module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire clknet_0_clk;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_1 _321_ (.A(net50),
    .X(_036_));
 sg13g2_buf_1 _322_ (.A(net42),
    .X(_037_));
 sg13g2_buf_1 _323_ (.A(_037_),
    .X(_038_));
 sg13g2_buf_1 _324_ (.A(\ctrl.state.out[2] ),
    .X(_039_));
 sg13g2_nor4_1 _325_ (.A(\dpath.a_lt_b$in1[7] ),
    .B(\dpath.a_lt_b$in1[6] ),
    .C(\dpath.a_lt_b$in1[5] ),
    .D(\dpath.a_lt_b$in1[0] ),
    .Y(_040_));
 sg13g2_nor4_1 _326_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(\dpath.a_lt_b$in1[3] ),
    .C(\dpath.a_lt_b$in1[2] ),
    .D(\dpath.a_lt_b$in1[1] ),
    .Y(_041_));
 sg13g2_nor4_1 _327_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(\dpath.a_lt_b$in1[14] ),
    .C(\dpath.a_lt_b$in1[13] ),
    .D(\dpath.a_lt_b$in1[8] ),
    .Y(_042_));
 sg13g2_buf_1 _328_ (.A(\dpath.a_lt_b$in1[9] ),
    .X(_043_));
 sg13g2_nor4_1 _329_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(\dpath.a_lt_b$in1[11] ),
    .C(\dpath.a_lt_b$in1[10] ),
    .D(net40),
    .Y(_044_));
 sg13g2_nand4_1 _330_ (.B(_041_),
    .C(_042_),
    .A(_040_),
    .Y(_045_),
    .D(_044_));
 sg13g2_a22oi_1 _331_ (.Y(_046_),
    .B1(net41),
    .B2(_045_),
    .A2(net47),
    .A1(net34));
 sg13g2_nor2_1 _332_ (.A(net48),
    .B(_046_),
    .Y(_002_));
 sg13g2_inv_1 _333_ (.Y(_047_),
    .A(net41));
 sg13g2_and3_1 _334_ (.X(net67),
    .A(_047_),
    .B(\ctrl.state.out[1] ),
    .C(_003_));
 sg13g2_nand2_1 _335_ (.Y(_048_),
    .A(net49),
    .B(net67));
 sg13g2_inv_1 _336_ (.Y(_049_),
    .A(net47));
 sg13g2_a21oi_1 _337_ (.A1(net34),
    .A2(_049_),
    .Y(_050_),
    .B1(net48));
 sg13g2_nand2_1 _338_ (.Y(_000_),
    .A(_048_),
    .B(_050_));
 sg13g2_buf_1 _339_ (.A(_047_),
    .X(_051_));
 sg13g2_nor2_1 _340_ (.A(net33),
    .B(_045_),
    .Y(_052_));
 sg13g2_a21oi_1 _341_ (.A1(\ctrl.state.out[1] ),
    .A2(_048_),
    .Y(_053_),
    .B1(_052_));
 sg13g2_nor2_1 _342_ (.A(net48),
    .B(_053_),
    .Y(_001_));
 sg13g2_xor2_1 _343_ (.B(\dpath.a_lt_b$in0[0] ),
    .A(\dpath.a_lt_b$in1[0] ),
    .X(net51));
 sg13g2_nand3b_1 _344_ (.B(net41),
    .C(_003_),
    .Y(_054_),
    .A_N(net50));
 sg13g2_inv_1 _345_ (.Y(_055_),
    .A(\dpath.a_lt_b$in0[0] ));
 sg13g2_xor2_1 _346_ (.B(\dpath.a_lt_b$in0[4] ),
    .A(\dpath.a_lt_b$in1[4] ),
    .X(_056_));
 sg13g2_xor2_1 _347_ (.B(\dpath.a_lt_b$in0[5] ),
    .A(\dpath.a_lt_b$in1[5] ),
    .X(_057_));
 sg13g2_nor2_1 _348_ (.A(_056_),
    .B(_057_),
    .Y(_058_));
 sg13g2_inv_1 _349_ (.Y(_059_),
    .A(\dpath.a_lt_b$in0[1] ));
 sg13g2_nor2b_1 _350_ (.A(\dpath.a_lt_b$in0[0] ),
    .B_N(\dpath.a_lt_b$in1[0] ),
    .Y(_060_));
 sg13g2_nand2_1 _351_ (.Y(_061_),
    .A(_059_),
    .B(_060_));
 sg13g2_o21ai_1 _352_ (.B1(\dpath.a_lt_b$in1[1] ),
    .Y(_062_),
    .A1(_059_),
    .A2(_060_));
 sg13g2_xor2_1 _353_ (.B(\dpath.a_lt_b$in0[2] ),
    .A(\dpath.a_lt_b$in1[2] ),
    .X(_063_));
 sg13g2_xor2_1 _354_ (.B(\dpath.a_lt_b$in0[3] ),
    .A(\dpath.a_lt_b$in1[3] ),
    .X(_064_));
 sg13g2_nor2_1 _355_ (.A(_063_),
    .B(_064_),
    .Y(_065_));
 sg13g2_nand4_1 _356_ (.B(_061_),
    .C(_062_),
    .A(_058_),
    .Y(_066_),
    .D(_065_));
 sg13g2_nor2b_1 _357_ (.A(\dpath.a_lt_b$in1[2] ),
    .B_N(\dpath.a_lt_b$in0[2] ),
    .Y(_067_));
 sg13g2_or2_1 _358_ (.X(_068_),
    .B(_067_),
    .A(\dpath.a_lt_b$in0[3] ));
 sg13g2_inv_1 _359_ (.Y(_069_),
    .A(\dpath.a_lt_b$in1[3] ));
 sg13g2_a21o_1 _360_ (.A2(_067_),
    .A1(\dpath.a_lt_b$in0[3] ),
    .B1(_069_),
    .X(_070_));
 sg13g2_nand3_1 _361_ (.B(_068_),
    .C(_070_),
    .A(_058_),
    .Y(_071_));
 sg13g2_nor2b_1 _362_ (.A(\dpath.a_lt_b$in1[7] ),
    .B_N(\dpath.a_lt_b$in0[7] ),
    .Y(_072_));
 sg13g2_inv_4 _363_ (.A(\dpath.a_lt_b$in0[5] ),
    .Y(_073_));
 sg13g2_nand2b_1 _364_ (.Y(_074_),
    .B(\dpath.a_lt_b$in0[4] ),
    .A_N(\dpath.a_lt_b$in1[4] ));
 sg13g2_nor2_1 _365_ (.A(_073_),
    .B(_074_),
    .Y(_075_));
 sg13g2_a21oi_1 _366_ (.A1(_073_),
    .A2(_074_),
    .Y(_076_),
    .B1(\dpath.a_lt_b$in1[5] ));
 sg13g2_nor4_1 _367_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(_072_),
    .C(_075_),
    .D(_076_),
    .Y(_077_));
 sg13g2_nand3_1 _368_ (.B(_071_),
    .C(_077_),
    .A(_066_),
    .Y(_078_));
 sg13g2_inv_1 _369_ (.Y(_079_),
    .A(\dpath.a_lt_b$in1[6] ));
 sg13g2_nor4_1 _370_ (.A(_079_),
    .B(_072_),
    .C(_075_),
    .D(_076_),
    .Y(_080_));
 sg13g2_nand3_1 _371_ (.B(_071_),
    .C(_080_),
    .A(_066_),
    .Y(_081_));
 sg13g2_nand2b_1 _372_ (.Y(_082_),
    .B(\dpath.a_lt_b$in1[6] ),
    .A_N(\dpath.a_lt_b$in0[6] ));
 sg13g2_nand2b_1 _373_ (.Y(_083_),
    .B(\dpath.a_lt_b$in1[7] ),
    .A_N(\dpath.a_lt_b$in0[7] ));
 sg13g2_o21ai_1 _374_ (.B1(_083_),
    .Y(_084_),
    .A1(_072_),
    .A2(_082_));
 sg13g2_inv_1 _375_ (.Y(_085_),
    .A(_084_));
 sg13g2_and3_1 _376_ (.X(_086_),
    .A(_078_),
    .B(_081_),
    .C(_085_));
 sg13g2_nand2b_2 _377_ (.Y(_087_),
    .B(\dpath.a_lt_b$in0[8] ),
    .A_N(\dpath.a_lt_b$in1[8] ));
 sg13g2_nand2b_1 _378_ (.Y(_088_),
    .B(\dpath.a_lt_b$in1[8] ),
    .A_N(\dpath.a_lt_b$in0[8] ));
 sg13g2_nand2_1 _379_ (.Y(_089_),
    .A(_087_),
    .B(_088_));
 sg13g2_xnor2_1 _380_ (.Y(_090_),
    .A(net40),
    .B(\dpath.a_lt_b$in0[9] ));
 sg13g2_buf_1 _381_ (.A(\dpath.a_lt_b$in0[11] ),
    .X(_091_));
 sg13g2_xnor2_1 _382_ (.Y(_092_),
    .A(\dpath.a_lt_b$in1[11] ),
    .B(_091_));
 sg13g2_xnor2_1 _383_ (.Y(_093_),
    .A(\dpath.a_lt_b$in1[10] ),
    .B(\dpath.a_lt_b$in0[10] ));
 sg13g2_nand3_1 _384_ (.B(_092_),
    .C(_093_),
    .A(_090_),
    .Y(_094_));
 sg13g2_nand2b_1 _385_ (.Y(_095_),
    .B(\dpath.a_lt_b$in0[12] ),
    .A_N(\dpath.a_lt_b$in1[12] ));
 sg13g2_nand2b_1 _386_ (.Y(_096_),
    .B(\dpath.a_lt_b$in1[12] ),
    .A_N(\dpath.a_lt_b$in0[12] ));
 sg13g2_and2_1 _387_ (.A(_095_),
    .B(_096_),
    .X(_097_));
 sg13g2_nand2b_2 _388_ (.Y(_098_),
    .B(_097_),
    .A_N(_094_));
 sg13g2_nand2b_1 _389_ (.Y(_099_),
    .B(\dpath.a_lt_b$in0[13] ),
    .A_N(\dpath.a_lt_b$in1[13] ));
 sg13g2_nand2b_1 _390_ (.Y(_100_),
    .B(\dpath.a_lt_b$in1[13] ),
    .A_N(\dpath.a_lt_b$in0[13] ));
 sg13g2_nand2_1 _391_ (.Y(_101_),
    .A(_099_),
    .B(_100_));
 sg13g2_nor3_1 _392_ (.A(_089_),
    .B(_098_),
    .C(_101_),
    .Y(_102_));
 sg13g2_nand2b_1 _393_ (.Y(_103_),
    .B(\dpath.a_lt_b$in0[15] ),
    .A_N(\dpath.a_lt_b$in1[15] ));
 sg13g2_nand2b_1 _394_ (.Y(_104_),
    .B(_103_),
    .A_N(\dpath.a_lt_b$in0[14] ));
 sg13g2_nand2_1 _395_ (.Y(_105_),
    .A(\dpath.a_lt_b$in1[14] ),
    .B(_103_));
 sg13g2_inv_1 _396_ (.Y(_106_),
    .A(\dpath.a_lt_b$in0[9] ));
 sg13g2_o21ai_1 _397_ (.B1(net40),
    .Y(_107_),
    .A1(_106_),
    .A2(_087_));
 sg13g2_inv_1 _398_ (.Y(_108_),
    .A(\dpath.a_lt_b$in0[10] ));
 sg13g2_inv_1 _399_ (.Y(_109_),
    .A(net39));
 sg13g2_a221oi_1 _400_ (.B2(_087_),
    .C1(_109_),
    .B1(_106_),
    .A1(\dpath.a_lt_b$in1[10] ),
    .Y(_110_),
    .A2(_108_));
 sg13g2_nand2b_1 _401_ (.Y(_111_),
    .B(\dpath.a_lt_b$in0[10] ),
    .A_N(\dpath.a_lt_b$in1[10] ));
 sg13g2_a21oi_1 _402_ (.A1(\dpath.a_lt_b$in1[11] ),
    .A2(_109_),
    .Y(_112_),
    .B1(_111_));
 sg13g2_a21oi_1 _403_ (.A1(_107_),
    .A2(_110_),
    .Y(_113_),
    .B1(_112_));
 sg13g2_inv_1 _404_ (.Y(_114_),
    .A(\dpath.a_lt_b$in1[11] ));
 sg13g2_a221oi_1 _405_ (.B2(_087_),
    .C1(\dpath.a_lt_b$in1[11] ),
    .B1(_106_),
    .A1(\dpath.a_lt_b$in1[10] ),
    .Y(_115_),
    .A2(_108_));
 sg13g2_a22oi_1 _406_ (.Y(_116_),
    .B1(_107_),
    .B2(_115_),
    .A2(net39),
    .A1(_114_));
 sg13g2_nand2_1 _407_ (.Y(_117_),
    .A(\dpath.a_lt_b$in0[12] ),
    .B(_100_));
 sg13g2_nand2b_1 _408_ (.Y(_118_),
    .B(_100_),
    .A_N(\dpath.a_lt_b$in1[12] ));
 sg13g2_a22oi_1 _409_ (.Y(_119_),
    .B1(_117_),
    .B2(_118_),
    .A2(_116_),
    .A1(_113_));
 sg13g2_nand2b_1 _410_ (.Y(_120_),
    .B(_100_),
    .A_N(_095_));
 sg13g2_nand3b_1 _411_ (.B(_120_),
    .C(_099_),
    .Y(_121_),
    .A_N(_119_));
 sg13g2_a221oi_1 _412_ (.B2(_105_),
    .C1(_121_),
    .B1(_104_),
    .A1(_086_),
    .Y(_122_),
    .A2(_102_));
 sg13g2_inv_1 _413_ (.Y(_123_),
    .A(\dpath.a_lt_b$in0[15] ));
 sg13g2_nor2_1 _414_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(_123_),
    .Y(_124_));
 sg13g2_nand2b_1 _415_ (.Y(_125_),
    .B(\dpath.a_lt_b$in1[14] ),
    .A_N(\dpath.a_lt_b$in0[14] ));
 sg13g2_nand2_1 _416_ (.Y(_126_),
    .A(\dpath.a_lt_b$in1[15] ),
    .B(_123_));
 sg13g2_o21ai_1 _417_ (.B1(_126_),
    .Y(_127_),
    .A1(_124_),
    .A2(_125_));
 sg13g2_nor3_1 _418_ (.A(_055_),
    .B(_122_),
    .C(_127_),
    .Y(_128_));
 sg13g2_xnor2_1 _419_ (.Y(_129_),
    .A(\dpath.a_lt_b$in1[0] ),
    .B(_128_));
 sg13g2_nor2_1 _420_ (.A(net42),
    .B(_055_),
    .Y(_130_));
 sg13g2_a22oi_1 _421_ (.Y(_131_),
    .B1(_130_),
    .B2(_051_),
    .A2(net8),
    .A1(_038_));
 sg13g2_o21ai_1 _422_ (.B1(_131_),
    .Y(_004_),
    .A1(_054_),
    .A2(_129_));
 sg13g2_nand4_1 _423_ (.B(_081_),
    .C(_085_),
    .A(_078_),
    .Y(_132_),
    .D(_088_));
 sg13g2_nand3_1 _424_ (.B(_087_),
    .C(_132_),
    .A(net40),
    .Y(_133_));
 sg13g2_a21oi_1 _425_ (.A1(_087_),
    .A2(_132_),
    .Y(_134_),
    .B1(net40));
 sg13g2_a21oi_1 _426_ (.A1(\dpath.a_lt_b$in0[9] ),
    .A2(_133_),
    .Y(_135_),
    .B1(_134_));
 sg13g2_xor2_1 _427_ (.B(_135_),
    .A(_093_),
    .X(_136_));
 sg13g2_inv_1 _428_ (.Y(_137_),
    .A(_003_));
 sg13g2_nor3_1 _429_ (.A(net50),
    .B(_047_),
    .C(_137_),
    .Y(_138_));
 sg13g2_nor2_2 _430_ (.A(_122_),
    .B(_127_),
    .Y(_139_));
 sg13g2_buf_1 _431_ (.A(_139_),
    .X(_140_));
 sg13g2_nand2_1 _432_ (.Y(_141_),
    .A(_138_),
    .B(net30));
 sg13g2_buf_1 _433_ (.A(net42),
    .X(_142_));
 sg13g2_or2_1 _434_ (.X(_143_),
    .B(_127_),
    .A(_122_));
 sg13g2_and2_1 _435_ (.A(\dpath.a_lt_b$in1[10] ),
    .B(net32),
    .X(_144_));
 sg13g2_buf_1 _436_ (.A(net42),
    .X(_145_));
 sg13g2_nor3_1 _437_ (.A(net36),
    .B(_108_),
    .C(net41),
    .Y(_146_));
 sg13g2_a221oi_1 _438_ (.B2(_144_),
    .C1(_146_),
    .B1(_143_),
    .A1(net37),
    .Y(_147_),
    .A2(net19));
 sg13g2_o21ai_1 _439_ (.B1(_147_),
    .Y(_005_),
    .A1(_136_),
    .A2(_141_));
 sg13g2_nand2_1 _440_ (.Y(_148_),
    .A(_114_),
    .B(net39));
 sg13g2_nor2b_1 _441_ (.A(\dpath.a_lt_b$in0[10] ),
    .B_N(\dpath.a_lt_b$in1[10] ),
    .Y(_149_));
 sg13g2_nand2b_1 _442_ (.Y(_150_),
    .B(\dpath.a_lt_b$in0[9] ),
    .A_N(net40));
 sg13g2_o21ai_1 _443_ (.B1(_111_),
    .Y(_151_),
    .A1(_149_),
    .A2(_150_));
 sg13g2_a221oi_1 _444_ (.B2(_132_),
    .C1(_149_),
    .B1(_087_),
    .A1(_043_),
    .Y(_152_),
    .A2(_106_));
 sg13g2_nor2_1 _445_ (.A(_151_),
    .B(_152_),
    .Y(_153_));
 sg13g2_or4_1 _446_ (.A(_054_),
    .B(_148_),
    .C(_143_),
    .D(_153_),
    .X(_154_));
 sg13g2_nor3_1 _447_ (.A(\dpath.a_lt_b$in1[11] ),
    .B(net39),
    .C(_054_),
    .Y(_155_));
 sg13g2_nand3_1 _448_ (.B(_153_),
    .C(_155_),
    .A(net30),
    .Y(_156_));
 sg13g2_nor2_1 _449_ (.A(net42),
    .B(_109_),
    .Y(_157_));
 sg13g2_a22oi_1 _450_ (.Y(_158_),
    .B1(_157_),
    .B2(_047_),
    .A2(net20),
    .A1(_036_));
 sg13g2_nor3_1 _451_ (.A(_114_),
    .B(net39),
    .C(_054_),
    .Y(_159_));
 sg13g2_o21ai_1 _452_ (.B1(_159_),
    .Y(_160_),
    .A1(_151_),
    .A2(_152_));
 sg13g2_nand3_1 _453_ (.B(net39),
    .C(_138_),
    .A(\dpath.a_lt_b$in1[11] ),
    .Y(_161_));
 sg13g2_or3_1 _454_ (.A(_151_),
    .B(_152_),
    .C(_161_),
    .X(_162_));
 sg13g2_nor2_1 _455_ (.A(_114_),
    .B(_054_),
    .Y(_163_));
 sg13g2_o21ai_1 _456_ (.B1(_163_),
    .Y(_164_),
    .A1(_122_),
    .A2(_127_));
 sg13g2_and4_1 _457_ (.A(_158_),
    .B(_160_),
    .C(_162_),
    .D(_164_),
    .X(_165_));
 sg13g2_nand3_1 _458_ (.B(_156_),
    .C(_165_),
    .A(_154_),
    .Y(_006_));
 sg13g2_buf_1 _459_ (.A(net32),
    .X(_166_));
 sg13g2_nor2_1 _460_ (.A(_094_),
    .B(_089_),
    .Y(_167_));
 sg13g2_nand2_1 _461_ (.Y(_168_),
    .A(_113_),
    .B(_116_));
 sg13g2_a21oi_1 _462_ (.A1(_086_),
    .A2(_167_),
    .Y(_169_),
    .B1(_168_));
 sg13g2_xnor2_1 _463_ (.Y(net54),
    .A(_169_),
    .B(_097_));
 sg13g2_mux2_1 _464_ (.A0(\dpath.a_lt_b$in1[12] ),
    .A1(net54),
    .S(net30),
    .X(_170_));
 sg13g2_inv_1 _465_ (.Y(_171_),
    .A(net21));
 sg13g2_buf_1 _466_ (.A(net42),
    .X(_172_));
 sg13g2_a21oi_1 _467_ (.A1(\dpath.a_lt_b$in0[12] ),
    .A2(net33),
    .Y(_173_),
    .B1(net35));
 sg13g2_a21oi_1 _468_ (.A1(net34),
    .A2(_171_),
    .Y(_174_),
    .B1(_173_));
 sg13g2_a21o_1 _469_ (.A2(_170_),
    .A1(net31),
    .B1(_174_),
    .X(_007_));
 sg13g2_and2_1 _470_ (.A(_087_),
    .B(_132_),
    .X(_175_));
 sg13g2_or3_1 _471_ (.A(_099_),
    .B(_098_),
    .C(_175_),
    .X(_176_));
 sg13g2_nor3_1 _472_ (.A(_054_),
    .B(_143_),
    .C(_176_),
    .Y(_177_));
 sg13g2_or3_1 _473_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(_098_),
    .C(_175_),
    .X(_178_));
 sg13g2_nand2_1 _474_ (.Y(_179_),
    .A(\dpath.a_lt_b$in1[13] ),
    .B(net32));
 sg13g2_a21oi_1 _475_ (.A1(_140_),
    .A2(_178_),
    .Y(_180_),
    .B1(_179_));
 sg13g2_nand2b_1 _476_ (.Y(_181_),
    .B(\dpath.a_lt_b$in0[13] ),
    .A_N(net42));
 sg13g2_nand2_1 _477_ (.Y(_182_),
    .A(net38),
    .B(net22));
 sg13g2_o21ai_1 _478_ (.B1(_182_),
    .Y(_183_),
    .A1(net41),
    .A2(_181_));
 sg13g2_and4_1 _479_ (.A(_078_),
    .B(_081_),
    .C(_085_),
    .D(_102_),
    .X(_184_));
 sg13g2_o21ai_1 _480_ (.B1(\dpath.a_lt_b$in0[14] ),
    .Y(_185_),
    .A1(_184_),
    .A2(_121_));
 sg13g2_nor3_1 _481_ (.A(\dpath.a_lt_b$in0[14] ),
    .B(_184_),
    .C(_121_),
    .Y(_186_));
 sg13g2_a21o_1 _482_ (.A2(_185_),
    .A1(\dpath.a_lt_b$in1[14] ),
    .B1(_186_),
    .X(_187_));
 sg13g2_a21oi_1 _483_ (.A1(net39),
    .A2(_151_),
    .Y(_188_),
    .B1(_114_));
 sg13g2_nor2_1 _484_ (.A(net39),
    .B(_151_),
    .Y(_189_));
 sg13g2_o21ai_1 _485_ (.B1(_095_),
    .Y(_190_),
    .A1(_188_),
    .A2(_189_));
 sg13g2_and2_1 _486_ (.A(_096_),
    .B(_190_),
    .X(_191_));
 sg13g2_nor2_1 _487_ (.A(_191_),
    .B(_101_),
    .Y(_192_));
 sg13g2_o21ai_1 _488_ (.B1(_192_),
    .Y(_193_),
    .A1(_098_),
    .A2(_175_));
 sg13g2_nand2_1 _489_ (.Y(_194_),
    .A(_191_),
    .B(_101_));
 sg13g2_nand2_1 _490_ (.Y(_195_),
    .A(net32),
    .B(_126_));
 sg13g2_a221oi_1 _491_ (.B2(_194_),
    .C1(_195_),
    .B1(_193_),
    .A1(_103_),
    .Y(_196_),
    .A2(_187_));
 sg13g2_or4_1 _492_ (.A(_177_),
    .B(_180_),
    .C(_183_),
    .D(_196_),
    .X(_008_));
 sg13g2_nor2_1 _493_ (.A(_184_),
    .B(_121_),
    .Y(_197_));
 sg13g2_xnor2_1 _494_ (.Y(_198_),
    .A(\dpath.a_lt_b$in1[14] ),
    .B(\dpath.a_lt_b$in0[14] ));
 sg13g2_xnor2_1 _495_ (.Y(net56),
    .A(_197_),
    .B(_198_));
 sg13g2_mux2_1 _496_ (.A0(\dpath.a_lt_b$in1[14] ),
    .A1(net56),
    .S(_140_),
    .X(_199_));
 sg13g2_inv_1 _497_ (.Y(_200_),
    .A(net24));
 sg13g2_a21oi_1 _498_ (.A1(\dpath.a_lt_b$in0[14] ),
    .A2(_051_),
    .Y(_201_),
    .B1(_172_));
 sg13g2_a21oi_1 _499_ (.A1(_038_),
    .A2(_200_),
    .Y(_202_),
    .B1(_201_));
 sg13g2_a21o_1 _500_ (.A2(_199_),
    .A1(_166_),
    .B1(_202_),
    .X(_009_));
 sg13g2_nand2_1 _501_ (.Y(_203_),
    .A(net32),
    .B(_124_));
 sg13g2_nand2_1 _502_ (.Y(_204_),
    .A(\dpath.a_lt_b$in1[15] ),
    .B(net32));
 sg13g2_mux2_1 _503_ (.A0(_203_),
    .A1(_204_),
    .S(_187_),
    .X(_205_));
 sg13g2_nor2b_1 _504_ (.A(\dpath.a_lt_b$in0[15] ),
    .B_N(\dpath.a_lt_b$in1[15] ),
    .Y(_206_));
 sg13g2_nor3_1 _505_ (.A(net36),
    .B(_123_),
    .C(net41),
    .Y(_207_));
 sg13g2_a221oi_1 _506_ (.B2(_206_),
    .C1(_207_),
    .B1(net32),
    .A1(net37),
    .Y(_208_),
    .A2(net25));
 sg13g2_nand2_1 _507_ (.Y(_010_),
    .A(_205_),
    .B(_208_));
 sg13g2_xnor2_1 _508_ (.Y(_209_),
    .A(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ));
 sg13g2_xnor2_1 _509_ (.Y(net58),
    .A(_060_),
    .B(_209_));
 sg13g2_mux2_1 _510_ (.A0(\dpath.a_lt_b$in1[1] ),
    .A1(net58),
    .S(net30),
    .X(_210_));
 sg13g2_nor3_1 _511_ (.A(net38),
    .B(_059_),
    .C(net41),
    .Y(_211_));
 sg13g2_a21o_1 _512_ (.A2(net9),
    .A1(net37),
    .B1(_211_),
    .X(_212_));
 sg13g2_a21o_1 _513_ (.A2(_210_),
    .A1(net31),
    .B1(_212_),
    .X(_011_));
 sg13g2_and2_1 _514_ (.A(_061_),
    .B(_062_),
    .X(_213_));
 sg13g2_xnor2_1 _515_ (.Y(net59),
    .A(_213_),
    .B(_063_));
 sg13g2_mux2_1 _516_ (.A0(\dpath.a_lt_b$in1[2] ),
    .A1(net59),
    .S(net30),
    .X(_214_));
 sg13g2_inv_1 _517_ (.Y(_215_),
    .A(net10));
 sg13g2_a21oi_1 _518_ (.A1(\dpath.a_lt_b$in0[2] ),
    .A2(net33),
    .Y(_216_),
    .B1(net35));
 sg13g2_a21oi_1 _519_ (.A1(net34),
    .A2(_215_),
    .Y(_217_),
    .B1(_216_));
 sg13g2_a21o_1 _520_ (.A2(_214_),
    .A1(net31),
    .B1(_217_),
    .X(_012_));
 sg13g2_inv_1 _521_ (.Y(_218_),
    .A(_213_));
 sg13g2_inv_1 _522_ (.Y(_219_),
    .A(\dpath.a_lt_b$in1[2] ));
 sg13g2_a21oi_1 _523_ (.A1(_219_),
    .A2(_213_),
    .Y(_220_),
    .B1(\dpath.a_lt_b$in0[2] ));
 sg13g2_a21oi_1 _524_ (.A1(\dpath.a_lt_b$in1[2] ),
    .A2(_218_),
    .Y(_221_),
    .B1(_220_));
 sg13g2_xnor2_1 _525_ (.Y(net60),
    .A(_064_),
    .B(_221_));
 sg13g2_mux2_1 _526_ (.A0(\dpath.a_lt_b$in1[3] ),
    .A1(net60),
    .S(net30),
    .X(_222_));
 sg13g2_inv_1 _527_ (.Y(_223_),
    .A(net11));
 sg13g2_a21oi_1 _528_ (.A1(\dpath.a_lt_b$in0[3] ),
    .A2(net33),
    .Y(_224_),
    .B1(net35));
 sg13g2_a21oi_1 _529_ (.A1(net34),
    .A2(_223_),
    .Y(_225_),
    .B1(_224_));
 sg13g2_a21o_1 _530_ (.A2(_222_),
    .A1(net31),
    .B1(_225_),
    .X(_013_));
 sg13g2_a22oi_1 _531_ (.Y(_226_),
    .B1(_213_),
    .B2(_065_),
    .A2(_070_),
    .A1(_068_));
 sg13g2_xor2_1 _532_ (.B(_226_),
    .A(_056_),
    .X(net61));
 sg13g2_mux2_1 _533_ (.A0(\dpath.a_lt_b$in1[4] ),
    .A1(net61),
    .S(net30),
    .X(_227_));
 sg13g2_inv_1 _534_ (.Y(_228_),
    .A(net13));
 sg13g2_a21oi_1 _535_ (.A1(\dpath.a_lt_b$in0[4] ),
    .A2(net33),
    .Y(_229_),
    .B1(net35));
 sg13g2_a21oi_1 _536_ (.A1(net34),
    .A2(_228_),
    .Y(_230_),
    .B1(_229_));
 sg13g2_a21o_1 _537_ (.A2(_227_),
    .A1(net31),
    .B1(_230_),
    .X(_014_));
 sg13g2_nand2_1 _538_ (.Y(_231_),
    .A(\dpath.a_lt_b$in1[4] ),
    .B(_226_));
 sg13g2_nor2_1 _539_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(_226_),
    .Y(_232_));
 sg13g2_a21oi_1 _540_ (.A1(\dpath.a_lt_b$in0[4] ),
    .A2(_231_),
    .Y(_233_),
    .B1(_232_));
 sg13g2_xor2_1 _541_ (.B(_233_),
    .A(_057_),
    .X(net62));
 sg13g2_mux2_1 _542_ (.A0(\dpath.a_lt_b$in1[5] ),
    .A1(net62),
    .S(net30),
    .X(_234_));
 sg13g2_nor3_1 _543_ (.A(net42),
    .B(_073_),
    .C(net41),
    .Y(_235_));
 sg13g2_a21o_1 _544_ (.A2(net14),
    .A1(net37),
    .B1(_235_),
    .X(_236_));
 sg13g2_a21o_1 _545_ (.A2(_234_),
    .A1(net31),
    .B1(_236_),
    .X(_015_));
 sg13g2_nor2_1 _546_ (.A(_075_),
    .B(_076_),
    .Y(_237_));
 sg13g2_and3_1 _547_ (.X(_238_),
    .A(_237_),
    .B(_066_),
    .C(_071_));
 sg13g2_xnor2_1 _548_ (.Y(_239_),
    .A(\dpath.a_lt_b$in1[6] ),
    .B(\dpath.a_lt_b$in0[6] ));
 sg13g2_xnor2_1 _549_ (.Y(net63),
    .A(_238_),
    .B(_239_));
 sg13g2_mux2_1 _550_ (.A0(\dpath.a_lt_b$in1[6] ),
    .A1(net63),
    .S(_139_),
    .X(_240_));
 sg13g2_inv_1 _551_ (.Y(_241_),
    .A(net15));
 sg13g2_a21oi_1 _552_ (.A1(\dpath.a_lt_b$in0[6] ),
    .A2(net33),
    .Y(_242_),
    .B1(net35));
 sg13g2_a21oi_1 _553_ (.A1(net34),
    .A2(_241_),
    .Y(_243_),
    .B1(_242_));
 sg13g2_a21o_1 _554_ (.A2(_240_),
    .A1(net31),
    .B1(_243_),
    .X(_016_));
 sg13g2_inv_1 _555_ (.Y(_244_),
    .A(\dpath.a_lt_b$in0[6] ));
 sg13g2_a21o_1 _556_ (.A2(_238_),
    .A1(_244_),
    .B1(\dpath.a_lt_b$in1[6] ),
    .X(_245_));
 sg13g2_o21ai_1 _557_ (.B1(_245_),
    .Y(_246_),
    .A1(_244_),
    .A2(_238_));
 sg13g2_nand2b_1 _558_ (.Y(_247_),
    .B(_083_),
    .A_N(_072_));
 sg13g2_xnor2_1 _559_ (.Y(net64),
    .A(_246_),
    .B(_247_));
 sg13g2_mux2_1 _560_ (.A0(\dpath.a_lt_b$in1[7] ),
    .A1(net64),
    .S(_139_),
    .X(_248_));
 sg13g2_inv_1 _561_ (.Y(_249_),
    .A(net16));
 sg13g2_a21oi_1 _562_ (.A1(\dpath.a_lt_b$in0[7] ),
    .A2(net33),
    .Y(_250_),
    .B1(net36));
 sg13g2_a21oi_1 _563_ (.A1(net34),
    .A2(_249_),
    .Y(_251_),
    .B1(_250_));
 sg13g2_a21o_1 _564_ (.A2(_248_),
    .A1(net31),
    .B1(_251_),
    .X(_017_));
 sg13g2_xnor2_1 _565_ (.Y(net65),
    .A(_086_),
    .B(_089_));
 sg13g2_mux2_1 _566_ (.A0(\dpath.a_lt_b$in1[8] ),
    .A1(net65),
    .S(_139_),
    .X(_252_));
 sg13g2_inv_1 _567_ (.Y(_253_),
    .A(net17));
 sg13g2_a21oi_1 _568_ (.A1(\dpath.a_lt_b$in0[8] ),
    .A2(net33),
    .Y(_254_),
    .B1(net36));
 sg13g2_a21oi_1 _569_ (.A1(net37),
    .A2(_253_),
    .Y(_255_),
    .B1(_254_));
 sg13g2_a21o_1 _570_ (.A2(_252_),
    .A1(_166_),
    .B1(_255_),
    .X(_018_));
 sg13g2_xnor2_1 _571_ (.Y(net66),
    .A(_090_),
    .B(_175_));
 sg13g2_mux2_1 _572_ (.A0(net40),
    .A1(net66),
    .S(_139_),
    .X(_256_));
 sg13g2_nor3_1 _573_ (.A(_036_),
    .B(_106_),
    .C(_039_),
    .Y(_257_));
 sg13g2_a21o_1 _574_ (.A2(net18),
    .A1(net35),
    .B1(_257_),
    .X(_258_));
 sg13g2_a21o_1 _575_ (.A2(_256_),
    .A1(net32),
    .B1(_258_),
    .X(_019_));
 sg13g2_a21o_1 _576_ (.A2(net1),
    .A1(_172_),
    .B1(_130_),
    .X(_259_));
 sg13g2_a21oi_2 _577_ (.B1(_137_),
    .Y(_260_),
    .A2(_143_),
    .A1(_039_));
 sg13g2_buf_8 _578_ (.A(_260_),
    .X(_261_));
 sg13g2_mux2_1 _579_ (.A0(_259_),
    .A1(\dpath.a_lt_b$in1[0] ),
    .S(net29),
    .X(_020_));
 sg13g2_nand2_1 _580_ (.Y(_262_),
    .A(net36),
    .B(net2));
 sg13g2_o21ai_1 _581_ (.B1(_262_),
    .Y(_263_),
    .A1(net37),
    .A2(_108_));
 sg13g2_mux2_1 _582_ (.A0(_263_),
    .A1(\dpath.a_lt_b$in1[10] ),
    .S(net29),
    .X(_021_));
 sg13g2_a21o_1 _583_ (.A2(net3),
    .A1(net35),
    .B1(_157_),
    .X(_264_));
 sg13g2_mux2_1 _584_ (.A0(_264_),
    .A1(\dpath.a_lt_b$in1[11] ),
    .S(net29),
    .X(_022_));
 sg13g2_mux2_1 _585_ (.A0(\dpath.a_lt_b$in0[12] ),
    .A1(net4),
    .S(_145_),
    .X(_265_));
 sg13g2_mux2_1 _586_ (.A0(_265_),
    .A1(\dpath.a_lt_b$in1[12] ),
    .S(net29),
    .X(_023_));
 sg13g2_nand2_1 _587_ (.Y(_266_),
    .A(net35),
    .B(net5));
 sg13g2_nand2_1 _588_ (.Y(_267_),
    .A(_181_),
    .B(_266_));
 sg13g2_mux2_1 _589_ (.A0(_267_),
    .A1(\dpath.a_lt_b$in1[13] ),
    .S(net29),
    .X(_024_));
 sg13g2_mux2_1 _590_ (.A0(\dpath.a_lt_b$in0[14] ),
    .A1(net6),
    .S(_037_),
    .X(_268_));
 sg13g2_mux2_1 _591_ (.A0(_268_),
    .A1(\dpath.a_lt_b$in1[14] ),
    .S(_261_),
    .X(_025_));
 sg13g2_nand2_1 _592_ (.Y(_269_),
    .A(net36),
    .B(net7));
 sg13g2_o21ai_1 _593_ (.B1(_269_),
    .Y(_270_),
    .A1(net37),
    .A2(_123_));
 sg13g2_mux2_1 _594_ (.A0(_270_),
    .A1(\dpath.a_lt_b$in1[15] ),
    .S(_261_),
    .X(_026_));
 sg13g2_nand2_1 _595_ (.Y(_271_),
    .A(net36),
    .B(net12));
 sg13g2_o21ai_1 _596_ (.B1(_271_),
    .Y(_272_),
    .A1(net37),
    .A2(_059_));
 sg13g2_mux2_1 _597_ (.A0(_272_),
    .A1(\dpath.a_lt_b$in1[1] ),
    .S(net29),
    .X(_027_));
 sg13g2_mux2_1 _598_ (.A0(\dpath.a_lt_b$in0[2] ),
    .A1(net23),
    .S(net38),
    .X(_273_));
 sg13g2_mux2_1 _599_ (.A0(_273_),
    .A1(\dpath.a_lt_b$in1[2] ),
    .S(net29),
    .X(_028_));
 sg13g2_mux2_1 _600_ (.A0(\dpath.a_lt_b$in0[3] ),
    .A1(net26),
    .S(net38),
    .X(_274_));
 sg13g2_mux2_1 _601_ (.A0(_274_),
    .A1(\dpath.a_lt_b$in1[3] ),
    .S(net29),
    .X(_029_));
 sg13g2_mux2_1 _602_ (.A0(\dpath.a_lt_b$in0[4] ),
    .A1(net27),
    .S(net38),
    .X(_275_));
 sg13g2_mux2_1 _603_ (.A0(_275_),
    .A1(\dpath.a_lt_b$in1[4] ),
    .S(_260_),
    .X(_030_));
 sg13g2_nand2_1 _604_ (.Y(_276_),
    .A(net36),
    .B(net28));
 sg13g2_o21ai_1 _605_ (.B1(_276_),
    .Y(_277_),
    .A1(_142_),
    .A2(_073_));
 sg13g2_mux2_1 _606_ (.A0(_277_),
    .A1(\dpath.a_lt_b$in1[5] ),
    .S(_260_),
    .X(_031_));
 sg13g2_mux2_1 _607_ (.A0(\dpath.a_lt_b$in0[6] ),
    .A1(net43),
    .S(net38),
    .X(_278_));
 sg13g2_mux2_1 _608_ (.A0(_278_),
    .A1(\dpath.a_lt_b$in1[6] ),
    .S(_260_),
    .X(_032_));
 sg13g2_mux2_1 _609_ (.A0(\dpath.a_lt_b$in0[7] ),
    .A1(net44),
    .S(net38),
    .X(_279_));
 sg13g2_mux2_1 _610_ (.A0(_279_),
    .A1(\dpath.a_lt_b$in1[7] ),
    .S(_260_),
    .X(_033_));
 sg13g2_mux2_1 _611_ (.A0(\dpath.a_lt_b$in0[8] ),
    .A1(net45),
    .S(net38),
    .X(_280_));
 sg13g2_mux2_1 _612_ (.A0(_280_),
    .A1(\dpath.a_lt_b$in1[8] ),
    .S(_260_),
    .X(_034_));
 sg13g2_nand2_1 _613_ (.Y(_281_),
    .A(_145_),
    .B(net46));
 sg13g2_o21ai_1 _614_ (.B1(_281_),
    .Y(_282_),
    .A1(_142_),
    .A2(_106_));
 sg13g2_mux2_1 _615_ (.A0(_282_),
    .A1(net40),
    .S(_260_),
    .X(_035_));
 sg13g2_inv_1 _616_ (.Y(net52),
    .A(_136_));
 sg13g2_xnor2_1 _617_ (.Y(net53),
    .A(_092_),
    .B(_153_));
 sg13g2_inv_1 _618_ (.Y(_283_),
    .A(_191_));
 sg13g2_o21ai_1 _619_ (.B1(_283_),
    .Y(_284_),
    .A1(_098_),
    .A2(_175_));
 sg13g2_xnor2_1 _620_ (.Y(net55),
    .A(_284_),
    .B(_101_));
 sg13g2_nor2_1 _621_ (.A(_124_),
    .B(_206_),
    .Y(_285_));
 sg13g2_xnor2_1 _622_ (.Y(net57),
    .A(_187_),
    .B(_285_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_dfrbp_1 \ctrl.state.out[0]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net68),
    .D(_000_),
    .Q_N(_003_),
    .Q(net50));
 sg13g2_dfrbp_1 \ctrl.state.out[1]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net69),
    .D(_001_),
    .Q_N(_319_),
    .Q(\ctrl.state.out[1] ));
 sg13g2_dfrbp_1 \ctrl.state.out[2]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net70),
    .D(_002_),
    .Q_N(_318_),
    .Q(\ctrl.state.out[2] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[0]$_DFFE_PP_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net71),
    .D(_004_),
    .Q_N(_317_),
    .Q(\dpath.a_lt_b$in0[0] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[10]$_DFFE_PP_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net72),
    .D(_005_),
    .Q_N(_316_),
    .Q(\dpath.a_lt_b$in0[10] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[11]$_DFFE_PP_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net73),
    .D(_006_),
    .Q_N(_315_),
    .Q(\dpath.a_lt_b$in0[11] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[12]$_DFFE_PP_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net74),
    .D(_007_),
    .Q_N(_314_),
    .Q(\dpath.a_lt_b$in0[12] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[13]$_DFFE_PP_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net75),
    .D(_008_),
    .Q_N(_313_),
    .Q(\dpath.a_lt_b$in0[13] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[14]$_DFFE_PP_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net76),
    .D(_009_),
    .Q_N(_312_),
    .Q(\dpath.a_lt_b$in0[14] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[15]$_DFFE_PP_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net77),
    .D(_010_),
    .Q_N(_311_),
    .Q(\dpath.a_lt_b$in0[15] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[1]$_DFFE_PP_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net78),
    .D(_011_),
    .Q_N(_310_),
    .Q(\dpath.a_lt_b$in0[1] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[2]$_DFFE_PP_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net79),
    .D(_012_),
    .Q_N(_309_),
    .Q(\dpath.a_lt_b$in0[2] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[3]$_DFFE_PP_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net80),
    .D(_013_),
    .Q_N(_308_),
    .Q(\dpath.a_lt_b$in0[3] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[4]$_DFFE_PP_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net81),
    .D(_014_),
    .Q_N(_307_),
    .Q(\dpath.a_lt_b$in0[4] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[5]$_DFFE_PP_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net82),
    .D(_015_),
    .Q_N(_306_),
    .Q(\dpath.a_lt_b$in0[5] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[6]$_DFFE_PP_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net83),
    .D(_016_),
    .Q_N(_305_),
    .Q(\dpath.a_lt_b$in0[6] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[7]$_DFFE_PP_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net84),
    .D(_017_),
    .Q_N(_304_),
    .Q(\dpath.a_lt_b$in0[7] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[8]$_DFFE_PP_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net85),
    .D(_018_),
    .Q_N(_303_),
    .Q(\dpath.a_lt_b$in0[8] ));
 sg13g2_dfrbp_1 \dpath.a_reg.out[9]$_DFFE_PP_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net86),
    .D(_019_),
    .Q_N(_302_),
    .Q(\dpath.a_lt_b$in0[9] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[0]$_DFFE_PP_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net87),
    .D(_020_),
    .Q_N(_301_),
    .Q(\dpath.a_lt_b$in1[0] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[10]$_DFFE_PP_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net88),
    .D(_021_),
    .Q_N(_300_),
    .Q(\dpath.a_lt_b$in1[10] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[11]$_DFFE_PP_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net89),
    .D(_022_),
    .Q_N(_299_),
    .Q(\dpath.a_lt_b$in1[11] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[12]$_DFFE_PP_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net90),
    .D(_023_),
    .Q_N(_298_),
    .Q(\dpath.a_lt_b$in1[12] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[13]$_DFFE_PP_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net91),
    .D(_024_),
    .Q_N(_297_),
    .Q(\dpath.a_lt_b$in1[13] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[14]$_DFFE_PP_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net92),
    .D(_025_),
    .Q_N(_296_),
    .Q(\dpath.a_lt_b$in1[14] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[15]$_DFFE_PP_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net93),
    .D(_026_),
    .Q_N(_295_),
    .Q(\dpath.a_lt_b$in1[15] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[1]$_DFFE_PP_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net94),
    .D(_027_),
    .Q_N(_294_),
    .Q(\dpath.a_lt_b$in1[1] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[2]$_DFFE_PP_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net95),
    .D(_028_),
    .Q_N(_293_),
    .Q(\dpath.a_lt_b$in1[2] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[3]$_DFFE_PP_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net96),
    .D(_029_),
    .Q_N(_292_),
    .Q(\dpath.a_lt_b$in1[3] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[4]$_DFFE_PP_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net97),
    .D(_030_),
    .Q_N(_291_),
    .Q(\dpath.a_lt_b$in1[4] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[5]$_DFFE_PP_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net98),
    .D(_031_),
    .Q_N(_290_),
    .Q(\dpath.a_lt_b$in1[5] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[6]$_DFFE_PP_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net99),
    .D(_032_),
    .Q_N(_289_),
    .Q(\dpath.a_lt_b$in1[6] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[7]$_DFFE_PP_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net100),
    .D(_033_),
    .Q_N(_288_),
    .Q(\dpath.a_lt_b$in1[7] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[8]$_DFFE_PP_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net101),
    .D(_034_),
    .Q_N(_287_),
    .Q(\dpath.a_lt_b$in1[8] ));
 sg13g2_dfrbp_1 \dpath.b_reg.out[9]$_DFFE_PP_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net102),
    .D(_035_),
    .Q_N(_286_),
    .Q(\dpath.a_lt_b$in1[9] ));
 sg13g2_buf_4 fanout29 (.X(net29),
    .A(_261_));
 sg13g2_buf_2 fanout30 (.A(_140_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_166_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_138_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_051_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_038_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_172_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_145_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_142_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_037_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_091_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_043_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_039_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_036_),
    .X(net42));
 sg13g2_buf_1 input1 (.A(req_msg[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(req_msg[10]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(req_msg[11]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(req_msg[12]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(req_msg[13]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(req_msg[14]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(req_msg[15]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(req_msg[16]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(req_msg[17]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(req_msg[18]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(req_msg[19]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(req_msg[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(req_msg[20]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(req_msg[21]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(req_msg[22]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(req_msg[23]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(req_msg[24]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(req_msg[25]),
    .X(net18));
 sg13g2_buf_1 input19 (.A(req_msg[26]),
    .X(net19));
 sg13g2_buf_1 input20 (.A(req_msg[27]),
    .X(net20));
 sg13g2_buf_1 input21 (.A(req_msg[28]),
    .X(net21));
 sg13g2_buf_1 input22 (.A(req_msg[29]),
    .X(net22));
 sg13g2_buf_1 input23 (.A(req_msg[2]),
    .X(net23));
 sg13g2_buf_1 input24 (.A(req_msg[30]),
    .X(net24));
 sg13g2_buf_1 input25 (.A(req_msg[31]),
    .X(net25));
 sg13g2_buf_1 input26 (.A(req_msg[3]),
    .X(net26));
 sg13g2_buf_1 input27 (.A(req_msg[4]),
    .X(net27));
 sg13g2_buf_1 input28 (.A(req_msg[5]),
    .X(net28));
 sg13g2_buf_1 input29 (.A(req_msg[6]),
    .X(net43));
 sg13g2_buf_1 input30 (.A(req_msg[7]),
    .X(net44));
 sg13g2_buf_1 input31 (.A(req_msg[8]),
    .X(net45));
 sg13g2_buf_1 input32 (.A(req_msg[9]),
    .X(net46));
 sg13g2_buf_1 input33 (.A(req_val),
    .X(net47));
 sg13g2_buf_1 input34 (.A(reset),
    .X(net48));
 sg13g2_buf_1 input35 (.A(resp_rdy),
    .X(net49));
 sg13g2_buf_1 output36 (.A(net50),
    .X(req_rdy));
 sg13g2_buf_1 output37 (.A(net51),
    .X(resp_msg[0]));
 sg13g2_buf_1 output38 (.A(net52),
    .X(resp_msg[10]));
 sg13g2_buf_1 output39 (.A(net53),
    .X(resp_msg[11]));
 sg13g2_buf_1 output40 (.A(net54),
    .X(resp_msg[12]));
 sg13g2_buf_1 output41 (.A(net55),
    .X(resp_msg[13]));
 sg13g2_buf_1 output42 (.A(net56),
    .X(resp_msg[14]));
 sg13g2_buf_1 output43 (.A(net57),
    .X(resp_msg[15]));
 sg13g2_buf_1 output44 (.A(net58),
    .X(resp_msg[1]));
 sg13g2_buf_1 output45 (.A(net59),
    .X(resp_msg[2]));
 sg13g2_buf_1 output46 (.A(net60),
    .X(resp_msg[3]));
 sg13g2_buf_1 output47 (.A(net61),
    .X(resp_msg[4]));
 sg13g2_buf_1 output48 (.A(net62),
    .X(resp_msg[5]));
 sg13g2_buf_1 output49 (.A(net63),
    .X(resp_msg[6]));
 sg13g2_buf_1 output50 (.A(net64),
    .X(resp_msg[7]));
 sg13g2_buf_1 output51 (.A(net65),
    .X(resp_msg[8]));
 sg13g2_buf_1 output52 (.A(net66),
    .X(resp_msg[9]));
 sg13g2_buf_1 output53 (.A(net67),
    .X(resp_val));
 sg13g2_tiehi \ctrl.state.out[0]$_DFF_P__54  (.L_HI(net68));
 sg13g2_tiehi \ctrl.state.out[1]$_DFF_P__55  (.L_HI(net69));
 sg13g2_tiehi \ctrl.state.out[2]$_DFF_P__56  (.L_HI(net70));
 sg13g2_tiehi \dpath.a_reg.out[0]$_DFFE_PP__57  (.L_HI(net71));
 sg13g2_tiehi \dpath.a_reg.out[10]$_DFFE_PP__58  (.L_HI(net72));
 sg13g2_tiehi \dpath.a_reg.out[11]$_DFFE_PP__59  (.L_HI(net73));
 sg13g2_tiehi \dpath.a_reg.out[12]$_DFFE_PP__60  (.L_HI(net74));
 sg13g2_tiehi \dpath.a_reg.out[13]$_DFFE_PP__61  (.L_HI(net75));
 sg13g2_tiehi \dpath.a_reg.out[14]$_DFFE_PP__62  (.L_HI(net76));
 sg13g2_tiehi \dpath.a_reg.out[15]$_DFFE_PP__63  (.L_HI(net77));
 sg13g2_tiehi \dpath.a_reg.out[1]$_DFFE_PP__64  (.L_HI(net78));
 sg13g2_tiehi \dpath.a_reg.out[2]$_DFFE_PP__65  (.L_HI(net79));
 sg13g2_tiehi \dpath.a_reg.out[3]$_DFFE_PP__66  (.L_HI(net80));
 sg13g2_tiehi \dpath.a_reg.out[4]$_DFFE_PP__67  (.L_HI(net81));
 sg13g2_tiehi \dpath.a_reg.out[5]$_DFFE_PP__68  (.L_HI(net82));
 sg13g2_tiehi \dpath.a_reg.out[6]$_DFFE_PP__69  (.L_HI(net83));
 sg13g2_tiehi \dpath.a_reg.out[7]$_DFFE_PP__70  (.L_HI(net84));
 sg13g2_tiehi \dpath.a_reg.out[8]$_DFFE_PP__71  (.L_HI(net85));
 sg13g2_tiehi \dpath.a_reg.out[9]$_DFFE_PP__72  (.L_HI(net86));
 sg13g2_tiehi \dpath.b_reg.out[0]$_DFFE_PP__73  (.L_HI(net87));
 sg13g2_tiehi \dpath.b_reg.out[10]$_DFFE_PP__74  (.L_HI(net88));
 sg13g2_tiehi \dpath.b_reg.out[11]$_DFFE_PP__75  (.L_HI(net89));
 sg13g2_tiehi \dpath.b_reg.out[12]$_DFFE_PP__76  (.L_HI(net90));
 sg13g2_tiehi \dpath.b_reg.out[13]$_DFFE_PP__77  (.L_HI(net91));
 sg13g2_tiehi \dpath.b_reg.out[14]$_DFFE_PP__78  (.L_HI(net92));
 sg13g2_tiehi \dpath.b_reg.out[15]$_DFFE_PP__79  (.L_HI(net93));
 sg13g2_tiehi \dpath.b_reg.out[1]$_DFFE_PP__80  (.L_HI(net94));
 sg13g2_tiehi \dpath.b_reg.out[2]$_DFFE_PP__81  (.L_HI(net95));
 sg13g2_tiehi \dpath.b_reg.out[3]$_DFFE_PP__82  (.L_HI(net96));
 sg13g2_tiehi \dpath.b_reg.out[4]$_DFFE_PP__83  (.L_HI(net97));
 sg13g2_tiehi \dpath.b_reg.out[5]$_DFFE_PP__84  (.L_HI(net98));
 sg13g2_tiehi \dpath.b_reg.out[6]$_DFFE_PP__85  (.L_HI(net99));
 sg13g2_tiehi \dpath.b_reg.out[7]$_DFFE_PP__86  (.L_HI(net100));
 sg13g2_tiehi \dpath.b_reg.out[8]$_DFFE_PP__87  (.L_HI(net101));
 sg13g2_tiehi \dpath.b_reg.out[9]$_DFFE_PP__88  (.L_HI(net102));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_4 FILLER_0_102 ();
 sg13g2_fill_1 FILLER_0_106 ();
 sg13g2_decap_4 FILLER_0_111 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_4 FILLER_0_130 ();
 sg13g2_decap_4 FILLER_0_138 ();
 sg13g2_decap_4 FILLER_0_146 ();
 sg13g2_decap_4 FILLER_0_154 ();
 sg13g2_fill_2 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_182 ();
 sg13g2_fill_2 FILLER_0_187 ();
 sg13g2_fill_2 FILLER_0_193 ();
 sg13g2_fill_1 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_fill_1 FILLER_0_326 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_4 FILLER_1_133 ();
 sg13g2_fill_1 FILLER_1_137 ();
 sg13g2_fill_1 FILLER_1_142 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_fill_1 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_173 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_208 ();
 sg13g2_decap_8 FILLER_1_215 ();
 sg13g2_decap_8 FILLER_1_222 ();
 sg13g2_decap_8 FILLER_1_229 ();
 sg13g2_decap_8 FILLER_1_236 ();
 sg13g2_decap_8 FILLER_1_243 ();
 sg13g2_decap_8 FILLER_1_250 ();
 sg13g2_decap_8 FILLER_1_257 ();
 sg13g2_decap_8 FILLER_1_264 ();
 sg13g2_decap_8 FILLER_1_271 ();
 sg13g2_decap_8 FILLER_1_278 ();
 sg13g2_decap_8 FILLER_1_285 ();
 sg13g2_decap_8 FILLER_1_292 ();
 sg13g2_decap_8 FILLER_1_299 ();
 sg13g2_decap_8 FILLER_1_306 ();
 sg13g2_decap_8 FILLER_1_313 ();
 sg13g2_decap_8 FILLER_1_320 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_4 FILLER_2_322 ();
 sg13g2_fill_1 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_4 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_4 FILLER_4_322 ();
 sg13g2_fill_1 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_4 FILLER_5_322 ();
 sg13g2_fill_1 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_4 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_4 FILLER_7_322 ();
 sg13g2_fill_1 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_4 FILLER_8_322 ();
 sg13g2_fill_1 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_4 FILLER_9_322 ();
 sg13g2_fill_1 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_4 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_decap_4 FILLER_10_122 ();
 sg13g2_decap_4 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_decap_8 FILLER_10_169 ();
 sg13g2_decap_4 FILLER_10_176 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_decap_8 FILLER_10_223 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_decap_8 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_251 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_4 FILLER_10_321 ();
 sg13g2_fill_2 FILLER_10_325 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_4 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_88 ();
 sg13g2_fill_1 FILLER_11_100 ();
 sg13g2_fill_1 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_229 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_271 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_121 ();
 sg13g2_fill_2 FILLER_12_145 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_fill_1 FILLER_12_165 ();
 sg13g2_fill_1 FILLER_12_176 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_201 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_fill_1 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_84 ();
 sg13g2_decap_4 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_124 ();
 sg13g2_fill_1 FILLER_13_128 ();
 sg13g2_fill_2 FILLER_13_159 ();
 sg13g2_fill_1 FILLER_13_175 ();
 sg13g2_fill_2 FILLER_13_202 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_244 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_decap_8 FILLER_13_279 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_314 ();
 sg13g2_decap_4 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_4 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_132 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_156 ();
 sg13g2_fill_2 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_16 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_4 FILLER_15_81 ();
 sg13g2_decap_4 FILLER_15_95 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_214 ();
 sg13g2_fill_2 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_fill_2 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_fill_1 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_fill_2 FILLER_16_200 ();
 sg13g2_decap_4 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_4 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_decap_4 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_fill_2 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_11 ();
 sg13g2_decap_8 FILLER_17_17 ();
 sg13g2_decap_8 FILLER_17_24 ();
 sg13g2_decap_8 FILLER_17_31 ();
 sg13g2_decap_8 FILLER_17_38 ();
 sg13g2_decap_8 FILLER_17_45 ();
 sg13g2_decap_8 FILLER_17_52 ();
 sg13g2_decap_8 FILLER_17_59 ();
 sg13g2_decap_8 FILLER_17_66 ();
 sg13g2_decap_8 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_80 ();
 sg13g2_fill_2 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_260 ();
 sg13g2_decap_8 FILLER_17_267 ();
 sg13g2_decap_4 FILLER_17_274 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_16 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_31 ();
 sg13g2_decap_8 FILLER_18_38 ();
 sg13g2_decap_8 FILLER_18_45 ();
 sg13g2_decap_8 FILLER_18_52 ();
 sg13g2_decap_8 FILLER_18_59 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_decap_8 FILLER_18_73 ();
 sg13g2_fill_2 FILLER_18_80 ();
 sg13g2_fill_1 FILLER_18_82 ();
 sg13g2_fill_1 FILLER_18_87 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_211 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_250 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_4 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_316 ();
 sg13g2_decap_4 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_4 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_4 FILLER_20_81 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_fill_2 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_4 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_25 ();
 sg13g2_decap_4 FILLER_21_30 ();
 sg13g2_fill_1 FILLER_21_34 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_4 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_decap_4 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_decap_4 FILLER_21_282 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_326 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_6 ();
 sg13g2_decap_4 FILLER_22_13 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_33 ();
 sg13g2_decap_8 FILLER_22_40 ();
 sg13g2_decap_8 FILLER_22_47 ();
 sg13g2_decap_8 FILLER_22_54 ();
 sg13g2_decap_8 FILLER_22_61 ();
 sg13g2_decap_8 FILLER_22_68 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_decap_8 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_fill_2 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_decap_4 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_153 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_164 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_272 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_4 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_15 ();
 sg13g2_decap_4 FILLER_25_22 ();
 sg13g2_decap_8 FILLER_25_30 ();
 sg13g2_decap_8 FILLER_25_37 ();
 sg13g2_decap_8 FILLER_25_44 ();
 sg13g2_decap_8 FILLER_25_51 ();
 sg13g2_decap_8 FILLER_25_58 ();
 sg13g2_decap_8 FILLER_25_65 ();
 sg13g2_decap_8 FILLER_25_72 ();
 sg13g2_decap_8 FILLER_25_79 ();
 sg13g2_decap_8 FILLER_25_86 ();
 sg13g2_decap_8 FILLER_25_93 ();
 sg13g2_decap_8 FILLER_25_104 ();
 sg13g2_fill_2 FILLER_25_111 ();
 sg13g2_fill_2 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_decap_8 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_fill_2 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_4 FILLER_26_321 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_decap_4 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_255 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_318 ();
 sg13g2_fill_2 FILLER_27_325 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_decap_8 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_decap_8 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_317 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_4 FILLER_29_112 ();
 sg13g2_decap_4 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_137 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_decap_8 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_306 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_decap_4 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_decap_4 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_227 ();
 sg13g2_decap_8 FILLER_30_234 ();
 sg13g2_decap_8 FILLER_30_241 ();
 sg13g2_decap_8 FILLER_30_248 ();
 sg13g2_decap_8 FILLER_30_255 ();
 sg13g2_decap_8 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_decap_8 FILLER_30_276 ();
 sg13g2_decap_8 FILLER_30_283 ();
 sg13g2_decap_8 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_4 FILLER_31_189 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_230 ();
 sg13g2_decap_8 FILLER_31_237 ();
 sg13g2_decap_8 FILLER_31_244 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_8 FILLER_31_258 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_314 ();
 sg13g2_decap_4 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_325 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_4 FILLER_32_322 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_4 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_4 FILLER_34_322 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_4 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_4 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_4 FILLER_37_322 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_4 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_140 ();
 sg13g2_fill_1 FILLER_39_142 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_4 FILLER_39_154 ();
 sg13g2_fill_2 FILLER_39_158 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_fill_2 FILLER_39_171 ();
 sg13g2_fill_1 FILLER_39_173 ();
 sg13g2_decap_8 FILLER_39_178 ();
 sg13g2_decap_8 FILLER_39_185 ();
 sg13g2_decap_8 FILLER_39_192 ();
 sg13g2_decap_8 FILLER_39_199 ();
 sg13g2_decap_8 FILLER_39_206 ();
 sg13g2_decap_8 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_227 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_decap_8 FILLER_39_241 ();
 sg13g2_decap_8 FILLER_39_248 ();
 sg13g2_decap_8 FILLER_39_255 ();
 sg13g2_decap_8 FILLER_39_262 ();
 sg13g2_decap_8 FILLER_39_269 ();
 sg13g2_decap_8 FILLER_39_276 ();
 sg13g2_decap_8 FILLER_39_283 ();
 sg13g2_decap_8 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_297 ();
 sg13g2_decap_8 FILLER_39_304 ();
 sg13g2_decap_8 FILLER_39_311 ();
 sg13g2_decap_8 FILLER_39_318 ();
 sg13g2_fill_2 FILLER_39_325 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_132 ();
 sg13g2_fill_1 FILLER_40_139 ();
 sg13g2_decap_8 FILLER_40_144 ();
 sg13g2_decap_8 FILLER_40_151 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_172 ();
 sg13g2_decap_8 FILLER_40_183 ();
 sg13g2_decap_8 FILLER_40_190 ();
 sg13g2_fill_1 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_206 ();
 sg13g2_fill_1 FILLER_40_208 ();
 sg13g2_fill_2 FILLER_40_213 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_decap_8 FILLER_40_233 ();
 sg13g2_decap_8 FILLER_40_240 ();
 sg13g2_decap_8 FILLER_40_247 ();
 sg13g2_decap_8 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_261 ();
 sg13g2_decap_8 FILLER_40_268 ();
 sg13g2_decap_8 FILLER_40_275 ();
 sg13g2_decap_8 FILLER_40_282 ();
 sg13g2_decap_8 FILLER_40_289 ();
 sg13g2_decap_8 FILLER_40_296 ();
 sg13g2_decap_8 FILLER_40_303 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_fill_2 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_326 ();
endmodule
