module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire net7;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire net291;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire net299;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire net308;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire net8;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire net356;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire net306;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire net437;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire clk_i_regs;
 wire \alu_adder_result_ex[0] ;
 wire \alu_adder_result_ex[10] ;
 wire \alu_adder_result_ex[11] ;
 wire \alu_adder_result_ex[12] ;
 wire \alu_adder_result_ex[13] ;
 wire \alu_adder_result_ex[14] ;
 wire \alu_adder_result_ex[15] ;
 wire \alu_adder_result_ex[16] ;
 wire \alu_adder_result_ex[17] ;
 wire \alu_adder_result_ex[18] ;
 wire \alu_adder_result_ex[19] ;
 wire \alu_adder_result_ex[1] ;
 wire \alu_adder_result_ex[20] ;
 wire \alu_adder_result_ex[21] ;
 wire \alu_adder_result_ex[22] ;
 wire \alu_adder_result_ex[23] ;
 wire \alu_adder_result_ex[24] ;
 wire \alu_adder_result_ex[25] ;
 wire \alu_adder_result_ex[26] ;
 wire \alu_adder_result_ex[27] ;
 wire \alu_adder_result_ex[28] ;
 wire \alu_adder_result_ex[29] ;
 wire \alu_adder_result_ex[2] ;
 wire \alu_adder_result_ex[30] ;
 wire net288;
 wire \alu_adder_result_ex[3] ;
 wire \alu_adder_result_ex[4] ;
 wire \alu_adder_result_ex[5] ;
 wire \alu_adder_result_ex[6] ;
 wire \alu_adder_result_ex[7] ;
 wire \alu_adder_result_ex[8] ;
 wire \alu_adder_result_ex[9] ;
 wire clk;
 wire core_busy_d;
 wire core_busy_q;
 wire \core_clock_gate_i.en_latch ;
 wire net146;
 wire \cs_registers_i.csr_depc_o[10] ;
 wire \cs_registers_i.csr_depc_o[11] ;
 wire \cs_registers_i.csr_depc_o[12] ;
 wire \cs_registers_i.csr_depc_o[13] ;
 wire \cs_registers_i.csr_depc_o[14] ;
 wire \cs_registers_i.csr_depc_o[15] ;
 wire \cs_registers_i.csr_depc_o[16] ;
 wire \cs_registers_i.csr_depc_o[17] ;
 wire \cs_registers_i.csr_depc_o[18] ;
 wire \cs_registers_i.csr_depc_o[19] ;
 wire \cs_registers_i.csr_depc_o[1] ;
 wire \cs_registers_i.csr_depc_o[20] ;
 wire \cs_registers_i.csr_depc_o[21] ;
 wire \cs_registers_i.csr_depc_o[22] ;
 wire \cs_registers_i.csr_depc_o[23] ;
 wire \cs_registers_i.csr_depc_o[24] ;
 wire \cs_registers_i.csr_depc_o[25] ;
 wire \cs_registers_i.csr_depc_o[26] ;
 wire \cs_registers_i.csr_depc_o[27] ;
 wire \cs_registers_i.csr_depc_o[28] ;
 wire \cs_registers_i.csr_depc_o[29] ;
 wire \cs_registers_i.csr_depc_o[2] ;
 wire \cs_registers_i.csr_depc_o[30] ;
 wire \cs_registers_i.csr_depc_o[31] ;
 wire \cs_registers_i.csr_depc_o[3] ;
 wire \cs_registers_i.csr_depc_o[4] ;
 wire \cs_registers_i.csr_depc_o[5] ;
 wire \cs_registers_i.csr_depc_o[6] ;
 wire \cs_registers_i.csr_depc_o[7] ;
 wire \cs_registers_i.csr_depc_o[8] ;
 wire \cs_registers_i.csr_depc_o[9] ;
 wire \cs_registers_i.csr_mepc_o[0] ;
 wire \cs_registers_i.csr_mepc_o[10] ;
 wire \cs_registers_i.csr_mepc_o[11] ;
 wire \cs_registers_i.csr_mepc_o[12] ;
 wire \cs_registers_i.csr_mepc_o[13] ;
 wire \cs_registers_i.csr_mepc_o[14] ;
 wire \cs_registers_i.csr_mepc_o[15] ;
 wire \cs_registers_i.csr_mepc_o[16] ;
 wire \cs_registers_i.csr_mepc_o[17] ;
 wire \cs_registers_i.csr_mepc_o[18] ;
 wire \cs_registers_i.csr_mepc_o[19] ;
 wire \cs_registers_i.csr_mepc_o[1] ;
 wire \cs_registers_i.csr_mepc_o[20] ;
 wire \cs_registers_i.csr_mepc_o[21] ;
 wire \cs_registers_i.csr_mepc_o[22] ;
 wire \cs_registers_i.csr_mepc_o[23] ;
 wire \cs_registers_i.csr_mepc_o[24] ;
 wire \cs_registers_i.csr_mepc_o[25] ;
 wire \cs_registers_i.csr_mepc_o[26] ;
 wire \cs_registers_i.csr_mepc_o[27] ;
 wire \cs_registers_i.csr_mepc_o[28] ;
 wire \cs_registers_i.csr_mepc_o[29] ;
 wire \cs_registers_i.csr_mepc_o[2] ;
 wire \cs_registers_i.csr_mepc_o[30] ;
 wire \cs_registers_i.csr_mepc_o[31] ;
 wire \cs_registers_i.csr_mepc_o[3] ;
 wire \cs_registers_i.csr_mepc_o[4] ;
 wire \cs_registers_i.csr_mepc_o[5] ;
 wire \cs_registers_i.csr_mepc_o[6] ;
 wire \cs_registers_i.csr_mepc_o[7] ;
 wire \cs_registers_i.csr_mepc_o[8] ;
 wire \cs_registers_i.csr_mepc_o[9] ;
 wire \cs_registers_i.csr_mstatus_mie_o ;
 wire \cs_registers_i.csr_mstatus_tw_o ;
 wire \cs_registers_i.csr_mtvec_o[10] ;
 wire \cs_registers_i.csr_mtvec_o[11] ;
 wire \cs_registers_i.csr_mtvec_o[12] ;
 wire \cs_registers_i.csr_mtvec_o[13] ;
 wire \cs_registers_i.csr_mtvec_o[14] ;
 wire \cs_registers_i.csr_mtvec_o[15] ;
 wire \cs_registers_i.csr_mtvec_o[16] ;
 wire \cs_registers_i.csr_mtvec_o[17] ;
 wire \cs_registers_i.csr_mtvec_o[18] ;
 wire \cs_registers_i.csr_mtvec_o[19] ;
 wire \cs_registers_i.csr_mtvec_o[20] ;
 wire \cs_registers_i.csr_mtvec_o[21] ;
 wire \cs_registers_i.csr_mtvec_o[22] ;
 wire \cs_registers_i.csr_mtvec_o[23] ;
 wire \cs_registers_i.csr_mtvec_o[24] ;
 wire \cs_registers_i.csr_mtvec_o[25] ;
 wire \cs_registers_i.csr_mtvec_o[26] ;
 wire \cs_registers_i.csr_mtvec_o[27] ;
 wire \cs_registers_i.csr_mtvec_o[28] ;
 wire \cs_registers_i.csr_mtvec_o[29] ;
 wire \cs_registers_i.csr_mtvec_o[30] ;
 wire \cs_registers_i.csr_mtvec_o[31] ;
 wire \cs_registers_i.csr_mtvec_o[8] ;
 wire \cs_registers_i.csr_mtvec_o[9] ;
 wire \cs_registers_i.dcsr_q[0] ;
 wire \cs_registers_i.dcsr_q[11] ;
 wire \cs_registers_i.dcsr_q[12] ;
 wire \cs_registers_i.dcsr_q[13] ;
 wire \cs_registers_i.dcsr_q[15] ;
 wire \cs_registers_i.dcsr_q[1] ;
 wire \cs_registers_i.dcsr_q[2] ;
 wire \cs_registers_i.dcsr_q[6] ;
 wire \cs_registers_i.dcsr_q[7] ;
 wire \cs_registers_i.dcsr_q[8] ;
 wire \cs_registers_i.debug_mode_i ;
 wire \cs_registers_i.dscratch0_q[0] ;
 wire \cs_registers_i.dscratch0_q[10] ;
 wire \cs_registers_i.dscratch0_q[11] ;
 wire \cs_registers_i.dscratch0_q[12] ;
 wire \cs_registers_i.dscratch0_q[13] ;
 wire \cs_registers_i.dscratch0_q[14] ;
 wire \cs_registers_i.dscratch0_q[15] ;
 wire \cs_registers_i.dscratch0_q[16] ;
 wire \cs_registers_i.dscratch0_q[17] ;
 wire \cs_registers_i.dscratch0_q[18] ;
 wire \cs_registers_i.dscratch0_q[19] ;
 wire \cs_registers_i.dscratch0_q[1] ;
 wire \cs_registers_i.dscratch0_q[20] ;
 wire \cs_registers_i.dscratch0_q[21] ;
 wire \cs_registers_i.dscratch0_q[22] ;
 wire \cs_registers_i.dscratch0_q[23] ;
 wire \cs_registers_i.dscratch0_q[24] ;
 wire \cs_registers_i.dscratch0_q[25] ;
 wire \cs_registers_i.dscratch0_q[26] ;
 wire \cs_registers_i.dscratch0_q[27] ;
 wire \cs_registers_i.dscratch0_q[28] ;
 wire \cs_registers_i.dscratch0_q[29] ;
 wire \cs_registers_i.dscratch0_q[2] ;
 wire \cs_registers_i.dscratch0_q[30] ;
 wire \cs_registers_i.dscratch0_q[31] ;
 wire \cs_registers_i.dscratch0_q[3] ;
 wire \cs_registers_i.dscratch0_q[4] ;
 wire \cs_registers_i.dscratch0_q[5] ;
 wire \cs_registers_i.dscratch0_q[6] ;
 wire \cs_registers_i.dscratch0_q[7] ;
 wire \cs_registers_i.dscratch0_q[8] ;
 wire \cs_registers_i.dscratch0_q[9] ;
 wire \cs_registers_i.dscratch1_q[0] ;
 wire \cs_registers_i.dscratch1_q[10] ;
 wire \cs_registers_i.dscratch1_q[11] ;
 wire \cs_registers_i.dscratch1_q[12] ;
 wire \cs_registers_i.dscratch1_q[13] ;
 wire \cs_registers_i.dscratch1_q[14] ;
 wire \cs_registers_i.dscratch1_q[15] ;
 wire \cs_registers_i.dscratch1_q[16] ;
 wire \cs_registers_i.dscratch1_q[17] ;
 wire \cs_registers_i.dscratch1_q[18] ;
 wire \cs_registers_i.dscratch1_q[19] ;
 wire \cs_registers_i.dscratch1_q[1] ;
 wire \cs_registers_i.dscratch1_q[20] ;
 wire \cs_registers_i.dscratch1_q[21] ;
 wire \cs_registers_i.dscratch1_q[22] ;
 wire \cs_registers_i.dscratch1_q[23] ;
 wire \cs_registers_i.dscratch1_q[24] ;
 wire \cs_registers_i.dscratch1_q[25] ;
 wire \cs_registers_i.dscratch1_q[26] ;
 wire \cs_registers_i.dscratch1_q[27] ;
 wire \cs_registers_i.dscratch1_q[28] ;
 wire \cs_registers_i.dscratch1_q[29] ;
 wire \cs_registers_i.dscratch1_q[2] ;
 wire \cs_registers_i.dscratch1_q[30] ;
 wire \cs_registers_i.dscratch1_q[31] ;
 wire \cs_registers_i.dscratch1_q[3] ;
 wire \cs_registers_i.dscratch1_q[4] ;
 wire \cs_registers_i.dscratch1_q[5] ;
 wire \cs_registers_i.dscratch1_q[6] ;
 wire \cs_registers_i.dscratch1_q[7] ;
 wire \cs_registers_i.dscratch1_q[8] ;
 wire \cs_registers_i.dscratch1_q[9] ;
 wire \cs_registers_i.mcause_q[0] ;
 wire \cs_registers_i.mcause_q[1] ;
 wire \cs_registers_i.mcause_q[2] ;
 wire \cs_registers_i.mcause_q[3] ;
 wire \cs_registers_i.mcause_q[4] ;
 wire \cs_registers_i.mcause_q[5] ;
 wire \cs_registers_i.mcountinhibit[0] ;
 wire \cs_registers_i.mcountinhibit[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter[11] ;
 wire \cs_registers_i.mcycle_counter_i.counter[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter[13] ;
 wire \cs_registers_i.mcycle_counter_i.counter[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter[15] ;
 wire \cs_registers_i.mcycle_counter_i.counter[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter[17] ;
 wire \cs_registers_i.mcycle_counter_i.counter[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter[19] ;
 wire \cs_registers_i.mcycle_counter_i.counter[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter[21] ;
 wire \cs_registers_i.mcycle_counter_i.counter[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter[23] ;
 wire \cs_registers_i.mcycle_counter_i.counter[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter[25] ;
 wire \cs_registers_i.mcycle_counter_i.counter[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter[27] ;
 wire \cs_registers_i.mcycle_counter_i.counter[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter[29] ;
 wire \cs_registers_i.mcycle_counter_i.counter[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter[31] ;
 wire \cs_registers_i.mcycle_counter_i.counter[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter[33] ;
 wire \cs_registers_i.mcycle_counter_i.counter[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter[35] ;
 wire \cs_registers_i.mcycle_counter_i.counter[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter[37] ;
 wire \cs_registers_i.mcycle_counter_i.counter[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter[39] ;
 wire \cs_registers_i.mcycle_counter_i.counter[3] ;
 wire \cs_registers_i.mcycle_counter_i.counter[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter[41] ;
 wire \cs_registers_i.mcycle_counter_i.counter[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter[43] ;
 wire \cs_registers_i.mcycle_counter_i.counter[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter[45] ;
 wire \cs_registers_i.mcycle_counter_i.counter[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter[47] ;
 wire \cs_registers_i.mcycle_counter_i.counter[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter[49] ;
 wire \cs_registers_i.mcycle_counter_i.counter[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter[51] ;
 wire \cs_registers_i.mcycle_counter_i.counter[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter[53] ;
 wire \cs_registers_i.mcycle_counter_i.counter[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter[55] ;
 wire \cs_registers_i.mcycle_counter_i.counter[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter[57] ;
 wire \cs_registers_i.mcycle_counter_i.counter[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter[59] ;
 wire \cs_registers_i.mcycle_counter_i.counter[5] ;
 wire \cs_registers_i.mcycle_counter_i.counter[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter[61] ;
 wire \cs_registers_i.mcycle_counter_i.counter[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter[63] ;
 wire \cs_registers_i.mcycle_counter_i.counter[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter[7] ;
 wire \cs_registers_i.mcycle_counter_i.counter[8] ;
 wire \cs_registers_i.mcycle_counter_i.counter[9] ;
 wire \cs_registers_i.mhpmcounter[2][0] ;
 wire \cs_registers_i.mhpmcounter[2][10] ;
 wire \cs_registers_i.mhpmcounter[2][11] ;
 wire \cs_registers_i.mhpmcounter[2][12] ;
 wire \cs_registers_i.mhpmcounter[2][13] ;
 wire \cs_registers_i.mhpmcounter[2][14] ;
 wire \cs_registers_i.mhpmcounter[2][15] ;
 wire \cs_registers_i.mhpmcounter[2][16] ;
 wire \cs_registers_i.mhpmcounter[2][17] ;
 wire \cs_registers_i.mhpmcounter[2][18] ;
 wire \cs_registers_i.mhpmcounter[2][19] ;
 wire \cs_registers_i.mhpmcounter[2][1] ;
 wire \cs_registers_i.mhpmcounter[2][20] ;
 wire \cs_registers_i.mhpmcounter[2][21] ;
 wire \cs_registers_i.mhpmcounter[2][22] ;
 wire \cs_registers_i.mhpmcounter[2][23] ;
 wire \cs_registers_i.mhpmcounter[2][24] ;
 wire \cs_registers_i.mhpmcounter[2][25] ;
 wire \cs_registers_i.mhpmcounter[2][26] ;
 wire \cs_registers_i.mhpmcounter[2][27] ;
 wire \cs_registers_i.mhpmcounter[2][28] ;
 wire \cs_registers_i.mhpmcounter[2][29] ;
 wire \cs_registers_i.mhpmcounter[2][2] ;
 wire \cs_registers_i.mhpmcounter[2][30] ;
 wire \cs_registers_i.mhpmcounter[2][31] ;
 wire \cs_registers_i.mhpmcounter[2][32] ;
 wire \cs_registers_i.mhpmcounter[2][33] ;
 wire \cs_registers_i.mhpmcounter[2][34] ;
 wire \cs_registers_i.mhpmcounter[2][35] ;
 wire \cs_registers_i.mhpmcounter[2][36] ;
 wire \cs_registers_i.mhpmcounter[2][37] ;
 wire \cs_registers_i.mhpmcounter[2][38] ;
 wire \cs_registers_i.mhpmcounter[2][39] ;
 wire \cs_registers_i.mhpmcounter[2][3] ;
 wire \cs_registers_i.mhpmcounter[2][40] ;
 wire \cs_registers_i.mhpmcounter[2][41] ;
 wire \cs_registers_i.mhpmcounter[2][42] ;
 wire \cs_registers_i.mhpmcounter[2][43] ;
 wire \cs_registers_i.mhpmcounter[2][44] ;
 wire \cs_registers_i.mhpmcounter[2][45] ;
 wire \cs_registers_i.mhpmcounter[2][46] ;
 wire \cs_registers_i.mhpmcounter[2][47] ;
 wire \cs_registers_i.mhpmcounter[2][48] ;
 wire \cs_registers_i.mhpmcounter[2][49] ;
 wire \cs_registers_i.mhpmcounter[2][4] ;
 wire \cs_registers_i.mhpmcounter[2][50] ;
 wire \cs_registers_i.mhpmcounter[2][51] ;
 wire \cs_registers_i.mhpmcounter[2][52] ;
 wire \cs_registers_i.mhpmcounter[2][53] ;
 wire \cs_registers_i.mhpmcounter[2][54] ;
 wire \cs_registers_i.mhpmcounter[2][55] ;
 wire \cs_registers_i.mhpmcounter[2][56] ;
 wire \cs_registers_i.mhpmcounter[2][57] ;
 wire \cs_registers_i.mhpmcounter[2][58] ;
 wire \cs_registers_i.mhpmcounter[2][59] ;
 wire \cs_registers_i.mhpmcounter[2][5] ;
 wire \cs_registers_i.mhpmcounter[2][60] ;
 wire \cs_registers_i.mhpmcounter[2][61] ;
 wire \cs_registers_i.mhpmcounter[2][62] ;
 wire \cs_registers_i.mhpmcounter[2][63] ;
 wire \cs_registers_i.mhpmcounter[2][6] ;
 wire \cs_registers_i.mhpmcounter[2][7] ;
 wire \cs_registers_i.mhpmcounter[2][8] ;
 wire \cs_registers_i.mhpmcounter[2][9] ;
 wire \cs_registers_i.mie_q[0] ;
 wire \cs_registers_i.mie_q[10] ;
 wire \cs_registers_i.mie_q[11] ;
 wire \cs_registers_i.mie_q[12] ;
 wire \cs_registers_i.mie_q[13] ;
 wire \cs_registers_i.mie_q[14] ;
 wire \cs_registers_i.mie_q[15] ;
 wire \cs_registers_i.mie_q[16] ;
 wire \cs_registers_i.mie_q[17] ;
 wire \cs_registers_i.mie_q[1] ;
 wire \cs_registers_i.mie_q[2] ;
 wire \cs_registers_i.mie_q[3] ;
 wire \cs_registers_i.mie_q[4] ;
 wire \cs_registers_i.mie_q[5] ;
 wire \cs_registers_i.mie_q[6] ;
 wire \cs_registers_i.mie_q[7] ;
 wire \cs_registers_i.mie_q[8] ;
 wire \cs_registers_i.mie_q[9] ;
 wire \cs_registers_i.mscratch_q[0] ;
 wire \cs_registers_i.mscratch_q[10] ;
 wire \cs_registers_i.mscratch_q[11] ;
 wire \cs_registers_i.mscratch_q[12] ;
 wire \cs_registers_i.mscratch_q[13] ;
 wire \cs_registers_i.mscratch_q[14] ;
 wire \cs_registers_i.mscratch_q[15] ;
 wire \cs_registers_i.mscratch_q[16] ;
 wire \cs_registers_i.mscratch_q[17] ;
 wire \cs_registers_i.mscratch_q[18] ;
 wire \cs_registers_i.mscratch_q[19] ;
 wire \cs_registers_i.mscratch_q[1] ;
 wire \cs_registers_i.mscratch_q[20] ;
 wire \cs_registers_i.mscratch_q[21] ;
 wire \cs_registers_i.mscratch_q[22] ;
 wire \cs_registers_i.mscratch_q[23] ;
 wire \cs_registers_i.mscratch_q[24] ;
 wire \cs_registers_i.mscratch_q[25] ;
 wire \cs_registers_i.mscratch_q[26] ;
 wire \cs_registers_i.mscratch_q[27] ;
 wire \cs_registers_i.mscratch_q[28] ;
 wire \cs_registers_i.mscratch_q[29] ;
 wire \cs_registers_i.mscratch_q[2] ;
 wire \cs_registers_i.mscratch_q[30] ;
 wire \cs_registers_i.mscratch_q[31] ;
 wire \cs_registers_i.mscratch_q[3] ;
 wire \cs_registers_i.mscratch_q[4] ;
 wire \cs_registers_i.mscratch_q[5] ;
 wire \cs_registers_i.mscratch_q[6] ;
 wire \cs_registers_i.mscratch_q[7] ;
 wire \cs_registers_i.mscratch_q[8] ;
 wire \cs_registers_i.mscratch_q[9] ;
 wire \cs_registers_i.mstack_cause_q[0] ;
 wire \cs_registers_i.mstack_cause_q[1] ;
 wire \cs_registers_i.mstack_cause_q[2] ;
 wire \cs_registers_i.mstack_cause_q[3] ;
 wire \cs_registers_i.mstack_cause_q[4] ;
 wire \cs_registers_i.mstack_cause_q[5] ;
 wire \cs_registers_i.mstack_d[0] ;
 wire \cs_registers_i.mstack_d[1] ;
 wire \cs_registers_i.mstack_d[2] ;
 wire \cs_registers_i.mstack_epc_q[0] ;
 wire \cs_registers_i.mstack_epc_q[10] ;
 wire \cs_registers_i.mstack_epc_q[11] ;
 wire \cs_registers_i.mstack_epc_q[12] ;
 wire \cs_registers_i.mstack_epc_q[13] ;
 wire \cs_registers_i.mstack_epc_q[14] ;
 wire \cs_registers_i.mstack_epc_q[15] ;
 wire \cs_registers_i.mstack_epc_q[16] ;
 wire \cs_registers_i.mstack_epc_q[17] ;
 wire \cs_registers_i.mstack_epc_q[18] ;
 wire \cs_registers_i.mstack_epc_q[19] ;
 wire \cs_registers_i.mstack_epc_q[1] ;
 wire \cs_registers_i.mstack_epc_q[20] ;
 wire \cs_registers_i.mstack_epc_q[21] ;
 wire \cs_registers_i.mstack_epc_q[22] ;
 wire \cs_registers_i.mstack_epc_q[23] ;
 wire \cs_registers_i.mstack_epc_q[24] ;
 wire \cs_registers_i.mstack_epc_q[25] ;
 wire \cs_registers_i.mstack_epc_q[26] ;
 wire \cs_registers_i.mstack_epc_q[27] ;
 wire \cs_registers_i.mstack_epc_q[28] ;
 wire \cs_registers_i.mstack_epc_q[29] ;
 wire \cs_registers_i.mstack_epc_q[2] ;
 wire \cs_registers_i.mstack_epc_q[30] ;
 wire \cs_registers_i.mstack_epc_q[31] ;
 wire \cs_registers_i.mstack_epc_q[3] ;
 wire \cs_registers_i.mstack_epc_q[4] ;
 wire \cs_registers_i.mstack_epc_q[5] ;
 wire \cs_registers_i.mstack_epc_q[6] ;
 wire \cs_registers_i.mstack_epc_q[7] ;
 wire \cs_registers_i.mstack_epc_q[8] ;
 wire \cs_registers_i.mstack_epc_q[9] ;
 wire \cs_registers_i.mstack_q[0] ;
 wire \cs_registers_i.mstack_q[1] ;
 wire \cs_registers_i.mstack_q[2] ;
 wire \cs_registers_i.mstatus_q[1] ;
 wire \cs_registers_i.mtval_q[0] ;
 wire \cs_registers_i.mtval_q[10] ;
 wire \cs_registers_i.mtval_q[11] ;
 wire \cs_registers_i.mtval_q[12] ;
 wire \cs_registers_i.mtval_q[13] ;
 wire \cs_registers_i.mtval_q[14] ;
 wire \cs_registers_i.mtval_q[15] ;
 wire \cs_registers_i.mtval_q[16] ;
 wire \cs_registers_i.mtval_q[17] ;
 wire \cs_registers_i.mtval_q[18] ;
 wire \cs_registers_i.mtval_q[19] ;
 wire \cs_registers_i.mtval_q[1] ;
 wire \cs_registers_i.mtval_q[20] ;
 wire \cs_registers_i.mtval_q[21] ;
 wire \cs_registers_i.mtval_q[22] ;
 wire \cs_registers_i.mtval_q[23] ;
 wire \cs_registers_i.mtval_q[24] ;
 wire \cs_registers_i.mtval_q[25] ;
 wire \cs_registers_i.mtval_q[26] ;
 wire \cs_registers_i.mtval_q[27] ;
 wire \cs_registers_i.mtval_q[28] ;
 wire \cs_registers_i.mtval_q[29] ;
 wire \cs_registers_i.mtval_q[2] ;
 wire \cs_registers_i.mtval_q[30] ;
 wire \cs_registers_i.mtval_q[31] ;
 wire \cs_registers_i.mtval_q[3] ;
 wire \cs_registers_i.mtval_q[4] ;
 wire \cs_registers_i.mtval_q[5] ;
 wire \cs_registers_i.mtval_q[6] ;
 wire \cs_registers_i.mtval_q[7] ;
 wire \cs_registers_i.mtval_q[8] ;
 wire \cs_registers_i.mtval_q[9] ;
 wire \cs_registers_i.nmi_mode_i ;
 wire \cs_registers_i.pc_id_i[10] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[12] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[14] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[16] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[18] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[20] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[22] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[24] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[26] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[28] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[30] ;
 wire \cs_registers_i.pc_id_i[31] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[4] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[6] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[8] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[10] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[12] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[14] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[16] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[18] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[1] ;
 wire \cs_registers_i.pc_if_i[20] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[22] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[24] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[26] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[28] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[30] ;
 wire \cs_registers_i.pc_if_i[31] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[4] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[6] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[8] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_lvl_q[0] ;
 wire \cs_registers_i.priv_lvl_q[1] ;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ;
 wire fetch_enable_q;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[4] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[4] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1000] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1001] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1002] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1003] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1004] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1005] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1006] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1007] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1008] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1009] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[100] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1010] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1011] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1012] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1013] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1014] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1015] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1016] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1017] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1018] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1019] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[101] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1020] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1021] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1022] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1023] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[102] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[103] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[104] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[105] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[106] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[107] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[108] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[109] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[110] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[111] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[112] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[113] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[114] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[115] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[116] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[117] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[118] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[119] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[120] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[121] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[122] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[123] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[124] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[125] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[126] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[127] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[128] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[129] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[130] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[131] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[132] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[133] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[134] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[135] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[136] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[137] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[138] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[139] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[140] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[141] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[142] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[143] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[144] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[145] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[146] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[147] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[148] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[149] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[150] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[151] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[152] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[153] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[154] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[155] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[156] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[157] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[158] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[159] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[160] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[161] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[162] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[163] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[164] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[165] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[166] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[167] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[168] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[169] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[170] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[171] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[172] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[173] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[174] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[175] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[176] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[177] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[178] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[179] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[180] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[181] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[182] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[183] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[184] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[185] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[186] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[187] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[188] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[189] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[190] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[191] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[192] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[193] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[194] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[195] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[196] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[197] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[198] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[199] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[200] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[201] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[202] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[203] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[204] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[205] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[206] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[207] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[208] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[209] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[210] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[211] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[212] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[213] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[214] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[215] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[216] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[217] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[218] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[219] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[220] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[221] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[222] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[223] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[224] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[225] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[226] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[227] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[228] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[229] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[230] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[231] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[232] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[233] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[234] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[235] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[236] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[237] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[238] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[239] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[240] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[241] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[242] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[243] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[244] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[245] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[246] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[247] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[248] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[249] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[250] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[251] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[252] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[253] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[254] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[255] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[256] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[257] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[258] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[259] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[260] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[261] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[262] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[263] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[264] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[265] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[266] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[267] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[268] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[269] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[270] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[271] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[272] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[273] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[274] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[275] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[276] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[277] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[278] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[279] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[280] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[281] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[282] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[283] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[284] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[285] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[286] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[287] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[288] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[289] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[290] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[291] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[292] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[293] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[294] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[295] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[296] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[297] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[298] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[299] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[300] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[301] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[302] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[303] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[304] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[305] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[306] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[307] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[308] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[309] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[310] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[311] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[312] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[313] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[314] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[315] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[316] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[317] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[318] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[319] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[320] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[321] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[322] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[323] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[324] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[325] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[326] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[327] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[328] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[329] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[32] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[330] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[331] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[332] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[333] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[334] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[335] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[336] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[337] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[338] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[339] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[33] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[340] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[341] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[342] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[343] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[344] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[345] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[346] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[347] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[348] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[349] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[34] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[350] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[351] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[352] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[353] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[354] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[355] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[356] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[357] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[358] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[359] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[35] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[360] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[361] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[362] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[363] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[364] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[365] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[366] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[367] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[368] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[369] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[36] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[370] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[371] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[372] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[373] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[374] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[375] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[376] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[377] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[378] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[379] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[37] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[380] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[381] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[382] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[383] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[384] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[385] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[386] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[387] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[388] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[389] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[38] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[390] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[391] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[392] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[393] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[394] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[395] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[396] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[397] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[398] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[399] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[39] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[400] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[401] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[402] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[403] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[404] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[405] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[406] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[407] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[408] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[409] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[40] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[410] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[411] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[412] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[413] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[414] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[415] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[416] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[417] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[418] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[419] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[41] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[420] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[421] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[422] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[423] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[424] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[425] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[426] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[427] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[428] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[429] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[42] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[430] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[431] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[432] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[433] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[434] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[435] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[436] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[437] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[438] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[439] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[43] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[440] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[441] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[442] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[443] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[444] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[445] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[446] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[447] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[448] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[449] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[44] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[450] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[451] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[452] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[453] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[454] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[455] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[456] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[457] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[458] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[459] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[45] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[460] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[461] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[462] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[463] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[464] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[465] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[466] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[467] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[468] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[469] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[46] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[470] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[471] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[472] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[473] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[474] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[475] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[476] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[477] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[478] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[479] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[47] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[480] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[481] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[482] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[483] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[484] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[485] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[486] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[487] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[488] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[489] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[48] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[490] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[491] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[492] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[493] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[494] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[495] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[496] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[497] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[498] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[499] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[49] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[500] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[501] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[502] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[503] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[504] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[505] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[506] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[507] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[508] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[509] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[50] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[510] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[511] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[512] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[513] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[514] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[515] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[516] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[517] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[518] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[519] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[51] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[520] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[521] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[522] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[523] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[524] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[525] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[526] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[527] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[528] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[529] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[52] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[530] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[531] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[532] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[533] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[534] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[535] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[536] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[537] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[538] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[539] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[53] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[540] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[541] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[542] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[543] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[544] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[545] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[546] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[547] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[548] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[549] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[54] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[550] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[551] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[552] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[553] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[554] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[555] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[556] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[557] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[558] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[559] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[55] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[560] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[561] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[562] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[563] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[564] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[565] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[566] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[567] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[568] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[569] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[56] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[570] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[571] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[572] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[573] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[574] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[575] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[576] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[577] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[578] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[579] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[57] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[580] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[581] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[582] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[583] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[584] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[585] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[586] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[587] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[588] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[589] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[58] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[590] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[591] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[592] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[593] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[594] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[595] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[596] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[597] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[598] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[599] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[59] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[600] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[601] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[602] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[603] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[604] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[605] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[606] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[607] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[608] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[609] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[60] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[610] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[611] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[612] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[613] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[614] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[615] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[616] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[617] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[618] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[619] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[61] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[620] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[621] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[622] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[623] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[624] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[625] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[626] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[627] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[628] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[629] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[62] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[630] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[631] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[632] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[633] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[634] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[635] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[636] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[637] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[638] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[639] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[63] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[640] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[641] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[642] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[643] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[644] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[645] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[646] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[647] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[648] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[649] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[64] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[650] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[651] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[652] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[653] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[654] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[655] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[656] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[657] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[658] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[659] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[65] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[660] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[661] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[662] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[663] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[664] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[665] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[666] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[667] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[668] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[669] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[66] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[670] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[671] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[672] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[673] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[674] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[675] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[676] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[677] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[678] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[679] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[67] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[680] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[681] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[682] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[683] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[684] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[685] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[686] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[687] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[688] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[689] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[68] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[690] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[691] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[692] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[693] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[694] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[695] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[696] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[697] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[698] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[699] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[69] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[700] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[701] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[702] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[703] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[704] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[705] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[706] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[707] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[708] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[709] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[70] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[710] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[711] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[712] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[713] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[714] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[715] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[716] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[717] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[718] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[719] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[71] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[720] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[721] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[722] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[723] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[724] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[725] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[726] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[727] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[728] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[729] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[72] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[730] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[731] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[732] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[733] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[734] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[735] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[736] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[737] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[738] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[739] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[73] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[740] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[741] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[742] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[743] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[744] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[745] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[746] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[747] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[748] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[749] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[74] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[750] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[751] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[752] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[753] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[754] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[755] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[756] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[757] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[758] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[759] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[75] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[760] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[761] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[762] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[763] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[764] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[765] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[766] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[767] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[768] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[769] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[76] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[770] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[771] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[772] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[773] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[774] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[775] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[776] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[777] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[778] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[779] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[77] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[780] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[781] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[782] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[783] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[784] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[785] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[786] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[787] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[788] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[789] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[78] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[790] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[791] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[792] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[793] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[794] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[795] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[796] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[797] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[798] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[799] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[79] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[800] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[801] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[802] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[803] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[804] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[805] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[806] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[807] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[808] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[809] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[80] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[810] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[811] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[812] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[813] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[814] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[815] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[816] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[817] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[818] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[819] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[81] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[820] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[821] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[822] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[823] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[824] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[825] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[826] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[827] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[828] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[829] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[82] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[830] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[831] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[832] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[833] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[834] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[835] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[836] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[837] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[838] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[839] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[83] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[840] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[841] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[842] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[843] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[844] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[845] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[846] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[847] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[848] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[849] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[84] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[850] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[851] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[852] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[853] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[854] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[855] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[856] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[857] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[858] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[859] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[85] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[860] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[861] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[862] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[863] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[864] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[865] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[866] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[867] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[868] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[869] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[86] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[870] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[871] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[872] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[873] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[874] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[875] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[876] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[877] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[878] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[879] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[87] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[880] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[881] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[882] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[883] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[884] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[885] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[886] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[887] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[888] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[889] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[88] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[890] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[891] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[892] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[893] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[894] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[895] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[896] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[897] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[898] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[899] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[89] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[900] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[901] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[902] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[903] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[904] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[905] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[906] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[907] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[908] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[909] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[90] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[910] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[911] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[912] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[913] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[914] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[915] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[916] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[917] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[918] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[919] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[91] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[920] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[921] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[922] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[923] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[924] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[925] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[926] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[927] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[928] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[929] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[92] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[930] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[931] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[932] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[933] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[934] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[935] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[936] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[937] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[938] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[939] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[93] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[940] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[941] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[942] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[943] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[944] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[945] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[946] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[947] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[948] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[949] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[94] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[950] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[951] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[952] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[953] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[954] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[955] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[956] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[957] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[958] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[959] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[95] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[960] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[961] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[962] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[963] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[964] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[965] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[966] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[967] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[968] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[969] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[96] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[970] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[971] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[972] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[973] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[974] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[975] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[976] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[977] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[978] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[979] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[97] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[980] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[981] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[982] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[983] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[984] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[985] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[986] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[987] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[988] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[989] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[98] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[990] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[991] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[992] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[993] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[994] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[995] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[996] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[997] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[998] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[999] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[99] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[4] ;
 wire \id_stage_i.branch_set ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[0] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[1] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[2] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[3] ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_compressed_i[0] ;
 wire \id_stage_i.controller_i.instr_compressed_i[10] ;
 wire \id_stage_i.controller_i.instr_compressed_i[11] ;
 wire \id_stage_i.controller_i.instr_compressed_i[12] ;
 wire \id_stage_i.controller_i.instr_compressed_i[13] ;
 wire \id_stage_i.controller_i.instr_compressed_i[14] ;
 wire \id_stage_i.controller_i.instr_compressed_i[15] ;
 wire \id_stage_i.controller_i.instr_compressed_i[1] ;
 wire \id_stage_i.controller_i.instr_compressed_i[2] ;
 wire \id_stage_i.controller_i.instr_compressed_i[3] ;
 wire \id_stage_i.controller_i.instr_compressed_i[4] ;
 wire \id_stage_i.controller_i.instr_compressed_i[5] ;
 wire \id_stage_i.controller_i.instr_compressed_i[6] ;
 wire \id_stage_i.controller_i.instr_compressed_i[7] ;
 wire \id_stage_i.controller_i.instr_compressed_i[8] ;
 wire \id_stage_i.controller_i.instr_compressed_i[9] ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_i[0] ;
 wire \id_stage_i.controller_i.instr_i[12] ;
 wire \id_stage_i.controller_i.instr_i[13] ;
 wire \id_stage_i.controller_i.instr_i[14] ;
 wire \id_stage_i.controller_i.instr_i[1] ;
 wire \id_stage_i.controller_i.instr_i[25] ;
 wire \id_stage_i.controller_i.instr_i[26] ;
 wire \id_stage_i.controller_i.instr_i[27] ;
 wire \id_stage_i.controller_i.instr_i[28] ;
 wire \id_stage_i.controller_i.instr_i[29] ;
 wire \id_stage_i.controller_i.instr_i[2] ;
 wire \id_stage_i.controller_i.instr_i[30] ;
 wire \id_stage_i.controller_i.instr_i[31] ;
 wire \id_stage_i.controller_i.instr_i[3] ;
 wire \id_stage_i.controller_i.instr_i[4] ;
 wire \id_stage_i.controller_i.instr_i[5] ;
 wire \id_stage_i.controller_i.instr_i[6] ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.load_err_d ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[0] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[10] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[11] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[12] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[13] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[14] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[15] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[16] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[17] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[18] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[19] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[1] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[20] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[21] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[22] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[23] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[24] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[25] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[26] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[27] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[28] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[29] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[2] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[30] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[31] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[3] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[4] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[5] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[6] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[7] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[8] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[9] ;
 wire \id_stage_i.controller_i.store_err_d ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_type_q[1] ;
 wire \load_store_unit_i.data_type_q[2] ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.ls_fsm_cs[0] ;
 wire \load_store_unit_i.ls_fsm_cs[1] ;
 wire \load_store_unit_i.ls_fsm_cs[2] ;
 wire \load_store_unit_i.lsu_err_q ;
 wire \load_store_unit_i.rdata_offset_q[0] ;
 wire \load_store_unit_i.rdata_offset_q[1] ;
 wire \load_store_unit_i.rdata_q[10] ;
 wire \load_store_unit_i.rdata_q[11] ;
 wire \load_store_unit_i.rdata_q[12] ;
 wire \load_store_unit_i.rdata_q[13] ;
 wire \load_store_unit_i.rdata_q[14] ;
 wire \load_store_unit_i.rdata_q[15] ;
 wire \load_store_unit_i.rdata_q[16] ;
 wire \load_store_unit_i.rdata_q[17] ;
 wire \load_store_unit_i.rdata_q[18] ;
 wire \load_store_unit_i.rdata_q[19] ;
 wire \load_store_unit_i.rdata_q[20] ;
 wire \load_store_unit_i.rdata_q[21] ;
 wire \load_store_unit_i.rdata_q[22] ;
 wire \load_store_unit_i.rdata_q[23] ;
 wire \load_store_unit_i.rdata_q[24] ;
 wire \load_store_unit_i.rdata_q[25] ;
 wire \load_store_unit_i.rdata_q[26] ;
 wire \load_store_unit_i.rdata_q[27] ;
 wire \load_store_unit_i.rdata_q[28] ;
 wire \load_store_unit_i.rdata_q[29] ;
 wire \load_store_unit_i.rdata_q[30] ;
 wire \load_store_unit_i.rdata_q[31] ;
 wire \load_store_unit_i.rdata_q[8] ;
 wire \load_store_unit_i.rdata_q[9] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_leaf_0_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_6_clk_i_regs;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_13_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_18_clk_i_regs;
 wire clknet_leaf_19_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_23_clk_i_regs;
 wire clknet_leaf_24_clk_i_regs;
 wire clknet_leaf_25_clk_i_regs;
 wire clknet_leaf_26_clk_i_regs;
 wire clknet_leaf_27_clk_i_regs;
 wire clknet_leaf_28_clk_i_regs;
 wire clknet_leaf_29_clk_i_regs;
 wire clknet_leaf_30_clk_i_regs;
 wire clknet_leaf_31_clk_i_regs;
 wire clknet_leaf_32_clk_i_regs;
 wire clknet_leaf_33_clk_i_regs;
 wire clknet_leaf_34_clk_i_regs;
 wire clknet_leaf_35_clk_i_regs;
 wire clknet_leaf_36_clk_i_regs;
 wire clknet_leaf_37_clk_i_regs;
 wire clknet_leaf_38_clk_i_regs;
 wire clknet_leaf_39_clk_i_regs;
 wire clknet_leaf_40_clk_i_regs;
 wire clknet_leaf_41_clk_i_regs;
 wire clknet_leaf_42_clk_i_regs;
 wire clknet_leaf_43_clk_i_regs;
 wire clknet_leaf_44_clk_i_regs;
 wire clknet_leaf_45_clk_i_regs;
 wire clknet_leaf_46_clk_i_regs;
 wire clknet_leaf_47_clk_i_regs;
 wire clknet_leaf_48_clk_i_regs;
 wire clknet_leaf_49_clk_i_regs;
 wire clknet_leaf_50_clk_i_regs;
 wire clknet_leaf_51_clk_i_regs;
 wire clknet_leaf_52_clk_i_regs;
 wire clknet_leaf_53_clk_i_regs;
 wire clknet_leaf_54_clk_i_regs;
 wire clknet_leaf_55_clk_i_regs;
 wire clknet_leaf_56_clk_i_regs;
 wire clknet_leaf_57_clk_i_regs;
 wire clknet_leaf_58_clk_i_regs;
 wire clknet_leaf_59_clk_i_regs;
 wire clknet_leaf_60_clk_i_regs;
 wire clknet_leaf_61_clk_i_regs;
 wire clknet_leaf_62_clk_i_regs;
 wire clknet_leaf_63_clk_i_regs;
 wire clknet_leaf_64_clk_i_regs;
 wire clknet_leaf_65_clk_i_regs;
 wire clknet_leaf_66_clk_i_regs;
 wire clknet_leaf_67_clk_i_regs;
 wire clknet_leaf_68_clk_i_regs;
 wire clknet_leaf_69_clk_i_regs;
 wire clknet_leaf_70_clk_i_regs;
 wire clknet_leaf_71_clk_i_regs;
 wire clknet_leaf_72_clk_i_regs;
 wire clknet_leaf_73_clk_i_regs;
 wire clknet_leaf_74_clk_i_regs;
 wire clknet_leaf_75_clk_i_regs;
 wire clknet_leaf_76_clk_i_regs;
 wire clknet_leaf_77_clk_i_regs;
 wire clknet_leaf_78_clk_i_regs;
 wire clknet_leaf_79_clk_i_regs;
 wire clknet_leaf_80_clk_i_regs;
 wire clknet_leaf_81_clk_i_regs;
 wire clknet_leaf_82_clk_i_regs;
 wire clknet_leaf_83_clk_i_regs;
 wire clknet_leaf_84_clk_i_regs;
 wire clknet_leaf_85_clk_i_regs;
 wire clknet_leaf_86_clk_i_regs;
 wire clknet_leaf_87_clk_i_regs;
 wire clknet_leaf_88_clk_i_regs;
 wire clknet_leaf_89_clk_i_regs;
 wire clknet_leaf_90_clk_i_regs;
 wire clknet_leaf_91_clk_i_regs;
 wire clknet_leaf_92_clk_i_regs;
 wire clknet_leaf_93_clk_i_regs;
 wire clknet_leaf_94_clk_i_regs;
 wire clknet_leaf_95_clk_i_regs;
 wire clknet_leaf_96_clk_i_regs;
 wire clknet_leaf_97_clk_i_regs;
 wire clknet_leaf_98_clk_i_regs;
 wire clknet_leaf_99_clk_i_regs;
 wire clknet_leaf_100_clk_i_regs;
 wire clknet_leaf_101_clk_i_regs;
 wire clknet_leaf_102_clk_i_regs;
 wire clknet_leaf_103_clk_i_regs;
 wire clknet_leaf_104_clk_i_regs;
 wire clknet_leaf_105_clk_i_regs;
 wire clknet_leaf_106_clk_i_regs;
 wire clknet_leaf_107_clk_i_regs;
 wire clknet_leaf_108_clk_i_regs;
 wire clknet_leaf_109_clk_i_regs;
 wire clknet_leaf_110_clk_i_regs;
 wire clknet_leaf_111_clk_i_regs;
 wire clknet_leaf_112_clk_i_regs;
 wire clknet_leaf_113_clk_i_regs;
 wire clknet_leaf_114_clk_i_regs;
 wire clknet_leaf_115_clk_i_regs;
 wire clknet_leaf_116_clk_i_regs;
 wire clknet_leaf_117_clk_i_regs;
 wire clknet_leaf_118_clk_i_regs;
 wire clknet_leaf_119_clk_i_regs;
 wire clknet_leaf_120_clk_i_regs;
 wire clknet_leaf_121_clk_i_regs;
 wire clknet_leaf_122_clk_i_regs;
 wire clknet_leaf_123_clk_i_regs;
 wire clknet_leaf_124_clk_i_regs;
 wire clknet_leaf_125_clk_i_regs;
 wire clknet_leaf_126_clk_i_regs;
 wire clknet_leaf_127_clk_i_regs;
 wire clknet_leaf_128_clk_i_regs;
 wire clknet_leaf_129_clk_i_regs;
 wire clknet_leaf_130_clk_i_regs;
 wire clknet_leaf_131_clk_i_regs;
 wire clknet_leaf_132_clk_i_regs;
 wire clknet_leaf_133_clk_i_regs;
 wire clknet_leaf_134_clk_i_regs;
 wire clknet_leaf_135_clk_i_regs;
 wire clknet_leaf_136_clk_i_regs;
 wire clknet_leaf_137_clk_i_regs;
 wire clknet_0_clk_i_regs;
 wire clknet_4_0_0_clk_i_regs;
 wire clknet_4_1_0_clk_i_regs;
 wire clknet_4_2_0_clk_i_regs;
 wire clknet_4_3_0_clk_i_regs;
 wire clknet_4_4_0_clk_i_regs;
 wire clknet_4_5_0_clk_i_regs;
 wire clknet_4_6_0_clk_i_regs;
 wire clknet_4_7_0_clk_i_regs;
 wire clknet_4_8_0_clk_i_regs;
 wire clknet_4_9_0_clk_i_regs;
 wire clknet_4_10_0_clk_i_regs;
 wire clknet_4_11_0_clk_i_regs;
 wire clknet_4_12_0_clk_i_regs;
 wire clknet_4_13_0_clk_i_regs;
 wire clknet_4_14_0_clk_i_regs;
 wire clknet_4_15_0_clk_i_regs;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire delaynet_0_core_clock;
 wire delaynet_1_core_clock;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net289;
 wire net290;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net307;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net358;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net599;
 wire net629;
 wire net630;
 wire net631;
 wire net313;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net357;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net386;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net435;
 wire net438;
 wire net439;
 wire net450;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;

 BUF_X8 _16515_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .Z(_10699_));
 BUF_X16 _16516_ (.A(_10699_),
    .Z(_10700_));
 BUF_X32 _16517_ (.A(_10700_),
    .Z(_10701_));
 BUF_X32 _16518_ (.A(_10701_),
    .Z(_10702_));
 BUF_X32 _16519_ (.A(_10702_),
    .Z(_10703_));
 BUF_X32 _16520_ (.A(_10703_),
    .Z(_10704_));
 BUF_X8 _16521_ (.A(_10704_),
    .Z(_10705_));
 MUX2_X1 _16522_ (.A(_00163_),
    .B(_00165_),
    .S(_10705_),
    .Z(_10706_));
 MUX2_X1 _16523_ (.A(_00164_),
    .B(_00166_),
    .S(_10705_),
    .Z(_10707_));
 BUF_X4 _16524_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(_10708_));
 BUF_X8 _16525_ (.A(_10708_),
    .Z(_10709_));
 BUF_X4 _16526_ (.A(_10709_),
    .Z(_10710_));
 BUF_X8 _16527_ (.A(_10710_),
    .Z(_10711_));
 BUF_X4 _16528_ (.A(_10711_),
    .Z(_10712_));
 MUX2_X1 _16529_ (.A(_10706_),
    .B(_10707_),
    .S(_10712_),
    .Z(_10713_));
 MUX2_X1 _16530_ (.A(_00155_),
    .B(_00157_),
    .S(_10705_),
    .Z(_10714_));
 MUX2_X1 _16531_ (.A(_00156_),
    .B(_00158_),
    .S(_10705_),
    .Z(_10715_));
 MUX2_X1 _16532_ (.A(_10714_),
    .B(_10715_),
    .S(_10712_),
    .Z(_10716_));
 BUF_X4 _16533_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(_10717_));
 INV_X8 _16534_ (.A(_10717_),
    .ZN(_10718_));
 BUF_X4 _16535_ (.A(_10718_),
    .Z(_10719_));
 MUX2_X1 _16536_ (.A(_10713_),
    .B(_10716_),
    .S(_10719_),
    .Z(_10720_));
 MUX2_X1 _16537_ (.A(_00167_),
    .B(_00169_),
    .S(_10705_),
    .Z(_10721_));
 MUX2_X1 _16538_ (.A(_00168_),
    .B(_00170_),
    .S(_10705_),
    .Z(_10722_));
 MUX2_X1 _16539_ (.A(_10721_),
    .B(_10722_),
    .S(_10712_),
    .Z(_10723_));
 MUX2_X1 _16540_ (.A(_00159_),
    .B(_00161_),
    .S(_10705_),
    .Z(_10724_));
 MUX2_X1 _16541_ (.A(_00160_),
    .B(_00162_),
    .S(_10705_),
    .Z(_10725_));
 MUX2_X1 _16542_ (.A(_10724_),
    .B(_10725_),
    .S(_10712_),
    .Z(_10726_));
 MUX2_X1 _16543_ (.A(_10723_),
    .B(_10726_),
    .S(_10719_),
    .Z(_10727_));
 BUF_X4 _16544_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(_10728_));
 BUF_X4 _16545_ (.A(_10728_),
    .Z(_10729_));
 BUF_X4 _16546_ (.A(_10729_),
    .Z(_10730_));
 BUF_X4 _16547_ (.A(_10730_),
    .Z(_10731_));
 MUX2_X1 _16548_ (.A(_10720_),
    .B(_10727_),
    .S(_10731_),
    .Z(_10732_));
 BUF_X4 _16549_ (.A(_10728_),
    .Z(_10733_));
 INV_X1 _16550_ (.A(_10733_),
    .ZN(_10734_));
 BUF_X8 _16551_ (.A(_10734_),
    .Z(_10735_));
 BUF_X8 _16552_ (.A(_10735_),
    .Z(_10736_));
 BUF_X8 _16553_ (.A(_10704_),
    .Z(_10737_));
 MUX2_X1 _16554_ (.A(_00151_),
    .B(_00153_),
    .S(_10737_),
    .Z(_10738_));
 MUX2_X1 _16555_ (.A(_00152_),
    .B(_00154_),
    .S(_10737_),
    .Z(_10739_));
 MUX2_X1 _16556_ (.A(_10738_),
    .B(_10739_),
    .S(_10711_),
    .Z(_10740_));
 MUX2_X1 _16557_ (.A(_00143_),
    .B(_00145_),
    .S(_10737_),
    .Z(_10741_));
 MUX2_X1 _16558_ (.A(_00144_),
    .B(_00146_),
    .S(_10737_),
    .Z(_10742_));
 MUX2_X1 _16559_ (.A(_10741_),
    .B(_10742_),
    .S(_10711_),
    .Z(_10743_));
 MUX2_X1 _16560_ (.A(_10740_),
    .B(_10743_),
    .S(_10719_),
    .Z(_10744_));
 NOR2_X1 _16561_ (.A1(_10736_),
    .A2(_10744_),
    .ZN(_10745_));
 BUF_X8 _16562_ (.A(_10717_),
    .Z(_10746_));
 BUF_X4 _16563_ (.A(_10746_),
    .Z(_10747_));
 BUF_X8 _16564_ (.A(_10704_),
    .Z(_10748_));
 NOR2_X1 _16565_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .A2(_10748_),
    .ZN(_10749_));
 BUF_X32 _16566_ (.A(_10704_),
    .Z(_10750_));
 AOI21_X1 _16567_ (.A(_10749_),
    .B1(net379),
    .B2(_00142_),
    .ZN(_10751_));
 NOR2_X1 _16568_ (.A1(_10712_),
    .A2(_00141_),
    .ZN(_10752_));
 AOI221_X2 _16569_ (.A(_10747_),
    .B1(_10751_),
    .B2(_10712_),
    .C1(_10752_),
    .C2(net379),
    .ZN(_10753_));
 MUX2_X1 _16570_ (.A(_00147_),
    .B(_00149_),
    .S(net379),
    .Z(_10754_));
 MUX2_X1 _16571_ (.A(_00148_),
    .B(_00150_),
    .S(net379),
    .Z(_10755_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 MUX2_X1 _16573_ (.A(_10754_),
    .B(_10755_),
    .S(_10711_),
    .Z(_10757_));
 BUF_X8 _16574_ (.A(_10747_),
    .Z(_10758_));
 AOI21_X1 _16575_ (.A(_10753_),
    .B1(_10757_),
    .B2(_10758_),
    .ZN(_10759_));
 AOI21_X1 _16576_ (.A(_10745_),
    .B1(_10759_),
    .B2(_10736_),
    .ZN(_10760_));
 BUF_X8 _16577_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .Z(_10761_));
 INV_X1 _16578_ (.A(_10761_),
    .ZN(_10762_));
 BUF_X4 _16579_ (.A(_10762_),
    .Z(_10763_));
 BUF_X8 _16580_ (.A(_10763_),
    .Z(_10764_));
 MUX2_X2 _16581_ (.A(_10732_),
    .B(_10760_),
    .S(_10764_),
    .Z(_10765_));
 INV_X1 _16582_ (.A(_16486_),
    .ZN(_10766_));
 BUF_X2 _16583_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .Z(_10767_));
 CLKBUF_X3 _16584_ (.A(_00171_),
    .Z(_10768_));
 AND2_X1 _16585_ (.A1(_10767_),
    .A2(_10768_),
    .ZN(_10769_));
 MUX2_X2 _16586_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(_10768_),
    .S(_10767_),
    .Z(_10770_));
 BUF_X4 _16587_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .Z(_10771_));
 INV_X2 _16588_ (.A(_10771_),
    .ZN(_10772_));
 AOI22_X4 _16589_ (.A1(_10766_),
    .A2(_10769_),
    .B1(_10770_),
    .B2(_10772_),
    .ZN(_10773_));
 BUF_X4 _16590_ (.A(_10773_),
    .Z(_10774_));
 BUF_X1 rebuffer17 (.A(\id_stage_i.controller_i.instr_i[14] ),
    .Z(net291));
 BUF_X8 _16592_ (.A(\id_stage_i.controller_i.instr_i[14] ),
    .Z(_10776_));
 BUF_X4 _16593_ (.A(\id_stage_i.controller_i.instr_i[4] ),
    .Z(_10777_));
 BUF_X4 _16594_ (.A(_10777_),
    .Z(_10778_));
 BUF_X4 _16595_ (.A(\id_stage_i.controller_i.instr_i[6] ),
    .Z(_10779_));
 OR2_X4 _16596_ (.A1(_10778_),
    .A2(_10779_),
    .ZN(_10780_));
 NOR2_X4 _16597_ (.A1(_10777_),
    .A2(_00172_),
    .ZN(_10781_));
 INV_X2 _16598_ (.A(_10779_),
    .ZN(_10782_));
 OAI22_X2 _16599_ (.A1(net303),
    .A2(_10780_),
    .B1(_10781_),
    .B2(_10782_),
    .ZN(_10783_));
 BUF_X8 _16600_ (.A(\id_stage_i.controller_i.instr_i[5] ),
    .Z(_10784_));
 BUF_X4 _16601_ (.A(_10784_),
    .Z(_10785_));
 BUF_X4 _16602_ (.A(\id_stage_i.controller_i.instr_i[1] ),
    .Z(_10786_));
 BUF_X4 _16603_ (.A(\id_stage_i.controller_i.instr_i[0] ),
    .Z(_10787_));
 AND2_X2 _16604_ (.A1(_10786_),
    .A2(_10787_),
    .ZN(_10788_));
 BUF_X8 _16605_ (.A(_10788_),
    .Z(_10789_));
 BUF_X8 _16606_ (.A(\id_stage_i.controller_i.instr_i[2] ),
    .Z(_10790_));
 NOR2_X4 _16607_ (.A1(_10790_),
    .A2(\id_stage_i.controller_i.instr_i[3] ),
    .ZN(_10791_));
 NAND3_X1 _16608_ (.A1(_10785_),
    .A2(_10789_),
    .A3(_10791_),
    .ZN(_10792_));
 BUF_X2 _16609_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .Z(_10793_));
 BUF_X4 _16610_ (.A(_10793_),
    .Z(_10794_));
 BUF_X4 _16611_ (.A(\id_stage_i.id_fsm_q ),
    .Z(_10795_));
 INV_X4 _16612_ (.A(_10795_),
    .ZN(_10796_));
 AOI21_X4 _16613_ (.A(_10790_),
    .B1(_10794_),
    .B2(_10796_),
    .ZN(_10797_));
 BUF_X4 _16614_ (.A(\id_stage_i.controller_i.instr_i[3] ),
    .Z(_10798_));
 INV_X8 _16615_ (.A(_10784_),
    .ZN(_10799_));
 OR2_X4 _16616_ (.A1(_10777_),
    .A2(_00172_),
    .ZN(_10800_));
 NAND2_X4 _16617_ (.A1(net310),
    .A2(net308),
    .ZN(_10801_));
 BUF_X8 _16618_ (.A(_10801_),
    .Z(_10802_));
 NOR4_X4 _16619_ (.A1(_10798_),
    .A2(_10799_),
    .A3(_10800_),
    .A4(_10802_),
    .ZN(_10803_));
 AOI211_X2 _16620_ (.A(_10783_),
    .B(_10792_),
    .C1(_10797_),
    .C2(_10803_),
    .ZN(_10804_));
 NAND2_X4 _16621_ (.A1(_10774_),
    .A2(_10804_),
    .ZN(_10805_));
 OR2_X1 _16622_ (.A1(_10765_),
    .A2(_10805_),
    .ZN(_10806_));
 INV_X4 _16623_ (.A(_10798_),
    .ZN(_10807_));
 NAND4_X4 _16624_ (.A1(_10807_),
    .A2(_10785_),
    .A3(_10781_),
    .A4(_10789_),
    .ZN(_10808_));
 INV_X4 _16625_ (.A(_10790_),
    .ZN(_10809_));
 INV_X4 _16626_ (.A(_10793_),
    .ZN(_10810_));
 OAI21_X2 _16627_ (.A(_10809_),
    .B1(_10810_),
    .B2(_10795_),
    .ZN(_10811_));
 NAND4_X4 _16628_ (.A1(_10807_),
    .A2(_10778_),
    .A3(_10782_),
    .A4(_10789_),
    .ZN(_10812_));
 OAI221_X2 _16629_ (.A(_10773_),
    .B1(_10808_),
    .B2(_10811_),
    .C1(_10812_),
    .C2(_10809_),
    .ZN(_10813_));
 BUF_X4 _16630_ (.A(_10813_),
    .Z(_10814_));
 NAND2_X1 _16631_ (.A1(_10772_),
    .A2(_10770_),
    .ZN(_10815_));
 NAND2_X2 _16632_ (.A1(_10767_),
    .A2(_10768_),
    .ZN(_10816_));
 OAI21_X4 _16633_ (.A(_10815_),
    .B1(_10816_),
    .B2(_16486_),
    .ZN(_10817_));
 BUF_X4 _16634_ (.A(_10817_),
    .Z(_10818_));
 BUF_X4 _16635_ (.A(_10818_),
    .Z(_10819_));
 NOR2_X4 _16636_ (.A1(_10777_),
    .A2(\id_stage_i.controller_i.instr_i[6] ),
    .ZN(_10820_));
 NAND4_X4 _16637_ (.A1(_10785_),
    .A2(_10820_),
    .A3(_10789_),
    .A4(_10791_),
    .ZN(_10821_));
 OAI22_X4 _16638_ (.A1(_10809_),
    .A2(_10812_),
    .B1(_10821_),
    .B2(_10776_),
    .ZN(_10822_));
 NAND2_X4 _16639_ (.A1(_10784_),
    .A2(_10781_),
    .ZN(_10823_));
 NOR2_X4 _16640_ (.A1(_10810_),
    .A2(_10795_),
    .ZN(_10824_));
 BUF_X4 _16641_ (.A(\id_stage_i.controller_i.instr_i[13] ),
    .Z(_10825_));
 INV_X4 _16642_ (.A(_10825_),
    .ZN(_10826_));
 BUF_X1 rebuffer25 (.A(_10879_),
    .Z(net299));
 BUF_X4 _16644_ (.A(\id_stage_i.controller_i.instr_i[12] ),
    .Z(_10828_));
 CLKBUF_X3 _16645_ (.A(_00173_),
    .Z(_10829_));
 NAND3_X4 _16646_ (.A1(_10826_),
    .A2(_10828_),
    .A3(_10829_),
    .ZN(_10830_));
 NAND3_X4 _16647_ (.A1(_10798_),
    .A2(_10799_),
    .A3(_10820_),
    .ZN(_10831_));
 OAI22_X4 _16648_ (.A1(_10823_),
    .A2(_10824_),
    .B1(_10830_),
    .B2(_10831_),
    .ZN(_10832_));
 AND3_X1 _16649_ (.A1(net310),
    .A2(net308),
    .A3(_10790_),
    .ZN(_10833_));
 BUF_X4 _16650_ (.A(_10833_),
    .Z(_10834_));
 AOI21_X2 _16651_ (.A(_10822_),
    .B1(_10832_),
    .B2(_10834_),
    .ZN(_10835_));
 CLKBUF_X3 _16652_ (.A(_10835_),
    .Z(_10836_));
 OAI21_X1 _16653_ (.A(net379),
    .B1(_10819_),
    .B2(_10836_),
    .ZN(_10837_));
 BUF_X4 _16654_ (.A(_10774_),
    .Z(_10838_));
 INV_X2 _16655_ (.A(_10778_),
    .ZN(_10839_));
 NOR4_X4 _16656_ (.A1(_10802_),
    .A2(_10839_),
    .A3(_10779_),
    .A4(_10798_),
    .ZN(_10840_));
 OR2_X2 _16657_ (.A1(\id_stage_i.controller_i.instr_i[2] ),
    .A2(\id_stage_i.controller_i.instr_i[3] ),
    .ZN(_10841_));
 BUF_X8 _16658_ (.A(_10841_),
    .Z(_10842_));
 NOR4_X4 _16659_ (.A1(_10799_),
    .A2(_10780_),
    .A3(_10802_),
    .A4(_10842_),
    .ZN(_10843_));
 INV_X4 _16660_ (.A(net293),
    .ZN(_10844_));
 AOI22_X4 _16661_ (.A1(_10790_),
    .A2(net367),
    .B1(_10843_),
    .B2(_10844_),
    .ZN(_10845_));
 NOR2_X4 _16662_ (.A1(_10799_),
    .A2(_10800_),
    .ZN(_10846_));
 NAND2_X4 _16663_ (.A1(_10793_),
    .A2(_10796_),
    .ZN(_10847_));
 INV_X1 _16664_ (.A(\id_stage_i.controller_i.instr_i[12] ),
    .ZN(_10848_));
 BUF_X4 _16665_ (.A(_10848_),
    .Z(_10849_));
 INV_X4 _16666_ (.A(_10829_),
    .ZN(_10850_));
 NOR3_X4 _16667_ (.A1(_10825_),
    .A2(_10849_),
    .A3(_10850_),
    .ZN(_10851_));
 NOR3_X4 _16668_ (.A1(_10807_),
    .A2(_10785_),
    .A3(_10780_),
    .ZN(_10852_));
 AOI22_X4 _16669_ (.A1(_10846_),
    .A2(_10847_),
    .B1(_10851_),
    .B2(_10852_),
    .ZN(_10853_));
 NAND3_X4 _16670_ (.A1(net311),
    .A2(net309),
    .A3(_10790_),
    .ZN(_10854_));
 OAI21_X4 _16671_ (.A(_10845_),
    .B1(_10853_),
    .B2(_10854_),
    .ZN(_10855_));
 NAND3_X2 _16672_ (.A1(_10807_),
    .A2(_10794_),
    .A3(_10796_),
    .ZN(_10856_));
 AOI22_X4 _16673_ (.A1(_10851_),
    .A2(_10852_),
    .B1(_10856_),
    .B2(_10846_),
    .ZN(_10857_));
 OAI21_X2 _16674_ (.A(_10773_),
    .B1(_10854_),
    .B2(_10857_),
    .ZN(_10858_));
 CLKBUF_X3 _16675_ (.A(_10858_),
    .Z(_10859_));
 NAND4_X1 _16676_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_10838_),
    .A3(_10855_),
    .A4(_10859_),
    .ZN(_10860_));
 AOI21_X1 _16677_ (.A(_10814_),
    .B1(_10837_),
    .B2(_10860_),
    .ZN(_10861_));
 BUF_X4 _16678_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .Z(_10862_));
 INV_X4 _16679_ (.A(_10862_),
    .ZN(_10863_));
 AOI22_X4 _16680_ (.A1(_10803_),
    .A2(_10797_),
    .B1(_10840_),
    .B2(_10790_),
    .ZN(_10864_));
 AND2_X1 _16681_ (.A1(_10773_),
    .A2(_10864_),
    .ZN(_10865_));
 XNOR2_X2 _16682_ (.A(_10865_),
    .B(_10835_),
    .ZN(_10866_));
 NOR3_X1 _16683_ (.A1(_10863_),
    .A2(_10859_),
    .A3(_10866_),
    .ZN(_10867_));
 OAI21_X1 _16684_ (.A(_10805_),
    .B1(_10861_),
    .B2(_10867_),
    .ZN(_10868_));
 AND2_X4 _16685_ (.A1(_10806_),
    .A2(_10868_),
    .ZN(_16236_));
 INV_X2 _16686_ (.A(_16236_),
    .ZN(_16247_));
 BUF_X4 _16687_ (.A(\id_stage_i.controller_i.instr_i[26] ),
    .Z(_10869_));
 NOR3_X4 _16688_ (.A1(_10842_),
    .A2(_10801_),
    .A3(_10799_),
    .ZN(_10870_));
 NOR2_X4 _16689_ (.A1(_10839_),
    .A2(_10779_),
    .ZN(_10871_));
 NAND2_X4 _16690_ (.A1(net297),
    .A2(_10871_),
    .ZN(_10872_));
 BUF_X4 _16691_ (.A(\id_stage_i.controller_i.instr_i[27] ),
    .Z(_10873_));
 NOR2_X1 _16692_ (.A1(\id_stage_i.controller_i.instr_i[25] ),
    .A2(_10873_),
    .ZN(_10874_));
 BUF_X4 _16693_ (.A(\id_stage_i.controller_i.instr_i[29] ),
    .Z(_10875_));
 BUF_X4 _16694_ (.A(\id_stage_i.controller_i.instr_i[28] ),
    .Z(_10876_));
 NOR2_X2 _16695_ (.A1(_10875_),
    .A2(_10876_),
    .ZN(_10877_));
 CLKBUF_X3 _16696_ (.A(\id_stage_i.controller_i.instr_i[31] ),
    .Z(_10878_));
 NOR2_X4 _16697_ (.A1(_10878_),
    .A2(\id_stage_i.controller_i.instr_i[26] ),
    .ZN(_10879_));
 AND3_X1 _16698_ (.A1(_10874_),
    .A2(_10877_),
    .A3(_10879_),
    .ZN(_10880_));
 BUF_X8 _16699_ (.A(_10825_),
    .Z(_10881_));
 BUF_X8 _16700_ (.A(_10881_),
    .Z(_10882_));
 CLKBUF_X2 _16701_ (.A(\id_stage_i.controller_i.instr_i[30] ),
    .Z(_10883_));
 BUF_X4 _16702_ (.A(_10883_),
    .Z(_10884_));
 NOR2_X2 _16703_ (.A1(_10776_),
    .A2(net412),
    .ZN(_10885_));
 AND2_X1 _16704_ (.A1(_10884_),
    .A2(_10885_),
    .ZN(_10886_));
 AND2_X4 _16705_ (.A1(net292),
    .A2(\id_stage_i.controller_i.instr_i[12] ),
    .ZN(_10887_));
 INV_X2 _16706_ (.A(_10883_),
    .ZN(_10888_));
 AOI21_X1 _16707_ (.A(_10886_),
    .B1(_10887_),
    .B2(_10888_),
    .ZN(_10889_));
 NAND2_X1 _16708_ (.A1(_10882_),
    .A2(_10849_),
    .ZN(_10890_));
 OAI22_X1 _16709_ (.A1(_10882_),
    .A2(_10889_),
    .B1(_10890_),
    .B2(_10884_),
    .ZN(_10891_));
 NAND2_X1 _16710_ (.A1(_10880_),
    .A2(_10891_),
    .ZN(_10892_));
 NAND2_X4 _16711_ (.A1(_10789_),
    .A2(_10791_),
    .ZN(_10893_));
 AND3_X4 _16712_ (.A1(_10825_),
    .A2(_10829_),
    .A3(_10887_),
    .ZN(_10894_));
 INV_X1 _16713_ (.A(_00176_),
    .ZN(_10895_));
 AOI211_X2 _16714_ (.A(_10825_),
    .B(_10895_),
    .C1(_10848_),
    .C2(net291),
    .ZN(_10896_));
 NOR2_X4 _16715_ (.A1(_10784_),
    .A2(\id_stage_i.controller_i.instr_i[6] ),
    .ZN(_10897_));
 NAND2_X4 _16716_ (.A1(_10777_),
    .A2(_10897_),
    .ZN(_10898_));
 OR4_X4 _16717_ (.A1(_10893_),
    .A2(_10894_),
    .A3(_10896_),
    .A4(_10898_),
    .ZN(_10899_));
 BUF_X2 _16718_ (.A(_00174_),
    .Z(_10900_));
 NOR3_X4 _16719_ (.A1(_10876_),
    .A2(_10875_),
    .A3(_10873_),
    .ZN(_10901_));
 AND2_X1 _16720_ (.A1(_10900_),
    .A2(_10901_),
    .ZN(_10902_));
 NOR3_X4 _16721_ (.A1(_10849_),
    .A2(_10825_),
    .A3(_10844_),
    .ZN(_10903_));
 NAND2_X2 _16722_ (.A1(_10902_),
    .A2(_10903_),
    .ZN(_10904_));
 OAI33_X1 _16723_ (.A1(_10869_),
    .A2(_10872_),
    .A3(_10892_),
    .B1(_10899_),
    .B2(_10904_),
    .B3(_10884_),
    .ZN(_10905_));
 INV_X1 _16724_ (.A(_10905_),
    .ZN(_10906_));
 NOR4_X4 _16725_ (.A1(_10893_),
    .A2(_10894_),
    .A3(_10896_),
    .A4(_10898_),
    .ZN(_10907_));
 NAND3_X1 _16726_ (.A1(_10882_),
    .A2(_10849_),
    .A3(_10907_),
    .ZN(_10908_));
 NOR4_X4 _16727_ (.A1(_10801_),
    .A2(_10800_),
    .A3(_10842_),
    .A4(_10799_),
    .ZN(_10909_));
 NAND2_X4 _16728_ (.A1(_10909_),
    .A2(_10824_),
    .ZN(_10910_));
 OAI21_X2 _16729_ (.A(_10908_),
    .B1(_10910_),
    .B2(_10882_),
    .ZN(_10911_));
 BUF_X4 _16730_ (.A(_10844_),
    .Z(_10912_));
 BUF_X4 _16731_ (.A(_10912_),
    .Z(_10913_));
 BUF_X4 _16732_ (.A(_10828_),
    .Z(_10914_));
 OAI21_X1 _16733_ (.A(_10913_),
    .B1(_10914_),
    .B2(_10850_),
    .ZN(_10915_));
 NAND2_X1 _16734_ (.A1(_10911_),
    .A2(_10915_),
    .ZN(_10916_));
 AND2_X4 _16735_ (.A1(_10906_),
    .A2(_10916_),
    .ZN(_15759_));
 INV_X1 _16736_ (.A(_15759_),
    .ZN(_15766_));
 BUF_X4 _16737_ (.A(_10829_),
    .Z(_10917_));
 NAND2_X2 _16738_ (.A1(_10900_),
    .A2(net295),
    .ZN(_10918_));
 OAI21_X1 _16739_ (.A(_10826_),
    .B1(_10917_),
    .B2(_10918_),
    .ZN(_10919_));
 AOI21_X1 _16740_ (.A(_10913_),
    .B1(_10914_),
    .B2(_10919_),
    .ZN(_10920_));
 BUF_X16 _16741_ (.A(_10776_),
    .Z(_10921_));
 BUF_X16 _16742_ (.A(_10921_),
    .Z(_10922_));
 BUF_X16 _16743_ (.A(_10922_),
    .Z(_10923_));
 BUF_X8 _16744_ (.A(_10923_),
    .Z(_10924_));
 OAI21_X1 _16745_ (.A(_10914_),
    .B1(_10917_),
    .B2(_10882_),
    .ZN(_10925_));
 NOR2_X1 _16746_ (.A1(_10924_),
    .A2(_10925_),
    .ZN(_10926_));
 OAI21_X1 _16747_ (.A(_10907_),
    .B1(_10920_),
    .B2(_10926_),
    .ZN(_10927_));
 NOR2_X2 _16748_ (.A1(_10881_),
    .A2(_10850_),
    .ZN(_10928_));
 NAND4_X2 _16749_ (.A1(_10798_),
    .A2(_10799_),
    .A3(_10820_),
    .A4(_10834_),
    .ZN(_10929_));
 OR2_X1 _16750_ (.A1(_10928_),
    .A2(_10929_),
    .ZN(_10930_));
 NAND2_X1 _16751_ (.A1(_10807_),
    .A2(_10789_),
    .ZN(_10931_));
 OAI21_X2 _16752_ (.A(_10782_),
    .B1(_10778_),
    .B2(_10809_),
    .ZN(_10932_));
 AOI21_X4 _16753_ (.A(_10931_),
    .B1(_10823_),
    .B2(_10932_),
    .ZN(_10933_));
 NAND2_X1 _16754_ (.A1(_10798_),
    .A2(_10839_),
    .ZN(_10934_));
 INV_X1 _16755_ (.A(_00172_),
    .ZN(_10935_));
 AOI21_X2 _16756_ (.A(_10897_),
    .B1(_10935_),
    .B2(_10784_),
    .ZN(_10936_));
 NOR3_X4 _16757_ (.A1(_10854_),
    .A2(_10934_),
    .A3(_10936_),
    .ZN(_10937_));
 OAI21_X1 _16758_ (.A(_10930_),
    .B1(_10933_),
    .B2(_10937_),
    .ZN(_10938_));
 NAND2_X2 _16759_ (.A1(_10826_),
    .A2(_10828_),
    .ZN(_10939_));
 NAND2_X1 _16760_ (.A1(_10939_),
    .A2(_10890_),
    .ZN(_10940_));
 AOI21_X1 _16761_ (.A(_10851_),
    .B1(_10940_),
    .B2(_10924_),
    .ZN(_10941_));
 NAND4_X4 _16762_ (.A1(_10784_),
    .A2(_10781_),
    .A3(_10789_),
    .A4(_10791_),
    .ZN(_10942_));
 NOR2_X4 _16763_ (.A1(_10847_),
    .A2(_10942_),
    .ZN(_10943_));
 NAND2_X1 _16764_ (.A1(_10879_),
    .A2(_10901_),
    .ZN(_10944_));
 BUF_X4 _16765_ (.A(\id_stage_i.controller_i.instr_i[25] ),
    .Z(_10945_));
 NOR2_X1 _16766_ (.A1(_10881_),
    .A2(_10945_),
    .ZN(_10946_));
 OAI21_X1 _16767_ (.A(_10946_),
    .B1(_10828_),
    .B2(_10844_),
    .ZN(_10947_));
 NOR2_X1 _16768_ (.A1(_10776_),
    .A2(_10849_),
    .ZN(_10948_));
 INV_X1 _16769_ (.A(_10945_),
    .ZN(_10949_));
 AOI221_X2 _16770_ (.A(_10944_),
    .B1(_10947_),
    .B2(_10884_),
    .C1(_10948_),
    .C2(_10949_),
    .ZN(_10950_));
 NOR2_X2 _16771_ (.A1(_10921_),
    .A2(_10881_),
    .ZN(_10951_));
 MUX2_X2 _16772_ (.A(_10923_),
    .B(_10951_),
    .S(_10828_),
    .Z(_10952_));
 NAND3_X2 _16773_ (.A1(_10888_),
    .A2(_10880_),
    .A3(_10952_),
    .ZN(_10953_));
 NAND3_X2 _16774_ (.A1(_00177_),
    .A2(_10950_),
    .A3(_10953_),
    .ZN(_10954_));
 AND2_X4 _16775_ (.A1(net297),
    .A2(_10871_),
    .ZN(_10955_));
 AOI221_X2 _16776_ (.A(_10938_),
    .B1(_10941_),
    .B2(_10943_),
    .C1(_10954_),
    .C2(_10955_),
    .ZN(_10956_));
 NAND2_X2 _16777_ (.A1(_10927_),
    .A2(_10956_),
    .ZN(_15760_));
 INV_X1 _16778_ (.A(_15760_),
    .ZN(_15763_));
 BUF_X4 _16779_ (.A(_10819_),
    .Z(_10957_));
 BUF_X4 _16780_ (.A(_10819_),
    .Z(_10958_));
 NOR3_X4 _16781_ (.A1(_10798_),
    .A2(_10810_),
    .A3(_10795_),
    .ZN(_10959_));
 NOR2_X1 _16782_ (.A1(_10790_),
    .A2(_10807_),
    .ZN(_10960_));
 NOR4_X2 _16783_ (.A1(_10802_),
    .A2(_10823_),
    .A3(_10959_),
    .A4(_10960_),
    .ZN(_10961_));
 NAND3_X4 _16784_ (.A1(_10778_),
    .A2(_10785_),
    .A3(_10779_),
    .ZN(_10962_));
 NAND2_X1 _16785_ (.A1(_10778_),
    .A2(_10784_),
    .ZN(_10963_));
 AOI211_X2 _16786_ (.A(_10802_),
    .B(_10842_),
    .C1(_10963_),
    .C2(_10779_),
    .ZN(_10964_));
 NOR4_X2 _16787_ (.A1(_10807_),
    .A2(_10785_),
    .A3(_10780_),
    .A4(_10854_),
    .ZN(_10965_));
 OAI33_X1 _16788_ (.A1(_10917_),
    .A2(_10893_),
    .A3(_10962_),
    .B1(_10964_),
    .B2(_10965_),
    .B3(_10803_),
    .ZN(_10966_));
 NOR2_X4 _16789_ (.A1(_10881_),
    .A2(_10828_),
    .ZN(_10967_));
 AND2_X1 _16790_ (.A1(_10917_),
    .A2(_10967_),
    .ZN(_10968_));
 OAI22_X2 _16791_ (.A1(_10798_),
    .A2(_10898_),
    .B1(_10968_),
    .B2(_10831_),
    .ZN(_10969_));
 AOI211_X2 _16792_ (.A(_10961_),
    .B(_10966_),
    .C1(_10834_),
    .C2(_10969_),
    .ZN(_10970_));
 NOR3_X4 _16793_ (.A1(_10802_),
    .A2(_10842_),
    .A3(_10962_),
    .ZN(_10971_));
 NAND2_X4 _16794_ (.A1(_10917_),
    .A2(_10967_),
    .ZN(_10972_));
 NAND2_X4 _16795_ (.A1(_10971_),
    .A2(_10972_),
    .ZN(_10973_));
 NOR3_X4 _16796_ (.A1(_10958_),
    .A2(_10970_),
    .A3(_10973_),
    .ZN(_10974_));
 INV_X2 _16797_ (.A(_00183_),
    .ZN(_10975_));
 AOI22_X2 _16798_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(_10957_),
    .B1(_10974_),
    .B2(_10975_),
    .ZN(_10976_));
 OR2_X2 _16799_ (.A1(_10818_),
    .A2(_10970_),
    .ZN(_10977_));
 BUF_X4 _16800_ (.A(_10977_),
    .Z(_10978_));
 INV_X2 _16801_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .ZN(_10979_));
 BUF_X8 _16802_ (.A(_10979_),
    .Z(_10980_));
 BUF_X8 _16803_ (.A(_10980_),
    .Z(_10981_));
 BUF_X8 _16804_ (.A(_10981_),
    .Z(_10982_));
 BUF_X8 _16805_ (.A(_10982_),
    .Z(_10983_));
 CLKBUF_X3 _16806_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .Z(_10984_));
 BUF_X4 _16807_ (.A(_10984_),
    .Z(_10985_));
 BUF_X8 _16808_ (.A(_10985_),
    .Z(_10986_));
 BUF_X8 _16809_ (.A(_10986_),
    .Z(_10987_));
 BUF_X4 _16810_ (.A(_10987_),
    .Z(_10988_));
 BUF_X4 _16811_ (.A(_10988_),
    .Z(_10989_));
 BUF_X2 _16812_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .Z(_10990_));
 INV_X2 _16813_ (.A(_10990_),
    .ZN(_10991_));
 BUF_X8 _16814_ (.A(_10991_),
    .Z(_10992_));
 BUF_X4 _16815_ (.A(_10992_),
    .Z(_10993_));
 BUF_X8 _16816_ (.A(_10993_),
    .Z(_10994_));
 BUF_X8 _16817_ (.A(_10994_),
    .Z(_10995_));
 BUF_X2 _16818_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .Z(_10996_));
 BUF_X8 _16819_ (.A(_10996_),
    .Z(_10997_));
 BUF_X8 _16820_ (.A(_10997_),
    .Z(_10998_));
 BUF_X8 _16821_ (.A(_10998_),
    .Z(_10999_));
 BUF_X4 _16822_ (.A(_10999_),
    .Z(_11000_));
 BUF_X8 _16823_ (.A(_11000_),
    .Z(_11001_));
 BUF_X4 _16824_ (.A(_11001_),
    .Z(_11002_));
 BUF_X2 _16825_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(_11003_));
 BUF_X8 _16826_ (.A(_11003_),
    .Z(_11004_));
 BUF_X4 _16827_ (.A(_11004_),
    .Z(_11005_));
 BUF_X4 _16828_ (.A(_11005_),
    .Z(_11006_));
 BUF_X4 _16829_ (.A(_11006_),
    .Z(_11007_));
 BUF_X4 _16830_ (.A(_11007_),
    .Z(_11008_));
 MUX2_X1 _16831_ (.A(_00147_),
    .B(_00149_),
    .S(_11008_),
    .Z(_11009_));
 NOR2_X1 _16832_ (.A1(_11002_),
    .A2(_11009_),
    .ZN(_11010_));
 INV_X2 _16833_ (.A(_10997_),
    .ZN(_11011_));
 BUF_X4 _16834_ (.A(_11011_),
    .Z(_11012_));
 BUF_X4 _16835_ (.A(_11012_),
    .Z(_11013_));
 BUF_X8 _16836_ (.A(_11004_),
    .Z(_11014_));
 BUF_X4 _16837_ (.A(_11014_),
    .Z(_11015_));
 BUF_X4 _16838_ (.A(_11015_),
    .Z(_11016_));
 BUF_X4 _16839_ (.A(_11016_),
    .Z(_11017_));
 MUX2_X1 _16840_ (.A(_00148_),
    .B(_00150_),
    .S(_11017_),
    .Z(_11018_));
 NOR2_X1 _16841_ (.A1(_11013_),
    .A2(_11018_),
    .ZN(_11019_));
 NOR3_X1 _16842_ (.A1(_10995_),
    .A2(_11010_),
    .A3(_11019_),
    .ZN(_11020_));
 BUF_X4 _16843_ (.A(_10990_),
    .Z(_11021_));
 BUF_X4 _16844_ (.A(_11021_),
    .Z(_11022_));
 NOR2_X1 _16845_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .A2(_11007_),
    .ZN(_11023_));
 AOI21_X1 _16846_ (.A(_11023_),
    .B1(_11017_),
    .B2(_00142_),
    .ZN(_11024_));
 BUF_X8 _16847_ (.A(_10997_),
    .Z(_11025_));
 BUF_X4 _16848_ (.A(_11025_),
    .Z(_11026_));
 BUF_X4 _16849_ (.A(_11026_),
    .Z(_11027_));
 BUF_X8 _16850_ (.A(_11027_),
    .Z(_11028_));
 INV_X2 _16851_ (.A(_11003_),
    .ZN(_11029_));
 NOR2_X4 _16852_ (.A1(_10996_),
    .A2(_11029_),
    .ZN(_11030_));
 BUF_X4 _16853_ (.A(_11030_),
    .Z(_11031_));
 BUF_X4 _16854_ (.A(_11031_),
    .Z(_11032_));
 INV_X1 _16855_ (.A(_00141_),
    .ZN(_11033_));
 AOI221_X2 _16856_ (.A(_11022_),
    .B1(_11024_),
    .B2(_11028_),
    .C1(_11032_),
    .C2(_11033_),
    .ZN(_11034_));
 NOR3_X2 _16857_ (.A1(_10989_),
    .A2(_11020_),
    .A3(_11034_),
    .ZN(_11035_));
 INV_X4 _16858_ (.A(_10985_),
    .ZN(_11036_));
 BUF_X4 _16859_ (.A(_11036_),
    .Z(_11037_));
 BUF_X8 _16860_ (.A(_11037_),
    .Z(_11038_));
 MUX2_X1 _16861_ (.A(_00151_),
    .B(_00153_),
    .S(_11016_),
    .Z(_11039_));
 MUX2_X1 _16862_ (.A(_00152_),
    .B(_00154_),
    .S(_11016_),
    .Z(_11040_));
 BUF_X8 _16863_ (.A(_11025_),
    .Z(_11041_));
 BUF_X8 _16864_ (.A(_11041_),
    .Z(_11042_));
 BUF_X8 _16865_ (.A(_11042_),
    .Z(_11043_));
 MUX2_X1 _16866_ (.A(_11039_),
    .B(_11040_),
    .S(_11043_),
    .Z(_11044_));
 MUX2_X1 _16867_ (.A(_00143_),
    .B(_00145_),
    .S(_11016_),
    .Z(_11045_));
 MUX2_X1 _16868_ (.A(_00144_),
    .B(_00146_),
    .S(_11016_),
    .Z(_11046_));
 MUX2_X1 _16869_ (.A(_11045_),
    .B(_11046_),
    .S(_11043_),
    .Z(_11047_));
 MUX2_X1 _16870_ (.A(_11044_),
    .B(_11047_),
    .S(_10994_),
    .Z(_11048_));
 NOR2_X2 _16871_ (.A1(_11038_),
    .A2(_11048_),
    .ZN(_11049_));
 OAI21_X4 _16872_ (.A(_10983_),
    .B1(_11035_),
    .B2(_11049_),
    .ZN(_11050_));
 BUF_X8 _16873_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .Z(_11051_));
 BUF_X8 _16874_ (.A(_11051_),
    .Z(_11052_));
 BUF_X8 _16875_ (.A(_11052_),
    .Z(_11053_));
 BUF_X8 _16876_ (.A(_11053_),
    .Z(_11054_));
 BUF_X8 _16877_ (.A(_11022_),
    .Z(_11055_));
 BUF_X4 _16878_ (.A(_11055_),
    .Z(_11056_));
 BUF_X8 _16879_ (.A(_10986_),
    .Z(_11057_));
 BUF_X8 _16880_ (.A(_11057_),
    .Z(_11058_));
 BUF_X8 _16881_ (.A(_11025_),
    .Z(_11059_));
 BUF_X4 _16882_ (.A(_11059_),
    .Z(_11060_));
 BUF_X4 _16883_ (.A(_11060_),
    .Z(_11061_));
 MUX2_X1 _16884_ (.A(_00165_),
    .B(_00166_),
    .S(_11061_),
    .Z(_11062_));
 BUF_X4 _16885_ (.A(_11003_),
    .Z(_11063_));
 BUF_X4 _16886_ (.A(_11063_),
    .Z(_11064_));
 BUF_X4 _16887_ (.A(_11064_),
    .Z(_11065_));
 BUF_X4 _16888_ (.A(_11065_),
    .Z(_11066_));
 BUF_X4 _16889_ (.A(_11066_),
    .Z(_11067_));
 BUF_X4 _16890_ (.A(_11067_),
    .Z(_11068_));
 BUF_X4 _16891_ (.A(_11068_),
    .Z(_11069_));
 AOI21_X2 _16892_ (.A(_11058_),
    .B1(_11062_),
    .B2(_11069_),
    .ZN(_11070_));
 MUX2_X1 _16893_ (.A(_00163_),
    .B(_00164_),
    .S(_11028_),
    .Z(_11071_));
 INV_X1 _16894_ (.A(_11071_),
    .ZN(_11072_));
 BUF_X4 _16895_ (.A(_11037_),
    .Z(_11073_));
 BUF_X4 _16896_ (.A(_11059_),
    .Z(_11074_));
 BUF_X8 _16897_ (.A(_11074_),
    .Z(_11075_));
 MUX2_X1 _16898_ (.A(_00169_),
    .B(_00170_),
    .S(_11075_),
    .Z(_11076_));
 AOI21_X2 _16899_ (.A(_11073_),
    .B1(_11076_),
    .B2(_11069_),
    .ZN(_11077_));
 MUX2_X1 _16900_ (.A(_00167_),
    .B(_00168_),
    .S(_11028_),
    .Z(_11078_));
 INV_X1 _16901_ (.A(_11078_),
    .ZN(_11079_));
 AOI22_X2 _16902_ (.A1(_11070_),
    .A2(_11072_),
    .B1(_11077_),
    .B2(_11079_),
    .ZN(_11080_));
 BUF_X8 _16903_ (.A(_11068_),
    .Z(_11081_));
 OAI21_X1 _16904_ (.A(_11081_),
    .B1(_11070_),
    .B2(_11077_),
    .ZN(_11082_));
 NAND3_X2 _16905_ (.A1(_11056_),
    .A2(_11080_),
    .A3(_11082_),
    .ZN(_11083_));
 NOR2_X2 _16906_ (.A1(_11036_),
    .A2(_11022_),
    .ZN(_11084_));
 BUF_X8 _16907_ (.A(_11084_),
    .Z(_11085_));
 MUX2_X1 _16908_ (.A(_00159_),
    .B(_00161_),
    .S(_11017_),
    .Z(_11086_));
 MUX2_X1 _16909_ (.A(_00160_),
    .B(_00162_),
    .S(_11017_),
    .Z(_11087_));
 BUF_X4 _16910_ (.A(_11043_),
    .Z(_11088_));
 MUX2_X1 _16911_ (.A(_11086_),
    .B(_11087_),
    .S(_11088_),
    .Z(_11089_));
 NOR3_X4 _16912_ (.A1(_11004_),
    .A2(_10985_),
    .A3(_10990_),
    .ZN(_11090_));
 BUF_X8 _16913_ (.A(_11090_),
    .Z(_11091_));
 BUF_X8 _16914_ (.A(_10998_),
    .Z(_11092_));
 BUF_X8 _16915_ (.A(_11092_),
    .Z(_11093_));
 BUF_X4 _16916_ (.A(_11093_),
    .Z(_11094_));
 MUX2_X1 _16917_ (.A(_00155_),
    .B(_00156_),
    .S(_11094_),
    .Z(_11095_));
 BUF_X4 _16918_ (.A(_11014_),
    .Z(_11096_));
 BUF_X4 _16919_ (.A(_11096_),
    .Z(_11097_));
 NOR2_X1 _16920_ (.A1(_10985_),
    .A2(_11021_),
    .ZN(_11098_));
 AND2_X2 _16921_ (.A1(_11097_),
    .A2(_11098_),
    .ZN(_11099_));
 BUF_X8 _16922_ (.A(_11099_),
    .Z(_11100_));
 MUX2_X1 _16923_ (.A(_00157_),
    .B(_00158_),
    .S(_11001_),
    .Z(_11101_));
 AOI222_X2 _16924_ (.A1(_11085_),
    .A2(_11089_),
    .B1(_11091_),
    .B2(_11095_),
    .C1(_11100_),
    .C2(_11101_),
    .ZN(_11102_));
 NAND3_X4 _16925_ (.A1(_11054_),
    .A2(_11083_),
    .A3(_11102_),
    .ZN(_11103_));
 AND3_X1 _16926_ (.A1(_10978_),
    .A2(_11050_),
    .A3(_11103_),
    .ZN(_11104_));
 OAI21_X1 _16927_ (.A(_10773_),
    .B1(_10928_),
    .B2(_10929_),
    .ZN(_11105_));
 AND3_X1 _16928_ (.A1(_10807_),
    .A2(_10778_),
    .A3(_10897_),
    .ZN(_11106_));
 NOR3_X1 _16929_ (.A1(_10807_),
    .A2(_10799_),
    .A3(_10800_),
    .ZN(_11107_));
 OAI21_X1 _16930_ (.A(_10834_),
    .B1(_11106_),
    .B2(_11107_),
    .ZN(_11108_));
 NOR3_X1 _16931_ (.A1(_10803_),
    .A2(_10965_),
    .A3(_10964_),
    .ZN(_11109_));
 AOI221_X2 _16932_ (.A(_11105_),
    .B1(_11108_),
    .B2(_11109_),
    .C1(_10850_),
    .C2(_10971_),
    .ZN(_11110_));
 CLKBUF_X3 _16933_ (.A(_11110_),
    .Z(_11111_));
 CLKBUF_X3 _16934_ (.A(_11111_),
    .Z(_11112_));
 CLKBUF_X3 _16935_ (.A(_11112_),
    .Z(_11113_));
 BUF_X4 _16936_ (.A(_10977_),
    .Z(_11114_));
 BUF_X4 _16937_ (.A(_11114_),
    .Z(_11115_));
 BUF_X2 _16938_ (.A(\cs_registers_i.pc_id_i[1] ),
    .Z(_11116_));
 OAI21_X2 _16939_ (.A(_11113_),
    .B1(_11115_),
    .B2(_11116_),
    .ZN(_11117_));
 OAI21_X4 _16940_ (.A(_10976_),
    .B1(_11104_),
    .B2(_11117_),
    .ZN(_16246_));
 INV_X1 _16941_ (.A(_16246_),
    .ZN(_16250_));
 OAI211_X2 _16942_ (.A(_10838_),
    .B(_10864_),
    .C1(_10854_),
    .C2(_10857_),
    .ZN(_11118_));
 AOI22_X4 _16943_ (.A1(_10844_),
    .A2(_10820_),
    .B1(_10800_),
    .B2(_10779_),
    .ZN(_11119_));
 OAI211_X4 _16944_ (.A(_11119_),
    .B(net297),
    .C1(_10811_),
    .C2(_10808_),
    .ZN(_11120_));
 BUF_X4 _16945_ (.A(_11120_),
    .Z(_11121_));
 NAND2_X2 _16946_ (.A1(_10774_),
    .A2(_11121_),
    .ZN(_11122_));
 NOR2_X1 _16947_ (.A1(_11118_),
    .A2(_11122_),
    .ZN(_11123_));
 OAI21_X1 _16948_ (.A(_10711_),
    .B1(_10819_),
    .B2(_10836_),
    .ZN(_11124_));
 NAND2_X1 _16949_ (.A1(_10838_),
    .A2(_10855_),
    .ZN(_11125_));
 OAI21_X2 _16950_ (.A(_11124_),
    .B1(_11125_),
    .B2(_00216_),
    .ZN(_11126_));
 MUX2_X1 _16951_ (.A(_00200_),
    .B(_00202_),
    .S(net379),
    .Z(_11127_));
 NOR2_X1 _16952_ (.A1(_10711_),
    .A2(_11127_),
    .ZN(_11128_));
 INV_X8 _16953_ (.A(_10708_),
    .ZN(_11129_));
 BUF_X4 _16954_ (.A(_11129_),
    .Z(_11130_));
 MUX2_X1 _16955_ (.A(_00201_),
    .B(_00203_),
    .S(net379),
    .Z(_11131_));
 NOR2_X1 _16956_ (.A1(_11130_),
    .A2(_11131_),
    .ZN(_11132_));
 NOR3_X1 _16957_ (.A1(_10764_),
    .A2(_11128_),
    .A3(_11132_),
    .ZN(_11133_));
 BUF_X8 _16958_ (.A(_10761_),
    .Z(_11134_));
 INV_X1 _16959_ (.A(_00186_),
    .ZN(_11135_));
 INV_X4 _16960_ (.A(net375),
    .ZN(_11136_));
 NOR2_X4 _16961_ (.A1(_10709_),
    .A2(_11136_),
    .ZN(_11137_));
 NOR2_X1 _16962_ (.A1(net379),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .ZN(_11138_));
 AOI21_X1 _16963_ (.A(_11138_),
    .B1(_00187_),
    .B2(net379),
    .ZN(_11139_));
 AOI221_X2 _16964_ (.A(_11134_),
    .B1(_11135_),
    .B2(_11137_),
    .C1(_11139_),
    .C2(_10711_),
    .ZN(_11140_));
 NOR3_X1 _16965_ (.A1(_10731_),
    .A2(_11133_),
    .A3(_11140_),
    .ZN(_11141_));
 MUX2_X1 _16966_ (.A(_00204_),
    .B(_00206_),
    .S(_10737_),
    .Z(_11142_));
 MUX2_X1 _16967_ (.A(_00205_),
    .B(_00207_),
    .S(_10737_),
    .Z(_11143_));
 MUX2_X1 _16968_ (.A(_11142_),
    .B(_11143_),
    .S(_10711_),
    .Z(_11144_));
 MUX2_X1 _16969_ (.A(_00188_),
    .B(_00190_),
    .S(_10737_),
    .Z(_11145_));
 MUX2_X1 _16970_ (.A(_00189_),
    .B(_00191_),
    .S(_10737_),
    .Z(_11146_));
 MUX2_X1 _16971_ (.A(_11145_),
    .B(_11146_),
    .S(_10711_),
    .Z(_11147_));
 MUX2_X1 _16972_ (.A(_11144_),
    .B(_11147_),
    .S(_10764_),
    .Z(_11148_));
 NOR2_X2 _16973_ (.A1(_10736_),
    .A2(_11148_),
    .ZN(_11149_));
 NOR3_X2 _16974_ (.A1(_10758_),
    .A2(_11141_),
    .A3(_11149_),
    .ZN(_11150_));
 MUX2_X1 _16975_ (.A(_00208_),
    .B(_00210_),
    .S(_10748_),
    .Z(_11151_));
 MUX2_X1 _16976_ (.A(_00209_),
    .B(_00211_),
    .S(_10748_),
    .Z(_11152_));
 MUX2_X1 _16977_ (.A(_11151_),
    .B(_11152_),
    .S(_10712_),
    .Z(_11153_));
 MUX2_X1 _16978_ (.A(_00192_),
    .B(_00194_),
    .S(_10748_),
    .Z(_11154_));
 MUX2_X1 _16979_ (.A(_00193_),
    .B(_00195_),
    .S(_10748_),
    .Z(_11155_));
 MUX2_X1 _16980_ (.A(_11154_),
    .B(_11155_),
    .S(_10712_),
    .Z(_11156_));
 MUX2_X1 _16981_ (.A(_11153_),
    .B(_11156_),
    .S(_10764_),
    .Z(_11157_));
 MUX2_X1 _16982_ (.A(_00212_),
    .B(_00214_),
    .S(_10748_),
    .Z(_11158_));
 MUX2_X1 _16983_ (.A(_00213_),
    .B(_00215_),
    .S(_10748_),
    .Z(_11159_));
 MUX2_X1 _16984_ (.A(_11158_),
    .B(_11159_),
    .S(_10712_),
    .Z(_11160_));
 MUX2_X1 _16985_ (.A(_00196_),
    .B(_00198_),
    .S(_10748_),
    .Z(_11161_));
 MUX2_X1 _16986_ (.A(_00197_),
    .B(_00199_),
    .S(_10748_),
    .Z(_11162_));
 MUX2_X1 _16987_ (.A(_11161_),
    .B(_11162_),
    .S(_10712_),
    .Z(_11163_));
 MUX2_X1 _16988_ (.A(_11160_),
    .B(_11163_),
    .S(_10764_),
    .Z(_11164_));
 MUX2_X1 _16989_ (.A(_11157_),
    .B(_11164_),
    .S(_10731_),
    .Z(_11165_));
 AOI21_X4 _16990_ (.A(_11150_),
    .B1(_10758_),
    .B2(_11165_),
    .ZN(_11166_));
 NOR2_X4 _16991_ (.A1(_10818_),
    .A2(_11120_),
    .ZN(_11167_));
 BUF_X8 _16992_ (.A(_11167_),
    .Z(_11168_));
 AOI22_X4 _16993_ (.A1(_11123_),
    .A2(_11126_),
    .B1(_11166_),
    .B2(_11168_),
    .ZN(_11169_));
 INV_X2 _16994_ (.A(_11169_),
    .ZN(_11170_));
 CLKBUF_X3 _16995_ (.A(_11170_),
    .Z(_11171_));
 BUF_X4 _16996_ (.A(_11171_),
    .Z(_16242_));
 BUF_X4 _16997_ (.A(_11169_),
    .Z(_11172_));
 BUF_X8 _16998_ (.A(_11172_),
    .Z(_11173_));
 BUF_X1 rebuffer32 (.A(_10893_),
    .Z(net306));
 BUF_X4 _17000_ (.A(_11037_),
    .Z(_11174_));
 MUX2_X1 _17001_ (.A(_00214_),
    .B(_00215_),
    .S(_11028_),
    .Z(_11175_));
 AOI21_X1 _17002_ (.A(_11174_),
    .B1(_11175_),
    .B2(_11081_),
    .ZN(_11176_));
 BUF_X4 _17003_ (.A(_11057_),
    .Z(_11177_));
 MUX2_X1 _17004_ (.A(_00210_),
    .B(_00211_),
    .S(_11028_),
    .Z(_11178_));
 AOI21_X1 _17005_ (.A(_11177_),
    .B1(_11178_),
    .B2(_11069_),
    .ZN(_11179_));
 OAI21_X1 _17006_ (.A(_11081_),
    .B1(_11176_),
    .B2(_11179_),
    .ZN(_11180_));
 NAND2_X1 _17007_ (.A1(_11013_),
    .A2(_00208_),
    .ZN(_11181_));
 NAND2_X1 _17008_ (.A1(_11002_),
    .A2(_00209_),
    .ZN(_11182_));
 NAND3_X1 _17009_ (.A1(_11179_),
    .A2(_11181_),
    .A3(_11182_),
    .ZN(_11183_));
 NAND2_X1 _17010_ (.A1(_11013_),
    .A2(_00212_),
    .ZN(_11184_));
 NAND2_X1 _17011_ (.A1(_11002_),
    .A2(_00213_),
    .ZN(_11185_));
 NAND3_X1 _17012_ (.A1(_11176_),
    .A2(_11184_),
    .A3(_11185_),
    .ZN(_11186_));
 NAND4_X2 _17013_ (.A1(_11056_),
    .A2(_11180_),
    .A3(_11183_),
    .A4(_11186_),
    .ZN(_11187_));
 BUF_X4 _17014_ (.A(_11067_),
    .Z(_11188_));
 MUX2_X1 _17015_ (.A(_00204_),
    .B(_00206_),
    .S(_11188_),
    .Z(_11189_));
 MUX2_X1 _17016_ (.A(_00205_),
    .B(_00207_),
    .S(_11188_),
    .Z(_11190_));
 MUX2_X1 _17017_ (.A(_11189_),
    .B(_11190_),
    .S(_11002_),
    .Z(_11191_));
 MUX2_X1 _17018_ (.A(_00200_),
    .B(_00201_),
    .S(_11088_),
    .Z(_11192_));
 MUX2_X1 _17019_ (.A(_00202_),
    .B(_00203_),
    .S(_11094_),
    .Z(_11193_));
 AOI222_X2 _17020_ (.A1(_11191_),
    .A2(_11085_),
    .B1(_11192_),
    .B2(_11091_),
    .C1(_11193_),
    .C2(_11100_),
    .ZN(_11194_));
 NAND3_X4 _17021_ (.A1(_11054_),
    .A2(_11187_),
    .A3(_11194_),
    .ZN(_11195_));
 MUX2_X1 _17022_ (.A(_00192_),
    .B(_00194_),
    .S(_11067_),
    .Z(_11196_));
 MUX2_X1 _17023_ (.A(_00193_),
    .B(_00195_),
    .S(_11067_),
    .Z(_11197_));
 MUX2_X1 _17024_ (.A(_11196_),
    .B(_11197_),
    .S(_11001_),
    .Z(_11198_));
 NOR2_X1 _17025_ (.A1(_11008_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .ZN(_11199_));
 AOI21_X1 _17026_ (.A(_11199_),
    .B1(_00187_),
    .B2(_11068_),
    .ZN(_11200_));
 AOI22_X1 _17027_ (.A1(_11135_),
    .A2(_11032_),
    .B1(_11200_),
    .B2(_11088_),
    .ZN(_11201_));
 MUX2_X1 _17028_ (.A(_11198_),
    .B(_11201_),
    .S(_10994_),
    .Z(_11202_));
 MUX2_X1 _17029_ (.A(_00196_),
    .B(_00198_),
    .S(_11067_),
    .Z(_11203_));
 MUX2_X1 _17030_ (.A(_00197_),
    .B(_00199_),
    .S(_11067_),
    .Z(_11204_));
 MUX2_X1 _17031_ (.A(_11203_),
    .B(_11204_),
    .S(_11001_),
    .Z(_11205_));
 MUX2_X1 _17032_ (.A(_00188_),
    .B(_00190_),
    .S(_11067_),
    .Z(_11206_));
 BUF_X4 _17033_ (.A(_11064_),
    .Z(_11207_));
 BUF_X4 _17034_ (.A(_11207_),
    .Z(_11208_));
 BUF_X4 _17035_ (.A(_11208_),
    .Z(_11209_));
 MUX2_X1 _17036_ (.A(_00189_),
    .B(_00191_),
    .S(_11209_),
    .Z(_11210_));
 MUX2_X1 _17037_ (.A(_11206_),
    .B(_11210_),
    .S(_11001_),
    .Z(_11211_));
 MUX2_X1 _17038_ (.A(_11205_),
    .B(_11211_),
    .S(_10994_),
    .Z(_11212_));
 MUX2_X2 _17039_ (.A(_11202_),
    .B(_11212_),
    .S(_10989_),
    .Z(_11213_));
 OAI211_X2 _17040_ (.A(_11113_),
    .B(_11195_),
    .C1(_11213_),
    .C2(_11054_),
    .ZN(_11214_));
 NOR2_X4 _17041_ (.A1(_10818_),
    .A2(_10970_),
    .ZN(_11215_));
 INV_X1 _17042_ (.A(_11111_),
    .ZN(_11216_));
 INV_X1 _17043_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .ZN(_11217_));
 AOI21_X2 _17044_ (.A(_11215_),
    .B1(_11216_),
    .B2(_11217_),
    .ZN(_11218_));
 NOR2_X1 _17045_ (.A1(_00184_),
    .A2(_11113_),
    .ZN(_11219_));
 AOI22_X4 _17046_ (.A1(_11214_),
    .A2(_11218_),
    .B1(_11219_),
    .B2(_10974_),
    .ZN(_16239_));
 BUF_X4 _17047_ (.A(_15774_),
    .Z(_11220_));
 XOR2_X2 _17048_ (.A(_14467_),
    .B(_11220_),
    .Z(\alu_adder_result_ex[1] ));
 INV_X4 _17049_ (.A(\alu_adder_result_ex[1] ),
    .ZN(_16491_));
 CLKBUF_X3 _17050_ (.A(_10819_),
    .Z(_11221_));
 NAND2_X1 _17051_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(_11221_),
    .ZN(_11222_));
 BUF_X4 _17052_ (.A(_11037_),
    .Z(_11223_));
 BUF_X4 _17053_ (.A(_11064_),
    .Z(_11224_));
 MUX2_X1 _17054_ (.A(_00228_),
    .B(_00230_),
    .S(_11224_),
    .Z(_11225_));
 MUX2_X1 _17055_ (.A(_00229_),
    .B(_00231_),
    .S(_11224_),
    .Z(_11226_));
 BUF_X8 _17056_ (.A(_11025_),
    .Z(_11227_));
 MUX2_X1 _17057_ (.A(_11225_),
    .B(_11226_),
    .S(_11227_),
    .Z(_11228_));
 MUX2_X1 _17058_ (.A(_00220_),
    .B(_00222_),
    .S(_11224_),
    .Z(_11229_));
 MUX2_X1 _17059_ (.A(_00221_),
    .B(_00223_),
    .S(_11065_),
    .Z(_11230_));
 MUX2_X1 _17060_ (.A(_11229_),
    .B(_11230_),
    .S(_11227_),
    .Z(_11231_));
 BUF_X4 _17061_ (.A(_10992_),
    .Z(_11232_));
 MUX2_X1 _17062_ (.A(_11228_),
    .B(_11231_),
    .S(_11232_),
    .Z(_11233_));
 NOR2_X1 _17063_ (.A1(_11223_),
    .A2(_11233_),
    .ZN(_11234_));
 BUF_X4 _17064_ (.A(_11021_),
    .Z(_11235_));
 INV_X1 _17065_ (.A(_00218_),
    .ZN(_11236_));
 NOR2_X1 _17066_ (.A1(_11006_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .ZN(_11237_));
 BUF_X4 _17067_ (.A(_11003_),
    .Z(_11238_));
 BUF_X4 _17068_ (.A(_11238_),
    .Z(_11239_));
 BUF_X4 _17069_ (.A(_11239_),
    .Z(_11240_));
 BUF_X4 _17070_ (.A(_11240_),
    .Z(_11241_));
 AOI21_X1 _17071_ (.A(_11237_),
    .B1(_00219_),
    .B2(_11241_),
    .ZN(_11242_));
 AOI221_X2 _17072_ (.A(_11235_),
    .B1(_11236_),
    .B2(_11031_),
    .C1(_11242_),
    .C2(_11042_),
    .ZN(_11243_));
 BUF_X4 _17073_ (.A(_11238_),
    .Z(_11244_));
 BUF_X4 _17074_ (.A(_11244_),
    .Z(_11245_));
 BUF_X4 _17075_ (.A(_11245_),
    .Z(_11246_));
 MUX2_X1 _17076_ (.A(_00224_),
    .B(_00226_),
    .S(_11246_),
    .Z(_11247_));
 MUX2_X1 _17077_ (.A(_00225_),
    .B(_00227_),
    .S(_11246_),
    .Z(_11248_));
 MUX2_X1 _17078_ (.A(_11247_),
    .B(_11248_),
    .S(_11075_),
    .Z(_11249_));
 AOI21_X1 _17079_ (.A(_11243_),
    .B1(_11249_),
    .B2(_11022_),
    .ZN(_11250_));
 AOI21_X2 _17080_ (.A(_11234_),
    .B1(_11250_),
    .B2(_11038_),
    .ZN(_11251_));
 BUF_X4 _17081_ (.A(_11022_),
    .Z(_11252_));
 MUX2_X1 _17082_ (.A(_00242_),
    .B(_00243_),
    .S(_11041_),
    .Z(_11253_));
 BUF_X4 _17083_ (.A(_11241_),
    .Z(_11254_));
 AOI21_X2 _17084_ (.A(_10986_),
    .B1(_11253_),
    .B2(_11254_),
    .ZN(_11255_));
 BUF_X4 _17085_ (.A(_10998_),
    .Z(_11256_));
 MUX2_X1 _17086_ (.A(_00246_),
    .B(_00247_),
    .S(_11256_),
    .Z(_11257_));
 AOI21_X2 _17087_ (.A(_11036_),
    .B1(_11257_),
    .B2(_11008_),
    .ZN(_11258_));
 OAI21_X1 _17088_ (.A(_11068_),
    .B1(_11255_),
    .B2(_11258_),
    .ZN(_11259_));
 BUF_X4 _17089_ (.A(_11059_),
    .Z(_11260_));
 MUX2_X1 _17090_ (.A(_00244_),
    .B(_00245_),
    .S(_11260_),
    .Z(_11261_));
 INV_X1 _17091_ (.A(_11261_),
    .ZN(_11262_));
 MUX2_X1 _17092_ (.A(_00240_),
    .B(_00241_),
    .S(_11092_),
    .Z(_11263_));
 INV_X1 _17093_ (.A(_11263_),
    .ZN(_11264_));
 AOI22_X2 _17094_ (.A1(_11258_),
    .A2(_11262_),
    .B1(_11264_),
    .B2(_11255_),
    .ZN(_11265_));
 NAND3_X2 _17095_ (.A1(_11252_),
    .A2(_11259_),
    .A3(_11265_),
    .ZN(_11266_));
 MUX2_X1 _17096_ (.A(_00236_),
    .B(_00238_),
    .S(_11066_),
    .Z(_11267_));
 MUX2_X1 _17097_ (.A(_00237_),
    .B(_00239_),
    .S(_11066_),
    .Z(_11268_));
 BUF_X4 _17098_ (.A(_11227_),
    .Z(_11269_));
 MUX2_X1 _17099_ (.A(_11267_),
    .B(_11268_),
    .S(_11269_),
    .Z(_11270_));
 BUF_X4 _17100_ (.A(_11041_),
    .Z(_11271_));
 MUX2_X1 _17101_ (.A(_00234_),
    .B(_00235_),
    .S(_11271_),
    .Z(_11272_));
 MUX2_X1 _17102_ (.A(_00232_),
    .B(_00233_),
    .S(_11260_),
    .Z(_11273_));
 AOI222_X2 _17103_ (.A1(_11084_),
    .A2(_11270_),
    .B1(_11272_),
    .B2(_11099_),
    .C1(_11273_),
    .C2(_11090_),
    .ZN(_11274_));
 NAND2_X1 _17104_ (.A1(_11266_),
    .A2(_11274_),
    .ZN(_11275_));
 MUX2_X2 _17105_ (.A(_11251_),
    .B(_11275_),
    .S(_11053_),
    .Z(_11276_));
 NAND2_X2 _17106_ (.A1(_10977_),
    .A2(_11111_),
    .ZN(_11277_));
 BUF_X4 _17107_ (.A(_11277_),
    .Z(_11278_));
 NAND2_X1 _17108_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_11112_),
    .ZN(_11279_));
 OAI221_X2 _17109_ (.A(_11222_),
    .B1(_11276_),
    .B2(_11278_),
    .C1(_11279_),
    .C2(_11114_),
    .ZN(_16333_));
 INV_X1 _17110_ (.A(_16333_),
    .ZN(_16337_));
 OR3_X4 _17111_ (.A1(_10802_),
    .A2(_10842_),
    .A3(_10962_),
    .ZN(_11280_));
 NOR2_X2 _17112_ (.A1(_11280_),
    .A2(_10968_),
    .ZN(_11281_));
 BUF_X4 _17113_ (.A(_11281_),
    .Z(_11282_));
 NOR2_X1 _17114_ (.A1(_10928_),
    .A2(_10929_),
    .ZN(_11283_));
 NOR3_X1 _17115_ (.A1(_10809_),
    .A2(_10808_),
    .A3(_10968_),
    .ZN(_11284_));
 OR3_X2 _17116_ (.A1(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .A2(_11283_),
    .A3(_11284_),
    .ZN(_11285_));
 NAND3_X2 _17117_ (.A1(_10874_),
    .A2(_10877_),
    .A3(_10879_),
    .ZN(_11286_));
 NAND2_X1 _17118_ (.A1(net329),
    .A2(_10888_),
    .ZN(_11287_));
 NOR3_X1 _17119_ (.A1(_10921_),
    .A2(_11286_),
    .A3(_11287_),
    .ZN(_11288_));
 NOR3_X2 _17120_ (.A1(_10872_),
    .A2(net305),
    .A3(_11288_),
    .ZN(_11289_));
 OAI21_X1 _17121_ (.A(_10849_),
    .B1(_10912_),
    .B2(_10785_),
    .ZN(_11290_));
 AOI22_X2 _17122_ (.A1(_10785_),
    .A2(_10850_),
    .B1(_11290_),
    .B2(_10881_),
    .ZN(_11291_));
 OAI33_X1 _17123_ (.A1(_10921_),
    .A2(_00175_),
    .A3(_10823_),
    .B1(_11291_),
    .B2(_10778_),
    .B3(_10779_),
    .ZN(_11292_));
 NOR2_X4 _17124_ (.A1(_10802_),
    .A2(_10842_),
    .ZN(_11293_));
 AOI211_X2 _17125_ (.A(_11285_),
    .B(_11289_),
    .C1(_11292_),
    .C2(_11293_),
    .ZN(_11294_));
 NOR2_X2 _17126_ (.A1(_10945_),
    .A2(_10869_),
    .ZN(_11295_));
 NAND4_X2 _17127_ (.A1(_10900_),
    .A2(_00177_),
    .A3(_10901_),
    .A4(_11295_),
    .ZN(_11296_));
 NAND4_X2 _17128_ (.A1(_10888_),
    .A2(_10900_),
    .A3(net294),
    .A4(_11295_),
    .ZN(_11297_));
 AOI22_X4 _17129_ (.A1(_10903_),
    .A2(_11296_),
    .B1(_11297_),
    .B2(_10917_),
    .ZN(_11298_));
 NOR4_X4 _17130_ (.A1(_10893_),
    .A2(_10939_),
    .A3(_10898_),
    .A4(_11298_),
    .ZN(_11299_));
 NOR2_X1 _17131_ (.A1(_11280_),
    .A2(_10967_),
    .ZN(_11300_));
 NOR3_X2 _17132_ (.A1(_10937_),
    .A2(_10933_),
    .A3(_11300_),
    .ZN(_11301_));
 NOR4_X4 _17133_ (.A1(_10761_),
    .A2(_10945_),
    .A3(_10873_),
    .A4(_10884_),
    .ZN(_11302_));
 AND4_X2 _17134_ (.A1(_10761_),
    .A2(_10945_),
    .A3(_10873_),
    .A4(_10884_),
    .ZN(_11303_));
 OAI21_X4 _17135_ (.A(net300),
    .B1(_11302_),
    .B2(_11303_),
    .ZN(_11304_));
 NAND3_X4 _17136_ (.A1(_11011_),
    .A2(_00180_),
    .A3(_11090_),
    .ZN(_11305_));
 BUF_X4 _17137_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .Z(_11306_));
 INV_X4 _17138_ (.A(_11306_),
    .ZN(_11307_));
 BUF_X4 _17139_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .Z(_11308_));
 BUF_X4 _17140_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .Z(_11309_));
 CLKBUF_X3 _17141_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .Z(_11310_));
 NOR3_X4 _17142_ (.A1(_11308_),
    .A2(_11309_),
    .A3(_11310_),
    .ZN(_11311_));
 NAND4_X2 _17143_ (.A1(_10917_),
    .A2(_10863_),
    .A3(_11307_),
    .A4(_11311_),
    .ZN(_11312_));
 NOR4_X2 _17144_ (.A1(_11280_),
    .A2(_11304_),
    .A3(_11305_),
    .A4(_11312_),
    .ZN(_11313_));
 INV_X1 _17145_ (.A(_10875_),
    .ZN(_11314_));
 BUF_X4 _17146_ (.A(_10709_),
    .Z(_11315_));
 BUF_X4 _17147_ (.A(_11315_),
    .Z(_11316_));
 NAND3_X4 _17148_ (.A1(_11316_),
    .A2(_10730_),
    .A3(_10876_),
    .ZN(_11317_));
 OAI21_X1 _17149_ (.A(_11317_),
    .B1(_10876_),
    .B2(_10730_),
    .ZN(_11318_));
 AND2_X2 _17150_ (.A1(net300),
    .A2(_11302_),
    .ZN(_11319_));
 NOR2_X2 _17151_ (.A1(_10748_),
    .A2(_10746_),
    .ZN(_11320_));
 AND4_X1 _17152_ (.A1(_11314_),
    .A2(_11318_),
    .A3(_11319_),
    .A4(_11320_),
    .ZN(_11321_));
 OR2_X2 _17153_ (.A1(_10730_),
    .A2(_10746_),
    .ZN(_11322_));
 NAND2_X2 _17154_ (.A1(_10875_),
    .A2(_10876_),
    .ZN(_11323_));
 NOR4_X4 _17155_ (.A1(_10711_),
    .A2(_11136_),
    .A3(_11322_),
    .A4(_11323_),
    .ZN(_11324_));
 OAI21_X2 _17156_ (.A(_11313_),
    .B1(_11321_),
    .B2(_11324_),
    .ZN(_11325_));
 AOI21_X4 _17157_ (.A(_11299_),
    .B1(_11301_),
    .B2(_11325_),
    .ZN(_11326_));
 AND3_X1 _17158_ (.A1(_11282_),
    .A2(_11294_),
    .A3(_11326_),
    .ZN(_11327_));
 BUF_X4 _17159_ (.A(_11327_),
    .Z(_11328_));
 BUF_X4 _17160_ (.A(_11328_),
    .Z(_11329_));
 NAND2_X2 _17161_ (.A1(_16242_),
    .A2(_11329_),
    .ZN(_15919_));
 NAND2_X2 _17162_ (.A1(_16247_),
    .A2(_11329_),
    .ZN(_15913_));
 INV_X1 _17163_ (.A(_15913_),
    .ZN(_15916_));
 INV_X1 _17164_ (.A(_11309_),
    .ZN(_11330_));
 NOR3_X2 _17165_ (.A1(_11330_),
    .A2(_10859_),
    .A3(_10866_),
    .ZN(_11331_));
 NAND2_X1 _17166_ (.A1(_11120_),
    .A2(_10865_),
    .ZN(_11332_));
 NAND4_X2 _17167_ (.A1(_00278_),
    .A2(_10773_),
    .A3(_10855_),
    .A4(_10858_),
    .ZN(_11333_));
 OAI21_X1 _17168_ (.A(_10731_),
    .B1(_10818_),
    .B2(_10836_),
    .ZN(_11334_));
 AOI21_X1 _17169_ (.A(_11332_),
    .B1(_11333_),
    .B2(_11334_),
    .ZN(_11335_));
 MUX2_X1 _17170_ (.A(_00274_),
    .B(_00276_),
    .S(_10699_),
    .Z(_11336_));
 MUX2_X1 _17171_ (.A(_00275_),
    .B(_00277_),
    .S(_10699_),
    .Z(_11337_));
 MUX2_X1 _17172_ (.A(_11336_),
    .B(_11337_),
    .S(_10708_),
    .Z(_11338_));
 MUX2_X1 _17173_ (.A(_00258_),
    .B(_00260_),
    .S(_10699_),
    .Z(_11339_));
 MUX2_X1 _17174_ (.A(_00259_),
    .B(_00261_),
    .S(_10700_),
    .Z(_11340_));
 MUX2_X1 _17175_ (.A(_11339_),
    .B(_11340_),
    .S(_10708_),
    .Z(_11341_));
 MUX2_X1 _17176_ (.A(_11338_),
    .B(_11341_),
    .S(_10762_),
    .Z(_11342_));
 AND3_X1 _17177_ (.A1(_10729_),
    .A2(_10717_),
    .A3(_11342_),
    .ZN(_11343_));
 NOR2_X2 _17178_ (.A1(_10734_),
    .A2(_10717_),
    .ZN(_11344_));
 MUX2_X1 _17179_ (.A(_00266_),
    .B(_00268_),
    .S(_10700_),
    .Z(_11345_));
 MUX2_X1 _17180_ (.A(_00267_),
    .B(_00269_),
    .S(_10700_),
    .Z(_11346_));
 MUX2_X1 _17181_ (.A(_11345_),
    .B(_11346_),
    .S(_10708_),
    .Z(_11347_));
 MUX2_X1 _17182_ (.A(_00250_),
    .B(_00252_),
    .S(net375),
    .Z(_11348_));
 MUX2_X1 _17183_ (.A(_00251_),
    .B(_00253_),
    .S(net375),
    .Z(_11349_));
 MUX2_X1 _17184_ (.A(_11348_),
    .B(_11349_),
    .S(_10708_),
    .Z(_11350_));
 MUX2_X1 _17185_ (.A(_11347_),
    .B(_11350_),
    .S(_10762_),
    .Z(_11351_));
 BUF_X4 _17186_ (.A(_10701_),
    .Z(_11352_));
 NAND2_X2 _17187_ (.A1(_11129_),
    .A2(_11352_),
    .ZN(_11353_));
 BUF_X8 _17188_ (.A(_10700_),
    .Z(_11354_));
 BUF_X4 _17189_ (.A(_11354_),
    .Z(_11355_));
 NAND2_X1 _17190_ (.A1(_11355_),
    .A2(_00249_),
    .ZN(_11356_));
 BUF_X4 _17191_ (.A(_11354_),
    .Z(_11357_));
 OAI21_X1 _17192_ (.A(_11356_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .B2(_11357_),
    .ZN(_11358_));
 OAI221_X2 _17193_ (.A(_10763_),
    .B1(_00248_),
    .B2(_11353_),
    .C1(_11358_),
    .C2(_11129_),
    .ZN(_11359_));
 MUX2_X1 _17194_ (.A(_00262_),
    .B(_00264_),
    .S(net375),
    .Z(_11360_));
 MUX2_X1 _17195_ (.A(_00263_),
    .B(_00265_),
    .S(net375),
    .Z(_11361_));
 MUX2_X1 _17196_ (.A(_11360_),
    .B(_11361_),
    .S(_10708_),
    .Z(_11362_));
 AOI21_X1 _17197_ (.A(_10717_),
    .B1(_10761_),
    .B2(_11362_),
    .ZN(_11363_));
 AOI21_X1 _17198_ (.A(_10729_),
    .B1(_11359_),
    .B2(_11363_),
    .ZN(_11364_));
 MUX2_X1 _17199_ (.A(_00270_),
    .B(_00272_),
    .S(_10701_),
    .Z(_11365_));
 MUX2_X1 _17200_ (.A(_00271_),
    .B(_00273_),
    .S(_10701_),
    .Z(_11366_));
 MUX2_X1 _17201_ (.A(_11365_),
    .B(_11366_),
    .S(_10709_),
    .Z(_11367_));
 NAND2_X1 _17202_ (.A1(_10761_),
    .A2(_11367_),
    .ZN(_11368_));
 MUX2_X1 _17203_ (.A(_00254_),
    .B(_00256_),
    .S(_10701_),
    .Z(_11369_));
 MUX2_X1 _17204_ (.A(_00255_),
    .B(_00257_),
    .S(_10701_),
    .Z(_11370_));
 MUX2_X1 _17205_ (.A(_11369_),
    .B(_11370_),
    .S(_10708_),
    .Z(_11371_));
 NAND2_X1 _17206_ (.A1(_10763_),
    .A2(_11371_),
    .ZN(_11372_));
 NAND3_X1 _17207_ (.A1(_10717_),
    .A2(_11368_),
    .A3(_11372_),
    .ZN(_11373_));
 AOI221_X2 _17208_ (.A(_11343_),
    .B1(_11344_),
    .B2(_11351_),
    .C1(_11364_),
    .C2(_11373_),
    .ZN(_11374_));
 BUF_X4 _17209_ (.A(_11374_),
    .Z(_11375_));
 AND2_X1 _17210_ (.A1(_10804_),
    .A2(_11375_),
    .ZN(_11376_));
 OR4_X1 _17211_ (.A1(_10818_),
    .A2(_11331_),
    .A3(_11335_),
    .A4(_11376_),
    .ZN(_11377_));
 BUF_X8 _17212_ (.A(_11377_),
    .Z(_16253_));
 INV_X4 _17213_ (.A(_16253_),
    .ZN(_11378_));
 BUF_X8 _17214_ (.A(_11378_),
    .Z(_11379_));
 BUF_X1 rebuffer146 (.A(\alu_adder_result_ex[15] ),
    .Z(net437));
 NAND3_X4 _17216_ (.A1(_11129_),
    .A2(_10729_),
    .A3(_10718_),
    .ZN(_11380_));
 MUX2_X1 _17217_ (.A(_00281_),
    .B(_00283_),
    .S(_11357_),
    .Z(_11381_));
 INV_X1 _17218_ (.A(_11381_),
    .ZN(_11382_));
 NAND3_X4 _17219_ (.A1(_10709_),
    .A2(_10733_),
    .A3(_10718_),
    .ZN(_11383_));
 MUX2_X1 _17220_ (.A(_00282_),
    .B(_00284_),
    .S(_11357_),
    .Z(_11384_));
 INV_X1 _17221_ (.A(_11384_),
    .ZN(_11385_));
 OAI22_X4 _17222_ (.A1(_11380_),
    .A2(_11382_),
    .B1(_11383_),
    .B2(_11385_),
    .ZN(_11386_));
 BUF_X4 _17223_ (.A(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(_11387_));
 NOR2_X2 _17224_ (.A1(_11387_),
    .A2(_10717_),
    .ZN(_11388_));
 NOR2_X4 _17225_ (.A1(_10761_),
    .A2(_11388_),
    .ZN(_11389_));
 NOR2_X4 _17226_ (.A1(_11129_),
    .A2(_10761_),
    .ZN(_11390_));
 NOR2_X1 _17227_ (.A1(net380),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .ZN(_11391_));
 AOI21_X1 _17228_ (.A(_11391_),
    .B1(_00280_),
    .B2(_11357_),
    .ZN(_11392_));
 NOR3_X4 _17229_ (.A1(_10708_),
    .A2(_11136_),
    .A3(_10761_),
    .ZN(_11393_));
 INV_X1 _17230_ (.A(_00279_),
    .ZN(_11394_));
 AOI221_X2 _17231_ (.A(_11389_),
    .B1(_11390_),
    .B2(_11392_),
    .C1(_11393_),
    .C2(_11394_),
    .ZN(_11395_));
 CLKBUF_X3 _17232_ (.A(_11387_),
    .Z(_11396_));
 MUX2_X1 _17233_ (.A(_00286_),
    .B(_00290_),
    .S(_11396_),
    .Z(_11397_));
 MUX2_X1 _17234_ (.A(_00288_),
    .B(_00292_),
    .S(_11396_),
    .Z(_11398_));
 BUF_X4 _17235_ (.A(_11354_),
    .Z(_11399_));
 BUF_X4 _17236_ (.A(_11399_),
    .Z(_11400_));
 MUX2_X1 _17237_ (.A(_11397_),
    .B(_11398_),
    .S(_11400_),
    .Z(_11401_));
 MUX2_X1 _17238_ (.A(_00285_),
    .B(_00289_),
    .S(_11396_),
    .Z(_11402_));
 MUX2_X1 _17239_ (.A(_00287_),
    .B(_00291_),
    .S(_11396_),
    .Z(_11403_));
 MUX2_X1 _17240_ (.A(_11402_),
    .B(_11403_),
    .S(_11400_),
    .Z(_11404_));
 BUF_X4 _17241_ (.A(_11129_),
    .Z(_11405_));
 MUX2_X1 _17242_ (.A(_11401_),
    .B(_11404_),
    .S(_11405_),
    .Z(_11406_));
 NOR3_X4 _17243_ (.A1(_11386_),
    .A2(_11395_),
    .A3(_11406_),
    .ZN(_11407_));
 NAND2_X4 _17244_ (.A1(_10717_),
    .A2(_10761_),
    .ZN(_11408_));
 MUX2_X1 _17245_ (.A(_00305_),
    .B(_00307_),
    .S(_11352_),
    .Z(_11409_));
 MUX2_X1 _17246_ (.A(_00306_),
    .B(_00308_),
    .S(_11352_),
    .Z(_11410_));
 MUX2_X1 _17247_ (.A(_11409_),
    .B(_11410_),
    .S(_11315_),
    .Z(_11411_));
 MUX2_X1 _17248_ (.A(_00301_),
    .B(_00303_),
    .S(_11352_),
    .Z(_11412_));
 MUX2_X1 _17249_ (.A(_00302_),
    .B(_00304_),
    .S(_11352_),
    .Z(_11413_));
 MUX2_X1 _17250_ (.A(_11412_),
    .B(_11413_),
    .S(_11315_),
    .Z(_11414_));
 MUX2_X1 _17251_ (.A(_11411_),
    .B(_11414_),
    .S(_10735_),
    .Z(_11415_));
 NOR2_X2 _17252_ (.A1(_11408_),
    .A2(_11415_),
    .ZN(_11416_));
 MUX2_X1 _17253_ (.A(_00294_),
    .B(_00298_),
    .S(_11396_),
    .Z(_11417_));
 MUX2_X1 _17254_ (.A(_00296_),
    .B(_00300_),
    .S(_11396_),
    .Z(_11418_));
 MUX2_X1 _17255_ (.A(_11417_),
    .B(_11418_),
    .S(_11400_),
    .Z(_11419_));
 MUX2_X1 _17256_ (.A(_00293_),
    .B(_00297_),
    .S(_11396_),
    .Z(_11420_));
 MUX2_X1 _17257_ (.A(_00295_),
    .B(_00299_),
    .S(_11396_),
    .Z(_11421_));
 MUX2_X1 _17258_ (.A(_11420_),
    .B(_11421_),
    .S(_11400_),
    .Z(_11422_));
 MUX2_X1 _17259_ (.A(_11419_),
    .B(_11422_),
    .S(_11405_),
    .Z(_11423_));
 NAND2_X4 _17260_ (.A1(_10718_),
    .A2(_11134_),
    .ZN(_11424_));
 NOR2_X2 _17261_ (.A1(_11423_),
    .A2(_11424_),
    .ZN(_11425_));
 NOR3_X4 _17262_ (.A1(_10746_),
    .A2(_11386_),
    .A3(_11395_),
    .ZN(_11426_));
 OR4_X4 _17263_ (.A1(_11407_),
    .A2(_11416_),
    .A3(_11425_),
    .A4(_11426_),
    .ZN(_11427_));
 INV_X1 _17264_ (.A(_11308_),
    .ZN(_11428_));
 NOR3_X1 _17265_ (.A1(_11428_),
    .A2(_10859_),
    .A3(_10866_),
    .ZN(_11429_));
 OAI21_X1 _17266_ (.A(_10865_),
    .B1(_10836_),
    .B2(_10818_),
    .ZN(_11430_));
 MUX2_X1 _17267_ (.A(_10719_),
    .B(_00139_),
    .S(_10858_),
    .Z(_11431_));
 OAI21_X1 _17268_ (.A(_11121_),
    .B1(_11430_),
    .B2(_11431_),
    .ZN(_11432_));
 OAI221_X2 _17269_ (.A(_10774_),
    .B1(_11121_),
    .B2(_11427_),
    .C1(_11429_),
    .C2(_11432_),
    .ZN(_11433_));
 BUF_X4 _17270_ (.A(_11433_),
    .Z(_11434_));
 INV_X1 _17271_ (.A(_11434_),
    .ZN(_11435_));
 BUF_X4 _17272_ (.A(_11435_),
    .Z(_16262_));
 BUF_X4 _17273_ (.A(_11434_),
    .Z(_16266_));
 BUF_X4 _17274_ (.A(_10728_),
    .Z(_11436_));
 MUX2_X1 _17275_ (.A(_00324_),
    .B(_00328_),
    .S(_11436_),
    .Z(_11437_));
 MUX2_X1 _17276_ (.A(_00326_),
    .B(_00330_),
    .S(_11436_),
    .Z(_11438_));
 BUF_X4 _17277_ (.A(_11357_),
    .Z(_11439_));
 MUX2_X1 _17278_ (.A(_11437_),
    .B(_11438_),
    .S(_11439_),
    .Z(_11440_));
 MUX2_X1 _17279_ (.A(_00323_),
    .B(_00327_),
    .S(_11436_),
    .Z(_11441_));
 MUX2_X1 _17280_ (.A(_00325_),
    .B(_00329_),
    .S(_11436_),
    .Z(_11442_));
 MUX2_X1 _17281_ (.A(_11441_),
    .B(_11442_),
    .S(_11439_),
    .Z(_11443_));
 MUX2_X1 _17282_ (.A(_11440_),
    .B(_11443_),
    .S(_11130_),
    .Z(_11444_));
 MUX2_X1 _17283_ (.A(_00335_),
    .B(_00337_),
    .S(_11399_),
    .Z(_11445_));
 MUX2_X1 _17284_ (.A(_00336_),
    .B(_00338_),
    .S(_11399_),
    .Z(_11446_));
 MUX2_X1 _17285_ (.A(_11445_),
    .B(_11446_),
    .S(_10710_),
    .Z(_11447_));
 MUX2_X1 _17286_ (.A(_00331_),
    .B(_00333_),
    .S(_11399_),
    .Z(_11448_));
 MUX2_X1 _17287_ (.A(_00332_),
    .B(_00334_),
    .S(_11399_),
    .Z(_11449_));
 MUX2_X1 _17288_ (.A(_11448_),
    .B(_11449_),
    .S(_10710_),
    .Z(_11450_));
 MUX2_X1 _17289_ (.A(_11447_),
    .B(_11450_),
    .S(_10735_),
    .Z(_11451_));
 MUX2_X2 _17290_ (.A(_11444_),
    .B(_11451_),
    .S(_10747_),
    .Z(_11452_));
 MUX2_X1 _17291_ (.A(_00319_),
    .B(_00321_),
    .S(_11439_),
    .Z(_11453_));
 MUX2_X1 _17292_ (.A(_00320_),
    .B(_00322_),
    .S(_11439_),
    .Z(_11454_));
 MUX2_X1 _17293_ (.A(_11453_),
    .B(_11454_),
    .S(_11316_),
    .Z(_11455_));
 NAND2_X1 _17294_ (.A1(_10747_),
    .A2(_11455_),
    .ZN(_11456_));
 MUX2_X1 _17295_ (.A(_00311_),
    .B(_00313_),
    .S(_11439_),
    .Z(_11457_));
 MUX2_X1 _17296_ (.A(_00312_),
    .B(_00314_),
    .S(_11439_),
    .Z(_11458_));
 MUX2_X1 _17297_ (.A(_11457_),
    .B(_11458_),
    .S(_11316_),
    .Z(_11459_));
 NAND2_X1 _17298_ (.A1(_10719_),
    .A2(_11459_),
    .ZN(_11460_));
 NAND3_X1 _17299_ (.A1(_10731_),
    .A2(_11456_),
    .A3(_11460_),
    .ZN(_11461_));
 NAND2_X1 _17300_ (.A1(net378),
    .A2(_00310_),
    .ZN(_11462_));
 OAI21_X1 _17301_ (.A(_11462_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B2(_10705_),
    .ZN(_11463_));
 OAI221_X2 _17302_ (.A(_10718_),
    .B1(_00309_),
    .B2(_11353_),
    .C1(_11463_),
    .C2(_11130_),
    .ZN(_11464_));
 MUX2_X1 _17303_ (.A(_00315_),
    .B(_00317_),
    .S(_11400_),
    .Z(_11465_));
 MUX2_X1 _17304_ (.A(_00316_),
    .B(_00318_),
    .S(_11400_),
    .Z(_11466_));
 MUX2_X1 _17305_ (.A(_11465_),
    .B(_11466_),
    .S(_11316_),
    .Z(_11467_));
 AOI21_X1 _17306_ (.A(_10730_),
    .B1(_10746_),
    .B2(_11467_),
    .ZN(_11468_));
 AOI21_X2 _17307_ (.A(_11134_),
    .B1(_11464_),
    .B2(_11468_),
    .ZN(_11469_));
 AOI22_X4 _17308_ (.A1(_11452_),
    .A2(_11134_),
    .B1(_11461_),
    .B2(_11469_),
    .ZN(_11470_));
 INV_X1 _17309_ (.A(_11310_),
    .ZN(_11471_));
 NOR3_X1 _17310_ (.A1(_11471_),
    .A2(_10859_),
    .A3(_10866_),
    .ZN(_11472_));
 MUX2_X1 _17311_ (.A(_10764_),
    .B(_00138_),
    .S(_10859_),
    .Z(_11473_));
 OAI21_X1 _17312_ (.A(_11121_),
    .B1(_11430_),
    .B2(_11473_),
    .ZN(_11474_));
 OAI221_X2 _17313_ (.A(_10774_),
    .B1(_11121_),
    .B2(_11470_),
    .C1(_11472_),
    .C2(_11474_),
    .ZN(_11475_));
 BUF_X4 _17314_ (.A(_11475_),
    .Z(_11476_));
 INV_X4 _17315_ (.A(_11476_),
    .ZN(_11477_));
 BUF_X4 _17316_ (.A(_11477_),
    .Z(_16270_));
 BUF_X4 _17317_ (.A(_11476_),
    .Z(_11478_));
 BUF_X4 _17318_ (.A(_11478_),
    .Z(_16274_));
 NAND3_X4 _17319_ (.A1(_11281_),
    .A2(_11294_),
    .A3(_11326_),
    .ZN(_11479_));
 OAI21_X1 _17320_ (.A(_10838_),
    .B1(_11121_),
    .B2(_11470_),
    .ZN(_11480_));
 AOI21_X4 _17321_ (.A(_10814_),
    .B1(_10855_),
    .B2(_10773_),
    .ZN(_11481_));
 INV_X1 _17322_ (.A(_00138_),
    .ZN(_11482_));
 MUX2_X1 _17323_ (.A(_11134_),
    .B(_11482_),
    .S(_10859_),
    .Z(_11483_));
 AOI21_X1 _17324_ (.A(_10804_),
    .B1(_11481_),
    .B2(_11483_),
    .ZN(_11484_));
 OAI22_X4 _17325_ (.A1(_10830_),
    .A2(_10831_),
    .B1(_10959_),
    .B2(_10823_),
    .ZN(_11485_));
 AOI21_X4 _17326_ (.A(_10817_),
    .B1(_10834_),
    .B2(_11485_),
    .ZN(_11486_));
 XNOR2_X2 _17327_ (.A(_10814_),
    .B(_10836_),
    .ZN(_11487_));
 NAND3_X1 _17328_ (.A1(_11310_),
    .A2(_11486_),
    .A3(_11487_),
    .ZN(_11488_));
 AOI211_X2 _17329_ (.A(_11479_),
    .B(_11480_),
    .C1(_11484_),
    .C2(_11488_),
    .ZN(_15909_));
 CLKBUF_X3 _17330_ (.A(_15920_),
    .Z(_11489_));
 BUF_X4 _17331_ (.A(_11489_),
    .Z(_11490_));
 OAI21_X4 _17332_ (.A(_11328_),
    .B1(_16253_),
    .B2(_16262_),
    .ZN(_11491_));
 BUF_X4 _17333_ (.A(_11491_),
    .Z(_11492_));
 NAND2_X4 _17334_ (.A1(_11490_),
    .A2(_11492_),
    .ZN(_11493_));
 INV_X2 _17335_ (.A(_11493_),
    .ZN(_15908_));
 MUX2_X1 _17336_ (.A(_00354_),
    .B(_00358_),
    .S(_10729_),
    .Z(_11494_));
 MUX2_X1 _17337_ (.A(_00356_),
    .B(_00360_),
    .S(_10729_),
    .Z(_11495_));
 MUX2_X1 _17338_ (.A(_11494_),
    .B(_11495_),
    .S(_10737_),
    .Z(_11496_));
 MUX2_X1 _17339_ (.A(_00353_),
    .B(_00357_),
    .S(_10730_),
    .Z(_11497_));
 MUX2_X1 _17340_ (.A(_00355_),
    .B(_00359_),
    .S(_10730_),
    .Z(_11498_));
 MUX2_X1 _17341_ (.A(_11497_),
    .B(_11498_),
    .S(_10737_),
    .Z(_11499_));
 MUX2_X1 _17342_ (.A(_11496_),
    .B(_11499_),
    .S(_11130_),
    .Z(_11500_));
 BUF_X4 _17343_ (.A(_10702_),
    .Z(_11501_));
 BUF_X4 _17344_ (.A(_11501_),
    .Z(_11502_));
 MUX2_X1 _17345_ (.A(_00365_),
    .B(_00367_),
    .S(_11502_),
    .Z(_11503_));
 MUX2_X1 _17346_ (.A(_00366_),
    .B(_00368_),
    .S(_11502_),
    .Z(_11504_));
 MUX2_X1 _17347_ (.A(_11503_),
    .B(_11504_),
    .S(_11316_),
    .Z(_11505_));
 MUX2_X1 _17348_ (.A(_00361_),
    .B(_00363_),
    .S(_11502_),
    .Z(_11506_));
 MUX2_X1 _17349_ (.A(_00362_),
    .B(_00364_),
    .S(_11502_),
    .Z(_11507_));
 MUX2_X1 _17350_ (.A(_11506_),
    .B(_11507_),
    .S(_10711_),
    .Z(_11508_));
 MUX2_X2 _17351_ (.A(_11505_),
    .B(_11508_),
    .S(_10736_),
    .Z(_11509_));
 OAI22_X4 _17352_ (.A1(_11424_),
    .A2(_11500_),
    .B1(_11509_),
    .B2(_11408_),
    .ZN(_11510_));
 MUX2_X1 _17353_ (.A(_00341_),
    .B(_00343_),
    .S(_11502_),
    .Z(_11511_));
 INV_X1 _17354_ (.A(_11511_),
    .ZN(_11512_));
 MUX2_X1 _17355_ (.A(_00342_),
    .B(_00344_),
    .S(_11502_),
    .Z(_11513_));
 INV_X1 _17356_ (.A(_11513_),
    .ZN(_11514_));
 OAI22_X2 _17357_ (.A1(_11380_),
    .A2(_11512_),
    .B1(_11514_),
    .B2(_11383_),
    .ZN(_11515_));
 NOR2_X1 _17358_ (.A1(net378),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .ZN(_11516_));
 AOI21_X1 _17359_ (.A(_11516_),
    .B1(_00340_),
    .B2(_10705_),
    .ZN(_11517_));
 NAND2_X1 _17360_ (.A1(_11390_),
    .A2(_11517_),
    .ZN(_11518_));
 INV_X1 _17361_ (.A(_00339_),
    .ZN(_11519_));
 AOI21_X1 _17362_ (.A(_11389_),
    .B1(_11393_),
    .B2(_11519_),
    .ZN(_11520_));
 MUX2_X1 _17363_ (.A(_00346_),
    .B(_00350_),
    .S(_10729_),
    .Z(_11521_));
 MUX2_X1 _17364_ (.A(_00348_),
    .B(_00352_),
    .S(_10729_),
    .Z(_11522_));
 MUX2_X1 _17365_ (.A(_11521_),
    .B(_11522_),
    .S(net378),
    .Z(_11523_));
 MUX2_X1 _17366_ (.A(_00345_),
    .B(_00349_),
    .S(_10729_),
    .Z(_11524_));
 MUX2_X1 _17367_ (.A(_00347_),
    .B(_00351_),
    .S(_10729_),
    .Z(_11525_));
 MUX2_X1 _17368_ (.A(_11524_),
    .B(_11525_),
    .S(net378),
    .Z(_11526_));
 MUX2_X1 _17369_ (.A(_11523_),
    .B(_11526_),
    .S(_11130_),
    .Z(_11527_));
 AOI221_X2 _17370_ (.A(_11515_),
    .B1(_11518_),
    .B2(_11520_),
    .C1(_11527_),
    .C2(_10747_),
    .ZN(_11528_));
 OAI21_X1 _17371_ (.A(_11167_),
    .B1(_11510_),
    .B2(_11528_),
    .ZN(_11529_));
 AOI211_X2 _17372_ (.A(_10817_),
    .B(_10814_),
    .C1(_10834_),
    .C2(_11485_),
    .ZN(_11530_));
 AOI211_X2 _17373_ (.A(_10817_),
    .B(_10822_),
    .C1(_10832_),
    .C2(_10834_),
    .ZN(_11531_));
 OAI21_X2 _17374_ (.A(_10805_),
    .B1(_11530_),
    .B2(_11531_),
    .ZN(_11532_));
 OAI21_X2 _17375_ (.A(_11529_),
    .B1(_11532_),
    .B2(_10949_),
    .ZN(_11533_));
 INV_X2 _17376_ (.A(_11533_),
    .ZN(_11534_));
 BUF_X4 _17377_ (.A(_11534_),
    .Z(_16282_));
 NAND2_X1 _17378_ (.A1(_10869_),
    .A2(_11120_),
    .ZN(_11535_));
 AOI211_X2 _17379_ (.A(_10858_),
    .B(_11535_),
    .C1(_10814_),
    .C2(_10855_),
    .ZN(_11536_));
 NOR3_X2 _17380_ (.A1(_00177_),
    .A2(_10804_),
    .A3(_11486_),
    .ZN(_11537_));
 MUX2_X1 _17381_ (.A(_00384_),
    .B(_00388_),
    .S(_10728_),
    .Z(_11538_));
 MUX2_X1 _17382_ (.A(_00386_),
    .B(_00390_),
    .S(_10728_),
    .Z(_11539_));
 MUX2_X1 _17383_ (.A(_11538_),
    .B(_11539_),
    .S(_11501_),
    .Z(_11540_));
 MUX2_X1 _17384_ (.A(_00383_),
    .B(_00387_),
    .S(_10728_),
    .Z(_11541_));
 MUX2_X1 _17385_ (.A(_00385_),
    .B(_00389_),
    .S(_10728_),
    .Z(_11542_));
 MUX2_X1 _17386_ (.A(_11541_),
    .B(_11542_),
    .S(_11501_),
    .Z(_11543_));
 MUX2_X1 _17387_ (.A(_11540_),
    .B(_11543_),
    .S(_11129_),
    .Z(_11544_));
 MUX2_X1 _17388_ (.A(_00395_),
    .B(_00397_),
    .S(_11354_),
    .Z(_11545_));
 MUX2_X1 _17389_ (.A(_00396_),
    .B(_00398_),
    .S(_11354_),
    .Z(_11546_));
 MUX2_X1 _17390_ (.A(_11545_),
    .B(_11546_),
    .S(_10709_),
    .Z(_11547_));
 MUX2_X1 _17391_ (.A(_00391_),
    .B(_00393_),
    .S(_11354_),
    .Z(_11548_));
 MUX2_X1 _17392_ (.A(_00392_),
    .B(_00394_),
    .S(_11354_),
    .Z(_11549_));
 MUX2_X1 _17393_ (.A(_11548_),
    .B(_11549_),
    .S(_10709_),
    .Z(_11550_));
 MUX2_X1 _17394_ (.A(_11547_),
    .B(_11550_),
    .S(_10735_),
    .Z(_11551_));
 MUX2_X1 _17395_ (.A(_11544_),
    .B(_11551_),
    .S(_10746_),
    .Z(_11552_));
 MUX2_X1 _17396_ (.A(_00379_),
    .B(_00381_),
    .S(_11501_),
    .Z(_11553_));
 MUX2_X1 _17397_ (.A(_00380_),
    .B(_00382_),
    .S(_11501_),
    .Z(_11554_));
 MUX2_X1 _17398_ (.A(_11553_),
    .B(_11554_),
    .S(_10710_),
    .Z(_11555_));
 NAND2_X1 _17399_ (.A1(_10746_),
    .A2(_11555_),
    .ZN(_11556_));
 MUX2_X1 _17400_ (.A(_00371_),
    .B(_00373_),
    .S(_11501_),
    .Z(_11557_));
 MUX2_X1 _17401_ (.A(_00372_),
    .B(_00374_),
    .S(_11501_),
    .Z(_11558_));
 MUX2_X1 _17402_ (.A(_11557_),
    .B(_11558_),
    .S(_10710_),
    .Z(_11559_));
 NAND2_X1 _17403_ (.A1(_10718_),
    .A2(_11559_),
    .ZN(_11560_));
 NAND3_X1 _17404_ (.A1(_10731_),
    .A2(_11556_),
    .A3(_11560_),
    .ZN(_11561_));
 NAND2_X1 _17405_ (.A1(_11502_),
    .A2(_00370_),
    .ZN(_11562_));
 OAI21_X1 _17406_ (.A(_11562_),
    .B1(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .B2(_10704_),
    .ZN(_11563_));
 OAI221_X2 _17407_ (.A(_10718_),
    .B1(_00369_),
    .B2(_11353_),
    .C1(_11563_),
    .C2(_11130_),
    .ZN(_11564_));
 MUX2_X1 _17408_ (.A(_00375_),
    .B(_00377_),
    .S(_11399_),
    .Z(_11565_));
 MUX2_X1 _17409_ (.A(_00376_),
    .B(_00378_),
    .S(_11399_),
    .Z(_11566_));
 MUX2_X1 _17410_ (.A(_11565_),
    .B(_11566_),
    .S(_10710_),
    .Z(_11567_));
 AOI21_X2 _17411_ (.A(_10730_),
    .B1(_10746_),
    .B2(_11567_),
    .ZN(_11568_));
 AOI21_X4 _17412_ (.A(_11134_),
    .B1(_11564_),
    .B2(_11568_),
    .ZN(_11569_));
 AOI22_X4 _17413_ (.A1(_11552_),
    .A2(_11134_),
    .B1(_11561_),
    .B2(_11569_),
    .ZN(_11570_));
 AOI221_X2 _17414_ (.A(_11536_),
    .B1(_11537_),
    .B2(_11481_),
    .C1(_11570_),
    .C2(_10804_),
    .ZN(_11571_));
 NOR2_X4 _17415_ (.A1(_10819_),
    .A2(net10),
    .ZN(_16286_));
 INV_X1 _17416_ (.A(_16286_),
    .ZN(_16290_));
 AND3_X1 _17417_ (.A1(_10873_),
    .A2(_10773_),
    .A3(_11120_),
    .ZN(_11572_));
 OAI21_X1 _17418_ (.A(_11572_),
    .B1(_11530_),
    .B2(_10836_),
    .ZN(_11573_));
 MUX2_X1 _17419_ (.A(_00414_),
    .B(_00418_),
    .S(_11436_),
    .Z(_11574_));
 MUX2_X1 _17420_ (.A(_00416_),
    .B(_00420_),
    .S(_11436_),
    .Z(_11575_));
 MUX2_X1 _17421_ (.A(_11574_),
    .B(_11575_),
    .S(_11439_),
    .Z(_11576_));
 MUX2_X1 _17422_ (.A(_00413_),
    .B(_00417_),
    .S(_11436_),
    .Z(_11577_));
 MUX2_X1 _17423_ (.A(_00415_),
    .B(_00419_),
    .S(_11436_),
    .Z(_11578_));
 MUX2_X1 _17424_ (.A(_11577_),
    .B(_11578_),
    .S(_11439_),
    .Z(_11579_));
 MUX2_X1 _17425_ (.A(_11576_),
    .B(_11579_),
    .S(_11130_),
    .Z(_11580_));
 MUX2_X1 _17426_ (.A(_00406_),
    .B(_00410_),
    .S(_10733_),
    .Z(_11581_));
 MUX2_X1 _17427_ (.A(_00408_),
    .B(_00412_),
    .S(_10733_),
    .Z(_11582_));
 MUX2_X1 _17428_ (.A(_11581_),
    .B(_11582_),
    .S(_11439_),
    .Z(_11583_));
 MUX2_X1 _17429_ (.A(_00405_),
    .B(_00409_),
    .S(_11436_),
    .Z(_11584_));
 MUX2_X1 _17430_ (.A(_00407_),
    .B(_00411_),
    .S(_11436_),
    .Z(_11585_));
 MUX2_X1 _17431_ (.A(_11584_),
    .B(_11585_),
    .S(_11439_),
    .Z(_11586_));
 MUX2_X1 _17432_ (.A(_11583_),
    .B(_11586_),
    .S(_11405_),
    .Z(_11587_));
 BUF_X4 _17433_ (.A(_11357_),
    .Z(_11588_));
 MUX2_X1 _17434_ (.A(_00401_),
    .B(_00403_),
    .S(_11588_),
    .Z(_11589_));
 INV_X1 _17435_ (.A(_11589_),
    .ZN(_11590_));
 MUX2_X1 _17436_ (.A(_00402_),
    .B(_00404_),
    .S(_11400_),
    .Z(_11591_));
 INV_X1 _17437_ (.A(_11591_),
    .ZN(_11592_));
 OAI22_X2 _17438_ (.A1(_11380_),
    .A2(_11590_),
    .B1(_11592_),
    .B2(_11383_),
    .ZN(_11593_));
 NOR2_X1 _17439_ (.A1(_11357_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .ZN(_11594_));
 AOI21_X1 _17440_ (.A(_11594_),
    .B1(_00400_),
    .B2(net377),
    .ZN(_11595_));
 INV_X1 _17441_ (.A(_00399_),
    .ZN(_11596_));
 AOI221_X2 _17442_ (.A(_11389_),
    .B1(_11390_),
    .B2(_11595_),
    .C1(_11393_),
    .C2(_11596_),
    .ZN(_11597_));
 OAI33_X1 _17443_ (.A1(_10747_),
    .A2(_10763_),
    .A3(_11580_),
    .B1(_11587_),
    .B2(_11593_),
    .B3(_11597_),
    .ZN(_11598_));
 MUX2_X1 _17444_ (.A(_00425_),
    .B(_00427_),
    .S(_11588_),
    .Z(_11599_));
 NOR2_X1 _17445_ (.A1(_11316_),
    .A2(_11599_),
    .ZN(_11600_));
 MUX2_X1 _17446_ (.A(_00426_),
    .B(_00428_),
    .S(_11400_),
    .Z(_11601_));
 NOR2_X1 _17447_ (.A1(_11130_),
    .A2(_11601_),
    .ZN(_11602_));
 NOR3_X1 _17448_ (.A1(_10735_),
    .A2(_11600_),
    .A3(_11602_),
    .ZN(_11603_));
 MUX2_X1 _17449_ (.A(_00421_),
    .B(_00423_),
    .S(_10703_),
    .Z(_11604_));
 NOR2_X1 _17450_ (.A1(_11316_),
    .A2(_11604_),
    .ZN(_11605_));
 MUX2_X1 _17451_ (.A(_00422_),
    .B(_00424_),
    .S(_10703_),
    .Z(_11606_));
 NOR2_X1 _17452_ (.A1(_11405_),
    .A2(_11606_),
    .ZN(_11607_));
 NOR3_X1 _17453_ (.A1(_10730_),
    .A2(_11605_),
    .A3(_11607_),
    .ZN(_11608_));
 OAI33_X1 _17454_ (.A1(_10747_),
    .A2(_11593_),
    .A3(_11597_),
    .B1(_11603_),
    .B2(_11608_),
    .B3(_11408_),
    .ZN(_11609_));
 OAI21_X1 _17455_ (.A(_11167_),
    .B1(_11598_),
    .B2(_11609_),
    .ZN(_11610_));
 AND2_X1 _17456_ (.A1(_11573_),
    .A2(_11610_),
    .ZN(_11611_));
 BUF_X4 _17457_ (.A(_11611_),
    .Z(_16298_));
 MUX2_X1 _17458_ (.A(_00431_),
    .B(_00433_),
    .S(_10703_),
    .Z(_11612_));
 INV_X1 _17459_ (.A(_11612_),
    .ZN(_11613_));
 BUF_X4 _17460_ (.A(_10702_),
    .Z(_11614_));
 MUX2_X1 _17461_ (.A(_00432_),
    .B(_00434_),
    .S(_11614_),
    .Z(_11615_));
 INV_X1 _17462_ (.A(_11615_),
    .ZN(_11616_));
 OAI22_X4 _17463_ (.A1(_11380_),
    .A2(_11613_),
    .B1(_11616_),
    .B2(_11383_),
    .ZN(_11617_));
 NOR2_X1 _17464_ (.A1(_11352_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .ZN(_11618_));
 AOI21_X1 _17465_ (.A(_11618_),
    .B1(_00430_),
    .B2(_11357_),
    .ZN(_11619_));
 INV_X1 _17466_ (.A(_00429_),
    .ZN(_11620_));
 AOI221_X2 _17467_ (.A(_11389_),
    .B1(_11390_),
    .B2(_11619_),
    .C1(_11393_),
    .C2(_11620_),
    .ZN(_11621_));
 CLKBUF_X3 _17468_ (.A(_10728_),
    .Z(_11622_));
 MUX2_X1 _17469_ (.A(_00436_),
    .B(_00440_),
    .S(_11622_),
    .Z(_11623_));
 MUX2_X1 _17470_ (.A(_00438_),
    .B(_00442_),
    .S(_11622_),
    .Z(_11624_));
 MUX2_X1 _17471_ (.A(_11623_),
    .B(_11624_),
    .S(_11588_),
    .Z(_11625_));
 MUX2_X1 _17472_ (.A(_00435_),
    .B(_00439_),
    .S(_10733_),
    .Z(_11626_));
 MUX2_X1 _17473_ (.A(_00437_),
    .B(_00441_),
    .S(_10733_),
    .Z(_11627_));
 MUX2_X1 _17474_ (.A(_11626_),
    .B(_11627_),
    .S(_11588_),
    .Z(_11628_));
 MUX2_X1 _17475_ (.A(_11625_),
    .B(_11628_),
    .S(_11405_),
    .Z(_11629_));
 NOR3_X4 _17476_ (.A1(_11617_),
    .A2(_11621_),
    .A3(_11629_),
    .ZN(_11630_));
 MUX2_X1 _17477_ (.A(_00455_),
    .B(_00457_),
    .S(_11355_),
    .Z(_11631_));
 MUX2_X1 _17478_ (.A(_00456_),
    .B(_00458_),
    .S(_11355_),
    .Z(_11632_));
 MUX2_X1 _17479_ (.A(_11631_),
    .B(_11632_),
    .S(_11315_),
    .Z(_11633_));
 MUX2_X1 _17480_ (.A(_00451_),
    .B(_00453_),
    .S(_11355_),
    .Z(_11634_));
 MUX2_X1 _17481_ (.A(_00452_),
    .B(_00454_),
    .S(_11355_),
    .Z(_11635_));
 MUX2_X1 _17482_ (.A(_11634_),
    .B(_11635_),
    .S(_11315_),
    .Z(_11636_));
 MUX2_X1 _17483_ (.A(_11633_),
    .B(_11636_),
    .S(_10735_),
    .Z(_11637_));
 NOR2_X2 _17484_ (.A1(_11408_),
    .A2(_11637_),
    .ZN(_11638_));
 MUX2_X1 _17485_ (.A(_00444_),
    .B(_00448_),
    .S(_11622_),
    .Z(_11639_));
 MUX2_X1 _17486_ (.A(_00446_),
    .B(_00450_),
    .S(_11622_),
    .Z(_11640_));
 MUX2_X1 _17487_ (.A(_11639_),
    .B(_11640_),
    .S(_11588_),
    .Z(_11641_));
 MUX2_X1 _17488_ (.A(_00443_),
    .B(_00447_),
    .S(_11622_),
    .Z(_11642_));
 MUX2_X1 _17489_ (.A(_00445_),
    .B(_00449_),
    .S(_11622_),
    .Z(_11643_));
 MUX2_X1 _17490_ (.A(_11642_),
    .B(_11643_),
    .S(_11588_),
    .Z(_11644_));
 MUX2_X1 _17491_ (.A(_11641_),
    .B(_11644_),
    .S(_11405_),
    .Z(_11645_));
 NOR2_X2 _17492_ (.A1(_11424_),
    .A2(_11645_),
    .ZN(_11646_));
 NOR3_X4 _17493_ (.A1(_10746_),
    .A2(_11617_),
    .A3(_11621_),
    .ZN(_11647_));
 OR4_X4 _17494_ (.A1(_11630_),
    .A2(_11638_),
    .A3(_11646_),
    .A4(_11647_),
    .ZN(_11648_));
 INV_X1 _17495_ (.A(_10876_),
    .ZN(_11649_));
 NOR2_X2 _17496_ (.A1(_11530_),
    .A2(_11531_),
    .ZN(_11650_));
 NOR2_X1 _17497_ (.A1(_11649_),
    .A2(_11650_),
    .ZN(_11651_));
 MUX2_X2 _17498_ (.A(_11648_),
    .B(_11651_),
    .S(_10805_),
    .Z(_16301_));
 INV_X1 _17499_ (.A(_16301_),
    .ZN(_16305_));
 MUX2_X1 _17500_ (.A(_00485_),
    .B(_00487_),
    .S(_10702_),
    .Z(_11652_));
 MUX2_X1 _17501_ (.A(_00486_),
    .B(_00488_),
    .S(net380),
    .Z(_11653_));
 MUX2_X1 _17502_ (.A(_11652_),
    .B(_11653_),
    .S(_10709_),
    .Z(_11654_));
 MUX2_X1 _17503_ (.A(_00481_),
    .B(_00483_),
    .S(_10702_),
    .Z(_11655_));
 MUX2_X1 _17504_ (.A(_00482_),
    .B(_00484_),
    .S(_10702_),
    .Z(_11656_));
 MUX2_X1 _17505_ (.A(_11655_),
    .B(_11656_),
    .S(_11315_),
    .Z(_11657_));
 MUX2_X1 _17506_ (.A(_11654_),
    .B(_11657_),
    .S(_10735_),
    .Z(_11658_));
 NOR2_X2 _17507_ (.A1(_11408_),
    .A2(_11658_),
    .ZN(_11659_));
 MUX2_X1 _17508_ (.A(_00466_),
    .B(_00470_),
    .S(_11622_),
    .Z(_11660_));
 MUX2_X1 _17509_ (.A(_00468_),
    .B(_00472_),
    .S(_11622_),
    .Z(_11661_));
 MUX2_X1 _17510_ (.A(_11660_),
    .B(_11661_),
    .S(_11588_),
    .Z(_11662_));
 MUX2_X1 _17511_ (.A(_00465_),
    .B(_00469_),
    .S(_11622_),
    .Z(_11663_));
 MUX2_X1 _17512_ (.A(_00467_),
    .B(_00471_),
    .S(_11622_),
    .Z(_11664_));
 MUX2_X1 _17513_ (.A(_11663_),
    .B(_11664_),
    .S(_11588_),
    .Z(_11665_));
 MUX2_X1 _17514_ (.A(_11662_),
    .B(_11665_),
    .S(_11405_),
    .Z(_11666_));
 INV_X1 _17515_ (.A(_11666_),
    .ZN(_11667_));
 MUX2_X1 _17516_ (.A(_00461_),
    .B(_00463_),
    .S(_10703_),
    .Z(_11668_));
 INV_X1 _17517_ (.A(_11668_),
    .ZN(_11669_));
 MUX2_X1 _17518_ (.A(_00462_),
    .B(_00464_),
    .S(_11614_),
    .Z(_11670_));
 INV_X1 _17519_ (.A(_11670_),
    .ZN(_11671_));
 OAI22_X2 _17520_ (.A1(_11380_),
    .A2(_11669_),
    .B1(_11671_),
    .B2(_11383_),
    .ZN(_11672_));
 NOR2_X1 _17521_ (.A1(_11352_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .ZN(_11673_));
 AOI21_X1 _17522_ (.A(_11673_),
    .B1(_00460_),
    .B2(_11357_),
    .ZN(_11674_));
 INV_X1 _17523_ (.A(_00459_),
    .ZN(_11675_));
 AOI221_X2 _17524_ (.A(_11389_),
    .B1(_11390_),
    .B2(_11674_),
    .C1(_11393_),
    .C2(_11675_),
    .ZN(_11676_));
 NOR2_X1 _17525_ (.A1(_11672_),
    .A2(_11676_),
    .ZN(_11677_));
 MUX2_X1 _17526_ (.A(_00474_),
    .B(_00478_),
    .S(_10728_),
    .Z(_11678_));
 MUX2_X1 _17527_ (.A(_00476_),
    .B(_00480_),
    .S(_10728_),
    .Z(_11679_));
 MUX2_X1 _17528_ (.A(_11678_),
    .B(_11679_),
    .S(net377),
    .Z(_11680_));
 MUX2_X1 _17529_ (.A(_00473_),
    .B(_00477_),
    .S(_11396_),
    .Z(_11681_));
 MUX2_X1 _17530_ (.A(_00475_),
    .B(_00479_),
    .S(_11396_),
    .Z(_11682_));
 MUX2_X1 _17531_ (.A(_11681_),
    .B(_11682_),
    .S(_11400_),
    .Z(_11683_));
 MUX2_X1 _17532_ (.A(_11680_),
    .B(_11683_),
    .S(_11405_),
    .Z(_11684_));
 OAI22_X2 _17533_ (.A1(_11672_),
    .A2(_11676_),
    .B1(_11684_),
    .B2(_10763_),
    .ZN(_11685_));
 AOI221_X2 _17534_ (.A(_11659_),
    .B1(_11667_),
    .B2(_11677_),
    .C1(_11685_),
    .C2(_10719_),
    .ZN(_11686_));
 OAI22_X4 _17535_ (.A1(_11314_),
    .A2(_11532_),
    .B1(_11686_),
    .B2(_10805_),
    .ZN(_16309_));
 INV_X2 _17536_ (.A(_16309_),
    .ZN(_16313_));
 OAI211_X2 _17537_ (.A(_10838_),
    .B(_10845_),
    .C1(_10853_),
    .C2(_10854_),
    .ZN(_11687_));
 AOI21_X2 _17538_ (.A(_11168_),
    .B1(_11118_),
    .B2(_11687_),
    .ZN(_11688_));
 MUX2_X1 _17539_ (.A(_00491_),
    .B(_00493_),
    .S(net380),
    .Z(_11689_));
 INV_X1 _17540_ (.A(_11689_),
    .ZN(_11690_));
 MUX2_X1 _17541_ (.A(_00492_),
    .B(_00494_),
    .S(_11354_),
    .Z(_11691_));
 INV_X1 _17542_ (.A(_11691_),
    .ZN(_11692_));
 OAI22_X4 _17543_ (.A1(_11380_),
    .A2(_11690_),
    .B1(_11692_),
    .B2(_11383_),
    .ZN(_11693_));
 NOR2_X1 _17544_ (.A1(net342),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .ZN(_11694_));
 AOI21_X2 _17545_ (.A(_11694_),
    .B1(_00490_),
    .B2(_11354_),
    .ZN(_11695_));
 INV_X1 _17546_ (.A(_00489_),
    .ZN(_11696_));
 AOI221_X2 _17547_ (.A(_11389_),
    .B1(_11390_),
    .B2(_11695_),
    .C1(_11393_),
    .C2(_11696_),
    .ZN(_11697_));
 MUX2_X1 _17548_ (.A(_00496_),
    .B(_00500_),
    .S(_11387_),
    .Z(_11698_));
 MUX2_X1 _17549_ (.A(_00498_),
    .B(_00502_),
    .S(_11387_),
    .Z(_11699_));
 MUX2_X1 _17550_ (.A(_11698_),
    .B(_11699_),
    .S(_11399_),
    .Z(_11700_));
 MUX2_X1 _17551_ (.A(_00495_),
    .B(_00499_),
    .S(_11387_),
    .Z(_11701_));
 MUX2_X1 _17552_ (.A(_00497_),
    .B(_00501_),
    .S(_11387_),
    .Z(_11702_));
 MUX2_X1 _17553_ (.A(_11701_),
    .B(_11702_),
    .S(_11399_),
    .Z(_11703_));
 MUX2_X1 _17554_ (.A(_11700_),
    .B(_11703_),
    .S(_11129_),
    .Z(_11704_));
 NOR3_X2 _17555_ (.A1(_11693_),
    .A2(_11697_),
    .A3(_11704_),
    .ZN(_11705_));
 MUX2_X1 _17556_ (.A(_00515_),
    .B(_00517_),
    .S(net342),
    .Z(_11706_));
 MUX2_X1 _17557_ (.A(_00516_),
    .B(_00518_),
    .S(net342),
    .Z(_11707_));
 MUX2_X1 _17558_ (.A(_11706_),
    .B(_11707_),
    .S(_10709_),
    .Z(_11708_));
 MUX2_X1 _17559_ (.A(_00511_),
    .B(_00513_),
    .S(net342),
    .Z(_11709_));
 MUX2_X1 _17560_ (.A(_00512_),
    .B(_00514_),
    .S(_11354_),
    .Z(_11710_));
 MUX2_X1 _17561_ (.A(_11709_),
    .B(_11710_),
    .S(_10709_),
    .Z(_11711_));
 MUX2_X1 _17562_ (.A(_11708_),
    .B(_11711_),
    .S(_10735_),
    .Z(_11712_));
 NOR2_X2 _17563_ (.A1(_11408_),
    .A2(_11712_),
    .ZN(_11713_));
 MUX2_X1 _17564_ (.A(_00504_),
    .B(_00508_),
    .S(_11387_),
    .Z(_11714_));
 MUX2_X1 _17565_ (.A(_00506_),
    .B(_00510_),
    .S(_11387_),
    .Z(_11715_));
 MUX2_X1 _17566_ (.A(_11714_),
    .B(_11715_),
    .S(_11355_),
    .Z(_11716_));
 MUX2_X1 _17567_ (.A(_00503_),
    .B(_00507_),
    .S(_11387_),
    .Z(_11717_));
 MUX2_X1 _17568_ (.A(_00505_),
    .B(_00509_),
    .S(_11387_),
    .Z(_11718_));
 MUX2_X1 _17569_ (.A(_11717_),
    .B(_11718_),
    .S(_11399_),
    .Z(_11719_));
 MUX2_X1 _17570_ (.A(_11716_),
    .B(_11719_),
    .S(_11129_),
    .Z(_11720_));
 NOR2_X2 _17571_ (.A1(_11424_),
    .A2(_11720_),
    .ZN(_11721_));
 NOR3_X2 _17572_ (.A1(_10746_),
    .A2(_11693_),
    .A3(_11697_),
    .ZN(_11722_));
 OR4_X2 _17573_ (.A1(_11705_),
    .A2(_11713_),
    .A3(_11721_),
    .A4(_11722_),
    .ZN(_11723_));
 BUF_X4 _17574_ (.A(_11723_),
    .Z(_11724_));
 AOI22_X4 _17575_ (.A1(_10884_),
    .A2(_11688_),
    .B1(_11724_),
    .B2(_11168_),
    .ZN(_16322_));
 NOR2_X1 _17576_ (.A1(_10818_),
    .A2(_10864_),
    .ZN(_11725_));
 AOI22_X2 _17577_ (.A1(_10774_),
    .A2(_10855_),
    .B1(_11725_),
    .B2(_11306_),
    .ZN(_11726_));
 INV_X1 _17578_ (.A(_10878_),
    .ZN(_11727_));
 MUX2_X1 _17579_ (.A(_11727_),
    .B(_00140_),
    .S(_10859_),
    .Z(_11728_));
 OAI21_X2 _17580_ (.A(_11726_),
    .B1(_11728_),
    .B2(_10814_),
    .ZN(_11729_));
 NOR2_X1 _17581_ (.A1(_10900_),
    .A2(_10814_),
    .ZN(_11730_));
 AOI211_X2 _17582_ (.A(_10818_),
    .B(_10836_),
    .C1(_11486_),
    .C2(_11730_),
    .ZN(_11731_));
 NOR2_X2 _17583_ (.A1(_11122_),
    .A2(_11731_),
    .ZN(_11732_));
 MUX2_X1 _17584_ (.A(_00534_),
    .B(_00538_),
    .S(_10733_),
    .Z(_11733_));
 MUX2_X1 _17585_ (.A(_00536_),
    .B(_00540_),
    .S(_10733_),
    .Z(_11734_));
 MUX2_X1 _17586_ (.A(_11733_),
    .B(_11734_),
    .S(_11588_),
    .Z(_11735_));
 MUX2_X1 _17587_ (.A(_00533_),
    .B(_00537_),
    .S(_10733_),
    .Z(_11736_));
 MUX2_X1 _17588_ (.A(_00535_),
    .B(_00539_),
    .S(_10733_),
    .Z(_11737_));
 MUX2_X1 _17589_ (.A(_11736_),
    .B(_11737_),
    .S(_11588_),
    .Z(_11738_));
 MUX2_X1 _17590_ (.A(_11735_),
    .B(_11738_),
    .S(_11405_),
    .Z(_11739_));
 NOR2_X2 _17591_ (.A1(_10747_),
    .A2(_11739_),
    .ZN(_11740_));
 MUX2_X1 _17592_ (.A(_00545_),
    .B(_00547_),
    .S(_11355_),
    .Z(_11741_));
 MUX2_X1 _17593_ (.A(_00546_),
    .B(_00548_),
    .S(_11355_),
    .Z(_11742_));
 MUX2_X1 _17594_ (.A(_11741_),
    .B(_11742_),
    .S(_11315_),
    .Z(_11743_));
 MUX2_X1 _17595_ (.A(_00541_),
    .B(_00543_),
    .S(_11355_),
    .Z(_11744_));
 MUX2_X1 _17596_ (.A(_00542_),
    .B(_00544_),
    .S(_11355_),
    .Z(_11745_));
 MUX2_X1 _17597_ (.A(_11744_),
    .B(_11745_),
    .S(_11315_),
    .Z(_11746_));
 MUX2_X1 _17598_ (.A(_11743_),
    .B(_11746_),
    .S(_10735_),
    .Z(_11747_));
 NOR2_X2 _17599_ (.A1(_10719_),
    .A2(_11747_),
    .ZN(_11748_));
 NOR3_X4 _17600_ (.A1(_10764_),
    .A2(_11740_),
    .A3(_11748_),
    .ZN(_11749_));
 MUX2_X1 _17601_ (.A(_00525_),
    .B(_00527_),
    .S(net377),
    .Z(_11750_));
 NOR2_X1 _17602_ (.A1(_11316_),
    .A2(_11750_),
    .ZN(_11751_));
 MUX2_X1 _17603_ (.A(_00526_),
    .B(_00528_),
    .S(_11614_),
    .Z(_11752_));
 NOR2_X1 _17604_ (.A1(_11405_),
    .A2(_11752_),
    .ZN(_11753_));
 NOR3_X2 _17605_ (.A1(_10718_),
    .A2(_11751_),
    .A3(_11753_),
    .ZN(_11754_));
 INV_X1 _17606_ (.A(_00519_),
    .ZN(_11755_));
 NOR2_X1 _17607_ (.A1(_11357_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .ZN(_11756_));
 AOI21_X2 _17608_ (.A(_11756_),
    .B1(_00520_),
    .B2(_11400_),
    .ZN(_11757_));
 AOI221_X2 _17609_ (.A(_10717_),
    .B1(_11755_),
    .B2(_11137_),
    .C1(_11757_),
    .C2(_10710_),
    .ZN(_11758_));
 NOR3_X2 _17610_ (.A1(_10730_),
    .A2(_11754_),
    .A3(_11758_),
    .ZN(_11759_));
 MUX2_X1 _17611_ (.A(_00529_),
    .B(_00531_),
    .S(net380),
    .Z(_11760_));
 MUX2_X1 _17612_ (.A(_00530_),
    .B(_00532_),
    .S(_11352_),
    .Z(_11761_));
 MUX2_X1 _17613_ (.A(_11760_),
    .B(_11761_),
    .S(_11315_),
    .Z(_11762_));
 MUX2_X1 _17614_ (.A(_00521_),
    .B(_00523_),
    .S(_11352_),
    .Z(_11763_));
 MUX2_X1 _17615_ (.A(_00522_),
    .B(_00524_),
    .S(_11352_),
    .Z(_11764_));
 MUX2_X1 _17616_ (.A(_11763_),
    .B(_11764_),
    .S(_11315_),
    .Z(_11765_));
 MUX2_X1 _17617_ (.A(_11762_),
    .B(_11765_),
    .S(_10718_),
    .Z(_11766_));
 NOR2_X2 _17618_ (.A1(_10735_),
    .A2(_11766_),
    .ZN(_11767_));
 NOR3_X4 _17619_ (.A1(_11134_),
    .A2(_11759_),
    .A3(_11767_),
    .ZN(_11768_));
 NOR2_X4 _17620_ (.A1(_11749_),
    .A2(_11768_),
    .ZN(_11769_));
 AOI22_X4 _17621_ (.A1(_11729_),
    .A2(_11732_),
    .B1(_11769_),
    .B2(_11167_),
    .ZN(_16330_));
 INV_X1 _17622_ (.A(_16330_),
    .ZN(_11770_));
 BUF_X4 _17623_ (.A(_11770_),
    .Z(_16326_));
 OR2_X1 _17624_ (.A1(_10826_),
    .A2(_11305_),
    .ZN(_11771_));
 NAND3_X2 _17625_ (.A1(_10914_),
    .A2(_10971_),
    .A3(_11771_),
    .ZN(_15924_));
 INV_X1 _17626_ (.A(_15924_),
    .ZN(_15931_));
 NAND3_X2 _17627_ (.A1(_10881_),
    .A2(_10971_),
    .A3(_11305_),
    .ZN(_11772_));
 BUF_X2 _17628_ (.A(_11772_),
    .Z(_15928_));
 NAND2_X1 _17629_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(_10957_),
    .ZN(_11773_));
 MUX2_X1 _17630_ (.A(_00541_),
    .B(_00543_),
    .S(_11096_),
    .Z(_11774_));
 MUX2_X1 _17631_ (.A(_00542_),
    .B(_00544_),
    .S(_11096_),
    .Z(_11775_));
 MUX2_X1 _17632_ (.A(_11774_),
    .B(_11775_),
    .S(_11271_),
    .Z(_11776_));
 MUX2_X1 _17633_ (.A(_00525_),
    .B(_00527_),
    .S(_11096_),
    .Z(_11777_));
 MUX2_X1 _17634_ (.A(_00526_),
    .B(_00528_),
    .S(_11096_),
    .Z(_11778_));
 MUX2_X1 _17635_ (.A(_11777_),
    .B(_11778_),
    .S(_11271_),
    .Z(_11779_));
 BUF_X4 _17636_ (.A(_10979_),
    .Z(_11780_));
 MUX2_X1 _17637_ (.A(_11776_),
    .B(_11779_),
    .S(_11780_),
    .Z(_11781_));
 NOR2_X1 _17638_ (.A1(_10988_),
    .A2(_11781_),
    .ZN(_11782_));
 BUF_X4 _17639_ (.A(_11239_),
    .Z(_11783_));
 MUX2_X1 _17640_ (.A(_00545_),
    .B(_00547_),
    .S(_11783_),
    .Z(_11784_));
 MUX2_X1 _17641_ (.A(_00546_),
    .B(_00548_),
    .S(_11783_),
    .Z(_11785_));
 MUX2_X1 _17642_ (.A(_11784_),
    .B(_11785_),
    .S(_11060_),
    .Z(_11786_));
 MUX2_X1 _17643_ (.A(_00529_),
    .B(_00531_),
    .S(_11783_),
    .Z(_11787_));
 MUX2_X1 _17644_ (.A(_00530_),
    .B(_00532_),
    .S(_11783_),
    .Z(_11788_));
 MUX2_X1 _17645_ (.A(_11787_),
    .B(_11788_),
    .S(_11060_),
    .Z(_11789_));
 MUX2_X1 _17646_ (.A(_11786_),
    .B(_11789_),
    .S(_11780_),
    .Z(_11790_));
 NOR2_X1 _17647_ (.A1(_11038_),
    .A2(_11790_),
    .ZN(_11791_));
 NOR3_X4 _17648_ (.A1(_10995_),
    .A2(_11782_),
    .A3(_11791_),
    .ZN(_11792_));
 MUX2_X1 _17649_ (.A(_00533_),
    .B(_00535_),
    .S(_11241_),
    .Z(_11793_));
 NOR2_X1 _17650_ (.A1(_11028_),
    .A2(_11793_),
    .ZN(_11794_));
 BUF_X4 _17651_ (.A(_11012_),
    .Z(_11795_));
 MUX2_X1 _17652_ (.A(_00534_),
    .B(_00536_),
    .S(_11246_),
    .Z(_11796_));
 NOR2_X1 _17653_ (.A1(_11795_),
    .A2(_11796_),
    .ZN(_11797_));
 NOR3_X1 _17654_ (.A1(_10981_),
    .A2(_11794_),
    .A3(_11797_),
    .ZN(_11798_));
 BUF_X4 _17655_ (.A(_11030_),
    .Z(_11799_));
 BUF_X4 _17656_ (.A(_11064_),
    .Z(_11800_));
 BUF_X4 _17657_ (.A(_11800_),
    .Z(_11801_));
 NOR2_X1 _17658_ (.A1(_11801_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .ZN(_11802_));
 AOI21_X1 _17659_ (.A(_11802_),
    .B1(_00520_),
    .B2(_11007_),
    .ZN(_11803_));
 BUF_X4 _17660_ (.A(_10998_),
    .Z(_11804_));
 BUF_X4 _17661_ (.A(_11804_),
    .Z(_11805_));
 AOI221_X2 _17662_ (.A(_11051_),
    .B1(_11755_),
    .B2(_11799_),
    .C1(_11803_),
    .C2(_11805_),
    .ZN(_11806_));
 NOR3_X2 _17663_ (.A1(_10988_),
    .A2(_11798_),
    .A3(_11806_),
    .ZN(_11807_));
 MUX2_X1 _17664_ (.A(_00537_),
    .B(_00539_),
    .S(_11240_),
    .Z(_11808_));
 MUX2_X1 _17665_ (.A(_00538_),
    .B(_00540_),
    .S(_11240_),
    .Z(_11809_));
 MUX2_X1 _17666_ (.A(_11808_),
    .B(_11809_),
    .S(_11260_),
    .Z(_11810_));
 MUX2_X1 _17667_ (.A(_00521_),
    .B(_00523_),
    .S(_11240_),
    .Z(_11811_));
 MUX2_X1 _17668_ (.A(_00522_),
    .B(_00524_),
    .S(_11240_),
    .Z(_11812_));
 MUX2_X1 _17669_ (.A(_11811_),
    .B(_11812_),
    .S(_11260_),
    .Z(_11813_));
 MUX2_X1 _17670_ (.A(_11810_),
    .B(_11813_),
    .S(_11780_),
    .Z(_11814_));
 NOR2_X1 _17671_ (.A1(_11174_),
    .A2(_11814_),
    .ZN(_11815_));
 NOR3_X4 _17672_ (.A1(_11055_),
    .A2(_11807_),
    .A3(_11815_),
    .ZN(_11816_));
 OR2_X1 _17673_ (.A1(_11792_),
    .A2(_11816_),
    .ZN(_11817_));
 BUF_X4 _17674_ (.A(_11277_),
    .Z(_11818_));
 NAND2_X1 _17675_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_11113_),
    .ZN(_11819_));
 OAI221_X2 _17676_ (.A(_11773_),
    .B1(_11817_),
    .B2(_11818_),
    .C1(_11819_),
    .C2(_11115_),
    .ZN(_16325_));
 INV_X2 _17677_ (.A(_16325_),
    .ZN(_16329_));
 INV_X1 _17678_ (.A(_16239_),
    .ZN(_16243_));
 NAND2_X1 _17679_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A2(_10957_),
    .ZN(_11820_));
 BUF_X4 _17680_ (.A(_11240_),
    .Z(_11821_));
 MUX2_X1 _17681_ (.A(_00274_),
    .B(_00276_),
    .S(_11821_),
    .Z(_11822_));
 MUX2_X1 _17682_ (.A(_00275_),
    .B(_00277_),
    .S(_11821_),
    .Z(_11823_));
 MUX2_X1 _17683_ (.A(_11822_),
    .B(_11823_),
    .S(_11075_),
    .Z(_11824_));
 MUX2_X1 _17684_ (.A(_00270_),
    .B(_00272_),
    .S(_11821_),
    .Z(_11825_));
 MUX2_X1 _17685_ (.A(_00271_),
    .B(_00273_),
    .S(_11821_),
    .Z(_11826_));
 MUX2_X1 _17686_ (.A(_11825_),
    .B(_11826_),
    .S(_11075_),
    .Z(_11827_));
 MUX2_X1 _17687_ (.A(_11824_),
    .B(_11827_),
    .S(_11073_),
    .Z(_11828_));
 MUX2_X1 _17688_ (.A(_00258_),
    .B(_00260_),
    .S(_11821_),
    .Z(_11829_));
 MUX2_X1 _17689_ (.A(_00259_),
    .B(_00261_),
    .S(_11821_),
    .Z(_11830_));
 MUX2_X1 _17690_ (.A(_11829_),
    .B(_11830_),
    .S(_11075_),
    .Z(_11831_));
 MUX2_X1 _17691_ (.A(_00254_),
    .B(_00256_),
    .S(_11821_),
    .Z(_11832_));
 MUX2_X1 _17692_ (.A(_00255_),
    .B(_00257_),
    .S(_11821_),
    .Z(_11833_));
 MUX2_X1 _17693_ (.A(_11832_),
    .B(_11833_),
    .S(_11075_),
    .Z(_11834_));
 MUX2_X1 _17694_ (.A(_11831_),
    .B(_11834_),
    .S(_11073_),
    .Z(_11835_));
 MUX2_X1 _17695_ (.A(_11828_),
    .B(_11835_),
    .S(_10982_),
    .Z(_11836_));
 NAND2_X2 _17696_ (.A1(_11056_),
    .A2(_11836_),
    .ZN(_11837_));
 BUF_X4 _17697_ (.A(_11037_),
    .Z(_11838_));
 MUX2_X1 _17698_ (.A(_00250_),
    .B(_00252_),
    .S(_11067_),
    .Z(_11839_));
 NOR2_X1 _17699_ (.A1(_11094_),
    .A2(_11839_),
    .ZN(_11840_));
 MUX2_X1 _17700_ (.A(_00251_),
    .B(_00253_),
    .S(_11067_),
    .Z(_11841_));
 NOR2_X1 _17701_ (.A1(_11013_),
    .A2(_11841_),
    .ZN(_11842_));
 NOR3_X1 _17702_ (.A1(_11838_),
    .A2(_11840_),
    .A3(_11842_),
    .ZN(_11843_));
 INV_X1 _17703_ (.A(_00248_),
    .ZN(_11844_));
 NOR2_X1 _17704_ (.A1(_11007_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .ZN(_11845_));
 AOI21_X1 _17705_ (.A(_11845_),
    .B1(_00249_),
    .B2(_11209_),
    .ZN(_11846_));
 AOI221_X2 _17706_ (.A(_11057_),
    .B1(_11844_),
    .B2(_11032_),
    .C1(_11846_),
    .C2(_11043_),
    .ZN(_11847_));
 NOR3_X1 _17707_ (.A1(_11053_),
    .A2(_11843_),
    .A3(_11847_),
    .ZN(_11848_));
 BUF_X4 _17708_ (.A(_11064_),
    .Z(_11849_));
 BUF_X4 _17709_ (.A(_11849_),
    .Z(_11850_));
 MUX2_X1 _17710_ (.A(_00266_),
    .B(_00268_),
    .S(_11850_),
    .Z(_11851_));
 MUX2_X1 _17711_ (.A(_00267_),
    .B(_00269_),
    .S(_11850_),
    .Z(_11852_));
 MUX2_X1 _17712_ (.A(_11851_),
    .B(_11852_),
    .S(_11000_),
    .Z(_11853_));
 MUX2_X1 _17713_ (.A(_00262_),
    .B(_00264_),
    .S(_11850_),
    .Z(_11854_));
 MUX2_X1 _17714_ (.A(_00263_),
    .B(_00265_),
    .S(_11850_),
    .Z(_11855_));
 MUX2_X1 _17715_ (.A(_11854_),
    .B(_11855_),
    .S(_11000_),
    .Z(_11856_));
 MUX2_X1 _17716_ (.A(_11853_),
    .B(_11856_),
    .S(_11037_),
    .Z(_11857_));
 NOR2_X1 _17717_ (.A1(_10982_),
    .A2(_11857_),
    .ZN(_11858_));
 OR3_X2 _17718_ (.A1(_11056_),
    .A2(_11848_),
    .A3(_11858_),
    .ZN(_11859_));
 AOI21_X1 _17719_ (.A(_11215_),
    .B1(_11837_),
    .B2(_11859_),
    .ZN(_11860_));
 OAI21_X1 _17720_ (.A(_11113_),
    .B1(_10978_),
    .B2(\cs_registers_i.pc_id_i[2] ),
    .ZN(_11861_));
 NAND2_X2 _17721_ (.A1(_11215_),
    .A2(_11282_),
    .ZN(_11862_));
 OAI221_X2 _17722_ (.A(_11820_),
    .B1(_11860_),
    .B2(_11861_),
    .C1(_11862_),
    .C2(_00182_),
    .ZN(_16254_));
 INV_X2 _17723_ (.A(_16254_),
    .ZN(_16258_));
 AND4_X4 _17724_ (.A1(_10945_),
    .A2(_10888_),
    .A3(net299),
    .A4(net296),
    .ZN(_11863_));
 NAND2_X4 _17725_ (.A1(_10955_),
    .A2(_11863_),
    .ZN(_11864_));
 BUF_X8 _17726_ (.A(_11864_),
    .Z(_11865_));
 NOR2_X2 _17727_ (.A1(_10881_),
    .A2(_10849_),
    .ZN(_11866_));
 INV_X1 _17728_ (.A(_00177_),
    .ZN(_11867_));
 AOI21_X1 _17729_ (.A(_11867_),
    .B1(_10883_),
    .B2(_10844_),
    .ZN(_11868_));
 NAND2_X1 _17730_ (.A1(_11866_),
    .A2(_11868_),
    .ZN(_11869_));
 NOR3_X2 _17731_ (.A1(_10872_),
    .A2(_11286_),
    .A3(_11869_),
    .ZN(_11870_));
 OAI33_X1 _17732_ (.A1(_10810_),
    .A2(_10795_),
    .A3(_10823_),
    .B1(_10894_),
    .B2(_10896_),
    .B3(_10898_),
    .ZN(_11871_));
 AND2_X1 _17733_ (.A1(_11293_),
    .A2(_11871_),
    .ZN(_11872_));
 OAI21_X2 _17734_ (.A(_10830_),
    .B1(_10899_),
    .B2(_10904_),
    .ZN(_11873_));
 AOI21_X4 _17735_ (.A(_11870_),
    .B1(_11872_),
    .B2(_11873_),
    .ZN(_11874_));
 NOR2_X2 _17736_ (.A1(net303),
    .A2(_10928_),
    .ZN(_11875_));
 OR2_X2 _17737_ (.A1(_10910_),
    .A2(_11875_),
    .ZN(_11876_));
 NOR2_X1 _17738_ (.A1(net303),
    .A2(_10826_),
    .ZN(_11877_));
 INV_X2 _17739_ (.A(_10869_),
    .ZN(_11878_));
 NAND3_X1 _17740_ (.A1(_10945_),
    .A2(_11878_),
    .A3(_10888_),
    .ZN(_11879_));
 AOI211_X2 _17741_ (.A(_11867_),
    .B(_10944_),
    .C1(_11877_),
    .C2(_11879_),
    .ZN(_11880_));
 OAI21_X1 _17742_ (.A(_10946_),
    .B1(_10885_),
    .B2(_10887_),
    .ZN(_11881_));
 NAND2_X1 _17743_ (.A1(_10883_),
    .A2(_11881_),
    .ZN(_11882_));
 AOI21_X4 _17744_ (.A(_10872_),
    .B1(_11880_),
    .B2(_11882_),
    .ZN(_11883_));
 AOI22_X2 _17745_ (.A1(_10881_),
    .A2(_10829_),
    .B1(_10918_),
    .B2(net413),
    .ZN(_11884_));
 OAI221_X2 _17746_ (.A(_10930_),
    .B1(_11884_),
    .B2(_10899_),
    .C1(_10937_),
    .C2(_10933_),
    .ZN(_11885_));
 NAND4_X1 _17747_ (.A1(_10778_),
    .A2(_10782_),
    .A3(_10789_),
    .A4(_10791_),
    .ZN(_11886_));
 OR4_X1 _17748_ (.A1(_10799_),
    .A2(_11286_),
    .A3(_11287_),
    .A4(_11886_),
    .ZN(_11887_));
 NAND2_X1 _17749_ (.A1(_10799_),
    .A2(net332),
    .ZN(_11888_));
 OR4_X1 _17750_ (.A1(_10894_),
    .A2(_10896_),
    .A3(_11886_),
    .A4(_11888_),
    .ZN(_11889_));
 NAND3_X1 _17751_ (.A1(_10910_),
    .A2(_11887_),
    .A3(_11889_),
    .ZN(_11890_));
 NAND3_X1 _17752_ (.A1(_10824_),
    .A2(_10830_),
    .A3(_10909_),
    .ZN(_11891_));
 NAND3_X1 _17753_ (.A1(net303),
    .A2(_10849_),
    .A3(_10850_),
    .ZN(_11892_));
 NAND3_X1 _17754_ (.A1(_10824_),
    .A2(_10909_),
    .A3(_11892_),
    .ZN(_11893_));
 AOI22_X2 _17755_ (.A1(_10844_),
    .A2(_11891_),
    .B1(_11893_),
    .B2(_10826_),
    .ZN(_11894_));
 AOI211_X2 _17756_ (.A(_11883_),
    .B(_11885_),
    .C1(_11890_),
    .C2(_11894_),
    .ZN(_11895_));
 NOR4_X4 _17757_ (.A1(_15764_),
    .A2(_11874_),
    .A3(_11876_),
    .A4(_11895_),
    .ZN(_11896_));
 BUF_X4 _17758_ (.A(_15767_),
    .Z(_11897_));
 OR3_X2 _17759_ (.A1(_10872_),
    .A2(_11286_),
    .A3(_11869_),
    .ZN(_11898_));
 NAND2_X2 _17760_ (.A1(_11293_),
    .A2(_11871_),
    .ZN(_11899_));
 NAND3_X2 _17761_ (.A1(_10776_),
    .A2(_10826_),
    .A3(net328),
    .ZN(_11900_));
 NOR2_X2 _17762_ (.A1(_10918_),
    .A2(_11900_),
    .ZN(_11901_));
 AOI21_X4 _17763_ (.A(_10851_),
    .B1(_10907_),
    .B2(_11901_),
    .ZN(_11902_));
 OAI21_X4 _17764_ (.A(_11898_),
    .B1(_11899_),
    .B2(_11902_),
    .ZN(_11903_));
 OAI22_X2 _17765_ (.A1(_10826_),
    .A2(_10850_),
    .B1(_10902_),
    .B2(_11900_),
    .ZN(_11904_));
 OR3_X1 _17766_ (.A1(_10854_),
    .A2(_10934_),
    .A3(_10936_),
    .ZN(_11905_));
 NOR2_X1 _17767_ (.A1(_10798_),
    .A2(_10802_),
    .ZN(_11906_));
 AOI21_X1 _17768_ (.A(_10779_),
    .B1(_10839_),
    .B2(_10790_),
    .ZN(_11907_));
 OAI21_X1 _17769_ (.A(_11906_),
    .B1(_10846_),
    .B2(_11907_),
    .ZN(_11908_));
 AOI221_X2 _17770_ (.A(_11283_),
    .B1(_11904_),
    .B2(_10907_),
    .C1(_11905_),
    .C2(_11908_),
    .ZN(_11909_));
 AND3_X1 _17771_ (.A1(_10910_),
    .A2(_11887_),
    .A3(_11889_),
    .ZN(_11910_));
 NOR3_X2 _17772_ (.A1(_10847_),
    .A2(_10851_),
    .A3(_10942_),
    .ZN(_11911_));
 AND3_X1 _17773_ (.A1(_10824_),
    .A2(_10909_),
    .A3(_11892_),
    .ZN(_11912_));
 OAI22_X4 _17774_ (.A1(net303),
    .A2(_11911_),
    .B1(_11912_),
    .B2(_10881_),
    .ZN(_11913_));
 AND2_X1 _17775_ (.A1(_11880_),
    .A2(_11882_),
    .ZN(_11914_));
 OAI221_X2 _17776_ (.A(_11909_),
    .B1(_11910_),
    .B2(_11913_),
    .C1(_11914_),
    .C2(_10872_),
    .ZN(_11915_));
 BUF_X4 _17777_ (.A(_11915_),
    .Z(_11916_));
 NOR4_X4 _17778_ (.A1(_11897_),
    .A2(_11903_),
    .A3(_11876_),
    .A4(_11916_),
    .ZN(_11917_));
 OR2_X2 _17779_ (.A1(_11896_),
    .A2(_11917_),
    .ZN(_11918_));
 NOR3_X2 _17780_ (.A1(_10847_),
    .A2(_10942_),
    .A3(_11875_),
    .ZN(_11919_));
 OR2_X2 _17781_ (.A1(_15762_),
    .A2(_11919_),
    .ZN(_11920_));
 BUF_X4 _17782_ (.A(_11895_),
    .Z(_11921_));
 AND2_X1 _17783_ (.A1(_10943_),
    .A2(_11875_),
    .ZN(_11922_));
 OAI33_X1 _17784_ (.A1(_11903_),
    .A2(_11920_),
    .A3(_11921_),
    .B1(_11922_),
    .B2(_11883_),
    .B3(_11885_),
    .ZN(_11923_));
 NOR3_X4 _17785_ (.A1(_10943_),
    .A2(_11883_),
    .A3(_11885_),
    .ZN(_11924_));
 OAI221_X2 _17786_ (.A(_11898_),
    .B1(_11899_),
    .B2(_11902_),
    .C1(_11910_),
    .C2(_11913_),
    .ZN(_11925_));
 CLKBUF_X3 _17787_ (.A(_15769_),
    .Z(_11926_));
 INV_X1 _17788_ (.A(_11926_),
    .ZN(_11927_));
 OAI21_X2 _17789_ (.A(_11924_),
    .B1(_11925_),
    .B2(_11927_),
    .ZN(_11928_));
 NAND2_X4 _17790_ (.A1(net9),
    .A2(_11928_),
    .ZN(_11929_));
 OAI21_X2 _17791_ (.A(_11865_),
    .B1(_11918_),
    .B2(_11929_),
    .ZN(_14464_));
 NAND2_X1 _17792_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(_10957_),
    .ZN(_11930_));
 BUF_X8 _17793_ (.A(_11052_),
    .Z(_11931_));
 MUX2_X1 _17794_ (.A(_00297_),
    .B(_00299_),
    .S(_11254_),
    .Z(_11932_));
 MUX2_X1 _17795_ (.A(_00298_),
    .B(_00300_),
    .S(_11254_),
    .Z(_11933_));
 MUX2_X1 _17796_ (.A(_11932_),
    .B(_11933_),
    .S(_11094_),
    .Z(_11934_));
 NAND2_X1 _17797_ (.A1(_11085_),
    .A2(_11934_),
    .ZN(_11935_));
 MUX2_X1 _17798_ (.A(_00295_),
    .B(_00296_),
    .S(_11094_),
    .Z(_11936_));
 MUX2_X1 _17799_ (.A(_00293_),
    .B(_00294_),
    .S(_11001_),
    .Z(_11937_));
 AOI22_X2 _17800_ (.A1(_11100_),
    .A2(_11936_),
    .B1(_11937_),
    .B2(_11091_),
    .ZN(_11938_));
 MUX2_X1 _17801_ (.A(_00307_),
    .B(_00308_),
    .S(_11027_),
    .Z(_11939_));
 AOI21_X1 _17802_ (.A(_11037_),
    .B1(_11939_),
    .B2(_11068_),
    .ZN(_11940_));
 MUX2_X1 _17803_ (.A(_00305_),
    .B(_00306_),
    .S(_11093_),
    .Z(_11941_));
 INV_X1 _17804_ (.A(_11941_),
    .ZN(_11942_));
 MUX2_X1 _17805_ (.A(_00303_),
    .B(_00304_),
    .S(_11271_),
    .Z(_11943_));
 AOI21_X1 _17806_ (.A(_11057_),
    .B1(_11943_),
    .B2(_11068_),
    .ZN(_11944_));
 MUX2_X1 _17807_ (.A(_00301_),
    .B(_00302_),
    .S(_11000_),
    .Z(_11945_));
 INV_X1 _17808_ (.A(_11945_),
    .ZN(_11946_));
 AOI22_X1 _17809_ (.A1(_11940_),
    .A2(_11942_),
    .B1(_11944_),
    .B2(_11946_),
    .ZN(_11947_));
 OAI21_X1 _17810_ (.A(_11081_),
    .B1(_11940_),
    .B2(_11944_),
    .ZN(_11948_));
 NAND3_X1 _17811_ (.A1(_11055_),
    .A2(_11947_),
    .A3(_11948_),
    .ZN(_11949_));
 NAND4_X2 _17812_ (.A1(_11931_),
    .A2(_11935_),
    .A3(_11938_),
    .A4(_11949_),
    .ZN(_11950_));
 MUX2_X1 _17813_ (.A(_00287_),
    .B(_00291_),
    .S(_10985_),
    .Z(_11951_));
 MUX2_X1 _17814_ (.A(_00288_),
    .B(_00292_),
    .S(_10985_),
    .Z(_11952_));
 MUX2_X1 _17815_ (.A(_11951_),
    .B(_11952_),
    .S(_11027_),
    .Z(_11953_));
 MUX2_X1 _17816_ (.A(_00285_),
    .B(_00289_),
    .S(_10985_),
    .Z(_11954_));
 MUX2_X1 _17817_ (.A(_00286_),
    .B(_00290_),
    .S(_10985_),
    .Z(_11955_));
 MUX2_X1 _17818_ (.A(_11954_),
    .B(_11955_),
    .S(_11027_),
    .Z(_11956_));
 MUX2_X1 _17819_ (.A(_11953_),
    .B(_11956_),
    .S(_11029_),
    .Z(_11957_));
 NOR2_X1 _17820_ (.A1(_10995_),
    .A2(_11957_),
    .ZN(_11958_));
 NOR2_X1 _17821_ (.A1(_11007_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .ZN(_11959_));
 AOI21_X1 _17822_ (.A(_11959_),
    .B1(_00280_),
    .B2(_11209_),
    .ZN(_11960_));
 AOI221_X1 _17823_ (.A(_10986_),
    .B1(_11394_),
    .B2(_11032_),
    .C1(_11960_),
    .C2(_11043_),
    .ZN(_11961_));
 MUX2_X1 _17824_ (.A(_00281_),
    .B(_00283_),
    .S(_11209_),
    .Z(_11962_));
 MUX2_X1 _17825_ (.A(_00282_),
    .B(_00284_),
    .S(_11209_),
    .Z(_11963_));
 MUX2_X1 _17826_ (.A(_11962_),
    .B(_11963_),
    .S(_11094_),
    .Z(_11964_));
 AOI21_X1 _17827_ (.A(_11961_),
    .B1(_11964_),
    .B2(_10988_),
    .ZN(_11965_));
 AOI21_X2 _17828_ (.A(_11958_),
    .B1(_11965_),
    .B2(_10995_),
    .ZN(_11966_));
 OAI21_X4 _17829_ (.A(_11950_),
    .B1(_11966_),
    .B2(_11931_),
    .ZN(_11967_));
 NOR2_X1 _17830_ (.A1(_11215_),
    .A2(_11967_),
    .ZN(_11968_));
 BUF_X2 _17831_ (.A(\cs_registers_i.pc_id_i[3] ),
    .Z(_11969_));
 OAI21_X1 _17832_ (.A(_11113_),
    .B1(_11115_),
    .B2(_11969_),
    .ZN(_11970_));
 OAI221_X2 _17833_ (.A(_11930_),
    .B1(_11968_),
    .B2(_11970_),
    .C1(_11862_),
    .C2(_00181_),
    .ZN(_11971_));
 BUF_X4 _17834_ (.A(_11971_),
    .Z(_16261_));
 INV_X1 _17835_ (.A(_16261_),
    .ZN(_16265_));
 NOR2_X1 _17836_ (.A1(_00180_),
    .A2(_11862_),
    .ZN(_11972_));
 NOR2_X2 _17837_ (.A1(_11215_),
    .A2(_11216_),
    .ZN(_11973_));
 MUX2_X1 _17838_ (.A(_00315_),
    .B(_00317_),
    .S(_11004_),
    .Z(_11974_));
 NOR2_X1 _17839_ (.A1(_10998_),
    .A2(_11974_),
    .ZN(_11975_));
 MUX2_X1 _17840_ (.A(_00316_),
    .B(_00318_),
    .S(_11004_),
    .Z(_11976_));
 NOR2_X1 _17841_ (.A1(_11011_),
    .A2(_11976_),
    .ZN(_11977_));
 NOR3_X1 _17842_ (.A1(_10992_),
    .A2(_11975_),
    .A3(_11977_),
    .ZN(_11978_));
 INV_X1 _17843_ (.A(_00309_),
    .ZN(_11979_));
 NOR2_X1 _17844_ (.A1(_11004_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .ZN(_11980_));
 AOI21_X1 _17845_ (.A(_11980_),
    .B1(_00310_),
    .B2(_11244_),
    .ZN(_11981_));
 AOI221_X1 _17846_ (.A(_11021_),
    .B1(_11979_),
    .B2(_11030_),
    .C1(_11981_),
    .C2(_11025_),
    .ZN(_11982_));
 NOR3_X1 _17847_ (.A1(_10986_),
    .A2(_11978_),
    .A3(_11982_),
    .ZN(_11983_));
 MUX2_X1 _17848_ (.A(_00319_),
    .B(_00321_),
    .S(_11063_),
    .Z(_11984_));
 MUX2_X1 _17849_ (.A(_00320_),
    .B(_00322_),
    .S(_11063_),
    .Z(_11985_));
 MUX2_X1 _17850_ (.A(_11984_),
    .B(_11985_),
    .S(_10997_),
    .Z(_11986_));
 MUX2_X1 _17851_ (.A(_00311_),
    .B(_00313_),
    .S(_11063_),
    .Z(_11987_));
 MUX2_X1 _17852_ (.A(_00312_),
    .B(_00314_),
    .S(_11063_),
    .Z(_11988_));
 MUX2_X1 _17853_ (.A(_11987_),
    .B(_11988_),
    .S(_10997_),
    .Z(_11989_));
 MUX2_X1 _17854_ (.A(_11986_),
    .B(_11989_),
    .S(_10992_),
    .Z(_11990_));
 NOR2_X1 _17855_ (.A1(_11036_),
    .A2(_11990_),
    .ZN(_11991_));
 NOR3_X2 _17856_ (.A1(_11052_),
    .A2(_11983_),
    .A3(_11991_),
    .ZN(_11992_));
 MUX2_X1 _17857_ (.A(_00331_),
    .B(_00333_),
    .S(_11063_),
    .Z(_11993_));
 MUX2_X1 _17858_ (.A(_00332_),
    .B(_00334_),
    .S(_11238_),
    .Z(_11994_));
 MUX2_X1 _17859_ (.A(_11993_),
    .B(_11994_),
    .S(_10997_),
    .Z(_11995_));
 MUX2_X1 _17860_ (.A(_00323_),
    .B(_00325_),
    .S(_11063_),
    .Z(_11996_));
 MUX2_X1 _17861_ (.A(_00324_),
    .B(_00326_),
    .S(_11238_),
    .Z(_11997_));
 MUX2_X1 _17862_ (.A(_11996_),
    .B(_11997_),
    .S(_10997_),
    .Z(_11998_));
 MUX2_X1 _17863_ (.A(_11995_),
    .B(_11998_),
    .S(_10992_),
    .Z(_11999_));
 MUX2_X1 _17864_ (.A(_00335_),
    .B(_00337_),
    .S(_11238_),
    .Z(_12000_));
 MUX2_X1 _17865_ (.A(_00336_),
    .B(_00338_),
    .S(_11238_),
    .Z(_12001_));
 MUX2_X1 _17866_ (.A(_12000_),
    .B(_12001_),
    .S(_10997_),
    .Z(_12002_));
 MUX2_X1 _17867_ (.A(_00327_),
    .B(_00329_),
    .S(_11238_),
    .Z(_12003_));
 MUX2_X1 _17868_ (.A(_00328_),
    .B(_00330_),
    .S(_11238_),
    .Z(_12004_));
 MUX2_X1 _17869_ (.A(_12003_),
    .B(_12004_),
    .S(_11025_),
    .Z(_12005_));
 MUX2_X1 _17870_ (.A(_12002_),
    .B(_12005_),
    .S(_10992_),
    .Z(_12006_));
 MUX2_X2 _17871_ (.A(_11999_),
    .B(_12006_),
    .S(_10986_),
    .Z(_12007_));
 AOI21_X4 _17872_ (.A(_11992_),
    .B1(_12007_),
    .B2(_11052_),
    .ZN(_12008_));
 AND2_X1 _17873_ (.A1(_11973_),
    .A2(_12008_),
    .ZN(_12009_));
 NAND2_X1 _17874_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .A2(_10819_),
    .ZN(_12010_));
 BUF_X1 _17875_ (.A(\cs_registers_i.pc_id_i[4] ),
    .Z(_12011_));
 NAND2_X1 _17876_ (.A1(_12011_),
    .A2(_11111_),
    .ZN(_12012_));
 OAI21_X1 _17877_ (.A(_12010_),
    .B1(_12012_),
    .B2(_10977_),
    .ZN(_12013_));
 OR3_X1 _17878_ (.A1(_11972_),
    .A2(_12009_),
    .A3(_12013_),
    .ZN(_12014_));
 CLKBUF_X3 _17879_ (.A(_12014_),
    .Z(_16269_));
 INV_X2 _17880_ (.A(_16269_),
    .ZN(_16273_));
 AND3_X1 _17881_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(_11215_),
    .A3(_11111_),
    .ZN(_12015_));
 MUX2_X1 _17882_ (.A(_00353_),
    .B(_00355_),
    .S(_11096_),
    .Z(_12016_));
 NOR2_X1 _17883_ (.A1(_11269_),
    .A2(_12016_),
    .ZN(_12017_));
 MUX2_X1 _17884_ (.A(_00354_),
    .B(_00356_),
    .S(_11783_),
    .Z(_12018_));
 NOR2_X1 _17885_ (.A1(_11012_),
    .A2(_12018_),
    .ZN(_12019_));
 NOR3_X1 _17886_ (.A1(_10980_),
    .A2(_12017_),
    .A3(_12019_),
    .ZN(_12020_));
 NOR2_X1 _17887_ (.A1(_11245_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .ZN(_12021_));
 AOI21_X1 _17888_ (.A(_12021_),
    .B1(_00340_),
    .B2(_11066_),
    .ZN(_12022_));
 AOI221_X1 _17889_ (.A(_11051_),
    .B1(_11519_),
    .B2(_11031_),
    .C1(_12022_),
    .C2(_11092_),
    .ZN(_12023_));
 NOR3_X1 _17890_ (.A1(_10987_),
    .A2(_12020_),
    .A3(_12023_),
    .ZN(_12024_));
 MUX2_X1 _17891_ (.A(_00357_),
    .B(_00359_),
    .S(_11239_),
    .Z(_12025_));
 MUX2_X1 _17892_ (.A(_00358_),
    .B(_00360_),
    .S(_11239_),
    .Z(_12026_));
 MUX2_X1 _17893_ (.A(_12025_),
    .B(_12026_),
    .S(_11059_),
    .Z(_12027_));
 MUX2_X1 _17894_ (.A(_00341_),
    .B(_00343_),
    .S(_11014_),
    .Z(_12028_));
 MUX2_X1 _17895_ (.A(_00342_),
    .B(_00344_),
    .S(_11014_),
    .Z(_12029_));
 MUX2_X1 _17896_ (.A(_12028_),
    .B(_12029_),
    .S(_11059_),
    .Z(_12030_));
 MUX2_X1 _17897_ (.A(_12027_),
    .B(_12030_),
    .S(_10980_),
    .Z(_12031_));
 NOR2_X1 _17898_ (.A1(_11037_),
    .A2(_12031_),
    .ZN(_12032_));
 NOR3_X2 _17899_ (.A1(_11252_),
    .A2(_12024_),
    .A3(_12032_),
    .ZN(_12033_));
 BUF_X4 _17900_ (.A(_11004_),
    .Z(_12034_));
 MUX2_X1 _17901_ (.A(_00361_),
    .B(_00363_),
    .S(_12034_),
    .Z(_12035_));
 MUX2_X1 _17902_ (.A(_00362_),
    .B(_00364_),
    .S(_12034_),
    .Z(_12036_));
 BUF_X4 _17903_ (.A(_11025_),
    .Z(_12037_));
 MUX2_X1 _17904_ (.A(_12035_),
    .B(_12036_),
    .S(_12037_),
    .Z(_12038_));
 MUX2_X1 _17905_ (.A(_00345_),
    .B(_00347_),
    .S(_12034_),
    .Z(_12039_));
 MUX2_X1 _17906_ (.A(_00346_),
    .B(_00348_),
    .S(_11224_),
    .Z(_12040_));
 MUX2_X1 _17907_ (.A(_12039_),
    .B(_12040_),
    .S(_12037_),
    .Z(_12041_));
 MUX2_X1 _17908_ (.A(_12038_),
    .B(_12041_),
    .S(_10980_),
    .Z(_12042_));
 MUX2_X1 _17909_ (.A(_00365_),
    .B(_00367_),
    .S(_12034_),
    .Z(_12043_));
 MUX2_X1 _17910_ (.A(_00366_),
    .B(_00368_),
    .S(_11224_),
    .Z(_12044_));
 MUX2_X1 _17911_ (.A(_12043_),
    .B(_12044_),
    .S(_12037_),
    .Z(_12045_));
 MUX2_X1 _17912_ (.A(_00349_),
    .B(_00351_),
    .S(_11224_),
    .Z(_12046_));
 MUX2_X1 _17913_ (.A(_00350_),
    .B(_00352_),
    .S(_11224_),
    .Z(_12047_));
 MUX2_X1 _17914_ (.A(_12046_),
    .B(_12047_),
    .S(_11227_),
    .Z(_12048_));
 MUX2_X1 _17915_ (.A(_12045_),
    .B(_12048_),
    .S(_10980_),
    .Z(_12049_));
 MUX2_X2 _17916_ (.A(_12042_),
    .B(_12049_),
    .S(_10987_),
    .Z(_12050_));
 AOI21_X4 _17917_ (.A(_12033_),
    .B1(_12050_),
    .B2(_11055_),
    .ZN(_12051_));
 AOI221_X2 _17918_ (.A(_12015_),
    .B1(_12051_),
    .B2(_11973_),
    .C1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .C2(_10958_),
    .ZN(_16281_));
 NAND2_X1 _17919_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(_10958_),
    .ZN(_12052_));
 MUX2_X1 _17920_ (.A(_00391_),
    .B(_00393_),
    .S(_11005_),
    .Z(_12053_));
 MUX2_X1 _17921_ (.A(_00392_),
    .B(_00394_),
    .S(_11005_),
    .Z(_12054_));
 MUX2_X1 _17922_ (.A(_12053_),
    .B(_12054_),
    .S(_12037_),
    .Z(_12055_));
 MUX2_X1 _17923_ (.A(_00383_),
    .B(_00385_),
    .S(_11005_),
    .Z(_12056_));
 MUX2_X1 _17924_ (.A(_00384_),
    .B(_00386_),
    .S(_12034_),
    .Z(_12057_));
 MUX2_X1 _17925_ (.A(_12056_),
    .B(_12057_),
    .S(_12037_),
    .Z(_12058_));
 MUX2_X1 _17926_ (.A(_12055_),
    .B(_12058_),
    .S(_11232_),
    .Z(_12059_));
 NOR2_X1 _17927_ (.A1(_11058_),
    .A2(_12059_),
    .ZN(_12060_));
 BUF_X4 _17928_ (.A(_11004_),
    .Z(_12061_));
 MUX2_X1 _17929_ (.A(_00395_),
    .B(_00397_),
    .S(_12061_),
    .Z(_12062_));
 MUX2_X1 _17930_ (.A(_00396_),
    .B(_00398_),
    .S(_12061_),
    .Z(_12063_));
 MUX2_X1 _17931_ (.A(_12062_),
    .B(_12063_),
    .S(_11026_),
    .Z(_12064_));
 MUX2_X1 _17932_ (.A(_00387_),
    .B(_00389_),
    .S(_12061_),
    .Z(_12065_));
 MUX2_X1 _17933_ (.A(_00388_),
    .B(_00390_),
    .S(_12061_),
    .Z(_12066_));
 MUX2_X1 _17934_ (.A(_12065_),
    .B(_12066_),
    .S(_11026_),
    .Z(_12067_));
 BUF_X4 _17935_ (.A(_10992_),
    .Z(_12068_));
 MUX2_X1 _17936_ (.A(_12064_),
    .B(_12067_),
    .S(_12068_),
    .Z(_12069_));
 NOR2_X1 _17937_ (.A1(_11073_),
    .A2(_12069_),
    .ZN(_12070_));
 NOR3_X4 _17938_ (.A1(_10981_),
    .A2(_12060_),
    .A3(_12070_),
    .ZN(_12071_));
 MUX2_X1 _17939_ (.A(_00375_),
    .B(_00377_),
    .S(_11015_),
    .Z(_12072_));
 NOR2_X1 _17940_ (.A1(_11000_),
    .A2(_12072_),
    .ZN(_12073_));
 MUX2_X1 _17941_ (.A(_00376_),
    .B(_00378_),
    .S(_11015_),
    .Z(_12074_));
 NOR2_X1 _17942_ (.A1(_11012_),
    .A2(_12074_),
    .ZN(_12075_));
 NOR3_X2 _17943_ (.A1(_10993_),
    .A2(_12073_),
    .A3(_12075_),
    .ZN(_12076_));
 INV_X1 _17944_ (.A(_00369_),
    .ZN(_12077_));
 NOR2_X1 _17945_ (.A1(_11240_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .ZN(_12078_));
 AOI21_X2 _17946_ (.A(_12078_),
    .B1(_00370_),
    .B2(_11801_),
    .ZN(_12079_));
 AOI221_X2 _17947_ (.A(_11021_),
    .B1(_12077_),
    .B2(_11031_),
    .C1(_12079_),
    .C2(_11074_),
    .ZN(_12080_));
 NOR3_X4 _17948_ (.A1(_10987_),
    .A2(_12076_),
    .A3(_12080_),
    .ZN(_12081_));
 MUX2_X1 _17949_ (.A(_00379_),
    .B(_00381_),
    .S(_11014_),
    .Z(_12082_));
 MUX2_X1 _17950_ (.A(_00380_),
    .B(_00382_),
    .S(_11014_),
    .Z(_12083_));
 MUX2_X1 _17951_ (.A(_12082_),
    .B(_12083_),
    .S(_11041_),
    .Z(_12084_));
 BUF_X4 _17952_ (.A(_11004_),
    .Z(_12085_));
 MUX2_X1 _17953_ (.A(_00371_),
    .B(_00373_),
    .S(_12085_),
    .Z(_12086_));
 MUX2_X1 _17954_ (.A(_00372_),
    .B(_00374_),
    .S(_12085_),
    .Z(_12087_));
 MUX2_X1 _17955_ (.A(_12086_),
    .B(_12087_),
    .S(_11041_),
    .Z(_12088_));
 MUX2_X1 _17956_ (.A(_12084_),
    .B(_12088_),
    .S(_12068_),
    .Z(_12089_));
 NOR2_X2 _17957_ (.A1(_11073_),
    .A2(_12089_),
    .ZN(_12090_));
 NOR3_X4 _17958_ (.A1(_11052_),
    .A2(_12081_),
    .A3(_12090_),
    .ZN(_12091_));
 OR2_X2 _17959_ (.A1(_12071_),
    .A2(_12091_),
    .ZN(_12092_));
 NAND2_X1 _17960_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(_11112_),
    .ZN(_12093_));
 OAI221_X1 _17961_ (.A(_12052_),
    .B1(_12092_),
    .B2(_11277_),
    .C1(_12093_),
    .C2(_11114_),
    .ZN(_12094_));
 CLKBUF_X3 _17962_ (.A(_12094_),
    .Z(_16285_));
 INV_X1 _17963_ (.A(_16285_),
    .ZN(_16289_));
 NAND2_X1 _17964_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(_11221_),
    .ZN(_12095_));
 MUX2_X1 _17965_ (.A(_00421_),
    .B(_00423_),
    .S(_11849_),
    .Z(_12096_));
 MUX2_X1 _17966_ (.A(_00422_),
    .B(_00424_),
    .S(_11849_),
    .Z(_12097_));
 BUF_X4 _17967_ (.A(_10998_),
    .Z(_12098_));
 MUX2_X1 _17968_ (.A(_12096_),
    .B(_12097_),
    .S(_12098_),
    .Z(_12099_));
 BUF_X4 _17969_ (.A(_11064_),
    .Z(_12100_));
 MUX2_X1 _17970_ (.A(_00413_),
    .B(_00415_),
    .S(_12100_),
    .Z(_12101_));
 MUX2_X1 _17971_ (.A(_00414_),
    .B(_00416_),
    .S(_12100_),
    .Z(_12102_));
 MUX2_X1 _17972_ (.A(_12101_),
    .B(_12102_),
    .S(_12098_),
    .Z(_12103_));
 BUF_X4 _17973_ (.A(_10992_),
    .Z(_12104_));
 MUX2_X1 _17974_ (.A(_12099_),
    .B(_12103_),
    .S(_12104_),
    .Z(_12105_));
 NOR2_X1 _17975_ (.A1(_11177_),
    .A2(_12105_),
    .ZN(_12106_));
 BUF_X4 _17976_ (.A(_11064_),
    .Z(_12107_));
 MUX2_X1 _17977_ (.A(_00425_),
    .B(_00427_),
    .S(_12107_),
    .Z(_12108_));
 MUX2_X1 _17978_ (.A(_00426_),
    .B(_00428_),
    .S(_12107_),
    .Z(_12109_));
 MUX2_X1 _17979_ (.A(_12108_),
    .B(_12109_),
    .S(_10999_),
    .Z(_12110_));
 MUX2_X1 _17980_ (.A(_00417_),
    .B(_00419_),
    .S(_12107_),
    .Z(_12111_));
 MUX2_X1 _17981_ (.A(_00418_),
    .B(_00420_),
    .S(_12107_),
    .Z(_12112_));
 MUX2_X1 _17982_ (.A(_12111_),
    .B(_12112_),
    .S(_10999_),
    .Z(_12113_));
 MUX2_X1 _17983_ (.A(_12110_),
    .B(_12113_),
    .S(_12104_),
    .Z(_12114_));
 NOR2_X1 _17984_ (.A1(_11838_),
    .A2(_12114_),
    .ZN(_12115_));
 NOR3_X4 _17985_ (.A1(_10982_),
    .A2(_12106_),
    .A3(_12115_),
    .ZN(_12116_));
 BUF_X4 _17986_ (.A(_12068_),
    .Z(_12117_));
 MUX2_X1 _17987_ (.A(_00405_),
    .B(_00407_),
    .S(_11066_),
    .Z(_12118_));
 NOR2_X1 _17988_ (.A1(_11093_),
    .A2(_12118_),
    .ZN(_12119_));
 MUX2_X1 _17989_ (.A(_00406_),
    .B(_00408_),
    .S(_11006_),
    .Z(_12120_));
 NOR2_X1 _17990_ (.A1(_11795_),
    .A2(_12120_),
    .ZN(_12121_));
 NOR3_X1 _17991_ (.A1(_12117_),
    .A2(_12119_),
    .A3(_12121_),
    .ZN(_12122_));
 NOR2_X1 _17992_ (.A1(_11015_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .ZN(_12123_));
 AOI21_X1 _17993_ (.A(_12123_),
    .B1(_00400_),
    .B2(_11246_),
    .ZN(_12124_));
 AOI221_X2 _17994_ (.A(_11235_),
    .B1(_11596_),
    .B2(_11031_),
    .C1(_12124_),
    .C2(_11271_),
    .ZN(_12125_));
 NOR3_X2 _17995_ (.A1(_11058_),
    .A2(_12122_),
    .A3(_12125_),
    .ZN(_12126_));
 MUX2_X1 _17996_ (.A(_00409_),
    .B(_00411_),
    .S(_11065_),
    .Z(_12127_));
 MUX2_X1 _17997_ (.A(_00410_),
    .B(_00412_),
    .S(_11065_),
    .Z(_12128_));
 MUX2_X1 _17998_ (.A(_12127_),
    .B(_12128_),
    .S(_11227_),
    .Z(_12129_));
 MUX2_X1 _17999_ (.A(_00401_),
    .B(_00403_),
    .S(_11065_),
    .Z(_12130_));
 MUX2_X1 _18000_ (.A(_00402_),
    .B(_00404_),
    .S(_11065_),
    .Z(_12131_));
 MUX2_X1 _18001_ (.A(_12130_),
    .B(_12131_),
    .S(_11227_),
    .Z(_12132_));
 MUX2_X1 _18002_ (.A(_12129_),
    .B(_12132_),
    .S(_11232_),
    .Z(_12133_));
 NOR2_X1 _18003_ (.A1(_11223_),
    .A2(_12133_),
    .ZN(_12134_));
 NOR3_X4 _18004_ (.A1(_11052_),
    .A2(_12126_),
    .A3(_12134_),
    .ZN(_12135_));
 OR2_X2 _18005_ (.A1(_12116_),
    .A2(_12135_),
    .ZN(_12136_));
 NAND2_X1 _18006_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_11112_),
    .ZN(_12137_));
 OAI221_X2 _18007_ (.A(_12095_),
    .B1(_12136_),
    .B2(_11278_),
    .C1(_12137_),
    .C2(_11114_),
    .ZN(_16293_));
 INV_X2 _18008_ (.A(_16293_),
    .ZN(_16297_));
 BUF_X4 _18009_ (.A(_15800_),
    .Z(_12138_));
 INV_X1 _18010_ (.A(_15795_),
    .ZN(_12139_));
 BUF_X4 _18011_ (.A(_15796_),
    .Z(_12140_));
 CLKBUF_X2 _18012_ (.A(_15791_),
    .Z(_12141_));
 BUF_X4 _18013_ (.A(_15792_),
    .Z(_12142_));
 BUF_X4 rebuffer34 (.A(_10787_),
    .Z(net308));
 OAI21_X1 _18015_ (.A(_12142_),
    .B1(_15787_),
    .B2(_15788_),
    .ZN(_12144_));
 INV_X1 _18016_ (.A(_12144_),
    .ZN(_12145_));
 OR2_X1 _18017_ (.A1(_15783_),
    .A2(_15787_),
    .ZN(_12146_));
 OR2_X1 _18018_ (.A1(_12141_),
    .A2(_12146_),
    .ZN(_12147_));
 BUF_X4 _18019_ (.A(_15784_),
    .Z(_12148_));
 INV_X1 _18020_ (.A(_15779_),
    .ZN(_12149_));
 AOI21_X4 _18021_ (.A(_15773_),
    .B1(_14467_),
    .B2(_11220_),
    .ZN(_12150_));
 BUF_X4 _18022_ (.A(_15780_),
    .Z(_12151_));
 INV_X2 _18023_ (.A(_12151_),
    .ZN(_12152_));
 OAI21_X4 _18024_ (.A(_12149_),
    .B1(_12150_),
    .B2(_12152_),
    .ZN(_12153_));
 AND2_X1 _18025_ (.A1(_12148_),
    .A2(_12153_),
    .ZN(_12154_));
 OAI221_X2 _18026_ (.A(_12140_),
    .B1(_12141_),
    .B2(_12145_),
    .C1(_12147_),
    .C2(_12154_),
    .ZN(_12155_));
 AND2_X1 _18027_ (.A1(_12139_),
    .A2(_12155_),
    .ZN(_12156_));
 XNOR2_X2 _18028_ (.A(_12138_),
    .B(_12156_),
    .ZN(\alu_adder_result_ex[7] ));
 INV_X1 _18029_ (.A(_12141_),
    .ZN(_12157_));
 INV_X1 _18030_ (.A(_15787_),
    .ZN(_12158_));
 AOI21_X1 _18031_ (.A(_15783_),
    .B1(_15779_),
    .B2(_12148_),
    .ZN(_12159_));
 INV_X1 _18032_ (.A(net347),
    .ZN(_12160_));
 OAI21_X1 _18033_ (.A(_12158_),
    .B1(_12159_),
    .B2(_12160_),
    .ZN(_12161_));
 NAND2_X1 _18034_ (.A1(_12142_),
    .A2(_12161_),
    .ZN(_12162_));
 NAND2_X1 _18035_ (.A1(_12157_),
    .A2(_12162_),
    .ZN(_12163_));
 NAND4_X4 _18036_ (.A1(net347),
    .A2(_12148_),
    .A3(_12151_),
    .A4(_12142_),
    .ZN(_12164_));
 AND3_X1 _18037_ (.A1(net298),
    .A2(_10871_),
    .A3(_11863_),
    .ZN(_12165_));
 AND2_X1 _18038_ (.A1(_15776_),
    .A2(_11220_),
    .ZN(_12166_));
 NAND2_X1 _18039_ (.A1(_12165_),
    .A2(_12166_),
    .ZN(_12167_));
 AOI21_X4 _18040_ (.A(_15773_),
    .B1(_15775_),
    .B2(_11220_),
    .ZN(_12168_));
 AOI21_X1 _18041_ (.A(_12164_),
    .B1(_12167_),
    .B2(_12168_),
    .ZN(_12169_));
 OAI21_X1 _18042_ (.A(_12140_),
    .B1(_12163_),
    .B2(_12169_),
    .ZN(_12170_));
 NAND2_X2 _18043_ (.A1(_15776_),
    .A2(_11220_),
    .ZN(_12171_));
 AOI21_X1 _18044_ (.A(_12164_),
    .B1(_12171_),
    .B2(_12168_),
    .ZN(_12172_));
 OR2_X1 _18045_ (.A1(_12163_),
    .A2(_12172_),
    .ZN(_12173_));
 OAI21_X1 _18046_ (.A(_12170_),
    .B1(_12173_),
    .B2(_12140_),
    .ZN(_12174_));
 AND2_X1 _18047_ (.A1(net9),
    .A2(_11928_),
    .ZN(_12175_));
 BUF_X4 _18048_ (.A(_12175_),
    .Z(_12176_));
 NOR2_X2 _18049_ (.A1(_11896_),
    .A2(_11917_),
    .ZN(_12177_));
 NOR2_X2 _18050_ (.A1(_12171_),
    .A2(_12164_),
    .ZN(_12178_));
 AND4_X1 _18051_ (.A1(_12140_),
    .A2(_12176_),
    .A3(_12177_),
    .A4(_12178_),
    .ZN(_12179_));
 NAND2_X1 _18052_ (.A1(_12176_),
    .A2(_12177_),
    .ZN(_12180_));
 NAND2_X1 _18053_ (.A1(_12168_),
    .A2(_12167_),
    .ZN(_12181_));
 NOR3_X1 _18054_ (.A1(_12140_),
    .A2(_12181_),
    .A3(_12163_),
    .ZN(_12182_));
 AOI211_X2 _18055_ (.A(_12174_),
    .B(_12179_),
    .C1(_12180_),
    .C2(_12182_),
    .ZN(\alu_adder_result_ex[6] ));
 NAND2_X1 _18056_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(_10958_),
    .ZN(_12183_));
 MUX2_X1 _18057_ (.A(_00451_),
    .B(_00453_),
    .S(_12100_),
    .Z(_12184_));
 MUX2_X1 _18058_ (.A(_00452_),
    .B(_00454_),
    .S(_12100_),
    .Z(_12185_));
 MUX2_X1 _18059_ (.A(_12184_),
    .B(_12185_),
    .S(_12098_),
    .Z(_12186_));
 MUX2_X1 _18060_ (.A(_00443_),
    .B(_00445_),
    .S(_12100_),
    .Z(_12187_));
 BUF_X4 _18061_ (.A(_11064_),
    .Z(_12188_));
 MUX2_X1 _18062_ (.A(_00444_),
    .B(_00446_),
    .S(_12188_),
    .Z(_12189_));
 MUX2_X1 _18063_ (.A(_12187_),
    .B(_12189_),
    .S(_11804_),
    .Z(_12190_));
 MUX2_X1 _18064_ (.A(_12186_),
    .B(_12190_),
    .S(_12104_),
    .Z(_12191_));
 MUX2_X1 _18065_ (.A(_00455_),
    .B(_00457_),
    .S(_12100_),
    .Z(_12192_));
 MUX2_X1 _18066_ (.A(_00456_),
    .B(_00458_),
    .S(_12188_),
    .Z(_12193_));
 MUX2_X1 _18067_ (.A(_12192_),
    .B(_12193_),
    .S(_11804_),
    .Z(_12194_));
 MUX2_X1 _18068_ (.A(_00447_),
    .B(_00449_),
    .S(_12100_),
    .Z(_12195_));
 MUX2_X1 _18069_ (.A(_00448_),
    .B(_00450_),
    .S(_12188_),
    .Z(_12196_));
 MUX2_X1 _18070_ (.A(_12195_),
    .B(_12196_),
    .S(_11804_),
    .Z(_12197_));
 MUX2_X1 _18071_ (.A(_12194_),
    .B(_12197_),
    .S(_12104_),
    .Z(_12198_));
 MUX2_X1 _18072_ (.A(_12191_),
    .B(_12198_),
    .S(_10987_),
    .Z(_12199_));
 BUF_X4 _18073_ (.A(_11064_),
    .Z(_12200_));
 MUX2_X1 _18074_ (.A(_00439_),
    .B(_00441_),
    .S(_12200_),
    .Z(_12201_));
 MUX2_X1 _18075_ (.A(_00440_),
    .B(_00442_),
    .S(_12200_),
    .Z(_12202_));
 MUX2_X1 _18076_ (.A(_12201_),
    .B(_12202_),
    .S(_10999_),
    .Z(_12203_));
 MUX2_X1 _18077_ (.A(_00431_),
    .B(_00433_),
    .S(_12200_),
    .Z(_12204_));
 MUX2_X1 _18078_ (.A(_00432_),
    .B(_00434_),
    .S(_12200_),
    .Z(_12205_));
 MUX2_X1 _18079_ (.A(_12204_),
    .B(_12205_),
    .S(_10999_),
    .Z(_12206_));
 MUX2_X1 _18080_ (.A(_12203_),
    .B(_12206_),
    .S(_11232_),
    .Z(_12207_));
 NOR2_X1 _18081_ (.A1(_11838_),
    .A2(_12207_),
    .ZN(_12208_));
 NOR2_X1 _18082_ (.A1(_11850_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .ZN(_12209_));
 AOI21_X1 _18083_ (.A(_12209_),
    .B1(_00430_),
    .B2(_11016_),
    .ZN(_12210_));
 AOI221_X1 _18084_ (.A(_11235_),
    .B1(_11620_),
    .B2(_11799_),
    .C1(_12210_),
    .C2(_11269_),
    .ZN(_12211_));
 MUX2_X1 _18085_ (.A(_00435_),
    .B(_00437_),
    .S(_11097_),
    .Z(_12212_));
 MUX2_X1 _18086_ (.A(_00436_),
    .B(_00438_),
    .S(_11097_),
    .Z(_12213_));
 MUX2_X1 _18087_ (.A(_12212_),
    .B(_12213_),
    .S(_11061_),
    .Z(_12214_));
 AOI21_X1 _18088_ (.A(_12211_),
    .B1(_12214_),
    .B2(_11252_),
    .ZN(_12215_));
 AOI21_X1 _18089_ (.A(_12208_),
    .B1(_12215_),
    .B2(_11038_),
    .ZN(_12216_));
 MUX2_X2 _18090_ (.A(_12199_),
    .B(_12216_),
    .S(_10982_),
    .Z(_12217_));
 CLKBUF_X2 _18091_ (.A(\cs_registers_i.pc_id_i[8] ),
    .Z(_12218_));
 CLKBUF_X3 _18092_ (.A(_11111_),
    .Z(_12219_));
 NAND2_X1 _18093_ (.A1(_12218_),
    .A2(_12219_),
    .ZN(_12220_));
 OAI221_X1 _18094_ (.A(_12183_),
    .B1(_12217_),
    .B2(_11278_),
    .C1(_12220_),
    .C2(_10978_),
    .ZN(_12221_));
 CLKBUF_X3 _18095_ (.A(_12221_),
    .Z(_16302_));
 INV_X1 _18096_ (.A(_16302_),
    .ZN(_16306_));
 NAND2_X1 _18097_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(_11221_),
    .ZN(_12222_));
 BUF_X4 _18098_ (.A(_11244_),
    .Z(_12223_));
 MUX2_X1 _18099_ (.A(_00481_),
    .B(_00483_),
    .S(_12223_),
    .Z(_12224_));
 MUX2_X1 _18100_ (.A(_00482_),
    .B(_00484_),
    .S(_12223_),
    .Z(_12225_));
 BUF_X8 _18101_ (.A(_11059_),
    .Z(_12226_));
 MUX2_X1 _18102_ (.A(_12224_),
    .B(_12225_),
    .S(_12226_),
    .Z(_12227_));
 MUX2_X1 _18103_ (.A(_00473_),
    .B(_00475_),
    .S(_12223_),
    .Z(_12228_));
 MUX2_X1 _18104_ (.A(_00474_),
    .B(_00476_),
    .S(_12223_),
    .Z(_12229_));
 MUX2_X1 _18105_ (.A(_12228_),
    .B(_12229_),
    .S(_12226_),
    .Z(_12230_));
 MUX2_X1 _18106_ (.A(_12227_),
    .B(_12230_),
    .S(_10993_),
    .Z(_12231_));
 NOR2_X1 _18107_ (.A1(_11177_),
    .A2(_12231_),
    .ZN(_12232_));
 MUX2_X1 _18108_ (.A(_00485_),
    .B(_00487_),
    .S(_11800_),
    .Z(_12233_));
 MUX2_X1 _18109_ (.A(_00486_),
    .B(_00488_),
    .S(_11800_),
    .Z(_12234_));
 MUX2_X1 _18110_ (.A(_12233_),
    .B(_12234_),
    .S(_11804_),
    .Z(_12235_));
 MUX2_X1 _18111_ (.A(_00477_),
    .B(_00479_),
    .S(_11800_),
    .Z(_12236_));
 MUX2_X1 _18112_ (.A(_00478_),
    .B(_00480_),
    .S(_11207_),
    .Z(_12237_));
 MUX2_X1 _18113_ (.A(_12236_),
    .B(_12237_),
    .S(_11092_),
    .Z(_12238_));
 MUX2_X1 _18114_ (.A(_12235_),
    .B(_12238_),
    .S(_10993_),
    .Z(_12239_));
 NOR2_X1 _18115_ (.A1(_11838_),
    .A2(_12239_),
    .ZN(_12240_));
 NOR3_X4 _18116_ (.A1(_10982_),
    .A2(_12232_),
    .A3(_12240_),
    .ZN(_12241_));
 MUX2_X1 _18117_ (.A(_00465_),
    .B(_00467_),
    .S(_11801_),
    .Z(_12242_));
 NOR2_X1 _18118_ (.A1(_11061_),
    .A2(_12242_),
    .ZN(_12243_));
 MUX2_X1 _18119_ (.A(_00466_),
    .B(_00468_),
    .S(_11850_),
    .Z(_12244_));
 NOR2_X1 _18120_ (.A1(_11795_),
    .A2(_12244_),
    .ZN(_12245_));
 NOR3_X1 _18121_ (.A1(_12117_),
    .A2(_12243_),
    .A3(_12245_),
    .ZN(_12246_));
 NOR2_X1 _18122_ (.A1(_11006_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .ZN(_12247_));
 AOI21_X1 _18123_ (.A(_12247_),
    .B1(_00460_),
    .B2(_11241_),
    .ZN(_12248_));
 AOI221_X2 _18124_ (.A(_11235_),
    .B1(_11675_),
    .B2(_11799_),
    .C1(_12248_),
    .C2(_11042_),
    .ZN(_12249_));
 NOR3_X2 _18125_ (.A1(_11058_),
    .A2(_12246_),
    .A3(_12249_),
    .ZN(_12250_));
 MUX2_X1 _18126_ (.A(_00469_),
    .B(_00471_),
    .S(_11849_),
    .Z(_12251_));
 MUX2_X1 _18127_ (.A(_00470_),
    .B(_00472_),
    .S(_12100_),
    .Z(_12252_));
 MUX2_X1 _18128_ (.A(_12251_),
    .B(_12252_),
    .S(_12098_),
    .Z(_12253_));
 MUX2_X1 _18129_ (.A(_00461_),
    .B(_00463_),
    .S(_12100_),
    .Z(_12254_));
 MUX2_X1 _18130_ (.A(_00462_),
    .B(_00464_),
    .S(_12100_),
    .Z(_12255_));
 MUX2_X1 _18131_ (.A(_12254_),
    .B(_12255_),
    .S(_12098_),
    .Z(_12256_));
 MUX2_X1 _18132_ (.A(_12253_),
    .B(_12256_),
    .S(_12104_),
    .Z(_12257_));
 NOR2_X1 _18133_ (.A1(_11838_),
    .A2(_12257_),
    .ZN(_12258_));
 NOR3_X4 _18134_ (.A1(_11053_),
    .A2(_12250_),
    .A3(_12258_),
    .ZN(_12259_));
 OR2_X2 _18135_ (.A1(_12241_),
    .A2(_12259_),
    .ZN(_12260_));
 BUF_X1 _18136_ (.A(\cs_registers_i.pc_id_i[9] ),
    .Z(_12261_));
 NAND2_X1 _18137_ (.A1(_12261_),
    .A2(_12219_),
    .ZN(_12262_));
 OAI221_X2 _18138_ (.A(_12222_),
    .B1(_12260_),
    .B2(_11818_),
    .C1(_12262_),
    .C2(_10978_),
    .ZN(_16310_));
 INV_X2 _18139_ (.A(_16310_),
    .ZN(_16314_));
 BUF_X2 _18140_ (.A(_15808_),
    .Z(_12263_));
 BUF_X1 _18141_ (.A(_15803_),
    .Z(_12264_));
 NOR3_X1 _18142_ (.A1(_12138_),
    .A2(_15799_),
    .A3(_12264_),
    .ZN(_12265_));
 NOR3_X1 _18143_ (.A1(_15795_),
    .A2(_15799_),
    .A3(_12264_),
    .ZN(_12266_));
 BUF_X4 _18144_ (.A(_15804_),
    .Z(_12267_));
 INV_X1 _18145_ (.A(_12267_),
    .ZN(_12268_));
 INV_X1 _18146_ (.A(_12264_),
    .ZN(_12269_));
 AOI221_X2 _18147_ (.A(_12265_),
    .B1(_12266_),
    .B2(_12155_),
    .C1(_12268_),
    .C2(_12269_),
    .ZN(_12270_));
 XNOR2_X2 _18148_ (.A(_12263_),
    .B(_12270_),
    .ZN(_12271_));
 INV_X4 _18149_ (.A(_12271_),
    .ZN(\alu_adder_result_ex[9] ));
 NAND2_X4 _18150_ (.A1(_12138_),
    .A2(_12140_),
    .ZN(_12272_));
 NOR3_X2 _18151_ (.A1(_12272_),
    .A2(_12171_),
    .A3(_12164_),
    .ZN(_12273_));
 NAND2_X1 _18152_ (.A1(_12267_),
    .A2(_12273_),
    .ZN(_12274_));
 NOR3_X2 _18153_ (.A1(net360),
    .A2(_11918_),
    .A3(_12274_),
    .ZN(_12275_));
 BUF_X4 _18154_ (.A(_12165_),
    .Z(_12276_));
 AOI21_X2 _18155_ (.A(_15799_),
    .B1(_15795_),
    .B2(_12138_),
    .ZN(_12277_));
 NOR2_X2 _18156_ (.A1(_12168_),
    .A2(_12164_),
    .ZN(_12278_));
 AOI211_X2 _18157_ (.A(_12141_),
    .B(_12278_),
    .C1(_12161_),
    .C2(_12142_),
    .ZN(_12279_));
 OAI21_X2 _18158_ (.A(_12277_),
    .B1(_12279_),
    .B2(_12272_),
    .ZN(_12280_));
 OR3_X1 _18159_ (.A1(_12267_),
    .A2(_12276_),
    .A3(_12280_),
    .ZN(_12281_));
 AOI21_X2 _18160_ (.A(_12281_),
    .B1(_12177_),
    .B2(_12176_),
    .ZN(_12282_));
 NAND2_X1 _18161_ (.A1(_12267_),
    .A2(_12280_),
    .ZN(_12283_));
 OR2_X1 _18162_ (.A1(_12267_),
    .A2(_12273_),
    .ZN(_12284_));
 OAI221_X2 _18163_ (.A(_12283_),
    .B1(_12284_),
    .B2(_12280_),
    .C1(_11865_),
    .C2(_12274_),
    .ZN(_12285_));
 OR3_X2 _18164_ (.A1(_12275_),
    .A2(_12282_),
    .A3(_12285_),
    .ZN(_12286_));
 INV_X4 _18165_ (.A(_12286_),
    .ZN(\alu_adder_result_ex[8] ));
 NAND2_X1 _18166_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(_11221_),
    .ZN(_12287_));
 MUX2_X1 _18167_ (.A(_00499_),
    .B(_00501_),
    .S(_12188_),
    .Z(_12288_));
 MUX2_X1 _18168_ (.A(_00500_),
    .B(_00502_),
    .S(_12188_),
    .Z(_12289_));
 MUX2_X1 _18169_ (.A(_12288_),
    .B(_12289_),
    .S(_11804_),
    .Z(_12290_));
 MUX2_X1 _18170_ (.A(_00491_),
    .B(_00493_),
    .S(_12188_),
    .Z(_12291_));
 MUX2_X1 _18171_ (.A(_00492_),
    .B(_00494_),
    .S(_12188_),
    .Z(_12292_));
 MUX2_X1 _18172_ (.A(_12291_),
    .B(_12292_),
    .S(_11804_),
    .Z(_12293_));
 MUX2_X1 _18173_ (.A(_12290_),
    .B(_12293_),
    .S(_12104_),
    .Z(_12294_));
 NOR2_X1 _18174_ (.A1(_11838_),
    .A2(_12294_),
    .ZN(_12295_));
 NOR2_X1 _18175_ (.A1(_11801_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .ZN(_12296_));
 BUF_X4 _18176_ (.A(_11015_),
    .Z(_12297_));
 AOI21_X1 _18177_ (.A(_12296_),
    .B1(_00490_),
    .B2(_12297_),
    .ZN(_12298_));
 AOI221_X2 _18178_ (.A(_11235_),
    .B1(_11696_),
    .B2(_11799_),
    .C1(_12298_),
    .C2(_11000_),
    .ZN(_12299_));
 MUX2_X1 _18179_ (.A(_00495_),
    .B(_00497_),
    .S(_11016_),
    .Z(_12300_));
 MUX2_X1 _18180_ (.A(_00496_),
    .B(_00498_),
    .S(_11016_),
    .Z(_12301_));
 MUX2_X1 _18181_ (.A(_12300_),
    .B(_12301_),
    .S(_11061_),
    .Z(_12302_));
 AOI21_X2 _18182_ (.A(_12299_),
    .B1(_12302_),
    .B2(_11252_),
    .ZN(_12303_));
 AOI21_X4 _18183_ (.A(_12295_),
    .B1(_12303_),
    .B2(_11038_),
    .ZN(_12304_));
 MUX2_X1 _18184_ (.A(_00517_),
    .B(_00518_),
    .S(_11256_),
    .Z(_12305_));
 AOI21_X1 _18185_ (.A(_11036_),
    .B1(_12305_),
    .B2(_11008_),
    .ZN(_12306_));
 MUX2_X1 _18186_ (.A(_00513_),
    .B(_00514_),
    .S(_11092_),
    .Z(_12307_));
 AOI21_X1 _18187_ (.A(_11057_),
    .B1(_12307_),
    .B2(_11068_),
    .ZN(_12308_));
 OAI21_X1 _18188_ (.A(_11069_),
    .B1(_12306_),
    .B2(_12308_),
    .ZN(_12309_));
 MUX2_X1 _18189_ (.A(_00511_),
    .B(_00512_),
    .S(_11042_),
    .Z(_12310_));
 INV_X1 _18190_ (.A(_12310_),
    .ZN(_12311_));
 MUX2_X1 _18191_ (.A(_00515_),
    .B(_00516_),
    .S(_11060_),
    .Z(_12312_));
 INV_X1 _18192_ (.A(_12312_),
    .ZN(_12313_));
 AOI22_X1 _18193_ (.A1(_12308_),
    .A2(_12311_),
    .B1(_12313_),
    .B2(_12306_),
    .ZN(_12314_));
 NAND3_X1 _18194_ (.A1(_11252_),
    .A2(_12309_),
    .A3(_12314_),
    .ZN(_12315_));
 MUX2_X1 _18195_ (.A(_00507_),
    .B(_00509_),
    .S(_11801_),
    .Z(_12316_));
 MUX2_X1 _18196_ (.A(_00508_),
    .B(_00510_),
    .S(_11801_),
    .Z(_12317_));
 MUX2_X1 _18197_ (.A(_12316_),
    .B(_12317_),
    .S(_11805_),
    .Z(_12318_));
 MUX2_X1 _18198_ (.A(_00505_),
    .B(_00506_),
    .S(_11269_),
    .Z(_12319_));
 MUX2_X1 _18199_ (.A(_00503_),
    .B(_00504_),
    .S(_11042_),
    .Z(_12320_));
 AOI222_X2 _18200_ (.A1(_11085_),
    .A2(_12318_),
    .B1(_12319_),
    .B2(_11100_),
    .C1(_12320_),
    .C2(_11091_),
    .ZN(_12321_));
 NAND2_X1 _18201_ (.A1(_12315_),
    .A2(_12321_),
    .ZN(_12322_));
 MUX2_X2 _18202_ (.A(_12304_),
    .B(_12322_),
    .S(_11931_),
    .Z(_12323_));
 NAND2_X1 _18203_ (.A1(\cs_registers_i.pc_id_i[10] ),
    .A2(_12219_),
    .ZN(_12324_));
 OAI221_X2 _18204_ (.A(_12287_),
    .B1(_12323_),
    .B2(_11818_),
    .C1(_12324_),
    .C2(_10978_),
    .ZN(_16317_));
 INV_X4 _18205_ (.A(_16317_),
    .ZN(_16321_));
 INV_X1 _18206_ (.A(_15816_),
    .ZN(_12325_));
 INV_X1 _18207_ (.A(_15807_),
    .ZN(_12326_));
 AOI21_X1 _18208_ (.A(_12264_),
    .B1(_15799_),
    .B2(_12267_),
    .ZN(_12327_));
 INV_X1 _18209_ (.A(_12263_),
    .ZN(_12328_));
 OAI21_X1 _18210_ (.A(_12326_),
    .B1(_12327_),
    .B2(_12328_),
    .ZN(_12329_));
 AOI21_X2 _18211_ (.A(_15811_),
    .B1(_12329_),
    .B2(_15812_),
    .ZN(_12330_));
 OR2_X1 _18212_ (.A1(_15812_),
    .A2(_15811_),
    .ZN(_12331_));
 NAND4_X1 _18213_ (.A1(_12138_),
    .A2(_12267_),
    .A3(_12263_),
    .A4(_12331_),
    .ZN(_12332_));
 OAI21_X2 _18214_ (.A(_12330_),
    .B1(_12332_),
    .B2(_12156_),
    .ZN(_12333_));
 XNOR2_X2 _18215_ (.A(_12333_),
    .B(_12325_),
    .ZN(\alu_adder_result_ex[11] ));
 OAI21_X1 _18216_ (.A(_12269_),
    .B1(_12277_),
    .B2(_12268_),
    .ZN(_12334_));
 AOI21_X1 _18217_ (.A(_15807_),
    .B1(_12334_),
    .B2(_12263_),
    .ZN(_12335_));
 NAND2_X1 _18218_ (.A1(_12267_),
    .A2(_12263_),
    .ZN(_12336_));
 NOR2_X1 _18219_ (.A1(_12272_),
    .A2(_12336_),
    .ZN(_12337_));
 OAI21_X2 _18220_ (.A(_12337_),
    .B1(_12169_),
    .B2(_12163_),
    .ZN(_12338_));
 NAND2_X2 _18221_ (.A1(_12335_),
    .A2(_12338_),
    .ZN(_12339_));
 NAND2_X2 _18222_ (.A1(_12178_),
    .A2(_12337_),
    .ZN(_12340_));
 NOR3_X4 _18223_ (.A1(_11896_),
    .A2(_11917_),
    .A3(_12340_),
    .ZN(_12341_));
 AOI21_X4 _18224_ (.A(_12339_),
    .B1(_12341_),
    .B2(_12176_),
    .ZN(_12342_));
 XNOR2_X2 _18225_ (.A(net349),
    .B(_12342_),
    .ZN(\alu_adder_result_ex[10] ));
 BUF_X8 _18226_ (.A(_11168_),
    .Z(_12343_));
 NAND2_X1 _18227_ (.A1(_10834_),
    .A2(_11485_),
    .ZN(_12344_));
 NAND4_X1 _18228_ (.A1(_10878_),
    .A2(_10774_),
    .A3(_10836_),
    .A4(_12344_),
    .ZN(_12345_));
 NAND4_X1 _18229_ (.A1(_10774_),
    .A2(_10855_),
    .A3(_11486_),
    .A4(_11730_),
    .ZN(_12346_));
 AND2_X1 _18230_ (.A1(_12345_),
    .A2(_12346_),
    .ZN(_12347_));
 BUF_X4 _18231_ (.A(_12347_),
    .Z(_12348_));
 NOR4_X2 _18232_ (.A1(_10809_),
    .A2(_10818_),
    .A3(_10802_),
    .A4(_10857_),
    .ZN(_12349_));
 MUX2_X1 _18233_ (.A(_11725_),
    .B(_12349_),
    .S(_10836_),
    .Z(_12350_));
 CLKBUF_X3 _18234_ (.A(_12350_),
    .Z(_12351_));
 NAND2_X1 _18235_ (.A1(_10828_),
    .A2(_12351_),
    .ZN(_12352_));
 AOI21_X2 _18236_ (.A(_12343_),
    .B1(_12348_),
    .B2(_12352_),
    .ZN(_12353_));
 BUF_X8 _18237_ (.A(_11134_),
    .Z(_12354_));
 BUF_X8 _18238_ (.A(_12354_),
    .Z(_12355_));
 BUF_X4 _18239_ (.A(_10731_),
    .Z(_12356_));
 BUF_X4 _18240_ (.A(_10719_),
    .Z(_12357_));
 BUF_X4 _18241_ (.A(_12357_),
    .Z(_12358_));
 BUF_X4 _18242_ (.A(_10711_),
    .Z(_12359_));
 BUF_X4 _18243_ (.A(_12359_),
    .Z(_12360_));
 BUF_X4 _18244_ (.A(_12360_),
    .Z(_12361_));
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 BUF_X8 _18246_ (.A(net341),
    .Z(_12363_));
 BUF_X8 _18247_ (.A(_12363_),
    .Z(_12364_));
 MUX2_X1 _18248_ (.A(_00224_),
    .B(_00226_),
    .S(_12364_),
    .Z(_12365_));
 NOR2_X1 _18249_ (.A1(_12361_),
    .A2(_12365_),
    .ZN(_12366_));
 BUF_X4 _18250_ (.A(_11130_),
    .Z(_12367_));
 BUF_X4 _18251_ (.A(_12367_),
    .Z(_12368_));
 MUX2_X1 _18252_ (.A(_00225_),
    .B(_00227_),
    .S(_12364_),
    .Z(_12369_));
 NOR2_X1 _18253_ (.A1(_12368_),
    .A2(_12369_),
    .ZN(_12370_));
 NOR3_X1 _18254_ (.A1(_12358_),
    .A2(_12366_),
    .A3(_12370_),
    .ZN(_12371_));
 BUF_X4 _18255_ (.A(_10758_),
    .Z(_12372_));
 BUF_X4 _18256_ (.A(_11137_),
    .Z(_12373_));
 BUF_X4 _18257_ (.A(_12373_),
    .Z(_12374_));
 NOR2_X1 _18258_ (.A1(_12364_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .ZN(_12375_));
 BUF_X32 _18259_ (.A(_10750_),
    .Z(_12376_));
 BUF_X4 _18260_ (.A(_12376_),
    .Z(_12377_));
 BUF_X4 _18261_ (.A(_12377_),
    .Z(_12378_));
 AOI21_X1 _18262_ (.A(_12375_),
    .B1(_00219_),
    .B2(_12378_),
    .ZN(_12379_));
 BUF_X4 _18263_ (.A(_12359_),
    .Z(_12380_));
 BUF_X4 _18264_ (.A(_12380_),
    .Z(_12381_));
 AOI221_X2 _18265_ (.A(_12372_),
    .B1(_11236_),
    .B2(_12374_),
    .C1(_12379_),
    .C2(_12381_),
    .ZN(_12382_));
 NOR3_X2 _18266_ (.A1(_12356_),
    .A2(_12371_),
    .A3(_12382_),
    .ZN(_12383_));
 BUF_X4 _18267_ (.A(_10736_),
    .Z(_12384_));
 BUF_X4 _18268_ (.A(net341),
    .Z(_12385_));
 MUX2_X1 _18269_ (.A(_00228_),
    .B(_00230_),
    .S(_12385_),
    .Z(_12386_));
 MUX2_X1 _18270_ (.A(_00229_),
    .B(_00231_),
    .S(_12385_),
    .Z(_12387_));
 BUF_X4 _18271_ (.A(_12359_),
    .Z(_12388_));
 MUX2_X1 _18272_ (.A(_12386_),
    .B(_12387_),
    .S(_12388_),
    .Z(_12389_));
 MUX2_X1 _18273_ (.A(_00220_),
    .B(_00222_),
    .S(_12385_),
    .Z(_12390_));
 MUX2_X1 _18274_ (.A(_00221_),
    .B(_00223_),
    .S(_12385_),
    .Z(_12391_));
 BUF_X4 _18275_ (.A(_12359_),
    .Z(_12392_));
 MUX2_X1 _18276_ (.A(_12390_),
    .B(_12391_),
    .S(_12392_),
    .Z(_12393_));
 BUF_X4 _18277_ (.A(_10719_),
    .Z(_12394_));
 MUX2_X1 _18278_ (.A(_12389_),
    .B(_12393_),
    .S(_12394_),
    .Z(_12395_));
 NOR2_X1 _18279_ (.A1(_12384_),
    .A2(_12395_),
    .ZN(_12396_));
 NOR3_X2 _18280_ (.A1(_12355_),
    .A2(_12383_),
    .A3(_12396_),
    .ZN(_12397_));
 BUF_X8 _18281_ (.A(_12376_),
    .Z(_12398_));
 MUX2_X1 _18282_ (.A(_00240_),
    .B(_00242_),
    .S(_12398_),
    .Z(_12399_));
 BUF_X8 _18283_ (.A(_10750_),
    .Z(_12400_));
 BUF_X8 _18284_ (.A(_12400_),
    .Z(_12401_));
 MUX2_X1 _18285_ (.A(_00241_),
    .B(_00243_),
    .S(_12401_),
    .Z(_12402_));
 BUF_X4 _18286_ (.A(_12359_),
    .Z(_12403_));
 MUX2_X1 _18287_ (.A(_12399_),
    .B(_12402_),
    .S(_12403_),
    .Z(_12404_));
 MUX2_X1 _18288_ (.A(_00232_),
    .B(_00234_),
    .S(_12398_),
    .Z(_12405_));
 MUX2_X1 _18289_ (.A(_00233_),
    .B(_00235_),
    .S(_12401_),
    .Z(_12406_));
 MUX2_X1 _18290_ (.A(_12405_),
    .B(_12406_),
    .S(_12403_),
    .Z(_12407_));
 BUF_X4 _18291_ (.A(_10719_),
    .Z(_12408_));
 BUF_X4 _18292_ (.A(_12408_),
    .Z(_12409_));
 MUX2_X1 _18293_ (.A(_12404_),
    .B(_12407_),
    .S(_12409_),
    .Z(_12410_));
 MUX2_X1 _18294_ (.A(_00244_),
    .B(_00246_),
    .S(_12401_),
    .Z(_12411_));
 MUX2_X1 _18295_ (.A(_00245_),
    .B(_00247_),
    .S(_12401_),
    .Z(_12412_));
 MUX2_X1 _18296_ (.A(_12411_),
    .B(_12412_),
    .S(_12403_),
    .Z(_12413_));
 MUX2_X1 _18297_ (.A(_00236_),
    .B(_00238_),
    .S(_12401_),
    .Z(_12414_));
 MUX2_X1 _18298_ (.A(_00237_),
    .B(_00239_),
    .S(_12401_),
    .Z(_12415_));
 MUX2_X1 _18299_ (.A(_12414_),
    .B(_12415_),
    .S(_12403_),
    .Z(_12416_));
 MUX2_X1 _18300_ (.A(_12413_),
    .B(_12416_),
    .S(_12409_),
    .Z(_12417_));
 MUX2_X1 _18301_ (.A(_12410_),
    .B(_12417_),
    .S(_12356_),
    .Z(_12418_));
 BUF_X8 _18302_ (.A(_12355_),
    .Z(_12419_));
 AOI21_X4 _18303_ (.A(_12397_),
    .B1(_12419_),
    .B2(_12418_),
    .ZN(_12420_));
 AOI21_X4 _18304_ (.A(_12353_),
    .B1(_12343_),
    .B2(_12420_),
    .ZN(_16338_));
 INV_X1 _18305_ (.A(_16338_),
    .ZN(_16334_));
 NAND2_X1 _18306_ (.A1(_10882_),
    .A2(_12351_),
    .ZN(_12421_));
 AOI21_X1 _18307_ (.A(_12343_),
    .B1(_12348_),
    .B2(_12421_),
    .ZN(_12422_));
 BUF_X4 _18308_ (.A(_10731_),
    .Z(_12423_));
 BUF_X8 _18309_ (.A(_12423_),
    .Z(_12424_));
 BUF_X4 _18310_ (.A(_12357_),
    .Z(_12425_));
 BUF_X4 _18311_ (.A(_12403_),
    .Z(_12426_));
 MUX2_X1 _18312_ (.A(_00575_),
    .B(_00577_),
    .S(_12378_),
    .Z(_12427_));
 NOR2_X1 _18313_ (.A1(_12426_),
    .A2(_12427_),
    .ZN(_12428_));
 MUX2_X1 _18314_ (.A(_00576_),
    .B(_00578_),
    .S(_12378_),
    .Z(_12429_));
 NOR2_X1 _18315_ (.A1(_12368_),
    .A2(_12429_),
    .ZN(_12430_));
 NOR3_X1 _18316_ (.A1(_12425_),
    .A2(_12428_),
    .A3(_12430_),
    .ZN(_12431_));
 BUF_X8 _18317_ (.A(_10758_),
    .Z(_12432_));
 INV_X1 _18318_ (.A(_00569_),
    .ZN(_12433_));
 BUF_X16 _18319_ (.A(_12376_),
    .Z(_12434_));
 BUF_X4 _18320_ (.A(_12434_),
    .Z(_12435_));
 NOR2_X1 _18321_ (.A1(_12435_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .ZN(_12436_));
 BUF_X4 _18322_ (.A(_12400_),
    .Z(_12437_));
 BUF_X4 _18323_ (.A(_12437_),
    .Z(_12438_));
 AOI21_X1 _18324_ (.A(_12436_),
    .B1(_00570_),
    .B2(_12438_),
    .ZN(_12439_));
 BUF_X4 _18325_ (.A(_12388_),
    .Z(_12440_));
 AOI221_X2 _18326_ (.A(_12432_),
    .B1(_12433_),
    .B2(_12374_),
    .C1(_12439_),
    .C2(_12440_),
    .ZN(_12441_));
 NOR3_X1 _18327_ (.A1(_12424_),
    .A2(_12431_),
    .A3(_12441_),
    .ZN(_12442_));
 MUX2_X1 _18328_ (.A(_00579_),
    .B(_00581_),
    .S(_12377_),
    .Z(_12443_));
 MUX2_X1 _18329_ (.A(_00580_),
    .B(_00582_),
    .S(_12398_),
    .Z(_12444_));
 BUF_X4 _18330_ (.A(_12359_),
    .Z(_12445_));
 MUX2_X1 _18331_ (.A(_12443_),
    .B(_12444_),
    .S(_12445_),
    .Z(_12446_));
 MUX2_X1 _18332_ (.A(_00571_),
    .B(_00573_),
    .S(_12398_),
    .Z(_12447_));
 MUX2_X1 _18333_ (.A(_00572_),
    .B(_00574_),
    .S(_12398_),
    .Z(_12448_));
 MUX2_X1 _18334_ (.A(_12447_),
    .B(_12448_),
    .S(_12445_),
    .Z(_12449_));
 BUF_X4 _18335_ (.A(_12408_),
    .Z(_12450_));
 MUX2_X1 _18336_ (.A(_12446_),
    .B(_12449_),
    .S(_12450_),
    .Z(_12451_));
 NOR2_X1 _18337_ (.A1(_12384_),
    .A2(_12451_),
    .ZN(_12452_));
 NOR3_X2 _18338_ (.A1(_12355_),
    .A2(_12442_),
    .A3(_12452_),
    .ZN(_12453_));
 BUF_X16 _18339_ (.A(_10750_),
    .Z(_12454_));
 BUF_X8 _18340_ (.A(_12454_),
    .Z(_12455_));
 MUX2_X1 _18341_ (.A(_00591_),
    .B(_00593_),
    .S(_12455_),
    .Z(_12456_));
 BUF_X4 _18342_ (.A(_12454_),
    .Z(_12457_));
 MUX2_X1 _18343_ (.A(_00592_),
    .B(_00594_),
    .S(_12457_),
    .Z(_12458_));
 BUF_X4 _18344_ (.A(_12380_),
    .Z(_12459_));
 MUX2_X1 _18345_ (.A(_12456_),
    .B(_12458_),
    .S(_12459_),
    .Z(_12460_));
 MUX2_X1 _18346_ (.A(_00583_),
    .B(_00585_),
    .S(_12457_),
    .Z(_12461_));
 MUX2_X1 _18347_ (.A(_00584_),
    .B(_00586_),
    .S(_12457_),
    .Z(_12462_));
 MUX2_X1 _18348_ (.A(_12461_),
    .B(_12462_),
    .S(_12459_),
    .Z(_12463_));
 MUX2_X1 _18349_ (.A(_12460_),
    .B(_12463_),
    .S(_12425_),
    .Z(_12464_));
 MUX2_X1 _18350_ (.A(_00595_),
    .B(_00597_),
    .S(_12457_),
    .Z(_12465_));
 MUX2_X1 _18351_ (.A(_00596_),
    .B(_00598_),
    .S(_12457_),
    .Z(_12466_));
 MUX2_X1 _18352_ (.A(_12465_),
    .B(_12466_),
    .S(_12459_),
    .Z(_12467_));
 MUX2_X1 _18353_ (.A(_00587_),
    .B(_00589_),
    .S(_12457_),
    .Z(_12468_));
 MUX2_X1 _18354_ (.A(_00588_),
    .B(_00590_),
    .S(_12364_),
    .Z(_12469_));
 MUX2_X1 _18355_ (.A(_12468_),
    .B(_12469_),
    .S(_12440_),
    .Z(_12470_));
 MUX2_X1 _18356_ (.A(_12467_),
    .B(_12470_),
    .S(_12425_),
    .Z(_12471_));
 MUX2_X1 _18357_ (.A(_12464_),
    .B(_12471_),
    .S(_12424_),
    .Z(_12472_));
 AOI21_X4 _18358_ (.A(_12453_),
    .B1(_12419_),
    .B2(_12472_),
    .ZN(_12473_));
 AOI21_X2 _18359_ (.A(_12422_),
    .B1(_12473_),
    .B2(_12343_),
    .ZN(_16341_));
 INV_X1 _18360_ (.A(_16341_),
    .ZN(_16345_));
 NAND2_X1 _18361_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(_11221_),
    .ZN(_12474_));
 MUX2_X1 _18362_ (.A(_00579_),
    .B(_00581_),
    .S(_11207_),
    .Z(_12475_));
 MUX2_X1 _18363_ (.A(_00580_),
    .B(_00582_),
    .S(_12223_),
    .Z(_12476_));
 MUX2_X1 _18364_ (.A(_12475_),
    .B(_12476_),
    .S(_11092_),
    .Z(_12477_));
 MUX2_X1 _18365_ (.A(_00571_),
    .B(_00573_),
    .S(_12223_),
    .Z(_12478_));
 MUX2_X1 _18366_ (.A(_00572_),
    .B(_00574_),
    .S(_12223_),
    .Z(_12479_));
 MUX2_X1 _18367_ (.A(_12478_),
    .B(_12479_),
    .S(_12226_),
    .Z(_12480_));
 MUX2_X1 _18368_ (.A(_12477_),
    .B(_12480_),
    .S(_10993_),
    .Z(_12481_));
 NOR2_X1 _18369_ (.A1(_11838_),
    .A2(_12481_),
    .ZN(_12482_));
 NOR2_X1 _18370_ (.A1(_11208_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .ZN(_12483_));
 AOI21_X1 _18371_ (.A(_12483_),
    .B1(_00570_),
    .B2(_11007_),
    .ZN(_12484_));
 AOI221_X1 _18372_ (.A(_11022_),
    .B1(_12433_),
    .B2(_11032_),
    .C1(_12484_),
    .C2(_11805_),
    .ZN(_12485_));
 MUX2_X1 _18373_ (.A(_00575_),
    .B(_00577_),
    .S(_12297_),
    .Z(_12486_));
 MUX2_X1 _18374_ (.A(_00576_),
    .B(_00578_),
    .S(_12297_),
    .Z(_12487_));
 MUX2_X1 _18375_ (.A(_12486_),
    .B(_12487_),
    .S(_11043_),
    .Z(_12488_));
 AOI21_X1 _18376_ (.A(_12485_),
    .B1(_12488_),
    .B2(_11252_),
    .ZN(_12489_));
 AOI21_X2 _18377_ (.A(_12482_),
    .B1(_12489_),
    .B2(_11038_),
    .ZN(_12490_));
 MUX2_X1 _18378_ (.A(_00597_),
    .B(_00598_),
    .S(_12098_),
    .Z(_12491_));
 AOI21_X1 _18379_ (.A(_11036_),
    .B1(_12491_),
    .B2(_11188_),
    .ZN(_12492_));
 MUX2_X1 _18380_ (.A(_00593_),
    .B(_00594_),
    .S(_11074_),
    .Z(_12493_));
 AOI21_X1 _18381_ (.A(_11057_),
    .B1(_12493_),
    .B2(_11068_),
    .ZN(_12494_));
 OAI21_X1 _18382_ (.A(_11069_),
    .B1(_12492_),
    .B2(_12494_),
    .ZN(_12495_));
 MUX2_X1 _18383_ (.A(_00591_),
    .B(_00592_),
    .S(_11042_),
    .Z(_12496_));
 INV_X1 _18384_ (.A(_12496_),
    .ZN(_12497_));
 MUX2_X1 _18385_ (.A(_00595_),
    .B(_00596_),
    .S(_11042_),
    .Z(_12498_));
 INV_X1 _18386_ (.A(_12498_),
    .ZN(_12499_));
 AOI22_X1 _18387_ (.A1(_12494_),
    .A2(_12497_),
    .B1(_12499_),
    .B2(_12492_),
    .ZN(_12500_));
 NAND3_X1 _18388_ (.A1(_11252_),
    .A2(_12495_),
    .A3(_12500_),
    .ZN(_12501_));
 BUF_X4 _18389_ (.A(_11244_),
    .Z(_12502_));
 BUF_X4 _18390_ (.A(_12502_),
    .Z(_12503_));
 MUX2_X1 _18391_ (.A(_00587_),
    .B(_00589_),
    .S(_12503_),
    .Z(_12504_));
 MUX2_X1 _18392_ (.A(_00588_),
    .B(_00590_),
    .S(_12503_),
    .Z(_12505_));
 MUX2_X1 _18393_ (.A(_12504_),
    .B(_12505_),
    .S(_11093_),
    .Z(_12506_));
 MUX2_X1 _18394_ (.A(_00583_),
    .B(_00584_),
    .S(_11000_),
    .Z(_12507_));
 MUX2_X1 _18395_ (.A(_00585_),
    .B(_00586_),
    .S(_11027_),
    .Z(_12508_));
 AOI222_X2 _18396_ (.A1(_11085_),
    .A2(_12506_),
    .B1(_12507_),
    .B2(_11091_),
    .C1(_12508_),
    .C2(_11100_),
    .ZN(_12509_));
 NAND2_X1 _18397_ (.A1(_12501_),
    .A2(_12509_),
    .ZN(_12510_));
 MUX2_X2 _18398_ (.A(_12490_),
    .B(_12510_),
    .S(_11931_),
    .Z(_12511_));
 BUF_X2 _18399_ (.A(\cs_registers_i.pc_id_i[13] ),
    .Z(_12512_));
 NAND2_X1 _18400_ (.A1(_12512_),
    .A2(_12219_),
    .ZN(_12513_));
 OAI221_X1 _18401_ (.A(_12474_),
    .B1(_12511_),
    .B2(_11818_),
    .C1(_12513_),
    .C2(_11115_),
    .ZN(_12514_));
 CLKBUF_X3 _18402_ (.A(_12514_),
    .Z(_16346_));
 INV_X2 _18403_ (.A(_16346_),
    .ZN(_16342_));
 BUF_X2 _18404_ (.A(_15824_),
    .Z(_12515_));
 INV_X4 _18405_ (.A(_12272_),
    .ZN(_12516_));
 AOI22_X4 _18406_ (.A1(_12138_),
    .A2(_15795_),
    .B1(_12516_),
    .B2(_12141_),
    .ZN(_12517_));
 NAND2_X2 _18407_ (.A1(_12145_),
    .A2(_12516_),
    .ZN(_12518_));
 AOI21_X4 _18408_ (.A(_12146_),
    .B1(_12153_),
    .B2(_12148_),
    .ZN(_12519_));
 OAI21_X4 _18409_ (.A(_12517_),
    .B1(_12519_),
    .B2(_12518_),
    .ZN(_12520_));
 BUF_X2 _18410_ (.A(_15820_),
    .Z(_12521_));
 INV_X2 _18411_ (.A(_12521_),
    .ZN(_12522_));
 NAND2_X2 _18412_ (.A1(_15812_),
    .A2(_15816_),
    .ZN(_12523_));
 NOR3_X1 _18413_ (.A1(_12522_),
    .A2(_12336_),
    .A3(_12523_),
    .ZN(_12524_));
 INV_X1 _18414_ (.A(_15815_),
    .ZN(_12525_));
 OAI21_X2 _18415_ (.A(_12525_),
    .B1(_12330_),
    .B2(_12325_),
    .ZN(_12526_));
 AOI221_X2 _18416_ (.A(_15819_),
    .B1(_12520_),
    .B2(_12524_),
    .C1(_12526_),
    .C2(_12521_),
    .ZN(_12527_));
 XNOR2_X2 _18417_ (.A(_12515_),
    .B(net275),
    .ZN(\alu_adder_result_ex[13] ));
 AOI21_X1 _18418_ (.A(_15815_),
    .B1(_15811_),
    .B2(_15816_),
    .ZN(_12528_));
 INV_X1 _18419_ (.A(_12523_),
    .ZN(_12529_));
 OAI21_X1 _18420_ (.A(_12529_),
    .B1(_15807_),
    .B2(_12263_),
    .ZN(_12530_));
 INV_X1 _18421_ (.A(_12528_),
    .ZN(_12531_));
 NOR3_X1 _18422_ (.A1(_12264_),
    .A2(_15807_),
    .A3(_12531_),
    .ZN(_12532_));
 AOI22_X1 _18423_ (.A1(_12528_),
    .A2(_12530_),
    .B1(_12532_),
    .B2(_12283_),
    .ZN(_12533_));
 NAND4_X2 _18424_ (.A1(_12267_),
    .A2(_12263_),
    .A3(_12273_),
    .A4(_12529_),
    .ZN(_12534_));
 NOR2_X1 _18425_ (.A1(_11864_),
    .A2(_12534_),
    .ZN(_12535_));
 OR2_X1 _18426_ (.A1(_12533_),
    .A2(_12535_),
    .ZN(_12536_));
 NOR3_X2 _18427_ (.A1(_11896_),
    .A2(_11917_),
    .A3(_12534_),
    .ZN(_12537_));
 AOI21_X4 _18428_ (.A(_12536_),
    .B1(_12537_),
    .B2(_12176_),
    .ZN(_12538_));
 XNOR2_X2 _18429_ (.A(_12521_),
    .B(_12538_),
    .ZN(\alu_adder_result_ex[12] ));
 NAND2_X1 _18430_ (.A1(_10924_),
    .A2(_12351_),
    .ZN(_12539_));
 AOI21_X1 _18431_ (.A(_11168_),
    .B1(_12348_),
    .B2(_12539_),
    .ZN(_12540_));
 MUX2_X1 _18432_ (.A(_00606_),
    .B(_00608_),
    .S(_12378_),
    .Z(_12541_));
 NOR2_X1 _18433_ (.A1(_12426_),
    .A2(_12541_),
    .ZN(_12542_));
 MUX2_X1 _18434_ (.A(_00607_),
    .B(_00609_),
    .S(_12435_),
    .Z(_12543_));
 NOR2_X1 _18435_ (.A1(_12368_),
    .A2(_12543_),
    .ZN(_12544_));
 NOR3_X1 _18436_ (.A1(_12425_),
    .A2(_12542_),
    .A3(_12544_),
    .ZN(_12545_));
 INV_X1 _18437_ (.A(_00600_),
    .ZN(_12546_));
 BUF_X4 _18438_ (.A(_12434_),
    .Z(_12547_));
 NOR2_X1 _18439_ (.A1(_12547_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .ZN(_12548_));
 AOI21_X1 _18440_ (.A(_12548_),
    .B1(_00601_),
    .B2(_12438_),
    .ZN(_12549_));
 AOI221_X2 _18441_ (.A(_12432_),
    .B1(_12546_),
    .B2(_12374_),
    .C1(_12549_),
    .C2(_12440_),
    .ZN(_12550_));
 NOR3_X1 _18442_ (.A1(_12356_),
    .A2(_12545_),
    .A3(_12550_),
    .ZN(_12551_));
 BUF_X4 _18443_ (.A(_12376_),
    .Z(_12552_));
 MUX2_X1 _18444_ (.A(_00610_),
    .B(_00612_),
    .S(_12552_),
    .Z(_12553_));
 MUX2_X1 _18445_ (.A(_00611_),
    .B(_00613_),
    .S(_12377_),
    .Z(_12554_));
 BUF_X4 _18446_ (.A(_12359_),
    .Z(_12555_));
 MUX2_X1 _18447_ (.A(_12553_),
    .B(_12554_),
    .S(_12555_),
    .Z(_12556_));
 MUX2_X1 _18448_ (.A(_00602_),
    .B(_00604_),
    .S(_12377_),
    .Z(_12557_));
 MUX2_X1 _18449_ (.A(_00603_),
    .B(_00605_),
    .S(_12377_),
    .Z(_12558_));
 MUX2_X1 _18450_ (.A(_12557_),
    .B(_12558_),
    .S(_12555_),
    .Z(_12559_));
 MUX2_X1 _18451_ (.A(_12556_),
    .B(_12559_),
    .S(_12450_),
    .Z(_12560_));
 NOR2_X1 _18452_ (.A1(_12384_),
    .A2(_12560_),
    .ZN(_12561_));
 NOR3_X2 _18453_ (.A1(_12355_),
    .A2(_12551_),
    .A3(_12561_),
    .ZN(_12562_));
 BUF_X32 _18454_ (.A(net341),
    .Z(_12563_));
 BUF_X8 _18455_ (.A(_12563_),
    .Z(_12564_));
 MUX2_X1 _18456_ (.A(_00622_),
    .B(_00624_),
    .S(_12564_),
    .Z(_12565_));
 MUX2_X1 _18457_ (.A(_00623_),
    .B(_00625_),
    .S(_12564_),
    .Z(_12566_));
 MUX2_X1 _18458_ (.A(_12565_),
    .B(_12566_),
    .S(_12381_),
    .Z(_12567_));
 MUX2_X1 _18459_ (.A(_00614_),
    .B(_00616_),
    .S(_12564_),
    .Z(_12568_));
 MUX2_X1 _18460_ (.A(_00615_),
    .B(_00617_),
    .S(_12455_),
    .Z(_12569_));
 MUX2_X1 _18461_ (.A(_12568_),
    .B(_12569_),
    .S(_12381_),
    .Z(_12570_));
 MUX2_X1 _18462_ (.A(_12567_),
    .B(_12570_),
    .S(_12358_),
    .Z(_12571_));
 MUX2_X1 _18463_ (.A(_00626_),
    .B(_00628_),
    .S(_12564_),
    .Z(_12572_));
 MUX2_X1 _18464_ (.A(_00627_),
    .B(_00629_),
    .S(_12455_),
    .Z(_12573_));
 MUX2_X1 _18465_ (.A(_12572_),
    .B(_12573_),
    .S(_12459_),
    .Z(_12574_));
 MUX2_X1 _18466_ (.A(_00618_),
    .B(_00620_),
    .S(_12455_),
    .Z(_12575_));
 MUX2_X1 _18467_ (.A(_00619_),
    .B(_00621_),
    .S(_12455_),
    .Z(_12576_));
 MUX2_X1 _18468_ (.A(_12575_),
    .B(_12576_),
    .S(_12459_),
    .Z(_12577_));
 MUX2_X1 _18469_ (.A(_12574_),
    .B(_12577_),
    .S(_12358_),
    .Z(_12578_));
 MUX2_X1 _18470_ (.A(_12571_),
    .B(_12578_),
    .S(_12424_),
    .Z(_12579_));
 AOI21_X4 _18471_ (.A(_12562_),
    .B1(_12419_),
    .B2(_12579_),
    .ZN(_12580_));
 AOI21_X4 _18472_ (.A(_12540_),
    .B1(_12580_),
    .B2(_12343_),
    .ZN(_16349_));
 INV_X1 _18473_ (.A(_16349_),
    .ZN(_16353_));
 NAND2_X1 _18474_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(_10958_),
    .ZN(_12581_));
 MUX2_X1 _18475_ (.A(_00622_),
    .B(_00624_),
    .S(_12107_),
    .Z(_12582_));
 MUX2_X1 _18476_ (.A(_00623_),
    .B(_00625_),
    .S(_12107_),
    .Z(_12583_));
 MUX2_X1 _18477_ (.A(_12582_),
    .B(_12583_),
    .S(_10999_),
    .Z(_12584_));
 MUX2_X1 _18478_ (.A(_00606_),
    .B(_00608_),
    .S(_11849_),
    .Z(_12585_));
 MUX2_X1 _18479_ (.A(_00607_),
    .B(_00609_),
    .S(_11849_),
    .Z(_12586_));
 MUX2_X1 _18480_ (.A(_12585_),
    .B(_12586_),
    .S(_10999_),
    .Z(_12587_));
 MUX2_X1 _18481_ (.A(_12584_),
    .B(_12587_),
    .S(_10980_),
    .Z(_12588_));
 NOR2_X1 _18482_ (.A1(_11058_),
    .A2(_12588_),
    .ZN(_12589_));
 MUX2_X1 _18483_ (.A(_00626_),
    .B(_00628_),
    .S(_12200_),
    .Z(_12590_));
 MUX2_X1 _18484_ (.A(_00627_),
    .B(_00629_),
    .S(_12200_),
    .Z(_12591_));
 MUX2_X1 _18485_ (.A(_12590_),
    .B(_12591_),
    .S(_11256_),
    .Z(_12592_));
 MUX2_X1 _18486_ (.A(_00610_),
    .B(_00612_),
    .S(_12200_),
    .Z(_12593_));
 MUX2_X1 _18487_ (.A(_00611_),
    .B(_00613_),
    .S(_12200_),
    .Z(_12594_));
 MUX2_X1 _18488_ (.A(_12593_),
    .B(_12594_),
    .S(_10999_),
    .Z(_12595_));
 MUX2_X1 _18489_ (.A(_12592_),
    .B(_12595_),
    .S(_10980_),
    .Z(_12596_));
 NOR2_X1 _18490_ (.A1(_11223_),
    .A2(_12596_),
    .ZN(_12597_));
 NOR3_X4 _18491_ (.A1(_10995_),
    .A2(_12589_),
    .A3(_12597_),
    .ZN(_12598_));
 MUX2_X1 _18492_ (.A(_00614_),
    .B(_00616_),
    .S(_11006_),
    .Z(_12599_));
 NOR2_X1 _18493_ (.A1(_11093_),
    .A2(_12599_),
    .ZN(_12600_));
 MUX2_X1 _18494_ (.A(_00615_),
    .B(_00617_),
    .S(_11006_),
    .Z(_12601_));
 NOR2_X1 _18495_ (.A1(_11012_),
    .A2(_12601_),
    .ZN(_12602_));
 NOR3_X1 _18496_ (.A1(_10981_),
    .A2(_12600_),
    .A3(_12602_),
    .ZN(_12603_));
 NOR2_X1 _18497_ (.A1(_11015_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .ZN(_12604_));
 AOI21_X1 _18498_ (.A(_12604_),
    .B1(_00601_),
    .B2(_12503_),
    .ZN(_12605_));
 AOI221_X2 _18499_ (.A(_11051_),
    .B1(_12546_),
    .B2(_11031_),
    .C1(_12605_),
    .C2(_11271_),
    .ZN(_12606_));
 NOR3_X2 _18500_ (.A1(_10987_),
    .A2(_12603_),
    .A3(_12606_),
    .ZN(_12607_));
 MUX2_X1 _18501_ (.A(_00618_),
    .B(_00620_),
    .S(_12034_),
    .Z(_12608_));
 MUX2_X1 _18502_ (.A(_00619_),
    .B(_00621_),
    .S(_11224_),
    .Z(_12609_));
 MUX2_X1 _18503_ (.A(_12608_),
    .B(_12609_),
    .S(_12037_),
    .Z(_12610_));
 MUX2_X1 _18504_ (.A(_00602_),
    .B(_00604_),
    .S(_11224_),
    .Z(_12611_));
 MUX2_X1 _18505_ (.A(_00603_),
    .B(_00605_),
    .S(_11224_),
    .Z(_12612_));
 MUX2_X1 _18506_ (.A(_12611_),
    .B(_12612_),
    .S(_11227_),
    .Z(_12613_));
 MUX2_X1 _18507_ (.A(_12610_),
    .B(_12613_),
    .S(_10980_),
    .Z(_12614_));
 NOR2_X1 _18508_ (.A1(_11223_),
    .A2(_12614_),
    .ZN(_12615_));
 NOR3_X4 _18509_ (.A1(_11055_),
    .A2(_12607_),
    .A3(_12615_),
    .ZN(_12616_));
 OR2_X2 _18510_ (.A1(_12598_),
    .A2(_12616_),
    .ZN(_12617_));
 BUF_X1 _18511_ (.A(\cs_registers_i.pc_id_i[14] ),
    .Z(_12618_));
 NAND2_X1 _18512_ (.A1(_12618_),
    .A2(_11112_),
    .ZN(_12619_));
 OAI221_X2 _18513_ (.A(_12581_),
    .B1(_12617_),
    .B2(_11278_),
    .C1(_12619_),
    .C2(_11114_),
    .ZN(_16354_));
 INV_X1 _18514_ (.A(_16354_),
    .ZN(_16350_));
 NAND2_X1 _18515_ (.A1(_11002_),
    .A2(_12351_),
    .ZN(_12620_));
 AOI21_X4 _18516_ (.A(_11168_),
    .B1(_12348_),
    .B2(_12620_),
    .ZN(_12621_));
 MUX2_X1 _18517_ (.A(_00637_),
    .B(_00639_),
    .S(_12378_),
    .Z(_12622_));
 NOR2_X1 _18518_ (.A1(_12426_),
    .A2(_12622_),
    .ZN(_12623_));
 MUX2_X1 _18519_ (.A(_00638_),
    .B(_00640_),
    .S(_12378_),
    .Z(_12624_));
 NOR2_X1 _18520_ (.A1(_12368_),
    .A2(_12624_),
    .ZN(_12625_));
 NOR3_X1 _18521_ (.A1(_12425_),
    .A2(_12623_),
    .A3(_12625_),
    .ZN(_12626_));
 INV_X1 _18522_ (.A(_00631_),
    .ZN(_12627_));
 NOR2_X1 _18523_ (.A1(_12435_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .ZN(_12628_));
 AOI21_X1 _18524_ (.A(_12628_),
    .B1(_00632_),
    .B2(_12438_),
    .ZN(_12629_));
 AOI221_X2 _18525_ (.A(_12432_),
    .B1(_12627_),
    .B2(_12374_),
    .C1(_12629_),
    .C2(_12440_),
    .ZN(_12630_));
 NOR3_X1 _18526_ (.A1(_12356_),
    .A2(_12626_),
    .A3(_12630_),
    .ZN(_12631_));
 MUX2_X1 _18527_ (.A(_00641_),
    .B(_00643_),
    .S(_12377_),
    .Z(_12632_));
 MUX2_X1 _18528_ (.A(_00642_),
    .B(_00644_),
    .S(_12377_),
    .Z(_12633_));
 MUX2_X1 _18529_ (.A(_12632_),
    .B(_12633_),
    .S(_12445_),
    .Z(_12634_));
 MUX2_X1 _18530_ (.A(_00633_),
    .B(_00635_),
    .S(_12377_),
    .Z(_12635_));
 MUX2_X1 _18531_ (.A(_00634_),
    .B(_00636_),
    .S(_12398_),
    .Z(_12636_));
 MUX2_X1 _18532_ (.A(_12635_),
    .B(_12636_),
    .S(_12445_),
    .Z(_12637_));
 MUX2_X1 _18533_ (.A(_12634_),
    .B(_12637_),
    .S(_12450_),
    .Z(_12638_));
 NOR2_X1 _18534_ (.A1(_12384_),
    .A2(_12638_),
    .ZN(_12639_));
 NOR3_X2 _18535_ (.A1(_12355_),
    .A2(_12631_),
    .A3(_12639_),
    .ZN(_12640_));
 MUX2_X1 _18536_ (.A(_00653_),
    .B(_00655_),
    .S(_12455_),
    .Z(_12641_));
 MUX2_X1 _18537_ (.A(_00654_),
    .B(_00656_),
    .S(_12455_),
    .Z(_12642_));
 MUX2_X1 _18538_ (.A(_12641_),
    .B(_12642_),
    .S(_12459_),
    .Z(_12643_));
 MUX2_X1 _18539_ (.A(_00645_),
    .B(_00647_),
    .S(_12455_),
    .Z(_12644_));
 MUX2_X1 _18540_ (.A(_00646_),
    .B(_00648_),
    .S(_12457_),
    .Z(_12645_));
 MUX2_X1 _18541_ (.A(_12644_),
    .B(_12645_),
    .S(_12459_),
    .Z(_12646_));
 MUX2_X1 _18542_ (.A(_12643_),
    .B(_12646_),
    .S(_12358_),
    .Z(_12647_));
 MUX2_X1 _18543_ (.A(_00657_),
    .B(_00659_),
    .S(_12457_),
    .Z(_12648_));
 MUX2_X1 _18544_ (.A(_00658_),
    .B(_00660_),
    .S(_12457_),
    .Z(_12649_));
 MUX2_X1 _18545_ (.A(_12648_),
    .B(_12649_),
    .S(_12459_),
    .Z(_12650_));
 MUX2_X1 _18546_ (.A(_00649_),
    .B(_00651_),
    .S(_12457_),
    .Z(_12651_));
 MUX2_X1 _18547_ (.A(_00650_),
    .B(_00652_),
    .S(_12364_),
    .Z(_12652_));
 MUX2_X1 _18548_ (.A(_12651_),
    .B(_12652_),
    .S(_12459_),
    .Z(_12653_));
 MUX2_X1 _18549_ (.A(_12650_),
    .B(_12653_),
    .S(_12425_),
    .Z(_12654_));
 MUX2_X1 _18550_ (.A(_12647_),
    .B(_12654_),
    .S(_12424_),
    .Z(_12655_));
 AOI21_X4 _18551_ (.A(_12640_),
    .B1(_12655_),
    .B2(_12419_),
    .ZN(_12656_));
 AOI21_X4 _18552_ (.A(_12621_),
    .B1(_12656_),
    .B2(_12343_),
    .ZN(_16357_));
 INV_X1 _18553_ (.A(_16357_),
    .ZN(_16361_));
 NAND2_X1 _18554_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(_11221_),
    .ZN(_12657_));
 MUX2_X1 _18555_ (.A(_00653_),
    .B(_00655_),
    .S(_11783_),
    .Z(_12658_));
 MUX2_X1 _18556_ (.A(_00654_),
    .B(_00656_),
    .S(_11783_),
    .Z(_12659_));
 MUX2_X1 _18557_ (.A(_12658_),
    .B(_12659_),
    .S(_11271_),
    .Z(_12660_));
 MUX2_X1 _18558_ (.A(_00645_),
    .B(_00647_),
    .S(_11096_),
    .Z(_12661_));
 MUX2_X1 _18559_ (.A(_00646_),
    .B(_00648_),
    .S(_11096_),
    .Z(_12662_));
 MUX2_X1 _18560_ (.A(_12661_),
    .B(_12662_),
    .S(_11271_),
    .Z(_12663_));
 MUX2_X1 _18561_ (.A(_12660_),
    .B(_12663_),
    .S(_12117_),
    .Z(_12664_));
 NOR2_X1 _18562_ (.A1(_10988_),
    .A2(_12664_),
    .ZN(_12665_));
 BUF_X4 _18563_ (.A(_11239_),
    .Z(_12666_));
 MUX2_X1 _18564_ (.A(_00657_),
    .B(_00659_),
    .S(_12666_),
    .Z(_12667_));
 MUX2_X1 _18565_ (.A(_00658_),
    .B(_00660_),
    .S(_12666_),
    .Z(_12668_));
 MUX2_X1 _18566_ (.A(_12667_),
    .B(_12668_),
    .S(_11060_),
    .Z(_12669_));
 MUX2_X1 _18567_ (.A(_00649_),
    .B(_00651_),
    .S(_11783_),
    .Z(_12670_));
 MUX2_X1 _18568_ (.A(_00650_),
    .B(_00652_),
    .S(_11783_),
    .Z(_12671_));
 MUX2_X1 _18569_ (.A(_12670_),
    .B(_12671_),
    .S(_11060_),
    .Z(_12672_));
 MUX2_X1 _18570_ (.A(_12669_),
    .B(_12672_),
    .S(_10993_),
    .Z(_12673_));
 NOR2_X1 _18571_ (.A1(_11174_),
    .A2(_12673_),
    .ZN(_12674_));
 NOR3_X4 _18572_ (.A1(_10982_),
    .A2(_12665_),
    .A3(_12674_),
    .ZN(_12675_));
 MUX2_X1 _18573_ (.A(_00637_),
    .B(_00639_),
    .S(_11821_),
    .Z(_12676_));
 NOR2_X1 _18574_ (.A1(_11043_),
    .A2(_12676_),
    .ZN(_12677_));
 MUX2_X1 _18575_ (.A(_00638_),
    .B(_00640_),
    .S(_11246_),
    .Z(_12678_));
 NOR2_X1 _18576_ (.A1(_11795_),
    .A2(_12678_),
    .ZN(_12679_));
 NOR3_X1 _18577_ (.A1(_12117_),
    .A2(_12677_),
    .A3(_12679_),
    .ZN(_12680_));
 NOR2_X1 _18578_ (.A1(_11801_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .ZN(_12681_));
 AOI21_X1 _18579_ (.A(_12681_),
    .B1(_00632_),
    .B2(_11007_),
    .ZN(_12682_));
 AOI221_X2 _18580_ (.A(_11235_),
    .B1(_12627_),
    .B2(_11799_),
    .C1(_12682_),
    .C2(_11000_),
    .ZN(_12683_));
 NOR3_X2 _18581_ (.A1(_11177_),
    .A2(_12680_),
    .A3(_12683_),
    .ZN(_12684_));
 BUF_X4 _18582_ (.A(_11239_),
    .Z(_12685_));
 MUX2_X1 _18583_ (.A(_00641_),
    .B(_00643_),
    .S(_12685_),
    .Z(_12686_));
 MUX2_X1 _18584_ (.A(_00642_),
    .B(_00644_),
    .S(_12685_),
    .Z(_12687_));
 MUX2_X1 _18585_ (.A(_12686_),
    .B(_12687_),
    .S(_11074_),
    .Z(_12688_));
 MUX2_X1 _18586_ (.A(_00633_),
    .B(_00635_),
    .S(_12685_),
    .Z(_12689_));
 MUX2_X1 _18587_ (.A(_00634_),
    .B(_00636_),
    .S(_12685_),
    .Z(_12690_));
 MUX2_X1 _18588_ (.A(_12689_),
    .B(_12690_),
    .S(_11260_),
    .Z(_12691_));
 MUX2_X1 _18589_ (.A(_12688_),
    .B(_12691_),
    .S(_10993_),
    .Z(_12692_));
 NOR2_X1 _18590_ (.A1(_11174_),
    .A2(_12692_),
    .ZN(_12693_));
 NOR3_X4 _18591_ (.A1(_11053_),
    .A2(_12684_),
    .A3(_12693_),
    .ZN(_12694_));
 OR2_X1 _18592_ (.A1(_12675_),
    .A2(_12694_),
    .ZN(_12695_));
 NAND2_X1 _18593_ (.A1(\cs_registers_i.pc_id_i[15] ),
    .A2(_12219_),
    .ZN(_12696_));
 OAI221_X2 _18594_ (.A(_12657_),
    .B1(_12695_),
    .B2(_11818_),
    .C1(_12696_),
    .C2(_11115_),
    .ZN(_12697_));
 BUF_X4 _18595_ (.A(_12697_),
    .Z(_16362_));
 INV_X1 _18596_ (.A(_16362_),
    .ZN(_16358_));
 BUF_X2 _18597_ (.A(_15832_),
    .Z(_12698_));
 INV_X1 _18598_ (.A(_15823_),
    .ZN(_12699_));
 INV_X1 _18599_ (.A(_12515_),
    .ZN(_12700_));
 OAI21_X1 _18600_ (.A(_12699_),
    .B1(net275),
    .B2(_12700_),
    .ZN(_12701_));
 BUF_X4 _18601_ (.A(_15828_),
    .Z(_12702_));
 AOI21_X2 _18602_ (.A(_15827_),
    .B1(_12701_),
    .B2(_12702_),
    .ZN(_12703_));
 XNOR2_X2 _18603_ (.A(_12703_),
    .B(_12698_),
    .ZN(\alu_adder_result_ex[15] ));
 NOR3_X2 _18604_ (.A1(_12522_),
    .A2(_12700_),
    .A3(_12523_),
    .ZN(_12704_));
 NOR2_X1 _18605_ (.A1(_12702_),
    .A2(_12704_),
    .ZN(_12705_));
 AOI21_X1 _18606_ (.A(_15819_),
    .B1(_12531_),
    .B2(_12521_),
    .ZN(_12706_));
 OAI21_X1 _18607_ (.A(_12699_),
    .B1(_12706_),
    .B2(_12700_),
    .ZN(_12707_));
 MUX2_X1 _18608_ (.A(_12705_),
    .B(_12702_),
    .S(_12707_),
    .Z(_12708_));
 OR2_X1 _18609_ (.A1(_12702_),
    .A2(_12707_),
    .ZN(_12709_));
 AOI211_X2 _18610_ (.A(_12339_),
    .B(_12709_),
    .C1(_12341_),
    .C2(_12176_),
    .ZN(_12710_));
 AND2_X1 _18611_ (.A1(_12702_),
    .A2(_12704_),
    .ZN(_12711_));
 AND2_X1 _18612_ (.A1(_12335_),
    .A2(_12338_),
    .ZN(_12712_));
 OR3_X2 _18613_ (.A1(_11896_),
    .A2(_11917_),
    .A3(_12340_),
    .ZN(_12713_));
 OAI21_X4 _18614_ (.A(_12712_),
    .B1(_12713_),
    .B2(net360),
    .ZN(_12714_));
 AOI211_X2 _18615_ (.A(_12708_),
    .B(_12710_),
    .C1(_12711_),
    .C2(_12714_),
    .ZN(\alu_adder_result_ex[14] ));
 NAND2_X1 _18616_ (.A1(_11081_),
    .A2(_12351_),
    .ZN(_12715_));
 AOI21_X2 _18617_ (.A(_11168_),
    .B1(_12348_),
    .B2(_12715_),
    .ZN(_12716_));
 MUX2_X1 _18618_ (.A(_00668_),
    .B(_00670_),
    .S(_12378_),
    .Z(_12717_));
 NOR2_X1 _18619_ (.A1(_12426_),
    .A2(_12717_),
    .ZN(_12718_));
 MUX2_X1 _18620_ (.A(_00669_),
    .B(_00671_),
    .S(_12435_),
    .Z(_12719_));
 NOR2_X1 _18621_ (.A1(_12368_),
    .A2(_12719_),
    .ZN(_12720_));
 NOR3_X1 _18622_ (.A1(_12425_),
    .A2(_12718_),
    .A3(_12720_),
    .ZN(_12721_));
 INV_X1 _18623_ (.A(_00662_),
    .ZN(_12722_));
 NOR2_X1 _18624_ (.A1(_12547_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .ZN(_12723_));
 AOI21_X1 _18625_ (.A(_12723_),
    .B1(_00663_),
    .B2(_12438_),
    .ZN(_12724_));
 AOI221_X2 _18626_ (.A(_12432_),
    .B1(_12722_),
    .B2(_12374_),
    .C1(_12724_),
    .C2(_12440_),
    .ZN(_12725_));
 NOR3_X1 _18627_ (.A1(_12356_),
    .A2(_12721_),
    .A3(_12725_),
    .ZN(_12726_));
 MUX2_X1 _18628_ (.A(_00672_),
    .B(_00674_),
    .S(_12552_),
    .Z(_12727_));
 MUX2_X1 _18629_ (.A(_00673_),
    .B(_00675_),
    .S(_12552_),
    .Z(_12728_));
 MUX2_X1 _18630_ (.A(_12727_),
    .B(_12728_),
    .S(_12555_),
    .Z(_12729_));
 MUX2_X1 _18631_ (.A(_00664_),
    .B(_00666_),
    .S(_12377_),
    .Z(_12730_));
 MUX2_X1 _18632_ (.A(_00665_),
    .B(_00667_),
    .S(_12377_),
    .Z(_12731_));
 MUX2_X1 _18633_ (.A(_12730_),
    .B(_12731_),
    .S(_12555_),
    .Z(_12732_));
 MUX2_X1 _18634_ (.A(_12729_),
    .B(_12732_),
    .S(_12450_),
    .Z(_12733_));
 NOR2_X2 _18635_ (.A1(_12384_),
    .A2(_12733_),
    .ZN(_12734_));
 NOR3_X2 _18636_ (.A1(_12355_),
    .A2(_12726_),
    .A3(_12734_),
    .ZN(_12735_));
 BUF_X8 _18637_ (.A(_12563_),
    .Z(_12736_));
 MUX2_X1 _18638_ (.A(_00684_),
    .B(_00686_),
    .S(_12736_),
    .Z(_12737_));
 MUX2_X1 _18639_ (.A(_00685_),
    .B(_00687_),
    .S(_12564_),
    .Z(_12738_));
 MUX2_X1 _18640_ (.A(_12737_),
    .B(_12738_),
    .S(_12381_),
    .Z(_12739_));
 MUX2_X1 _18641_ (.A(_00676_),
    .B(_00678_),
    .S(_12564_),
    .Z(_12740_));
 MUX2_X1 _18642_ (.A(_00677_),
    .B(_00679_),
    .S(_12564_),
    .Z(_12741_));
 MUX2_X1 _18643_ (.A(_12740_),
    .B(_12741_),
    .S(_12381_),
    .Z(_12742_));
 MUX2_X1 _18644_ (.A(_12739_),
    .B(_12742_),
    .S(_12358_),
    .Z(_12743_));
 MUX2_X1 _18645_ (.A(_00688_),
    .B(_00690_),
    .S(_12564_),
    .Z(_12744_));
 MUX2_X1 _18646_ (.A(_00689_),
    .B(_00691_),
    .S(_12564_),
    .Z(_12745_));
 MUX2_X1 _18647_ (.A(_12744_),
    .B(_12745_),
    .S(_12381_),
    .Z(_12746_));
 MUX2_X1 _18648_ (.A(_00680_),
    .B(_00682_),
    .S(_12564_),
    .Z(_12747_));
 MUX2_X1 _18649_ (.A(_00681_),
    .B(_00683_),
    .S(_12455_),
    .Z(_12748_));
 MUX2_X1 _18650_ (.A(_12747_),
    .B(_12748_),
    .S(_12459_),
    .Z(_12749_));
 MUX2_X1 _18651_ (.A(_12746_),
    .B(_12749_),
    .S(_12358_),
    .Z(_12750_));
 MUX2_X1 _18652_ (.A(_12743_),
    .B(_12750_),
    .S(_12424_),
    .Z(_12751_));
 AOI21_X4 _18653_ (.A(_12735_),
    .B1(_12419_),
    .B2(_12751_),
    .ZN(_12752_));
 AOI21_X4 _18654_ (.A(_12716_),
    .B1(net281),
    .B2(_12343_),
    .ZN(_16370_));
 INV_X1 _18655_ (.A(_16370_),
    .ZN(_16366_));
 NAND2_X1 _18656_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(_10957_),
    .ZN(_12753_));
 MUX2_X1 _18657_ (.A(_00676_),
    .B(_00677_),
    .S(_10998_),
    .Z(_12754_));
 NAND2_X1 _18658_ (.A1(_11090_),
    .A2(_12754_),
    .ZN(_12755_));
 MUX2_X1 _18659_ (.A(_00678_),
    .B(_00679_),
    .S(_11059_),
    .Z(_12756_));
 INV_X1 _18660_ (.A(_12756_),
    .ZN(_12757_));
 NAND2_X1 _18661_ (.A1(_11067_),
    .A2(_11098_),
    .ZN(_12758_));
 OAI21_X1 _18662_ (.A(_12755_),
    .B1(_12757_),
    .B2(_12758_),
    .ZN(_12759_));
 MUX2_X1 _18663_ (.A(_00684_),
    .B(_00686_),
    .S(_11800_),
    .Z(_12760_));
 MUX2_X1 _18664_ (.A(_00685_),
    .B(_00687_),
    .S(_11800_),
    .Z(_12761_));
 MUX2_X1 _18665_ (.A(_12760_),
    .B(_12761_),
    .S(_11804_),
    .Z(_12762_));
 NOR2_X1 _18666_ (.A1(_10986_),
    .A2(_12068_),
    .ZN(_12763_));
 MUX2_X1 _18667_ (.A(_00688_),
    .B(_00690_),
    .S(_11244_),
    .Z(_12764_));
 MUX2_X1 _18668_ (.A(_00689_),
    .B(_00691_),
    .S(_11244_),
    .Z(_12765_));
 MUX2_X1 _18669_ (.A(_12764_),
    .B(_12765_),
    .S(_10998_),
    .Z(_12766_));
 MUX2_X1 _18670_ (.A(_00680_),
    .B(_00682_),
    .S(_11244_),
    .Z(_12767_));
 MUX2_X1 _18671_ (.A(_00681_),
    .B(_00683_),
    .S(_11244_),
    .Z(_12768_));
 MUX2_X1 _18672_ (.A(_12767_),
    .B(_12768_),
    .S(_10998_),
    .Z(_12769_));
 MUX2_X1 _18673_ (.A(_12766_),
    .B(_12769_),
    .S(_10992_),
    .Z(_12770_));
 AOI221_X2 _18674_ (.A(_12759_),
    .B1(_12762_),
    .B2(_12763_),
    .C1(_12770_),
    .C2(_11057_),
    .ZN(_12771_));
 OR2_X1 _18675_ (.A1(_10982_),
    .A2(_12771_),
    .ZN(_12772_));
 MUX2_X1 _18676_ (.A(_00668_),
    .B(_00670_),
    .S(_12503_),
    .Z(_12773_));
 NOR2_X1 _18677_ (.A1(_11061_),
    .A2(_12773_),
    .ZN(_12774_));
 MUX2_X1 _18678_ (.A(_00669_),
    .B(_00671_),
    .S(_11208_),
    .Z(_12775_));
 NOR2_X1 _18679_ (.A1(_11795_),
    .A2(_12775_),
    .ZN(_12776_));
 NOR3_X1 _18680_ (.A1(_12117_),
    .A2(_12774_),
    .A3(_12776_),
    .ZN(_12777_));
 NOR2_X1 _18681_ (.A1(_11066_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .ZN(_12778_));
 AOI21_X1 _18682_ (.A(_12778_),
    .B1(_00663_),
    .B2(_11097_),
    .ZN(_12779_));
 AOI221_X1 _18683_ (.A(_11235_),
    .B1(_12722_),
    .B2(_11799_),
    .C1(_12779_),
    .C2(_11269_),
    .ZN(_12780_));
 OR3_X1 _18684_ (.A1(_11177_),
    .A2(_12777_),
    .A3(_12780_),
    .ZN(_12781_));
 MUX2_X1 _18685_ (.A(_00672_),
    .B(_00674_),
    .S(_11241_),
    .Z(_12782_));
 MUX2_X1 _18686_ (.A(_00673_),
    .B(_00675_),
    .S(_11241_),
    .Z(_12783_));
 MUX2_X1 _18687_ (.A(_12782_),
    .B(_12783_),
    .S(_11075_),
    .Z(_12784_));
 MUX2_X1 _18688_ (.A(_00664_),
    .B(_00666_),
    .S(_11241_),
    .Z(_12785_));
 MUX2_X1 _18689_ (.A(_00665_),
    .B(_00667_),
    .S(_11241_),
    .Z(_12786_));
 MUX2_X1 _18690_ (.A(_12785_),
    .B(_12786_),
    .S(_11075_),
    .Z(_12787_));
 MUX2_X1 _18691_ (.A(_12784_),
    .B(_12787_),
    .S(_10994_),
    .Z(_12788_));
 OAI21_X2 _18692_ (.A(_12781_),
    .B1(_12788_),
    .B2(_11038_),
    .ZN(_12789_));
 OAI21_X4 _18693_ (.A(_12772_),
    .B1(_12789_),
    .B2(_11931_),
    .ZN(_12790_));
 NAND2_X1 _18694_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(_12219_),
    .ZN(_12791_));
 OAI221_X2 _18695_ (.A(_12753_),
    .B1(_12790_),
    .B2(_11278_),
    .C1(_12791_),
    .C2(_10978_),
    .ZN(_16365_));
 INV_X2 _18696_ (.A(_16365_),
    .ZN(_16369_));
 MUX2_X1 _18697_ (.A(_00715_),
    .B(_00717_),
    .S(_12363_),
    .Z(_12792_));
 MUX2_X1 _18698_ (.A(_00716_),
    .B(_00718_),
    .S(_12363_),
    .Z(_12793_));
 MUX2_X1 _18699_ (.A(_12792_),
    .B(_12793_),
    .S(_12380_),
    .Z(_12794_));
 MUX2_X1 _18700_ (.A(_00707_),
    .B(_00709_),
    .S(_12363_),
    .Z(_12795_));
 MUX2_X1 _18701_ (.A(_00708_),
    .B(_00710_),
    .S(_12363_),
    .Z(_12796_));
 MUX2_X1 _18702_ (.A(_12795_),
    .B(_12796_),
    .S(_12380_),
    .Z(_12797_));
 MUX2_X1 _18703_ (.A(_12794_),
    .B(_12797_),
    .S(_12357_),
    .Z(_12798_));
 MUX2_X1 _18704_ (.A(_00719_),
    .B(_00721_),
    .S(_12363_),
    .Z(_12799_));
 MUX2_X1 _18705_ (.A(_00720_),
    .B(_00722_),
    .S(_12363_),
    .Z(_12800_));
 MUX2_X1 _18706_ (.A(_12799_),
    .B(_12800_),
    .S(_12388_),
    .Z(_12801_));
 MUX2_X1 _18707_ (.A(_00711_),
    .B(_00713_),
    .S(_12363_),
    .Z(_12802_));
 MUX2_X1 _18708_ (.A(_00712_),
    .B(_00714_),
    .S(_12363_),
    .Z(_12803_));
 MUX2_X1 _18709_ (.A(_12802_),
    .B(_12803_),
    .S(_12388_),
    .Z(_12804_));
 MUX2_X1 _18710_ (.A(_12801_),
    .B(_12804_),
    .S(_12357_),
    .Z(_12805_));
 MUX2_X1 _18711_ (.A(_12798_),
    .B(_12805_),
    .S(_12423_),
    .Z(_12806_));
 BUF_X4 _18712_ (.A(_10736_),
    .Z(_12807_));
 MUX2_X1 _18713_ (.A(_00703_),
    .B(_00705_),
    .S(_12454_),
    .Z(_12808_));
 MUX2_X1 _18714_ (.A(_00704_),
    .B(_00706_),
    .S(_12454_),
    .Z(_12809_));
 MUX2_X1 _18715_ (.A(_12808_),
    .B(_12809_),
    .S(_12380_),
    .Z(_12810_));
 MUX2_X1 _18716_ (.A(_00695_),
    .B(_00697_),
    .S(_12454_),
    .Z(_12811_));
 MUX2_X1 _18717_ (.A(_00696_),
    .B(_00698_),
    .S(_12454_),
    .Z(_12812_));
 MUX2_X1 _18718_ (.A(_12811_),
    .B(_12812_),
    .S(_12380_),
    .Z(_12813_));
 MUX2_X1 _18719_ (.A(_12810_),
    .B(_12813_),
    .S(_12357_),
    .Z(_12814_));
 NOR2_X2 _18720_ (.A1(_12807_),
    .A2(_12814_),
    .ZN(_12815_));
 INV_X1 _18721_ (.A(_00693_),
    .ZN(_12816_));
 NOR2_X1 _18722_ (.A1(_12455_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .ZN(_12817_));
 AOI21_X1 _18723_ (.A(_12817_),
    .B1(_00694_),
    .B2(_12378_),
    .ZN(_12818_));
 AOI221_X1 _18724_ (.A(_12372_),
    .B1(_12816_),
    .B2(_12374_),
    .C1(_12818_),
    .C2(_12403_),
    .ZN(_12819_));
 MUX2_X1 _18725_ (.A(_00699_),
    .B(_00701_),
    .S(_12435_),
    .Z(_12820_));
 MUX2_X1 _18726_ (.A(_00700_),
    .B(_00702_),
    .S(_12435_),
    .Z(_12821_));
 MUX2_X1 _18727_ (.A(_12820_),
    .B(_12821_),
    .S(_12361_),
    .Z(_12822_));
 AOI21_X1 _18728_ (.A(_12819_),
    .B1(_12822_),
    .B2(_12432_),
    .ZN(_12823_));
 AOI21_X2 _18729_ (.A(_12815_),
    .B1(_12823_),
    .B2(_12384_),
    .ZN(_12824_));
 MUX2_X2 _18730_ (.A(_12806_),
    .B(_12824_),
    .S(_10764_),
    .Z(_12825_));
 NOR2_X2 _18731_ (.A1(_10805_),
    .A2(_12825_),
    .ZN(_12826_));
 NAND2_X1 _18732_ (.A1(_10989_),
    .A2(_12351_),
    .ZN(_12827_));
 AOI21_X1 _18733_ (.A(_12343_),
    .B1(_12348_),
    .B2(_12827_),
    .ZN(_12828_));
 NOR2_X2 _18734_ (.A1(_12826_),
    .A2(_12828_),
    .ZN(_16378_));
 INV_X1 _18735_ (.A(_16378_),
    .ZN(_16374_));
 NAND2_X1 _18736_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(_10958_),
    .ZN(_12829_));
 MUX2_X1 _18737_ (.A(_00699_),
    .B(_00701_),
    .S(_11821_),
    .Z(_12830_));
 NOR2_X1 _18738_ (.A1(_11043_),
    .A2(_12830_),
    .ZN(_12831_));
 MUX2_X1 _18739_ (.A(_00700_),
    .B(_00702_),
    .S(_11246_),
    .Z(_12832_));
 NOR2_X1 _18740_ (.A1(_11795_),
    .A2(_12832_),
    .ZN(_12833_));
 NOR3_X1 _18741_ (.A1(_12117_),
    .A2(_12831_),
    .A3(_12833_),
    .ZN(_12834_));
 NOR2_X1 _18742_ (.A1(_11801_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .ZN(_12835_));
 AOI21_X1 _18743_ (.A(_12835_),
    .B1(_00694_),
    .B2(_12297_),
    .ZN(_12836_));
 AOI221_X1 _18744_ (.A(_11235_),
    .B1(_12816_),
    .B2(_11799_),
    .C1(_12836_),
    .C2(_11269_),
    .ZN(_12837_));
 OR3_X1 _18745_ (.A1(_11177_),
    .A2(_12834_),
    .A3(_12837_),
    .ZN(_12838_));
 MUX2_X1 _18746_ (.A(_00703_),
    .B(_00705_),
    .S(_12297_),
    .Z(_12839_));
 MUX2_X1 _18747_ (.A(_00704_),
    .B(_00706_),
    .S(_12297_),
    .Z(_12840_));
 MUX2_X1 _18748_ (.A(_12839_),
    .B(_12840_),
    .S(_11028_),
    .Z(_12841_));
 NAND2_X1 _18749_ (.A1(_11252_),
    .A2(_12841_),
    .ZN(_12842_));
 MUX2_X1 _18750_ (.A(_00695_),
    .B(_00697_),
    .S(_12297_),
    .Z(_12843_));
 MUX2_X1 _18751_ (.A(_00696_),
    .B(_00698_),
    .S(_12297_),
    .Z(_12844_));
 MUX2_X1 _18752_ (.A(_12843_),
    .B(_12844_),
    .S(_11043_),
    .Z(_12845_));
 NAND2_X1 _18753_ (.A1(_10994_),
    .A2(_12845_),
    .ZN(_12846_));
 NAND3_X2 _18754_ (.A1(_10988_),
    .A2(_12842_),
    .A3(_12846_),
    .ZN(_12847_));
 AOI21_X4 _18755_ (.A(_11931_),
    .B1(_12838_),
    .B2(_12847_),
    .ZN(_12848_));
 MUX2_X1 _18756_ (.A(_00711_),
    .B(_00713_),
    .S(_11850_),
    .Z(_12849_));
 MUX2_X1 _18757_ (.A(_00712_),
    .B(_00714_),
    .S(_11850_),
    .Z(_12850_));
 MUX2_X1 _18758_ (.A(_12849_),
    .B(_12850_),
    .S(_11805_),
    .Z(_12851_));
 MUX2_X1 _18759_ (.A(_00709_),
    .B(_00710_),
    .S(_11027_),
    .Z(_12852_));
 MUX2_X1 _18760_ (.A(_00707_),
    .B(_00708_),
    .S(_11042_),
    .Z(_12853_));
 AOI222_X2 _18761_ (.A1(_11085_),
    .A2(_12851_),
    .B1(_12852_),
    .B2(_11100_),
    .C1(_12853_),
    .C2(_11091_),
    .ZN(_12854_));
 NAND2_X1 _18762_ (.A1(_11053_),
    .A2(_12854_),
    .ZN(_12855_));
 MUX2_X1 _18763_ (.A(_00717_),
    .B(_00718_),
    .S(_11227_),
    .Z(_12856_));
 AOI21_X2 _18764_ (.A(_10986_),
    .B1(_12856_),
    .B2(_11008_),
    .ZN(_12857_));
 MUX2_X1 _18765_ (.A(_00721_),
    .B(_00722_),
    .S(_11041_),
    .Z(_12858_));
 AOI21_X2 _18766_ (.A(_11036_),
    .B1(_12858_),
    .B2(_11254_),
    .ZN(_12859_));
 OAI21_X2 _18767_ (.A(_11081_),
    .B1(_12857_),
    .B2(_12859_),
    .ZN(_12860_));
 MUX2_X1 _18768_ (.A(_00719_),
    .B(_00720_),
    .S(_11256_),
    .Z(_12861_));
 INV_X1 _18769_ (.A(_12861_),
    .ZN(_12862_));
 MUX2_X1 _18770_ (.A(_00715_),
    .B(_00716_),
    .S(_11271_),
    .Z(_12863_));
 INV_X1 _18771_ (.A(_12863_),
    .ZN(_12864_));
 AOI221_X2 _18772_ (.A(_12117_),
    .B1(_12859_),
    .B2(_12862_),
    .C1(_12864_),
    .C2(_12857_),
    .ZN(_12865_));
 AOI21_X4 _18773_ (.A(_12855_),
    .B1(_12860_),
    .B2(_12865_),
    .ZN(_12866_));
 NOR2_X2 _18774_ (.A1(_12848_),
    .A2(_12866_),
    .ZN(_12867_));
 CLKBUF_X2 _18775_ (.A(\cs_registers_i.pc_id_i[17] ),
    .Z(_12868_));
 NAND2_X1 _18776_ (.A1(_12868_),
    .A2(_11112_),
    .ZN(_12869_));
 OAI221_X1 _18777_ (.A(_12829_),
    .B1(_12867_),
    .B2(_11278_),
    .C1(_12869_),
    .C2(_10978_),
    .ZN(_12870_));
 CLKBUF_X3 _18778_ (.A(_12870_),
    .Z(_16373_));
 INV_X1 _18779_ (.A(_16373_),
    .ZN(_16377_));
 BUF_X2 _18780_ (.A(_15840_),
    .Z(_12871_));
 INV_X1 _18781_ (.A(_15831_),
    .ZN(_12872_));
 AOI21_X1 _18782_ (.A(_15827_),
    .B1(_15823_),
    .B2(_12702_),
    .ZN(_12873_));
 INV_X1 _18783_ (.A(_12698_),
    .ZN(_12874_));
 OAI21_X1 _18784_ (.A(_12872_),
    .B1(_12873_),
    .B2(_12874_),
    .ZN(_12875_));
 BUF_X4 _18785_ (.A(_15836_),
    .Z(_12876_));
 AOI21_X2 _18786_ (.A(_15835_),
    .B1(_12875_),
    .B2(_12876_),
    .ZN(_12877_));
 NAND4_X1 _18787_ (.A1(_12515_),
    .A2(_12702_),
    .A3(_12698_),
    .A4(_12876_),
    .ZN(_12878_));
 OR2_X1 _18788_ (.A1(net275),
    .A2(_12878_),
    .ZN(_12879_));
 AND2_X2 _18789_ (.A1(_12877_),
    .A2(_12879_),
    .ZN(_12880_));
 XOR2_X2 _18790_ (.A(_12871_),
    .B(_12880_),
    .Z(_12881_));
 INV_X4 _18791_ (.A(_12881_),
    .ZN(\alu_adder_result_ex[17] ));
 NAND3_X1 _18792_ (.A1(_12521_),
    .A2(_12515_),
    .A3(_12702_),
    .ZN(_12882_));
 OR2_X1 _18793_ (.A1(_12874_),
    .A2(_12882_),
    .ZN(_12883_));
 OR2_X1 _18794_ (.A1(_12876_),
    .A2(_12883_),
    .ZN(_12884_));
 AOI21_X1 _18795_ (.A(_15823_),
    .B1(_15819_),
    .B2(_12515_),
    .ZN(_12885_));
 INV_X1 _18796_ (.A(_12885_),
    .ZN(_12886_));
 AOI21_X2 _18797_ (.A(_15827_),
    .B1(_12886_),
    .B2(_12702_),
    .ZN(_12887_));
 NAND3_X1 _18798_ (.A1(_12876_),
    .A2(_12872_),
    .A3(_12887_),
    .ZN(_12888_));
 MUX2_X2 _18799_ (.A(_12884_),
    .B(_12888_),
    .S(_12538_),
    .Z(_12889_));
 AOI21_X1 _18800_ (.A(_12874_),
    .B1(_12887_),
    .B2(_12882_),
    .ZN(_12890_));
 OAI21_X1 _18801_ (.A(_12876_),
    .B1(_15831_),
    .B2(_12890_),
    .ZN(_12891_));
 INV_X1 _18802_ (.A(_12876_),
    .ZN(_12892_));
 INV_X1 _18803_ (.A(_12887_),
    .ZN(_12893_));
 AOI21_X1 _18804_ (.A(_15831_),
    .B1(_12893_),
    .B2(_12698_),
    .ZN(_12894_));
 NAND2_X1 _18805_ (.A1(_12892_),
    .A2(_12894_),
    .ZN(_12895_));
 NAND2_X2 _18806_ (.A1(_12891_),
    .A2(_12895_),
    .ZN(_12896_));
 NAND2_X4 _18807_ (.A1(_12889_),
    .A2(_12896_),
    .ZN(\alu_adder_result_ex[16] ));
 NAND2_X1 _18808_ (.A1(_11056_),
    .A2(_12351_),
    .ZN(_12897_));
 AOI21_X2 _18809_ (.A(_11168_),
    .B1(_12348_),
    .B2(_12897_),
    .ZN(_12898_));
 MUX2_X1 _18810_ (.A(_00730_),
    .B(_00732_),
    .S(_12435_),
    .Z(_12899_));
 NOR2_X1 _18811_ (.A1(_12426_),
    .A2(_12899_),
    .ZN(_12900_));
 MUX2_X1 _18812_ (.A(_00731_),
    .B(_00733_),
    .S(_12435_),
    .Z(_12901_));
 NOR2_X1 _18813_ (.A1(_12368_),
    .A2(_12901_),
    .ZN(_12902_));
 NOR3_X1 _18814_ (.A1(_12425_),
    .A2(_12900_),
    .A3(_12902_),
    .ZN(_12903_));
 INV_X1 _18815_ (.A(_00724_),
    .ZN(_12904_));
 NOR2_X1 _18816_ (.A1(_12364_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .ZN(_12905_));
 AOI21_X1 _18817_ (.A(_12905_),
    .B1(_00725_),
    .B2(_12438_),
    .ZN(_12906_));
 AOI221_X2 _18818_ (.A(_12372_),
    .B1(_12904_),
    .B2(_12374_),
    .C1(_12906_),
    .C2(_12440_),
    .ZN(_12907_));
 NOR3_X1 _18819_ (.A1(_12356_),
    .A2(_12903_),
    .A3(_12907_),
    .ZN(_12908_));
 MUX2_X1 _18820_ (.A(_00734_),
    .B(_00736_),
    .S(_12434_),
    .Z(_12909_));
 MUX2_X1 _18821_ (.A(_00735_),
    .B(_00737_),
    .S(_12552_),
    .Z(_12910_));
 BUF_X4 _18822_ (.A(_12359_),
    .Z(_12911_));
 MUX2_X1 _18823_ (.A(_12909_),
    .B(_12910_),
    .S(_12911_),
    .Z(_12912_));
 MUX2_X1 _18824_ (.A(_00726_),
    .B(_00728_),
    .S(_12552_),
    .Z(_12913_));
 MUX2_X1 _18825_ (.A(_00727_),
    .B(_00729_),
    .S(_12552_),
    .Z(_12914_));
 MUX2_X1 _18826_ (.A(_12913_),
    .B(_12914_),
    .S(_12911_),
    .Z(_12915_));
 MUX2_X1 _18827_ (.A(_12912_),
    .B(_12915_),
    .S(_12450_),
    .Z(_12916_));
 NOR2_X1 _18828_ (.A1(_12384_),
    .A2(_12916_),
    .ZN(_12917_));
 NOR3_X2 _18829_ (.A1(_12355_),
    .A2(_12908_),
    .A3(_12917_),
    .ZN(_12918_));
 BUF_X8 _18830_ (.A(net341),
    .Z(_12919_));
 BUF_X4 _18831_ (.A(_12919_),
    .Z(_12920_));
 MUX2_X1 _18832_ (.A(_00746_),
    .B(_00748_),
    .S(_12920_),
    .Z(_12921_));
 MUX2_X1 _18833_ (.A(_00747_),
    .B(_00749_),
    .S(_12920_),
    .Z(_12922_));
 MUX2_X1 _18834_ (.A(_12921_),
    .B(_12922_),
    .S(_12403_),
    .Z(_12923_));
 MUX2_X1 _18835_ (.A(_00738_),
    .B(_00740_),
    .S(_12920_),
    .Z(_12924_));
 MUX2_X1 _18836_ (.A(_00739_),
    .B(_00741_),
    .S(_12920_),
    .Z(_12925_));
 MUX2_X1 _18837_ (.A(_12924_),
    .B(_12925_),
    .S(_12403_),
    .Z(_12926_));
 MUX2_X1 _18838_ (.A(_12923_),
    .B(_12926_),
    .S(_12358_),
    .Z(_12927_));
 MUX2_X1 _18839_ (.A(_00750_),
    .B(_00752_),
    .S(_12920_),
    .Z(_12928_));
 MUX2_X1 _18840_ (.A(_00751_),
    .B(_00753_),
    .S(_12920_),
    .Z(_12929_));
 MUX2_X1 _18841_ (.A(_12928_),
    .B(_12929_),
    .S(_12403_),
    .Z(_12930_));
 MUX2_X1 _18842_ (.A(_00742_),
    .B(_00744_),
    .S(_12920_),
    .Z(_12931_));
 MUX2_X1 _18843_ (.A(_00743_),
    .B(_00745_),
    .S(_12920_),
    .Z(_12932_));
 MUX2_X1 _18844_ (.A(_12931_),
    .B(_12932_),
    .S(_12403_),
    .Z(_12933_));
 MUX2_X1 _18845_ (.A(_12930_),
    .B(_12933_),
    .S(_12358_),
    .Z(_12934_));
 MUX2_X1 _18846_ (.A(_12927_),
    .B(_12934_),
    .S(_12424_),
    .Z(_12935_));
 AOI21_X4 _18847_ (.A(_12918_),
    .B1(_12935_),
    .B2(_12419_),
    .ZN(_12936_));
 AOI21_X4 _18848_ (.A(_12898_),
    .B1(net286),
    .B2(_12343_),
    .ZN(_16386_));
 INV_X1 _18849_ (.A(_16386_),
    .ZN(_16382_));
 NAND2_X1 _18850_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(_11221_),
    .ZN(_12937_));
 MUX2_X1 _18851_ (.A(_00734_),
    .B(_00736_),
    .S(_11207_),
    .Z(_12938_));
 MUX2_X1 _18852_ (.A(_00735_),
    .B(_00737_),
    .S(_12223_),
    .Z(_12939_));
 MUX2_X1 _18853_ (.A(_12938_),
    .B(_12939_),
    .S(_12226_),
    .Z(_12940_));
 MUX2_X1 _18854_ (.A(_00726_),
    .B(_00728_),
    .S(_12223_),
    .Z(_12941_));
 MUX2_X1 _18855_ (.A(_00727_),
    .B(_00729_),
    .S(_12223_),
    .Z(_12942_));
 MUX2_X1 _18856_ (.A(_12941_),
    .B(_12942_),
    .S(_12226_),
    .Z(_12943_));
 MUX2_X1 _18857_ (.A(_12940_),
    .B(_12943_),
    .S(_10993_),
    .Z(_12944_));
 NOR2_X1 _18858_ (.A1(_11174_),
    .A2(_12944_),
    .ZN(_12945_));
 NOR2_X1 _18859_ (.A1(_11208_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .ZN(_12946_));
 AOI21_X1 _18860_ (.A(_12946_),
    .B1(_00725_),
    .B2(_11007_),
    .ZN(_12947_));
 AOI221_X1 _18861_ (.A(_11022_),
    .B1(_12904_),
    .B2(_11032_),
    .C1(_12947_),
    .C2(_11805_),
    .ZN(_12948_));
 MUX2_X1 _18862_ (.A(_00730_),
    .B(_00732_),
    .S(_12297_),
    .Z(_12949_));
 MUX2_X1 _18863_ (.A(_00731_),
    .B(_00733_),
    .S(_12297_),
    .Z(_12950_));
 MUX2_X1 _18864_ (.A(_12949_),
    .B(_12950_),
    .S(_11043_),
    .Z(_12951_));
 AOI21_X1 _18865_ (.A(_12948_),
    .B1(_12951_),
    .B2(_11252_),
    .ZN(_12952_));
 AOI21_X2 _18866_ (.A(_12945_),
    .B1(_12952_),
    .B2(_11038_),
    .ZN(_12953_));
 MUX2_X1 _18867_ (.A(_00748_),
    .B(_00749_),
    .S(_12098_),
    .Z(_12954_));
 AOI21_X1 _18868_ (.A(_10986_),
    .B1(_12954_),
    .B2(_11188_),
    .ZN(_12955_));
 MUX2_X1 _18869_ (.A(_00752_),
    .B(_00753_),
    .S(_11074_),
    .Z(_12956_));
 AOI21_X1 _18870_ (.A(_11037_),
    .B1(_12956_),
    .B2(_11068_),
    .ZN(_12957_));
 OAI21_X1 _18871_ (.A(_11069_),
    .B1(_12955_),
    .B2(_12957_),
    .ZN(_12958_));
 MUX2_X1 _18872_ (.A(_00750_),
    .B(_00751_),
    .S(_11042_),
    .Z(_12959_));
 INV_X1 _18873_ (.A(_12959_),
    .ZN(_12960_));
 MUX2_X1 _18874_ (.A(_00746_),
    .B(_00747_),
    .S(_11042_),
    .Z(_12961_));
 INV_X1 _18875_ (.A(_12961_),
    .ZN(_12962_));
 AOI22_X1 _18876_ (.A1(_12957_),
    .A2(_12960_),
    .B1(_12962_),
    .B2(_12955_),
    .ZN(_12963_));
 NAND3_X1 _18877_ (.A1(_11252_),
    .A2(_12958_),
    .A3(_12963_),
    .ZN(_12964_));
 MUX2_X1 _18878_ (.A(_00742_),
    .B(_00744_),
    .S(_12503_),
    .Z(_12965_));
 MUX2_X1 _18879_ (.A(_00743_),
    .B(_00745_),
    .S(_12503_),
    .Z(_12966_));
 MUX2_X1 _18880_ (.A(_12965_),
    .B(_12966_),
    .S(_11093_),
    .Z(_12967_));
 MUX2_X1 _18881_ (.A(_00738_),
    .B(_00739_),
    .S(_11000_),
    .Z(_12968_));
 MUX2_X1 _18882_ (.A(_00740_),
    .B(_00741_),
    .S(_11027_),
    .Z(_12969_));
 AOI222_X2 _18883_ (.A1(_11085_),
    .A2(_12967_),
    .B1(_12968_),
    .B2(_11091_),
    .C1(_12969_),
    .C2(_11100_),
    .ZN(_12970_));
 NAND2_X1 _18884_ (.A1(_12964_),
    .A2(_12970_),
    .ZN(_12971_));
 MUX2_X2 _18885_ (.A(_12953_),
    .B(_12971_),
    .S(_11931_),
    .Z(_12972_));
 BUF_X1 _18886_ (.A(\cs_registers_i.pc_id_i[18] ),
    .Z(_12973_));
 NAND2_X1 _18887_ (.A1(_12973_),
    .A2(_12219_),
    .ZN(_12974_));
 OAI221_X1 _18888_ (.A(_12937_),
    .B1(_12972_),
    .B2(_11818_),
    .C1(_12974_),
    .C2(_11115_),
    .ZN(_12975_));
 CLKBUF_X3 _18889_ (.A(_12975_),
    .Z(_16381_));
 INV_X2 _18890_ (.A(_16381_),
    .ZN(_16385_));
 NAND2_X1 _18891_ (.A1(_11054_),
    .A2(_12351_),
    .ZN(_12976_));
 AOI21_X2 _18892_ (.A(_11168_),
    .B1(_12348_),
    .B2(_12976_),
    .ZN(_12977_));
 MUX2_X1 _18893_ (.A(_00761_),
    .B(_00763_),
    .S(_12435_),
    .Z(_12978_));
 NOR2_X1 _18894_ (.A1(_12426_),
    .A2(_12978_),
    .ZN(_12979_));
 MUX2_X1 _18895_ (.A(_00762_),
    .B(_00764_),
    .S(_12435_),
    .Z(_12980_));
 NOR2_X1 _18896_ (.A1(_12368_),
    .A2(_12980_),
    .ZN(_12981_));
 NOR3_X1 _18897_ (.A1(_12425_),
    .A2(_12979_),
    .A3(_12981_),
    .ZN(_12982_));
 INV_X1 _18898_ (.A(_00755_),
    .ZN(_12983_));
 NOR2_X1 _18899_ (.A1(_12364_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .ZN(_12984_));
 AOI21_X1 _18900_ (.A(_12984_),
    .B1(_00756_),
    .B2(_12438_),
    .ZN(_12985_));
 AOI221_X2 _18901_ (.A(_12432_),
    .B1(_12983_),
    .B2(_12374_),
    .C1(_12985_),
    .C2(_12440_),
    .ZN(_12986_));
 NOR3_X2 _18902_ (.A1(_12356_),
    .A2(_12982_),
    .A3(_12986_),
    .ZN(_12987_));
 MUX2_X1 _18903_ (.A(_00765_),
    .B(_00767_),
    .S(_12552_),
    .Z(_12988_));
 MUX2_X1 _18904_ (.A(_00766_),
    .B(_00768_),
    .S(_12552_),
    .Z(_12989_));
 MUX2_X1 _18905_ (.A(_12988_),
    .B(_12989_),
    .S(_12555_),
    .Z(_12990_));
 MUX2_X1 _18906_ (.A(_00757_),
    .B(_00759_),
    .S(_12552_),
    .Z(_12991_));
 MUX2_X1 _18907_ (.A(_00758_),
    .B(_00760_),
    .S(_12552_),
    .Z(_12992_));
 MUX2_X1 _18908_ (.A(_12991_),
    .B(_12992_),
    .S(_12555_),
    .Z(_12993_));
 MUX2_X1 _18909_ (.A(_12990_),
    .B(_12993_),
    .S(_12450_),
    .Z(_12994_));
 NOR2_X1 _18910_ (.A1(_12384_),
    .A2(_12994_),
    .ZN(_12995_));
 NOR3_X2 _18911_ (.A1(_12355_),
    .A2(_12987_),
    .A3(_12995_),
    .ZN(_12996_));
 MUX2_X1 _18912_ (.A(_00777_),
    .B(_00779_),
    .S(_12437_),
    .Z(_12997_));
 MUX2_X1 _18913_ (.A(_00778_),
    .B(_00780_),
    .S(_12437_),
    .Z(_12998_));
 MUX2_X1 _18914_ (.A(_12997_),
    .B(_12998_),
    .S(_12381_),
    .Z(_12999_));
 MUX2_X1 _18915_ (.A(_00769_),
    .B(_00771_),
    .S(_12437_),
    .Z(_13000_));
 MUX2_X1 _18916_ (.A(_00770_),
    .B(_00772_),
    .S(_12437_),
    .Z(_13001_));
 MUX2_X1 _18917_ (.A(_13000_),
    .B(_13001_),
    .S(_12381_),
    .Z(_13002_));
 MUX2_X1 _18918_ (.A(_12999_),
    .B(_13002_),
    .S(_12358_),
    .Z(_13003_));
 MUX2_X1 _18919_ (.A(_00781_),
    .B(_00783_),
    .S(_12437_),
    .Z(_13004_));
 MUX2_X1 _18920_ (.A(_00782_),
    .B(_00784_),
    .S(_12437_),
    .Z(_13005_));
 MUX2_X1 _18921_ (.A(_13004_),
    .B(_13005_),
    .S(_12381_),
    .Z(_13006_));
 MUX2_X1 _18922_ (.A(_00773_),
    .B(_00775_),
    .S(_12437_),
    .Z(_13007_));
 MUX2_X1 _18923_ (.A(_00774_),
    .B(_00776_),
    .S(_12437_),
    .Z(_13008_));
 MUX2_X1 _18924_ (.A(_13007_),
    .B(_13008_),
    .S(_12381_),
    .Z(_13009_));
 MUX2_X1 _18925_ (.A(_13006_),
    .B(_13009_),
    .S(_12358_),
    .Z(_13010_));
 MUX2_X1 _18926_ (.A(_13003_),
    .B(_13010_),
    .S(_12424_),
    .Z(_13011_));
 AOI21_X4 _18927_ (.A(_12996_),
    .B1(_13011_),
    .B2(_12419_),
    .ZN(_13012_));
 AOI21_X4 _18928_ (.A(_12977_),
    .B1(net283),
    .B2(_12343_),
    .ZN(_16394_));
 INV_X1 _18929_ (.A(_16394_),
    .ZN(_16390_));
 NAND2_X1 _18930_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(_10958_),
    .ZN(_13013_));
 MUX2_X1 _18931_ (.A(_00777_),
    .B(_00779_),
    .S(_11245_),
    .Z(_13014_));
 MUX2_X1 _18932_ (.A(_00778_),
    .B(_00780_),
    .S(_11245_),
    .Z(_13015_));
 MUX2_X1 _18933_ (.A(_13014_),
    .B(_13015_),
    .S(_11074_),
    .Z(_13016_));
 MUX2_X1 _18934_ (.A(_00761_),
    .B(_00763_),
    .S(_11245_),
    .Z(_13017_));
 MUX2_X1 _18935_ (.A(_00762_),
    .B(_00764_),
    .S(_11245_),
    .Z(_13018_));
 MUX2_X1 _18936_ (.A(_13017_),
    .B(_13018_),
    .S(_11074_),
    .Z(_13019_));
 MUX2_X1 _18937_ (.A(_13016_),
    .B(_13019_),
    .S(_11780_),
    .Z(_13020_));
 NOR2_X1 _18938_ (.A1(_10988_),
    .A2(_13020_),
    .ZN(_13021_));
 MUX2_X1 _18939_ (.A(_00781_),
    .B(_00783_),
    .S(_12502_),
    .Z(_13022_));
 MUX2_X1 _18940_ (.A(_00782_),
    .B(_00784_),
    .S(_12502_),
    .Z(_13023_));
 MUX2_X1 _18941_ (.A(_13022_),
    .B(_13023_),
    .S(_12226_),
    .Z(_13024_));
 MUX2_X1 _18942_ (.A(_00765_),
    .B(_00767_),
    .S(_12502_),
    .Z(_13025_));
 MUX2_X1 _18943_ (.A(_00766_),
    .B(_00768_),
    .S(_12502_),
    .Z(_13026_));
 MUX2_X1 _18944_ (.A(_13025_),
    .B(_13026_),
    .S(_12226_),
    .Z(_13027_));
 MUX2_X1 _18945_ (.A(_13024_),
    .B(_13027_),
    .S(_11780_),
    .Z(_13028_));
 NOR2_X1 _18946_ (.A1(_11174_),
    .A2(_13028_),
    .ZN(_13029_));
 NOR3_X4 _18947_ (.A1(_10995_),
    .A2(_13021_),
    .A3(_13029_),
    .ZN(_13030_));
 MUX2_X1 _18948_ (.A(_00769_),
    .B(_00771_),
    .S(_11208_),
    .Z(_13031_));
 NOR2_X1 _18949_ (.A1(_11061_),
    .A2(_13031_),
    .ZN(_13032_));
 MUX2_X1 _18950_ (.A(_00770_),
    .B(_00772_),
    .S(_11801_),
    .Z(_13033_));
 NOR2_X1 _18951_ (.A1(_11795_),
    .A2(_13033_),
    .ZN(_13034_));
 NOR3_X1 _18952_ (.A1(_10981_),
    .A2(_13032_),
    .A3(_13034_),
    .ZN(_13035_));
 NOR2_X1 _18953_ (.A1(_11066_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .ZN(_13036_));
 AOI21_X1 _18954_ (.A(_13036_),
    .B1(_00756_),
    .B2(_11097_),
    .ZN(_13037_));
 AOI221_X2 _18955_ (.A(_11051_),
    .B1(_12983_),
    .B2(_11799_),
    .C1(_13037_),
    .C2(_11269_),
    .ZN(_13038_));
 NOR3_X2 _18956_ (.A1(_11177_),
    .A2(_13035_),
    .A3(_13038_),
    .ZN(_13039_));
 MUX2_X1 _18957_ (.A(_00773_),
    .B(_00775_),
    .S(_11800_),
    .Z(_13040_));
 MUX2_X1 _18958_ (.A(_00774_),
    .B(_00776_),
    .S(_11800_),
    .Z(_13041_));
 MUX2_X1 _18959_ (.A(_13040_),
    .B(_13041_),
    .S(_11092_),
    .Z(_13042_));
 MUX2_X1 _18960_ (.A(_00757_),
    .B(_00759_),
    .S(_11800_),
    .Z(_13043_));
 MUX2_X1 _18961_ (.A(_00758_),
    .B(_00760_),
    .S(_11207_),
    .Z(_13044_));
 MUX2_X1 _18962_ (.A(_13043_),
    .B(_13044_),
    .S(_11092_),
    .Z(_13045_));
 MUX2_X1 _18963_ (.A(_13042_),
    .B(_13045_),
    .S(_10980_),
    .Z(_13046_));
 NOR2_X1 _18964_ (.A1(_11838_),
    .A2(_13046_),
    .ZN(_13047_));
 NOR3_X4 _18965_ (.A1(_11055_),
    .A2(_13039_),
    .A3(_13047_),
    .ZN(_13048_));
 OR2_X2 _18966_ (.A1(_13030_),
    .A2(_13048_),
    .ZN(_13049_));
 NAND2_X1 _18967_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(_12219_),
    .ZN(_13050_));
 OAI221_X2 _18968_ (.A(_13013_),
    .B1(_13049_),
    .B2(_11278_),
    .C1(_13050_),
    .C2(_10978_),
    .ZN(_13051_));
 BUF_X4 _18969_ (.A(_13051_),
    .Z(_16389_));
 INV_X2 _18970_ (.A(_16389_),
    .ZN(_16393_));
 BUF_X2 _18971_ (.A(_15848_),
    .Z(_13052_));
 INV_X2 _18972_ (.A(_13052_),
    .ZN(_13053_));
 CLKBUF_X3 _18973_ (.A(_15844_),
    .Z(_13054_));
 AOI21_X2 _18974_ (.A(_15843_),
    .B1(_15839_),
    .B2(_13054_),
    .ZN(_13055_));
 NAND2_X1 _18975_ (.A1(_12871_),
    .A2(_13054_),
    .ZN(_13056_));
 OAI21_X2 _18976_ (.A(_13055_),
    .B1(_13056_),
    .B2(_12880_),
    .ZN(_13057_));
 XNOR2_X2 _18977_ (.A(_13057_),
    .B(_13053_),
    .ZN(\alu_adder_result_ex[19] ));
 AND4_X1 _18978_ (.A1(_12702_),
    .A2(_12698_),
    .A3(_12876_),
    .A4(_12871_),
    .ZN(_13058_));
 NAND2_X1 _18979_ (.A1(_12707_),
    .A2(_13058_),
    .ZN(_13059_));
 INV_X1 _18980_ (.A(_15835_),
    .ZN(_13060_));
 AOI21_X1 _18981_ (.A(_15831_),
    .B1(_15827_),
    .B2(_12698_),
    .ZN(_13061_));
 OAI21_X1 _18982_ (.A(_13060_),
    .B1(_13061_),
    .B2(_12892_),
    .ZN(_13062_));
 AOI21_X2 _18983_ (.A(_15839_),
    .B1(_13062_),
    .B2(_12871_),
    .ZN(_13063_));
 NAND2_X2 _18984_ (.A1(_13059_),
    .A2(_13063_),
    .ZN(_13064_));
 AND2_X2 _18985_ (.A1(_13054_),
    .A2(_13064_),
    .ZN(_13065_));
 AND2_X2 _18986_ (.A1(_12704_),
    .A2(_13058_),
    .ZN(_13066_));
 NOR3_X4 _18987_ (.A1(_13054_),
    .A2(_13064_),
    .A3(_13066_),
    .ZN(_13067_));
 NOR2_X1 _18988_ (.A1(_13054_),
    .A2(_13064_),
    .ZN(_13068_));
 AND2_X1 _18989_ (.A1(_13054_),
    .A2(_13066_),
    .ZN(_13069_));
 MUX2_X2 _18990_ (.A(_13068_),
    .B(_13069_),
    .S(_12714_),
    .Z(_13070_));
 NOR3_X4 _18991_ (.A1(_13065_),
    .A2(_13067_),
    .A3(_13070_),
    .ZN(\alu_adder_result_ex[18] ));
 NAND3_X1 _18992_ (.A1(_10878_),
    .A2(_10836_),
    .A3(_12349_),
    .ZN(_13071_));
 NAND3_X2 _18993_ (.A1(_11121_),
    .A2(_12348_),
    .A3(_13071_),
    .ZN(_13072_));
 BUF_X2 _18994_ (.A(_13072_),
    .Z(_13073_));
 NOR2_X2 _18995_ (.A1(_10864_),
    .A2(_11125_),
    .ZN(_13074_));
 CLKBUF_X3 _18996_ (.A(_13074_),
    .Z(_13075_));
 AOI21_X1 _18997_ (.A(_13073_),
    .B1(_13075_),
    .B2(_12426_),
    .ZN(_13076_));
 CLKBUF_X3 _18998_ (.A(_10838_),
    .Z(_13077_));
 CLKBUF_X3 _18999_ (.A(_11121_),
    .Z(_13078_));
 BUF_X4 _19000_ (.A(_12400_),
    .Z(_13079_));
 MUX2_X1 _19001_ (.A(_00792_),
    .B(_00794_),
    .S(_13079_),
    .Z(_13080_));
 NOR2_X1 _19002_ (.A1(_12440_),
    .A2(_13080_),
    .ZN(_13081_));
 MUX2_X1 _19003_ (.A(_00793_),
    .B(_00795_),
    .S(_13079_),
    .Z(_13082_));
 NOR2_X1 _19004_ (.A1(_12367_),
    .A2(_13082_),
    .ZN(_13083_));
 NOR3_X1 _19005_ (.A1(_12450_),
    .A2(_13081_),
    .A3(_13083_),
    .ZN(_13084_));
 INV_X1 _19006_ (.A(_00786_),
    .ZN(_13085_));
 NOR2_X1 _19007_ (.A1(_12398_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .ZN(_13086_));
 AOI21_X1 _19008_ (.A(_13086_),
    .B1(_00787_),
    .B2(_12364_),
    .ZN(_13087_));
 AOI221_X1 _19009_ (.A(_10758_),
    .B1(_13085_),
    .B2(_12373_),
    .C1(_13087_),
    .C2(_12555_),
    .ZN(_13088_));
 NOR3_X1 _19010_ (.A1(_12423_),
    .A2(_13084_),
    .A3(_13088_),
    .ZN(_13089_));
 MUX2_X1 _19011_ (.A(_00796_),
    .B(_00798_),
    .S(_12400_),
    .Z(_13090_));
 MUX2_X1 _19012_ (.A(_00797_),
    .B(_00799_),
    .S(_12400_),
    .Z(_13091_));
 BUF_X4 _19013_ (.A(_10711_),
    .Z(_13092_));
 MUX2_X1 _19014_ (.A(_13090_),
    .B(_13091_),
    .S(_13092_),
    .Z(_13093_));
 MUX2_X1 _19015_ (.A(_00788_),
    .B(_00790_),
    .S(_12400_),
    .Z(_13094_));
 MUX2_X1 _19016_ (.A(_00789_),
    .B(_00791_),
    .S(_12400_),
    .Z(_13095_));
 MUX2_X1 _19017_ (.A(_13094_),
    .B(_13095_),
    .S(_13092_),
    .Z(_13096_));
 MUX2_X1 _19018_ (.A(_13093_),
    .B(_13096_),
    .S(_12408_),
    .Z(_13097_));
 NOR2_X2 _19019_ (.A1(_10736_),
    .A2(_13097_),
    .ZN(_13098_));
 NOR3_X2 _19020_ (.A1(_12354_),
    .A2(_13089_),
    .A3(_13098_),
    .ZN(_13099_));
 MUX2_X1 _19021_ (.A(_00808_),
    .B(_00810_),
    .S(_12363_),
    .Z(_13100_));
 BUF_X8 _19022_ (.A(net341),
    .Z(_13101_));
 MUX2_X1 _19023_ (.A(_00809_),
    .B(_00811_),
    .S(_13101_),
    .Z(_13102_));
 MUX2_X1 _19024_ (.A(_13100_),
    .B(_13102_),
    .S(_12388_),
    .Z(_13103_));
 MUX2_X1 _19025_ (.A(_00800_),
    .B(_00802_),
    .S(_13101_),
    .Z(_13104_));
 MUX2_X1 _19026_ (.A(_00801_),
    .B(_00803_),
    .S(_13101_),
    .Z(_13105_));
 MUX2_X1 _19027_ (.A(_13104_),
    .B(_13105_),
    .S(_12388_),
    .Z(_13106_));
 MUX2_X1 _19028_ (.A(_13103_),
    .B(_13106_),
    .S(_12394_),
    .Z(_13107_));
 MUX2_X1 _19029_ (.A(_00812_),
    .B(_00814_),
    .S(_13101_),
    .Z(_13108_));
 MUX2_X1 _19030_ (.A(_00813_),
    .B(_00815_),
    .S(_13101_),
    .Z(_13109_));
 MUX2_X1 _19031_ (.A(_13108_),
    .B(_13109_),
    .S(_12388_),
    .Z(_13110_));
 MUX2_X1 _19032_ (.A(_00804_),
    .B(_00806_),
    .S(_13101_),
    .Z(_13111_));
 MUX2_X1 _19033_ (.A(_00805_),
    .B(_00807_),
    .S(_13101_),
    .Z(_13112_));
 MUX2_X1 _19034_ (.A(_13111_),
    .B(_13112_),
    .S(_12388_),
    .Z(_13113_));
 MUX2_X1 _19035_ (.A(_13110_),
    .B(_13113_),
    .S(_12394_),
    .Z(_13114_));
 BUF_X4 _19036_ (.A(_10731_),
    .Z(_13115_));
 MUX2_X1 _19037_ (.A(_13107_),
    .B(_13114_),
    .S(_13115_),
    .Z(_13116_));
 BUF_X8 _19038_ (.A(_12354_),
    .Z(_13117_));
 AOI21_X4 _19039_ (.A(_13099_),
    .B1(_13117_),
    .B2(_13116_),
    .ZN(_13118_));
 OAI21_X4 _19040_ (.A(_13077_),
    .B1(_13078_),
    .B2(net368),
    .ZN(_13119_));
 OR2_X4 _19041_ (.A1(_13076_),
    .A2(_13119_),
    .ZN(_16397_));
 INV_X1 _19042_ (.A(_16397_),
    .ZN(_16401_));
 NAND2_X1 _19043_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(_10957_),
    .ZN(_13120_));
 MUX2_X1 _19044_ (.A(_00808_),
    .B(_00810_),
    .S(_12666_),
    .Z(_13121_));
 MUX2_X1 _19045_ (.A(_00809_),
    .B(_00811_),
    .S(_12666_),
    .Z(_13122_));
 MUX2_X1 _19046_ (.A(_13121_),
    .B(_13122_),
    .S(_11260_),
    .Z(_13123_));
 MUX2_X1 _19047_ (.A(_00792_),
    .B(_00794_),
    .S(_12666_),
    .Z(_13124_));
 MUX2_X1 _19048_ (.A(_00793_),
    .B(_00795_),
    .S(_12666_),
    .Z(_13125_));
 MUX2_X1 _19049_ (.A(_13124_),
    .B(_13125_),
    .S(_11060_),
    .Z(_13126_));
 MUX2_X1 _19050_ (.A(_13123_),
    .B(_13126_),
    .S(_11780_),
    .Z(_13127_));
 NOR2_X1 _19051_ (.A1(_10988_),
    .A2(_13127_),
    .ZN(_13128_));
 MUX2_X1 _19052_ (.A(_00812_),
    .B(_00814_),
    .S(_12685_),
    .Z(_13129_));
 MUX2_X1 _19053_ (.A(_00813_),
    .B(_00815_),
    .S(_12685_),
    .Z(_13130_));
 MUX2_X1 _19054_ (.A(_13129_),
    .B(_13130_),
    .S(_11260_),
    .Z(_13131_));
 MUX2_X1 _19055_ (.A(_00796_),
    .B(_00798_),
    .S(_12685_),
    .Z(_13132_));
 MUX2_X1 _19056_ (.A(_00797_),
    .B(_00799_),
    .S(_11240_),
    .Z(_13133_));
 MUX2_X1 _19057_ (.A(_13132_),
    .B(_13133_),
    .S(_11260_),
    .Z(_13134_));
 MUX2_X1 _19058_ (.A(_13131_),
    .B(_13134_),
    .S(_11780_),
    .Z(_13135_));
 NOR2_X1 _19059_ (.A1(_11174_),
    .A2(_13135_),
    .ZN(_13136_));
 NOR3_X4 _19060_ (.A1(_10995_),
    .A2(_13128_),
    .A3(_13136_),
    .ZN(_13137_));
 MUX2_X1 _19061_ (.A(_00800_),
    .B(_00802_),
    .S(_11246_),
    .Z(_13138_));
 NOR2_X1 _19062_ (.A1(_11061_),
    .A2(_13138_),
    .ZN(_13139_));
 MUX2_X1 _19063_ (.A(_00801_),
    .B(_00803_),
    .S(_11208_),
    .Z(_13140_));
 NOR2_X1 _19064_ (.A1(_11795_),
    .A2(_13140_),
    .ZN(_13141_));
 NOR3_X1 _19065_ (.A1(_10981_),
    .A2(_13139_),
    .A3(_13141_),
    .ZN(_13142_));
 NOR2_X1 _19066_ (.A1(_11850_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .ZN(_13143_));
 AOI21_X1 _19067_ (.A(_13143_),
    .B1(_00787_),
    .B2(_11016_),
    .ZN(_13144_));
 AOI221_X2 _19068_ (.A(_11051_),
    .B1(_13085_),
    .B2(_11799_),
    .C1(_13144_),
    .C2(_11269_),
    .ZN(_13145_));
 NOR3_X2 _19069_ (.A1(_11177_),
    .A2(_13142_),
    .A3(_13145_),
    .ZN(_13146_));
 MUX2_X1 _19070_ (.A(_00804_),
    .B(_00806_),
    .S(_12502_),
    .Z(_13147_));
 MUX2_X1 _19071_ (.A(_00805_),
    .B(_00807_),
    .S(_12502_),
    .Z(_13148_));
 MUX2_X1 _19072_ (.A(_13147_),
    .B(_13148_),
    .S(_12226_),
    .Z(_13149_));
 MUX2_X1 _19073_ (.A(_00788_),
    .B(_00790_),
    .S(_12502_),
    .Z(_13150_));
 MUX2_X1 _19074_ (.A(_00789_),
    .B(_00791_),
    .S(_12502_),
    .Z(_13151_));
 MUX2_X1 _19075_ (.A(_13150_),
    .B(_13151_),
    .S(_12226_),
    .Z(_13152_));
 MUX2_X1 _19076_ (.A(_13149_),
    .B(_13152_),
    .S(_11780_),
    .Z(_13153_));
 NOR2_X1 _19077_ (.A1(_11174_),
    .A2(_13153_),
    .ZN(_13154_));
 NOR3_X4 _19078_ (.A1(_11055_),
    .A2(_13146_),
    .A3(_13154_),
    .ZN(_13155_));
 OR2_X2 _19079_ (.A1(_13137_),
    .A2(_13155_),
    .ZN(_13156_));
 NAND2_X1 _19080_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(_11113_),
    .ZN(_13157_));
 OAI221_X2 _19081_ (.A(_13120_),
    .B1(_13156_),
    .B2(_11818_),
    .C1(_13157_),
    .C2(_11115_),
    .ZN(_16402_));
 INV_X2 _19082_ (.A(_16402_),
    .ZN(_16398_));
 AOI21_X1 _19083_ (.A(_13073_),
    .B1(_13075_),
    .B2(_12438_),
    .ZN(_13158_));
 MUX2_X1 _19084_ (.A(_00823_),
    .B(_00825_),
    .S(_12736_),
    .Z(_13159_));
 NOR2_X1 _19085_ (.A1(_12440_),
    .A2(_13159_),
    .ZN(_13160_));
 MUX2_X1 _19086_ (.A(_00824_),
    .B(_00826_),
    .S(_13079_),
    .Z(_13161_));
 NOR2_X1 _19087_ (.A1(_12367_),
    .A2(_13161_),
    .ZN(_13162_));
 NOR3_X1 _19088_ (.A1(_12450_),
    .A2(_13160_),
    .A3(_13162_),
    .ZN(_13163_));
 INV_X1 _19089_ (.A(_00817_),
    .ZN(_13164_));
 NOR2_X1 _19090_ (.A1(_12398_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .ZN(_13165_));
 AOI21_X1 _19091_ (.A(_13165_),
    .B1(_00818_),
    .B2(_12364_),
    .ZN(_13166_));
 AOI221_X2 _19092_ (.A(_10758_),
    .B1(_13164_),
    .B2(_12373_),
    .C1(_13166_),
    .C2(_12555_),
    .ZN(_13167_));
 NOR3_X1 _19093_ (.A1(_12423_),
    .A2(_13163_),
    .A3(_13167_),
    .ZN(_13168_));
 MUX2_X1 _19094_ (.A(_00827_),
    .B(_00829_),
    .S(_12400_),
    .Z(_13169_));
 BUF_X4 _19095_ (.A(_10750_),
    .Z(_13170_));
 MUX2_X1 _19096_ (.A(_00828_),
    .B(_00830_),
    .S(_13170_),
    .Z(_13171_));
 MUX2_X1 _19097_ (.A(_13169_),
    .B(_13171_),
    .S(_13092_),
    .Z(_13172_));
 MUX2_X1 _19098_ (.A(_00819_),
    .B(_00821_),
    .S(_13170_),
    .Z(_13173_));
 MUX2_X1 _19099_ (.A(_00820_),
    .B(_00822_),
    .S(_12919_),
    .Z(_13174_));
 MUX2_X1 _19100_ (.A(_13173_),
    .B(_13174_),
    .S(_13092_),
    .Z(_13175_));
 MUX2_X1 _19101_ (.A(_13172_),
    .B(_13175_),
    .S(_12408_),
    .Z(_13176_));
 NOR2_X1 _19102_ (.A1(_10736_),
    .A2(_13176_),
    .ZN(_13177_));
 NOR3_X2 _19103_ (.A1(_12354_),
    .A2(_13168_),
    .A3(_13177_),
    .ZN(_13178_));
 MUX2_X1 _19104_ (.A(_00839_),
    .B(_00841_),
    .S(_12385_),
    .Z(_13179_));
 BUF_X32 _19105_ (.A(net374),
    .Z(_13180_));
 MUX2_X1 _19106_ (.A(_00840_),
    .B(_00842_),
    .S(_13180_),
    .Z(_13181_));
 MUX2_X1 _19107_ (.A(_13179_),
    .B(_13181_),
    .S(_12392_),
    .Z(_13182_));
 MUX2_X1 _19108_ (.A(_00831_),
    .B(_00833_),
    .S(_12385_),
    .Z(_13183_));
 BUF_X32 _19109_ (.A(net374),
    .Z(_13184_));
 MUX2_X1 _19110_ (.A(_00832_),
    .B(_00834_),
    .S(_13184_),
    .Z(_13185_));
 MUX2_X1 _19111_ (.A(_13183_),
    .B(_13185_),
    .S(_12392_),
    .Z(_13186_));
 MUX2_X1 _19112_ (.A(_13182_),
    .B(_13186_),
    .S(_12394_),
    .Z(_13187_));
 MUX2_X1 _19113_ (.A(_00843_),
    .B(_00845_),
    .S(_13180_),
    .Z(_13188_));
 MUX2_X1 _19114_ (.A(_00844_),
    .B(_00846_),
    .S(_13184_),
    .Z(_13189_));
 MUX2_X1 _19115_ (.A(_13188_),
    .B(_13189_),
    .S(_12392_),
    .Z(_13190_));
 MUX2_X1 _19116_ (.A(_00835_),
    .B(_00837_),
    .S(_13184_),
    .Z(_13191_));
 BUF_X16 _19117_ (.A(_12376_),
    .Z(_13192_));
 MUX2_X1 _19118_ (.A(_00836_),
    .B(_00838_),
    .S(_13192_),
    .Z(_13193_));
 BUF_X4 _19119_ (.A(_12359_),
    .Z(_13194_));
 MUX2_X1 _19120_ (.A(_13191_),
    .B(_13193_),
    .S(_13194_),
    .Z(_13195_));
 MUX2_X1 _19121_ (.A(_13190_),
    .B(_13195_),
    .S(_12394_),
    .Z(_13196_));
 MUX2_X1 _19122_ (.A(_13187_),
    .B(_13196_),
    .S(_13115_),
    .Z(_13197_));
 AOI21_X4 _19123_ (.A(_13178_),
    .B1(_13117_),
    .B2(_13197_),
    .ZN(_13198_));
 OAI21_X1 _19124_ (.A(_13077_),
    .B1(_13078_),
    .B2(_13198_),
    .ZN(_13199_));
 OR2_X1 _19125_ (.A1(_13158_),
    .A2(_13199_),
    .ZN(_16405_));
 INV_X1 _19126_ (.A(_16405_),
    .ZN(_16409_));
 NAND2_X1 _19127_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(_10958_),
    .ZN(_13200_));
 MUX2_X1 _19128_ (.A(_00839_),
    .B(_00841_),
    .S(_11245_),
    .Z(_13201_));
 MUX2_X1 _19129_ (.A(_00840_),
    .B(_00842_),
    .S(_12685_),
    .Z(_13202_));
 MUX2_X1 _19130_ (.A(_13201_),
    .B(_13202_),
    .S(_11074_),
    .Z(_13203_));
 MUX2_X1 _19131_ (.A(_00823_),
    .B(_00825_),
    .S(_12685_),
    .Z(_13204_));
 MUX2_X1 _19132_ (.A(_00824_),
    .B(_00826_),
    .S(_12685_),
    .Z(_13205_));
 MUX2_X1 _19133_ (.A(_13204_),
    .B(_13205_),
    .S(_11260_),
    .Z(_13206_));
 MUX2_X1 _19134_ (.A(_13203_),
    .B(_13206_),
    .S(_11780_),
    .Z(_13207_));
 NOR2_X1 _19135_ (.A1(_10988_),
    .A2(_13207_),
    .ZN(_13208_));
 MUX2_X1 _19136_ (.A(_00843_),
    .B(_00845_),
    .S(_12502_),
    .Z(_13209_));
 MUX2_X1 _19137_ (.A(_00844_),
    .B(_00846_),
    .S(_11245_),
    .Z(_13210_));
 MUX2_X1 _19138_ (.A(_13209_),
    .B(_13210_),
    .S(_12226_),
    .Z(_13211_));
 MUX2_X1 _19139_ (.A(_00827_),
    .B(_00829_),
    .S(_11245_),
    .Z(_13212_));
 MUX2_X1 _19140_ (.A(_00828_),
    .B(_00830_),
    .S(_11245_),
    .Z(_13213_));
 MUX2_X1 _19141_ (.A(_13212_),
    .B(_13213_),
    .S(_11074_),
    .Z(_13214_));
 MUX2_X1 _19142_ (.A(_13211_),
    .B(_13214_),
    .S(_11780_),
    .Z(_13215_));
 NOR2_X1 _19143_ (.A1(_11174_),
    .A2(_13215_),
    .ZN(_13216_));
 NOR3_X4 _19144_ (.A1(_10995_),
    .A2(_13208_),
    .A3(_13216_),
    .ZN(_13217_));
 MUX2_X1 _19145_ (.A(_00831_),
    .B(_00833_),
    .S(_11208_),
    .Z(_13218_));
 NOR2_X1 _19146_ (.A1(_11061_),
    .A2(_13218_),
    .ZN(_13219_));
 MUX2_X1 _19147_ (.A(_00832_),
    .B(_00834_),
    .S(_11801_),
    .Z(_13220_));
 NOR2_X1 _19148_ (.A1(_11795_),
    .A2(_13220_),
    .ZN(_13221_));
 NOR3_X1 _19149_ (.A1(_10981_),
    .A2(_13219_),
    .A3(_13221_),
    .ZN(_13222_));
 NOR2_X1 _19150_ (.A1(_11066_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .ZN(_13223_));
 AOI21_X1 _19151_ (.A(_13223_),
    .B1(_00818_),
    .B2(_11016_),
    .ZN(_13224_));
 AOI221_X2 _19152_ (.A(_11051_),
    .B1(_13164_),
    .B2(_11799_),
    .C1(_13224_),
    .C2(_11269_),
    .ZN(_13225_));
 NOR3_X2 _19153_ (.A1(_11177_),
    .A2(_13222_),
    .A3(_13225_),
    .ZN(_13226_));
 MUX2_X1 _19154_ (.A(_00835_),
    .B(_00837_),
    .S(_11207_),
    .Z(_13227_));
 MUX2_X1 _19155_ (.A(_00836_),
    .B(_00838_),
    .S(_11207_),
    .Z(_13228_));
 MUX2_X1 _19156_ (.A(_13227_),
    .B(_13228_),
    .S(_11092_),
    .Z(_13229_));
 MUX2_X1 _19157_ (.A(_00819_),
    .B(_00821_),
    .S(_11207_),
    .Z(_13230_));
 MUX2_X1 _19158_ (.A(_00820_),
    .B(_00822_),
    .S(_11207_),
    .Z(_13231_));
 MUX2_X1 _19159_ (.A(_13230_),
    .B(_13231_),
    .S(_11092_),
    .Z(_13232_));
 MUX2_X1 _19160_ (.A(_13229_),
    .B(_13232_),
    .S(_10980_),
    .Z(_13233_));
 NOR2_X1 _19161_ (.A1(_11838_),
    .A2(_13233_),
    .ZN(_13234_));
 NOR3_X4 _19162_ (.A1(_11055_),
    .A2(_13226_),
    .A3(_13234_),
    .ZN(_13235_));
 OR2_X2 _19163_ (.A1(_13217_),
    .A2(_13235_),
    .ZN(_13236_));
 BUF_X1 _19164_ (.A(\cs_registers_i.pc_id_i[21] ),
    .Z(_13237_));
 NAND2_X1 _19165_ (.A1(_13237_),
    .A2(_12219_),
    .ZN(_13238_));
 OAI221_X2 _19166_ (.A(_13200_),
    .B1(_13236_),
    .B2(_11278_),
    .C1(_13238_),
    .C2(_10978_),
    .ZN(_13239_));
 BUF_X4 _19167_ (.A(_13239_),
    .Z(_16410_));
 INV_X2 _19168_ (.A(_16410_),
    .ZN(_16406_));
 BUF_X2 _19169_ (.A(_15856_),
    .Z(_13240_));
 INV_X1 _19170_ (.A(_15847_),
    .ZN(_13241_));
 OAI21_X1 _19171_ (.A(_13241_),
    .B1(_13055_),
    .B2(_13053_),
    .ZN(_13242_));
 BUF_X4 _19172_ (.A(_15852_),
    .Z(_13243_));
 AOI21_X1 _19173_ (.A(_15851_),
    .B1(_13242_),
    .B2(_13243_),
    .ZN(_13244_));
 AND3_X4 _19174_ (.A1(_13054_),
    .A2(_13052_),
    .A3(_13243_),
    .ZN(_13245_));
 NAND2_X2 _19175_ (.A1(_12871_),
    .A2(_13245_),
    .ZN(_13246_));
 OAI21_X2 _19176_ (.A(_13244_),
    .B1(_13246_),
    .B2(_12877_),
    .ZN(_13247_));
 NAND2_X2 _19177_ (.A1(_13247_),
    .A2(_13240_),
    .ZN(_13248_));
 INV_X1 _19178_ (.A(_13240_),
    .ZN(_13249_));
 OR3_X4 _19179_ (.A1(_13249_),
    .A2(_12878_),
    .A3(_13246_),
    .ZN(_13250_));
 OAI21_X4 _19180_ (.A(_13248_),
    .B1(_13250_),
    .B2(net275),
    .ZN(_13251_));
 NOR3_X1 _19181_ (.A1(net275),
    .A2(_12878_),
    .A3(_13246_),
    .ZN(_13252_));
 NOR3_X2 _19182_ (.A1(_13240_),
    .A2(_13247_),
    .A3(_13252_),
    .ZN(_13253_));
 NOR2_X4 _19183_ (.A1(_13251_),
    .A2(_13253_),
    .ZN(\alu_adder_result_ex[21] ));
 AOI21_X1 _19184_ (.A(_15839_),
    .B1(_15835_),
    .B2(_12871_),
    .ZN(_13254_));
 INV_X1 _19185_ (.A(_13254_),
    .ZN(_13255_));
 AOI21_X2 _19186_ (.A(_15843_),
    .B1(_13255_),
    .B2(_13054_),
    .ZN(_13256_));
 NAND3_X1 _19187_ (.A1(_13243_),
    .A2(_13241_),
    .A3(_13256_),
    .ZN(_13257_));
 AND3_X1 _19188_ (.A1(_12876_),
    .A2(_12871_),
    .A3(_13054_),
    .ZN(_13258_));
 OAI21_X2 _19189_ (.A(_12894_),
    .B1(_12883_),
    .B2(_12538_),
    .ZN(_13259_));
 AOI21_X2 _19190_ (.A(_13257_),
    .B1(_13258_),
    .B2(_13259_),
    .ZN(_13260_));
 INV_X1 _19191_ (.A(_13243_),
    .ZN(_13261_));
 AND4_X1 _19192_ (.A1(_13052_),
    .A2(_13261_),
    .A3(_13259_),
    .A4(_13258_),
    .ZN(_13262_));
 NAND3_X1 _19193_ (.A1(_13053_),
    .A2(_13243_),
    .A3(_13241_),
    .ZN(_13263_));
 NAND2_X1 _19194_ (.A1(_13052_),
    .A2(_13261_),
    .ZN(_13264_));
 OAI221_X2 _19195_ (.A(_13263_),
    .B1(_13264_),
    .B2(_13256_),
    .C1(_13243_),
    .C2(_13241_),
    .ZN(_13265_));
 NOR3_X4 _19196_ (.A1(_13262_),
    .A2(_13260_),
    .A3(_13265_),
    .ZN(_13266_));
 INV_X4 _19197_ (.A(_13266_),
    .ZN(\alu_adder_result_ex[20] ));
 AOI21_X1 _19198_ (.A(_13073_),
    .B1(_13075_),
    .B2(_12424_),
    .ZN(_13267_));
 MUX2_X1 _19199_ (.A(_00854_),
    .B(_00856_),
    .S(_12736_),
    .Z(_13268_));
 NOR2_X1 _19200_ (.A1(_12361_),
    .A2(_13268_),
    .ZN(_13269_));
 MUX2_X1 _19201_ (.A(_00855_),
    .B(_00857_),
    .S(_12437_),
    .Z(_13270_));
 NOR2_X1 _19202_ (.A1(_12368_),
    .A2(_13270_),
    .ZN(_13271_));
 NOR3_X1 _19203_ (.A1(_12409_),
    .A2(_13269_),
    .A3(_13271_),
    .ZN(_13272_));
 INV_X1 _19204_ (.A(_00848_),
    .ZN(_13273_));
 NOR2_X1 _19205_ (.A1(_13079_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .ZN(_13274_));
 AOI21_X1 _19206_ (.A(_13274_),
    .B1(_00849_),
    .B2(_12547_),
    .ZN(_13275_));
 AOI221_X2 _19207_ (.A(_12372_),
    .B1(_13273_),
    .B2(_12374_),
    .C1(_13275_),
    .C2(_12445_),
    .ZN(_13276_));
 NOR3_X2 _19208_ (.A1(_13115_),
    .A2(_13272_),
    .A3(_13276_),
    .ZN(_13277_));
 BUF_X4 _19209_ (.A(net379),
    .Z(_13278_));
 MUX2_X1 _19210_ (.A(_00858_),
    .B(_00860_),
    .S(_13278_),
    .Z(_13279_));
 MUX2_X1 _19211_ (.A(_00859_),
    .B(_00861_),
    .S(_13278_),
    .Z(_13280_));
 BUF_X4 _19212_ (.A(_12359_),
    .Z(_13281_));
 MUX2_X1 _19213_ (.A(_13279_),
    .B(_13280_),
    .S(_13281_),
    .Z(_13282_));
 MUX2_X1 _19214_ (.A(_00850_),
    .B(_00852_),
    .S(_12563_),
    .Z(_13283_));
 MUX2_X1 _19215_ (.A(_00851_),
    .B(_00853_),
    .S(_12563_),
    .Z(_13284_));
 MUX2_X1 _19216_ (.A(_13283_),
    .B(_13284_),
    .S(_13281_),
    .Z(_13285_));
 MUX2_X1 _19217_ (.A(_13282_),
    .B(_13285_),
    .S(_12357_),
    .Z(_13286_));
 NOR2_X1 _19218_ (.A1(_12807_),
    .A2(_13286_),
    .ZN(_13287_));
 NOR3_X4 _19219_ (.A1(_12355_),
    .A2(_13277_),
    .A3(_13287_),
    .ZN(_13288_));
 BUF_X16 _19220_ (.A(net374),
    .Z(_13289_));
 MUX2_X1 _19221_ (.A(_00870_),
    .B(_00872_),
    .S(_13289_),
    .Z(_13290_));
 BUF_X16 _19222_ (.A(net374),
    .Z(_13291_));
 MUX2_X1 _19223_ (.A(_00871_),
    .B(_00873_),
    .S(_13291_),
    .Z(_13292_));
 MUX2_X1 _19224_ (.A(_13290_),
    .B(_13292_),
    .S(_12360_),
    .Z(_13293_));
 MUX2_X1 _19225_ (.A(_00862_),
    .B(_00864_),
    .S(_13291_),
    .Z(_13294_));
 MUX2_X1 _19226_ (.A(_00863_),
    .B(_00865_),
    .S(_13291_),
    .Z(_13295_));
 MUX2_X1 _19227_ (.A(_13294_),
    .B(_13295_),
    .S(_12911_),
    .Z(_13296_));
 BUF_X4 _19228_ (.A(_12408_),
    .Z(_13297_));
 MUX2_X1 _19229_ (.A(_13293_),
    .B(_13296_),
    .S(_13297_),
    .Z(_13298_));
 MUX2_X1 _19230_ (.A(_00874_),
    .B(_00876_),
    .S(_13291_),
    .Z(_13299_));
 MUX2_X1 _19231_ (.A(_00875_),
    .B(_00877_),
    .S(_12434_),
    .Z(_13300_));
 MUX2_X1 _19232_ (.A(_13299_),
    .B(_13300_),
    .S(_12911_),
    .Z(_13301_));
 MUX2_X1 _19233_ (.A(_00866_),
    .B(_00868_),
    .S(_12434_),
    .Z(_13302_));
 MUX2_X1 _19234_ (.A(_00867_),
    .B(_00869_),
    .S(_12434_),
    .Z(_13303_));
 MUX2_X1 _19235_ (.A(_13302_),
    .B(_13303_),
    .S(_12911_),
    .Z(_13304_));
 MUX2_X1 _19236_ (.A(_13301_),
    .B(_13304_),
    .S(_12450_),
    .Z(_13305_));
 MUX2_X1 _19237_ (.A(_13298_),
    .B(_13305_),
    .S(_12356_),
    .Z(_13306_));
 AOI21_X4 _19238_ (.A(_13288_),
    .B1(_13117_),
    .B2(_13306_),
    .ZN(_13307_));
 OAI21_X1 _19239_ (.A(_13077_),
    .B1(_13078_),
    .B2(_13307_),
    .ZN(_13308_));
 OR2_X1 _19240_ (.A1(_13267_),
    .A2(_13308_),
    .ZN(_16413_));
 INV_X1 _19241_ (.A(_16413_),
    .ZN(_16417_));
 NAND2_X1 _19242_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(_11221_),
    .ZN(_13309_));
 MUX2_X1 _19243_ (.A(_00870_),
    .B(_00872_),
    .S(_12107_),
    .Z(_13310_));
 MUX2_X1 _19244_ (.A(_00871_),
    .B(_00873_),
    .S(_12107_),
    .Z(_13311_));
 MUX2_X1 _19245_ (.A(_13310_),
    .B(_13311_),
    .S(_10999_),
    .Z(_13312_));
 MUX2_X1 _19246_ (.A(_00862_),
    .B(_00864_),
    .S(_12107_),
    .Z(_13313_));
 MUX2_X1 _19247_ (.A(_00863_),
    .B(_00865_),
    .S(_12107_),
    .Z(_13314_));
 MUX2_X1 _19248_ (.A(_13313_),
    .B(_13314_),
    .S(_10999_),
    .Z(_13315_));
 MUX2_X1 _19249_ (.A(_13312_),
    .B(_13315_),
    .S(_12104_),
    .Z(_13316_));
 NOR2_X2 _19250_ (.A1(_11058_),
    .A2(_13316_),
    .ZN(_13317_));
 BUF_X4 _19251_ (.A(_11064_),
    .Z(_13318_));
 MUX2_X1 _19252_ (.A(_00874_),
    .B(_00876_),
    .S(_13318_),
    .Z(_13319_));
 MUX2_X1 _19253_ (.A(_00875_),
    .B(_00877_),
    .S(_13318_),
    .Z(_13320_));
 MUX2_X1 _19254_ (.A(_13319_),
    .B(_13320_),
    .S(_11256_),
    .Z(_13321_));
 MUX2_X1 _19255_ (.A(_00866_),
    .B(_00868_),
    .S(_13318_),
    .Z(_13322_));
 MUX2_X1 _19256_ (.A(_00867_),
    .B(_00869_),
    .S(_13318_),
    .Z(_13323_));
 MUX2_X1 _19257_ (.A(_13322_),
    .B(_13323_),
    .S(_11256_),
    .Z(_13324_));
 MUX2_X1 _19258_ (.A(_13321_),
    .B(_13324_),
    .S(_11232_),
    .Z(_13325_));
 NOR2_X1 _19259_ (.A1(_11223_),
    .A2(_13325_),
    .ZN(_13326_));
 NOR3_X4 _19260_ (.A1(_10981_),
    .A2(_13317_),
    .A3(_13326_),
    .ZN(_13327_));
 MUX2_X1 _19261_ (.A(_00854_),
    .B(_00856_),
    .S(_11006_),
    .Z(_13328_));
 NOR2_X1 _19262_ (.A1(_11805_),
    .A2(_13328_),
    .ZN(_13329_));
 MUX2_X1 _19263_ (.A(_00855_),
    .B(_00857_),
    .S(_11006_),
    .Z(_13330_));
 NOR2_X1 _19264_ (.A1(_11012_),
    .A2(_13330_),
    .ZN(_13331_));
 NOR3_X1 _19265_ (.A1(_12117_),
    .A2(_13329_),
    .A3(_13331_),
    .ZN(_13332_));
 NOR2_X1 _19266_ (.A1(_11096_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .ZN(_13333_));
 AOI21_X1 _19267_ (.A(_13333_),
    .B1(_00849_),
    .B2(_12503_),
    .ZN(_13334_));
 AOI221_X2 _19268_ (.A(_11235_),
    .B1(_13273_),
    .B2(_11031_),
    .C1(_13334_),
    .C2(_11060_),
    .ZN(_13335_));
 NOR3_X2 _19269_ (.A1(_10987_),
    .A2(_13332_),
    .A3(_13335_),
    .ZN(_13336_));
 MUX2_X1 _19270_ (.A(_00858_),
    .B(_00860_),
    .S(_12034_),
    .Z(_13337_));
 MUX2_X1 _19271_ (.A(_00859_),
    .B(_00861_),
    .S(_12034_),
    .Z(_13338_));
 MUX2_X1 _19272_ (.A(_13337_),
    .B(_13338_),
    .S(_12037_),
    .Z(_13339_));
 MUX2_X1 _19273_ (.A(_00850_),
    .B(_00852_),
    .S(_12034_),
    .Z(_13340_));
 MUX2_X1 _19274_ (.A(_00851_),
    .B(_00853_),
    .S(_12034_),
    .Z(_13341_));
 MUX2_X1 _19275_ (.A(_13340_),
    .B(_13341_),
    .S(_12037_),
    .Z(_13342_));
 MUX2_X1 _19276_ (.A(_13339_),
    .B(_13342_),
    .S(_11232_),
    .Z(_13343_));
 NOR2_X1 _19277_ (.A1(_11223_),
    .A2(_13343_),
    .ZN(_13344_));
 NOR3_X4 _19278_ (.A1(_11052_),
    .A2(_13336_),
    .A3(_13344_),
    .ZN(_13345_));
 OR2_X2 _19279_ (.A1(_13327_),
    .A2(_13345_),
    .ZN(_13346_));
 CLKBUF_X2 _19280_ (.A(\cs_registers_i.pc_id_i[22] ),
    .Z(_13347_));
 NAND2_X1 _19281_ (.A1(_13347_),
    .A2(_11112_),
    .ZN(_13348_));
 OAI221_X2 _19282_ (.A(_13309_),
    .B1(_13346_),
    .B2(_11278_),
    .C1(_13348_),
    .C2(_11114_),
    .ZN(_16418_));
 INV_X1 _19283_ (.A(_16418_),
    .ZN(_16414_));
 AOI21_X1 _19284_ (.A(_13073_),
    .B1(_13075_),
    .B2(_12432_),
    .ZN(_13349_));
 MUX2_X1 _19285_ (.A(_00885_),
    .B(_00887_),
    .S(_12736_),
    .Z(_13350_));
 NOR2_X1 _19286_ (.A1(_12361_),
    .A2(_13350_),
    .ZN(_13351_));
 MUX2_X1 _19287_ (.A(_00886_),
    .B(_00888_),
    .S(_12920_),
    .Z(_13352_));
 NOR2_X1 _19288_ (.A1(_12368_),
    .A2(_13352_),
    .ZN(_13353_));
 NOR3_X1 _19289_ (.A1(_12409_),
    .A2(_13351_),
    .A3(_13353_),
    .ZN(_13354_));
 INV_X1 _19290_ (.A(_00879_),
    .ZN(_13355_));
 NOR2_X1 _19291_ (.A1(_13079_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .ZN(_13356_));
 AOI21_X1 _19292_ (.A(_13356_),
    .B1(_00880_),
    .B2(_12547_),
    .ZN(_13357_));
 AOI221_X1 _19293_ (.A(_12372_),
    .B1(_13355_),
    .B2(_12373_),
    .C1(_13357_),
    .C2(_12445_),
    .ZN(_13358_));
 NOR3_X1 _19294_ (.A1(_13115_),
    .A2(_13354_),
    .A3(_13358_),
    .ZN(_13359_));
 MUX2_X1 _19295_ (.A(_00889_),
    .B(_00891_),
    .S(_13278_),
    .Z(_13360_));
 MUX2_X1 _19296_ (.A(_00890_),
    .B(_00892_),
    .S(_13278_),
    .Z(_13361_));
 MUX2_X1 _19297_ (.A(_13360_),
    .B(_13361_),
    .S(_13281_),
    .Z(_13362_));
 MUX2_X1 _19298_ (.A(_00881_),
    .B(_00883_),
    .S(_13278_),
    .Z(_13363_));
 MUX2_X1 _19299_ (.A(_00882_),
    .B(_00884_),
    .S(_12563_),
    .Z(_13364_));
 MUX2_X1 _19300_ (.A(_13363_),
    .B(_13364_),
    .S(_13281_),
    .Z(_13365_));
 MUX2_X1 _19301_ (.A(_13362_),
    .B(_13365_),
    .S(_12357_),
    .Z(_13366_));
 NOR2_X1 _19302_ (.A1(_12807_),
    .A2(_13366_),
    .ZN(_13367_));
 NOR3_X2 _19303_ (.A1(_12355_),
    .A2(_13359_),
    .A3(_13367_),
    .ZN(_13368_));
 MUX2_X1 _19304_ (.A(_00901_),
    .B(_00903_),
    .S(_13289_),
    .Z(_13369_));
 MUX2_X1 _19305_ (.A(_00902_),
    .B(_00904_),
    .S(_13289_),
    .Z(_13370_));
 MUX2_X1 _19306_ (.A(_13369_),
    .B(_13370_),
    .S(_12360_),
    .Z(_13371_));
 MUX2_X1 _19307_ (.A(_00893_),
    .B(_00895_),
    .S(_13289_),
    .Z(_13372_));
 MUX2_X1 _19308_ (.A(_00894_),
    .B(_00896_),
    .S(_13291_),
    .Z(_13373_));
 MUX2_X1 _19309_ (.A(_13372_),
    .B(_13373_),
    .S(_12911_),
    .Z(_13374_));
 MUX2_X1 _19310_ (.A(_13371_),
    .B(_13374_),
    .S(_13297_),
    .Z(_13375_));
 MUX2_X1 _19311_ (.A(_00905_),
    .B(_00907_),
    .S(_13291_),
    .Z(_13376_));
 MUX2_X1 _19312_ (.A(_00906_),
    .B(_00908_),
    .S(_12434_),
    .Z(_13377_));
 MUX2_X1 _19313_ (.A(_13376_),
    .B(_13377_),
    .S(_12911_),
    .Z(_13378_));
 MUX2_X1 _19314_ (.A(_00897_),
    .B(_00899_),
    .S(_12434_),
    .Z(_13379_));
 MUX2_X1 _19315_ (.A(_00898_),
    .B(_00900_),
    .S(_12434_),
    .Z(_13380_));
 MUX2_X1 _19316_ (.A(_13379_),
    .B(_13380_),
    .S(_12911_),
    .Z(_13381_));
 MUX2_X1 _19317_ (.A(_13378_),
    .B(_13381_),
    .S(_12450_),
    .Z(_13382_));
 MUX2_X1 _19318_ (.A(_13375_),
    .B(_13382_),
    .S(_12356_),
    .Z(_13383_));
 AOI21_X4 _19319_ (.A(_13368_),
    .B1(_13117_),
    .B2(_13383_),
    .ZN(_13384_));
 OAI21_X2 _19320_ (.A(_13077_),
    .B1(_13078_),
    .B2(net350),
    .ZN(_13385_));
 OR2_X4 _19321_ (.A1(_13349_),
    .A2(_13385_),
    .ZN(_16426_));
 INV_X1 _19322_ (.A(_16426_),
    .ZN(_16422_));
 NAND2_X1 _19323_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(_10958_),
    .ZN(_13386_));
 MUX2_X1 _19324_ (.A(_00901_),
    .B(_00903_),
    .S(_12188_),
    .Z(_13387_));
 MUX2_X1 _19325_ (.A(_00902_),
    .B(_00904_),
    .S(_12188_),
    .Z(_13388_));
 MUX2_X1 _19326_ (.A(_13387_),
    .B(_13388_),
    .S(_11804_),
    .Z(_13389_));
 MUX2_X1 _19327_ (.A(_00893_),
    .B(_00895_),
    .S(_12188_),
    .Z(_13390_));
 MUX2_X1 _19328_ (.A(_00894_),
    .B(_00896_),
    .S(_11800_),
    .Z(_13391_));
 MUX2_X1 _19329_ (.A(_13390_),
    .B(_13391_),
    .S(_11804_),
    .Z(_13392_));
 MUX2_X1 _19330_ (.A(_13389_),
    .B(_13392_),
    .S(_12104_),
    .Z(_13393_));
 NOR2_X1 _19331_ (.A1(_11177_),
    .A2(_13393_),
    .ZN(_13394_));
 MUX2_X1 _19332_ (.A(_00905_),
    .B(_00907_),
    .S(_11849_),
    .Z(_13395_));
 MUX2_X1 _19333_ (.A(_00906_),
    .B(_00908_),
    .S(_11849_),
    .Z(_13396_));
 MUX2_X1 _19334_ (.A(_13395_),
    .B(_13396_),
    .S(_12098_),
    .Z(_13397_));
 MUX2_X1 _19335_ (.A(_00897_),
    .B(_00899_),
    .S(_11849_),
    .Z(_13398_));
 MUX2_X1 _19336_ (.A(_00898_),
    .B(_00900_),
    .S(_11849_),
    .Z(_13399_));
 MUX2_X1 _19337_ (.A(_13398_),
    .B(_13399_),
    .S(_12098_),
    .Z(_13400_));
 MUX2_X1 _19338_ (.A(_13397_),
    .B(_13400_),
    .S(_12104_),
    .Z(_13401_));
 NOR2_X2 _19339_ (.A1(_11838_),
    .A2(_13401_),
    .ZN(_13402_));
 NOR3_X4 _19340_ (.A1(_10982_),
    .A2(_13394_),
    .A3(_13402_),
    .ZN(_13403_));
 MUX2_X1 _19341_ (.A(_00885_),
    .B(_00887_),
    .S(_11066_),
    .Z(_13404_));
 NOR2_X1 _19342_ (.A1(_11075_),
    .A2(_13404_),
    .ZN(_13405_));
 MUX2_X1 _19343_ (.A(_00886_),
    .B(_00888_),
    .S(_11066_),
    .Z(_13406_));
 NOR2_X1 _19344_ (.A1(_11795_),
    .A2(_13406_),
    .ZN(_13407_));
 NOR3_X1 _19345_ (.A1(_12117_),
    .A2(_13405_),
    .A3(_13407_),
    .ZN(_13408_));
 NOR2_X1 _19346_ (.A1(_11015_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .ZN(_13409_));
 AOI21_X1 _19347_ (.A(_13409_),
    .B1(_00880_),
    .B2(_11246_),
    .ZN(_13410_));
 AOI221_X2 _19348_ (.A(_11235_),
    .B1(_13355_),
    .B2(_11031_),
    .C1(_13410_),
    .C2(_11271_),
    .ZN(_13411_));
 NOR3_X2 _19349_ (.A1(_11058_),
    .A2(_13408_),
    .A3(_13411_),
    .ZN(_13412_));
 MUX2_X1 _19350_ (.A(_00889_),
    .B(_00891_),
    .S(_13318_),
    .Z(_13413_));
 MUX2_X1 _19351_ (.A(_00890_),
    .B(_00892_),
    .S(_13318_),
    .Z(_13414_));
 MUX2_X1 _19352_ (.A(_13413_),
    .B(_13414_),
    .S(_11256_),
    .Z(_13415_));
 MUX2_X1 _19353_ (.A(_00881_),
    .B(_00883_),
    .S(_13318_),
    .Z(_13416_));
 MUX2_X1 _19354_ (.A(_00882_),
    .B(_00884_),
    .S(_13318_),
    .Z(_13417_));
 MUX2_X1 _19355_ (.A(_13416_),
    .B(_13417_),
    .S(_11256_),
    .Z(_13418_));
 MUX2_X1 _19356_ (.A(_13415_),
    .B(_13418_),
    .S(_11232_),
    .Z(_13419_));
 NOR2_X1 _19357_ (.A1(_11223_),
    .A2(_13419_),
    .ZN(_13420_));
 NOR3_X4 _19358_ (.A1(_11053_),
    .A2(_13412_),
    .A3(_13420_),
    .ZN(_13421_));
 OR2_X2 _19359_ (.A1(_13403_),
    .A2(_13421_),
    .ZN(_13422_));
 CLKBUF_X2 _19360_ (.A(\cs_registers_i.pc_id_i[23] ),
    .Z(_13423_));
 NAND2_X1 _19361_ (.A1(_13423_),
    .A2(_12219_),
    .ZN(_13424_));
 OAI221_X2 _19362_ (.A(_13386_),
    .B1(_13422_),
    .B2(_11818_),
    .C1(_13424_),
    .C2(_10978_),
    .ZN(_13425_));
 BUF_X4 _19363_ (.A(_13425_),
    .Z(_16421_));
 INV_X1 _19364_ (.A(_16421_),
    .ZN(_16425_));
 BUF_X1 rebuffer68 (.A(\alu_adder_result_ex[23] ),
    .Z(net356));
 BUF_X2 _19366_ (.A(_15859_),
    .Z(_13427_));
 OR2_X4 _19367_ (.A1(_13251_),
    .A2(_15855_),
    .ZN(_13428_));
 CLKBUF_X3 _19368_ (.A(_15860_),
    .Z(_13429_));
 AOI21_X4 _19369_ (.A(_13427_),
    .B1(_13428_),
    .B2(_13429_),
    .ZN(_13430_));
 XNOR2_X2 _19370_ (.A(_13430_),
    .B(_15864_),
    .ZN(\alu_adder_result_ex[23] ));
 INV_X1 _19371_ (.A(_15851_),
    .ZN(_13431_));
 AOI21_X1 _19372_ (.A(_15847_),
    .B1(_15843_),
    .B2(_13052_),
    .ZN(_13432_));
 OAI21_X1 _19373_ (.A(_13431_),
    .B1(_13432_),
    .B2(_13261_),
    .ZN(_13433_));
 AOI21_X2 _19374_ (.A(_15855_),
    .B1(_13433_),
    .B2(_13240_),
    .ZN(_13434_));
 NAND2_X1 _19375_ (.A1(_13240_),
    .A2(_13245_),
    .ZN(_13435_));
 AND2_X2 _19376_ (.A1(_13059_),
    .A2(_13063_),
    .ZN(_13436_));
 OAI21_X4 _19377_ (.A(_13434_),
    .B1(_13435_),
    .B2(_13436_),
    .ZN(_13437_));
 NAND2_X2 _19378_ (.A1(_13429_),
    .A2(_13437_),
    .ZN(_13438_));
 AND3_X2 _19379_ (.A1(_13240_),
    .A2(_13066_),
    .A3(_13245_),
    .ZN(_13439_));
 NAND2_X4 _19380_ (.A1(_13429_),
    .A2(_13439_),
    .ZN(_13440_));
 OAI21_X4 _19381_ (.A(_13438_),
    .B1(_12342_),
    .B2(_13440_),
    .ZN(_13441_));
 OR2_X1 _19382_ (.A1(_13429_),
    .A2(_13437_),
    .ZN(_13442_));
 AOI21_X2 _19383_ (.A(_13442_),
    .B1(_13439_),
    .B2(_12714_),
    .ZN(_13443_));
 NOR2_X4 _19384_ (.A1(_13441_),
    .A2(_13443_),
    .ZN(\alu_adder_result_ex[22] ));
 AOI21_X1 _19385_ (.A(_13073_),
    .B1(_13075_),
    .B2(_12419_),
    .ZN(_13444_));
 MUX2_X1 _19386_ (.A(_00916_),
    .B(_00918_),
    .S(_12736_),
    .Z(_13445_));
 NOR2_X1 _19387_ (.A1(_12361_),
    .A2(_13445_),
    .ZN(_13446_));
 MUX2_X1 _19388_ (.A(_00917_),
    .B(_00919_),
    .S(_13079_),
    .Z(_13447_));
 NOR2_X1 _19389_ (.A1(_12367_),
    .A2(_13447_),
    .ZN(_13448_));
 NOR3_X1 _19390_ (.A1(_12409_),
    .A2(_13446_),
    .A3(_13448_),
    .ZN(_13449_));
 INV_X1 _19391_ (.A(_00910_),
    .ZN(_13450_));
 NOR2_X1 _19392_ (.A1(_12398_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .ZN(_13451_));
 AOI21_X1 _19393_ (.A(_13451_),
    .B1(_00911_),
    .B2(_12547_),
    .ZN(_13452_));
 AOI221_X2 _19394_ (.A(_10758_),
    .B1(_13450_),
    .B2(_12373_),
    .C1(_13452_),
    .C2(_12555_),
    .ZN(_13453_));
 NOR3_X2 _19395_ (.A1(_12423_),
    .A2(_13449_),
    .A3(_13453_),
    .ZN(_13454_));
 MUX2_X1 _19396_ (.A(_00920_),
    .B(_00922_),
    .S(_12400_),
    .Z(_13455_));
 MUX2_X1 _19397_ (.A(_00921_),
    .B(_00923_),
    .S(_13170_),
    .Z(_13456_));
 MUX2_X1 _19398_ (.A(_13455_),
    .B(_13456_),
    .S(_13092_),
    .Z(_13457_));
 MUX2_X1 _19399_ (.A(_00912_),
    .B(_00914_),
    .S(_13170_),
    .Z(_13458_));
 MUX2_X1 _19400_ (.A(_00913_),
    .B(_00915_),
    .S(_12919_),
    .Z(_13459_));
 MUX2_X1 _19401_ (.A(_13458_),
    .B(_13459_),
    .S(_13281_),
    .Z(_13460_));
 MUX2_X1 _19402_ (.A(_13457_),
    .B(_13460_),
    .S(_12408_),
    .Z(_13461_));
 NOR2_X1 _19403_ (.A1(_12807_),
    .A2(_13461_),
    .ZN(_13462_));
 NOR3_X4 _19404_ (.A1(_12354_),
    .A2(_13454_),
    .A3(_13462_),
    .ZN(_13463_));
 MUX2_X1 _19405_ (.A(_00932_),
    .B(_00934_),
    .S(_12385_),
    .Z(_13464_));
 MUX2_X1 _19406_ (.A(_00933_),
    .B(_00935_),
    .S(_13180_),
    .Z(_13465_));
 MUX2_X1 _19407_ (.A(_13464_),
    .B(_13465_),
    .S(_12392_),
    .Z(_13466_));
 MUX2_X1 _19408_ (.A(_00924_),
    .B(_00926_),
    .S(_13180_),
    .Z(_13467_));
 MUX2_X1 _19409_ (.A(_00925_),
    .B(_00927_),
    .S(net344),
    .Z(_13468_));
 MUX2_X1 _19410_ (.A(_13467_),
    .B(_13468_),
    .S(_12392_),
    .Z(_13469_));
 MUX2_X1 _19411_ (.A(_13466_),
    .B(_13469_),
    .S(_12394_),
    .Z(_13470_));
 MUX2_X1 _19412_ (.A(_00936_),
    .B(_00938_),
    .S(_13180_),
    .Z(_13471_));
 BUF_X4 _19413_ (.A(net374),
    .Z(_13472_));
 MUX2_X1 _19414_ (.A(_00937_),
    .B(_00939_),
    .S(_13472_),
    .Z(_13473_));
 MUX2_X1 _19415_ (.A(_13471_),
    .B(_13473_),
    .S(_13194_),
    .Z(_13474_));
 MUX2_X1 _19416_ (.A(_00928_),
    .B(_00930_),
    .S(net344),
    .Z(_13475_));
 MUX2_X1 _19417_ (.A(_00929_),
    .B(_00931_),
    .S(_13192_),
    .Z(_13476_));
 MUX2_X1 _19418_ (.A(_13475_),
    .B(_13476_),
    .S(_13194_),
    .Z(_13477_));
 MUX2_X1 _19419_ (.A(_13474_),
    .B(_13477_),
    .S(_13297_),
    .Z(_13478_));
 MUX2_X1 _19420_ (.A(_13470_),
    .B(_13478_),
    .S(_13115_),
    .Z(_13479_));
 AOI21_X4 _19421_ (.A(_13463_),
    .B1(_13117_),
    .B2(_13479_),
    .ZN(_13480_));
 OAI21_X1 _19422_ (.A(_13077_),
    .B1(_13078_),
    .B2(_13480_),
    .ZN(_13481_));
 OR2_X1 _19423_ (.A1(_13444_),
    .A2(_13481_),
    .ZN(_16434_));
 INV_X1 _19424_ (.A(_16434_),
    .ZN(_16430_));
 NAND2_X1 _19425_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(_11221_),
    .ZN(_13482_));
 MUX2_X1 _19426_ (.A(_00932_),
    .B(_00934_),
    .S(_13318_),
    .Z(_13483_));
 MUX2_X1 _19427_ (.A(_00933_),
    .B(_00935_),
    .S(_13318_),
    .Z(_13484_));
 MUX2_X1 _19428_ (.A(_13483_),
    .B(_13484_),
    .S(_11256_),
    .Z(_13485_));
 MUX2_X1 _19429_ (.A(_00924_),
    .B(_00926_),
    .S(_12200_),
    .Z(_13486_));
 MUX2_X1 _19430_ (.A(_00925_),
    .B(_00927_),
    .S(_12200_),
    .Z(_13487_));
 MUX2_X1 _19431_ (.A(_13486_),
    .B(_13487_),
    .S(_11256_),
    .Z(_13488_));
 MUX2_X1 _19432_ (.A(_13485_),
    .B(_13488_),
    .S(_11232_),
    .Z(_13489_));
 NOR2_X2 _19433_ (.A1(_11058_),
    .A2(_13489_),
    .ZN(_13490_));
 MUX2_X1 _19434_ (.A(_00936_),
    .B(_00938_),
    .S(_11065_),
    .Z(_13491_));
 MUX2_X1 _19435_ (.A(_00937_),
    .B(_00939_),
    .S(_11065_),
    .Z(_13492_));
 MUX2_X1 _19436_ (.A(_13491_),
    .B(_13492_),
    .S(_11227_),
    .Z(_13493_));
 MUX2_X1 _19437_ (.A(_00928_),
    .B(_00930_),
    .S(_11065_),
    .Z(_13494_));
 MUX2_X1 _19438_ (.A(_00929_),
    .B(_00931_),
    .S(_11065_),
    .Z(_13495_));
 MUX2_X1 _19439_ (.A(_13494_),
    .B(_13495_),
    .S(_11227_),
    .Z(_13496_));
 MUX2_X1 _19440_ (.A(_13493_),
    .B(_13496_),
    .S(_11232_),
    .Z(_13497_));
 NOR2_X1 _19441_ (.A1(_11223_),
    .A2(_13497_),
    .ZN(_13498_));
 NOR3_X4 _19442_ (.A1(_10981_),
    .A2(_13490_),
    .A3(_13498_),
    .ZN(_13499_));
 MUX2_X1 _19443_ (.A(_00916_),
    .B(_00918_),
    .S(_11006_),
    .Z(_13500_));
 NOR2_X1 _19444_ (.A1(_11805_),
    .A2(_13500_),
    .ZN(_13501_));
 MUX2_X1 _19445_ (.A(_00917_),
    .B(_00919_),
    .S(_11015_),
    .Z(_13502_));
 NOR2_X1 _19446_ (.A1(_11012_),
    .A2(_13502_),
    .ZN(_13503_));
 NOR3_X1 _19447_ (.A1(_12117_),
    .A2(_13501_),
    .A3(_13503_),
    .ZN(_13504_));
 NOR2_X1 _19448_ (.A1(_11096_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .ZN(_13505_));
 AOI21_X1 _19449_ (.A(_13505_),
    .B1(_00911_),
    .B2(_11208_),
    .ZN(_13506_));
 AOI221_X2 _19450_ (.A(_11021_),
    .B1(_13450_),
    .B2(_11031_),
    .C1(_13506_),
    .C2(_11260_),
    .ZN(_13507_));
 NOR3_X2 _19451_ (.A1(_10987_),
    .A2(_13504_),
    .A3(_13507_),
    .ZN(_13508_));
 MUX2_X1 _19452_ (.A(_00920_),
    .B(_00922_),
    .S(_12061_),
    .Z(_13509_));
 MUX2_X1 _19453_ (.A(_00921_),
    .B(_00923_),
    .S(_12061_),
    .Z(_13510_));
 MUX2_X1 _19454_ (.A(_13509_),
    .B(_13510_),
    .S(_11026_),
    .Z(_13511_));
 MUX2_X1 _19455_ (.A(_00912_),
    .B(_00914_),
    .S(_11005_),
    .Z(_13512_));
 MUX2_X1 _19456_ (.A(_00913_),
    .B(_00915_),
    .S(_11005_),
    .Z(_13513_));
 MUX2_X1 _19457_ (.A(_13512_),
    .B(_13513_),
    .S(_11026_),
    .Z(_13514_));
 MUX2_X1 _19458_ (.A(_13511_),
    .B(_13514_),
    .S(_12068_),
    .Z(_13515_));
 NOR2_X2 _19459_ (.A1(_11223_),
    .A2(_13515_),
    .ZN(_13516_));
 NOR3_X4 _19460_ (.A1(_11052_),
    .A2(_13508_),
    .A3(_13516_),
    .ZN(_13517_));
 OR2_X4 _19461_ (.A1(_13499_),
    .A2(_13517_),
    .ZN(_13518_));
 NAND2_X1 _19462_ (.A1(\cs_registers_i.pc_id_i[24] ),
    .A2(_11112_),
    .ZN(_13519_));
 OAI221_X2 _19463_ (.A(_13482_),
    .B1(_13518_),
    .B2(_11278_),
    .C1(_13519_),
    .C2(_11114_),
    .ZN(_16429_));
 INV_X2 _19464_ (.A(_16429_),
    .ZN(_16433_));
 AOI21_X1 _19465_ (.A(_13073_),
    .B1(_13075_),
    .B2(_10945_),
    .ZN(_13520_));
 MUX2_X1 _19466_ (.A(_00963_),
    .B(_00965_),
    .S(_12454_),
    .Z(_13521_));
 MUX2_X1 _19467_ (.A(_00964_),
    .B(_00966_),
    .S(_12454_),
    .Z(_13522_));
 MUX2_X1 _19468_ (.A(_13521_),
    .B(_13522_),
    .S(_12380_),
    .Z(_13523_));
 MUX2_X1 _19469_ (.A(_00955_),
    .B(_00957_),
    .S(_12454_),
    .Z(_13524_));
 MUX2_X1 _19470_ (.A(_00956_),
    .B(_00958_),
    .S(_12454_),
    .Z(_13525_));
 MUX2_X1 _19471_ (.A(_13524_),
    .B(_13525_),
    .S(_12380_),
    .Z(_13526_));
 MUX2_X1 _19472_ (.A(_13523_),
    .B(_13526_),
    .S(_12357_),
    .Z(_13527_));
 NOR2_X1 _19473_ (.A1(_12356_),
    .A2(_13527_),
    .ZN(_13528_));
 MUX2_X1 _19474_ (.A(_00967_),
    .B(_00969_),
    .S(_12563_),
    .Z(_13529_));
 MUX2_X1 _19475_ (.A(_00968_),
    .B(_00970_),
    .S(_12563_),
    .Z(_13530_));
 MUX2_X1 _19476_ (.A(_13529_),
    .B(_13530_),
    .S(_12380_),
    .Z(_13531_));
 MUX2_X1 _19477_ (.A(_00959_),
    .B(_00961_),
    .S(_12563_),
    .Z(_13532_));
 MUX2_X1 _19478_ (.A(_00960_),
    .B(_00962_),
    .S(_12563_),
    .Z(_13533_));
 MUX2_X1 _19479_ (.A(_13532_),
    .B(_13533_),
    .S(_12380_),
    .Z(_13534_));
 MUX2_X1 _19480_ (.A(_13531_),
    .B(_13534_),
    .S(_12357_),
    .Z(_13535_));
 NOR2_X1 _19481_ (.A1(_12807_),
    .A2(_13535_),
    .ZN(_13536_));
 NOR3_X2 _19482_ (.A1(_10764_),
    .A2(_13528_),
    .A3(_13536_),
    .ZN(_13537_));
 MUX2_X1 _19483_ (.A(_00951_),
    .B(_00953_),
    .S(_13101_),
    .Z(_13538_));
 MUX2_X1 _19484_ (.A(_00952_),
    .B(_00954_),
    .S(_13101_),
    .Z(_13539_));
 MUX2_X1 _19485_ (.A(_13538_),
    .B(_13539_),
    .S(_12388_),
    .Z(_13540_));
 MUX2_X1 _19486_ (.A(_00943_),
    .B(_00945_),
    .S(_13101_),
    .Z(_13541_));
 MUX2_X1 _19487_ (.A(_00944_),
    .B(_00946_),
    .S(_12385_),
    .Z(_13542_));
 MUX2_X1 _19488_ (.A(_13541_),
    .B(_13542_),
    .S(_12388_),
    .Z(_13543_));
 MUX2_X1 _19489_ (.A(_13540_),
    .B(_13543_),
    .S(_12394_),
    .Z(_13544_));
 NOR2_X1 _19490_ (.A1(_12384_),
    .A2(_13544_),
    .ZN(_13545_));
 INV_X1 _19491_ (.A(_00941_),
    .ZN(_13546_));
 NOR2_X1 _19492_ (.A1(_12364_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .ZN(_13547_));
 AOI21_X1 _19493_ (.A(_13547_),
    .B1(_00942_),
    .B2(_12438_),
    .ZN(_13548_));
 AOI221_X2 _19494_ (.A(_12372_),
    .B1(_13546_),
    .B2(_12374_),
    .C1(_13548_),
    .C2(_12440_),
    .ZN(_13549_));
 MUX2_X1 _19495_ (.A(_00947_),
    .B(_00949_),
    .S(_12378_),
    .Z(_13550_));
 MUX2_X1 _19496_ (.A(_00948_),
    .B(_00950_),
    .S(_12378_),
    .Z(_13551_));
 MUX2_X1 _19497_ (.A(_13550_),
    .B(_13551_),
    .S(_12426_),
    .Z(_13552_));
 AOI21_X2 _19498_ (.A(_13549_),
    .B1(_13552_),
    .B2(_12432_),
    .ZN(_13553_));
 AOI21_X4 _19499_ (.A(_13545_),
    .B1(_13553_),
    .B2(_12384_),
    .ZN(_13554_));
 AOI21_X4 _19500_ (.A(_13537_),
    .B1(_13554_),
    .B2(_10764_),
    .ZN(_13555_));
 OAI21_X1 _19501_ (.A(_13077_),
    .B1(_13078_),
    .B2(_13555_),
    .ZN(_13556_));
 OR2_X2 _19502_ (.A1(_13520_),
    .A2(_13556_),
    .ZN(_16442_));
 INV_X1 _19503_ (.A(_16442_),
    .ZN(_16438_));
 NAND2_X1 _19504_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(_10958_),
    .ZN(_13557_));
 MUX2_X1 _19505_ (.A(_00963_),
    .B(_00965_),
    .S(_11005_),
    .Z(_13558_));
 MUX2_X1 _19506_ (.A(_00964_),
    .B(_00966_),
    .S(_11005_),
    .Z(_13559_));
 MUX2_X1 _19507_ (.A(_13558_),
    .B(_13559_),
    .S(_12037_),
    .Z(_13560_));
 MUX2_X1 _19508_ (.A(_00955_),
    .B(_00957_),
    .S(_11005_),
    .Z(_13561_));
 MUX2_X1 _19509_ (.A(_00956_),
    .B(_00958_),
    .S(_11005_),
    .Z(_13562_));
 MUX2_X1 _19510_ (.A(_13561_),
    .B(_13562_),
    .S(_12037_),
    .Z(_13563_));
 MUX2_X1 _19511_ (.A(_13560_),
    .B(_13563_),
    .S(_12068_),
    .Z(_13564_));
 NOR2_X1 _19512_ (.A1(_11058_),
    .A2(_13564_),
    .ZN(_13565_));
 MUX2_X1 _19513_ (.A(_00967_),
    .B(_00969_),
    .S(_12085_),
    .Z(_13566_));
 MUX2_X1 _19514_ (.A(_00968_),
    .B(_00970_),
    .S(_12061_),
    .Z(_13567_));
 MUX2_X1 _19515_ (.A(_13566_),
    .B(_13567_),
    .S(_11026_),
    .Z(_13568_));
 MUX2_X1 _19516_ (.A(_00959_),
    .B(_00961_),
    .S(_12061_),
    .Z(_13569_));
 MUX2_X1 _19517_ (.A(_00960_),
    .B(_00962_),
    .S(_12061_),
    .Z(_13570_));
 MUX2_X1 _19518_ (.A(_13569_),
    .B(_13570_),
    .S(_11026_),
    .Z(_13571_));
 MUX2_X1 _19519_ (.A(_13568_),
    .B(_13571_),
    .S(_12068_),
    .Z(_13572_));
 NOR2_X1 _19520_ (.A1(_11073_),
    .A2(_13572_),
    .ZN(_13573_));
 NOR3_X4 _19521_ (.A1(_10981_),
    .A2(_13565_),
    .A3(_13573_),
    .ZN(_13574_));
 MUX2_X1 _19522_ (.A(_00947_),
    .B(_00949_),
    .S(_11015_),
    .Z(_13575_));
 NOR2_X1 _19523_ (.A1(_11000_),
    .A2(_13575_),
    .ZN(_13576_));
 MUX2_X1 _19524_ (.A(_00948_),
    .B(_00950_),
    .S(_11015_),
    .Z(_13577_));
 NOR2_X1 _19525_ (.A1(_11012_),
    .A2(_13577_),
    .ZN(_13578_));
 NOR3_X1 _19526_ (.A1(_10993_),
    .A2(_13576_),
    .A3(_13578_),
    .ZN(_13579_));
 NOR2_X1 _19527_ (.A1(_11240_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .ZN(_13580_));
 AOI21_X1 _19528_ (.A(_13580_),
    .B1(_00942_),
    .B2(_11850_),
    .ZN(_13581_));
 AOI221_X2 _19529_ (.A(_11021_),
    .B1(_13546_),
    .B2(_11031_),
    .C1(_13581_),
    .C2(_11074_),
    .ZN(_13582_));
 NOR3_X2 _19530_ (.A1(_10987_),
    .A2(_13579_),
    .A3(_13582_),
    .ZN(_13583_));
 MUX2_X1 _19531_ (.A(_00951_),
    .B(_00953_),
    .S(_11014_),
    .Z(_13584_));
 MUX2_X1 _19532_ (.A(_00952_),
    .B(_00954_),
    .S(_11014_),
    .Z(_13585_));
 MUX2_X1 _19533_ (.A(_13584_),
    .B(_13585_),
    .S(_11041_),
    .Z(_13586_));
 MUX2_X1 _19534_ (.A(_00943_),
    .B(_00945_),
    .S(_11014_),
    .Z(_13587_));
 MUX2_X1 _19535_ (.A(_00944_),
    .B(_00946_),
    .S(_11014_),
    .Z(_13588_));
 MUX2_X1 _19536_ (.A(_13587_),
    .B(_13588_),
    .S(_11041_),
    .Z(_13589_));
 MUX2_X1 _19537_ (.A(_13586_),
    .B(_13589_),
    .S(_12068_),
    .Z(_13590_));
 NOR2_X2 _19538_ (.A1(_11073_),
    .A2(_13590_),
    .ZN(_13591_));
 NOR3_X4 _19539_ (.A1(_11052_),
    .A2(_13583_),
    .A3(_13591_),
    .ZN(_13592_));
 OR2_X2 _19540_ (.A1(_13574_),
    .A2(_13592_),
    .ZN(_13593_));
 NAND2_X1 _19541_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(_11112_),
    .ZN(_13594_));
 OAI221_X1 _19542_ (.A(_13557_),
    .B1(_13593_),
    .B2(_11277_),
    .C1(_13594_),
    .C2(_11114_),
    .ZN(_13595_));
 CLKBUF_X3 _19543_ (.A(_13595_),
    .Z(_16437_));
 INV_X1 _19544_ (.A(_16437_),
    .ZN(_16441_));
 BUF_X2 _19545_ (.A(_15863_),
    .Z(_13596_));
 AOI21_X2 _19546_ (.A(_15867_),
    .B1(_13596_),
    .B2(_15868_),
    .ZN(_13597_));
 NAND2_X1 _19547_ (.A1(_15864_),
    .A2(_15868_),
    .ZN(_13598_));
 NOR2_X1 _19548_ (.A1(_13429_),
    .A2(_13427_),
    .ZN(_13599_));
 OAI21_X2 _19549_ (.A(_13597_),
    .B1(_13598_),
    .B2(_13599_),
    .ZN(_13600_));
 NOR2_X1 _19550_ (.A1(_15855_),
    .A2(_13427_),
    .ZN(_13601_));
 NAND2_X1 _19551_ (.A1(_13597_),
    .A2(_13601_),
    .ZN(_13602_));
 OAI21_X4 _19552_ (.A(_13600_),
    .B1(_13602_),
    .B2(_13251_),
    .ZN(_13603_));
 XNOR2_X2 _19553_ (.A(_13603_),
    .B(_15872_),
    .ZN(\alu_adder_result_ex[25] ));
 INV_X2 _19554_ (.A(_15868_),
    .ZN(_13604_));
 NOR3_X1 _19555_ (.A1(_13604_),
    .A2(_13427_),
    .A3(_13596_),
    .ZN(_13605_));
 OAI211_X2 _19556_ (.A(_13438_),
    .B(_13605_),
    .C1(_13440_),
    .C2(_12342_),
    .ZN(_13606_));
 NOR3_X1 _19557_ (.A1(_15864_),
    .A2(_13604_),
    .A3(_13596_),
    .ZN(_13607_));
 AND2_X1 _19558_ (.A1(_15864_),
    .A2(_13604_),
    .ZN(_13608_));
 AOI221_X2 _19559_ (.A(_13607_),
    .B1(_13608_),
    .B2(_13427_),
    .C1(_13604_),
    .C2(_13596_),
    .ZN(_13609_));
 NAND2_X1 _19560_ (.A1(_15864_),
    .A2(_13604_),
    .ZN(_13610_));
 INV_X1 _19561_ (.A(_13440_),
    .ZN(_13611_));
 AOI22_X4 _19562_ (.A1(_13429_),
    .A2(_13437_),
    .B1(_12714_),
    .B2(_13611_),
    .ZN(_13612_));
 OAI211_X4 _19563_ (.A(_13606_),
    .B(_13609_),
    .C1(_13610_),
    .C2(_13612_),
    .ZN(\alu_adder_result_ex[24] ));
 AOI21_X1 _19564_ (.A(_13073_),
    .B1(_13075_),
    .B2(_10869_),
    .ZN(_13613_));
 MUX2_X1 _19565_ (.A(_00978_),
    .B(_00980_),
    .S(_12736_),
    .Z(_13614_));
 NOR2_X1 _19566_ (.A1(_12361_),
    .A2(_13614_),
    .ZN(_13615_));
 MUX2_X1 _19567_ (.A(_00979_),
    .B(_00981_),
    .S(_13079_),
    .Z(_13616_));
 NOR2_X1 _19568_ (.A1(_12367_),
    .A2(_13616_),
    .ZN(_13617_));
 NOR3_X1 _19569_ (.A1(_12409_),
    .A2(_13615_),
    .A3(_13617_),
    .ZN(_13618_));
 INV_X1 _19570_ (.A(_00972_),
    .ZN(_13619_));
 NOR2_X1 _19571_ (.A1(_12401_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .ZN(_13620_));
 AOI21_X1 _19572_ (.A(_13620_),
    .B1(_00973_),
    .B2(_12547_),
    .ZN(_13621_));
 AOI221_X1 _19573_ (.A(_12372_),
    .B1(_13619_),
    .B2(_12373_),
    .C1(_13621_),
    .C2(_12445_),
    .ZN(_13622_));
 NOR3_X1 _19574_ (.A1(_12423_),
    .A2(_13618_),
    .A3(_13622_),
    .ZN(_13623_));
 MUX2_X1 _19575_ (.A(_00982_),
    .B(_00984_),
    .S(_13170_),
    .Z(_13624_));
 MUX2_X1 _19576_ (.A(_00983_),
    .B(_00985_),
    .S(_13170_),
    .Z(_13625_));
 MUX2_X1 _19577_ (.A(_13624_),
    .B(_13625_),
    .S(_13092_),
    .Z(_13626_));
 MUX2_X1 _19578_ (.A(_00974_),
    .B(_00976_),
    .S(_12919_),
    .Z(_13627_));
 MUX2_X1 _19579_ (.A(_00975_),
    .B(_00977_),
    .S(_12919_),
    .Z(_13628_));
 MUX2_X1 _19580_ (.A(_13627_),
    .B(_13628_),
    .S(_13281_),
    .Z(_13629_));
 MUX2_X1 _19581_ (.A(_13626_),
    .B(_13629_),
    .S(_12408_),
    .Z(_13630_));
 NOR2_X1 _19582_ (.A1(_12807_),
    .A2(_13630_),
    .ZN(_13631_));
 NOR3_X2 _19583_ (.A1(_12354_),
    .A2(_13623_),
    .A3(_13631_),
    .ZN(_13632_));
 MUX2_X1 _19584_ (.A(_00994_),
    .B(_00996_),
    .S(_12385_),
    .Z(_13633_));
 MUX2_X1 _19585_ (.A(_00995_),
    .B(_00997_),
    .S(_13184_),
    .Z(_13634_));
 MUX2_X1 _19586_ (.A(_13633_),
    .B(_13634_),
    .S(_12392_),
    .Z(_13635_));
 MUX2_X1 _19587_ (.A(_00986_),
    .B(_00988_),
    .S(_13184_),
    .Z(_13636_));
 MUX2_X1 _19588_ (.A(_00987_),
    .B(_00989_),
    .S(_13472_),
    .Z(_13637_));
 MUX2_X1 _19589_ (.A(_13636_),
    .B(_13637_),
    .S(_13194_),
    .Z(_13638_));
 MUX2_X1 _19590_ (.A(_13635_),
    .B(_13638_),
    .S(_12394_),
    .Z(_13639_));
 MUX2_X1 _19591_ (.A(_00998_),
    .B(_01000_),
    .S(net344),
    .Z(_13640_));
 MUX2_X1 _19592_ (.A(_00999_),
    .B(_01001_),
    .S(_13192_),
    .Z(_13641_));
 MUX2_X1 _19593_ (.A(_13640_),
    .B(_13641_),
    .S(_13194_),
    .Z(_13642_));
 MUX2_X1 _19594_ (.A(_00990_),
    .B(_00992_),
    .S(_13472_),
    .Z(_13643_));
 MUX2_X1 _19595_ (.A(_00991_),
    .B(_00993_),
    .S(_13289_),
    .Z(_13644_));
 MUX2_X1 _19596_ (.A(_13643_),
    .B(_13644_),
    .S(_12360_),
    .Z(_13645_));
 MUX2_X1 _19597_ (.A(_13642_),
    .B(_13645_),
    .S(_13297_),
    .Z(_13646_));
 MUX2_X1 _19598_ (.A(_13639_),
    .B(_13646_),
    .S(_13115_),
    .Z(_13647_));
 AOI21_X4 _19599_ (.A(_13632_),
    .B1(_13647_),
    .B2(_13117_),
    .ZN(_13648_));
 OAI21_X1 _19600_ (.A(_13077_),
    .B1(_13078_),
    .B2(_13648_),
    .ZN(_13649_));
 OR2_X1 _19601_ (.A1(_13613_),
    .A2(_13649_),
    .ZN(_16450_));
 INV_X1 _19602_ (.A(_16450_),
    .ZN(_16446_));
 MUX2_X1 _19603_ (.A(_00978_),
    .B(_00980_),
    .S(_11097_),
    .Z(_13650_));
 NOR2_X1 _19604_ (.A1(_11028_),
    .A2(_13650_),
    .ZN(_13651_));
 MUX2_X1 _19605_ (.A(_00979_),
    .B(_00981_),
    .S(_11241_),
    .Z(_13652_));
 NOR2_X1 _19606_ (.A1(_11013_),
    .A2(_13652_),
    .ZN(_13653_));
 NOR3_X1 _19607_ (.A1(_10994_),
    .A2(_13651_),
    .A3(_13653_),
    .ZN(_13654_));
 NOR2_X1 _19608_ (.A1(_11246_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .ZN(_13655_));
 AOI21_X1 _19609_ (.A(_13655_),
    .B1(_00973_),
    .B2(_11007_),
    .ZN(_13656_));
 AOI221_X2 _19610_ (.A(_11022_),
    .B1(_13619_),
    .B2(_11032_),
    .C1(_13656_),
    .C2(_11805_),
    .ZN(_13657_));
 NOR3_X1 _19611_ (.A1(_10988_),
    .A2(_13654_),
    .A3(_13657_),
    .ZN(_13658_));
 MUX2_X1 _19612_ (.A(_00982_),
    .B(_00984_),
    .S(_12666_),
    .Z(_13659_));
 MUX2_X1 _19613_ (.A(_00983_),
    .B(_00985_),
    .S(_12666_),
    .Z(_13660_));
 MUX2_X1 _19614_ (.A(_13659_),
    .B(_13660_),
    .S(_11060_),
    .Z(_13661_));
 MUX2_X1 _19615_ (.A(_00974_),
    .B(_00976_),
    .S(_12666_),
    .Z(_13662_));
 MUX2_X1 _19616_ (.A(_00975_),
    .B(_00977_),
    .S(_11783_),
    .Z(_13663_));
 MUX2_X1 _19617_ (.A(_13662_),
    .B(_13663_),
    .S(_11060_),
    .Z(_13664_));
 MUX2_X1 _19618_ (.A(_13661_),
    .B(_13664_),
    .S(_10993_),
    .Z(_13665_));
 NOR2_X1 _19619_ (.A1(_11174_),
    .A2(_13665_),
    .ZN(_13666_));
 OAI21_X2 _19620_ (.A(_10982_),
    .B1(_13658_),
    .B2(_13666_),
    .ZN(_13667_));
 MUX2_X1 _19621_ (.A(_00990_),
    .B(_00992_),
    .S(_11208_),
    .Z(_13668_));
 MUX2_X1 _19622_ (.A(_00991_),
    .B(_00993_),
    .S(_11208_),
    .Z(_13669_));
 MUX2_X1 _19623_ (.A(_13668_),
    .B(_13669_),
    .S(_11093_),
    .Z(_13670_));
 MUX2_X1 _19624_ (.A(_00986_),
    .B(_00987_),
    .S(_11269_),
    .Z(_13671_));
 MUX2_X1 _19625_ (.A(_00988_),
    .B(_00989_),
    .S(_11027_),
    .Z(_13672_));
 AOI222_X2 _19626_ (.A1(_11085_),
    .A2(_13670_),
    .B1(_13671_),
    .B2(_11091_),
    .C1(_13672_),
    .C2(_11100_),
    .ZN(_13673_));
 NAND2_X1 _19627_ (.A1(_11053_),
    .A2(_13673_),
    .ZN(_13674_));
 MUX2_X1 _19628_ (.A(_01000_),
    .B(_01001_),
    .S(_11025_),
    .Z(_13675_));
 AOI21_X1 _19629_ (.A(_11036_),
    .B1(_13675_),
    .B2(_11007_),
    .ZN(_13676_));
 MUX2_X1 _19630_ (.A(_00996_),
    .B(_00997_),
    .S(_11025_),
    .Z(_13677_));
 AOI21_X1 _19631_ (.A(_10986_),
    .B1(_13677_),
    .B2(_11241_),
    .ZN(_13678_));
 OAI21_X1 _19632_ (.A(_11069_),
    .B1(_13676_),
    .B2(_13678_),
    .ZN(_13679_));
 MUX2_X1 _19633_ (.A(_00994_),
    .B(_00995_),
    .S(_10998_),
    .Z(_13680_));
 INV_X1 _19634_ (.A(_13680_),
    .ZN(_13681_));
 MUX2_X1 _19635_ (.A(_00998_),
    .B(_00999_),
    .S(_11059_),
    .Z(_13682_));
 INV_X1 _19636_ (.A(_13682_),
    .ZN(_13683_));
 AOI221_X1 _19637_ (.A(_11232_),
    .B1(_13678_),
    .B2(_13681_),
    .C1(_13683_),
    .C2(_13676_),
    .ZN(_13684_));
 AND2_X1 _19638_ (.A1(_13679_),
    .A2(_13684_),
    .ZN(_13685_));
 OAI21_X4 _19639_ (.A(_13667_),
    .B1(_13674_),
    .B2(_13685_),
    .ZN(_13686_));
 NAND2_X1 _19640_ (.A1(_11973_),
    .A2(_13686_),
    .ZN(_13687_));
 BUF_X2 _19641_ (.A(\cs_registers_i.pc_id_i[26] ),
    .Z(_13688_));
 NAND2_X1 _19642_ (.A1(_13688_),
    .A2(_11112_),
    .ZN(_13689_));
 INV_X1 _19643_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .ZN(_13690_));
 OAI221_X2 _19644_ (.A(_13687_),
    .B1(_13689_),
    .B2(_11114_),
    .C1(_10838_),
    .C2(_13690_),
    .ZN(_16445_));
 INV_X2 _19645_ (.A(_16445_),
    .ZN(_16449_));
 AOI21_X1 _19646_ (.A(_13073_),
    .B1(_13075_),
    .B2(_10873_),
    .ZN(_13691_));
 MUX2_X1 _19647_ (.A(_01009_),
    .B(_01011_),
    .S(_12736_),
    .Z(_13692_));
 NOR2_X1 _19648_ (.A1(_12361_),
    .A2(_13692_),
    .ZN(_13693_));
 MUX2_X1 _19649_ (.A(_01010_),
    .B(_01012_),
    .S(_12920_),
    .Z(_13694_));
 NOR2_X1 _19650_ (.A1(_12367_),
    .A2(_13694_),
    .ZN(_13695_));
 NOR3_X1 _19651_ (.A1(_12409_),
    .A2(_13693_),
    .A3(_13695_),
    .ZN(_13696_));
 INV_X1 _19652_ (.A(_01003_),
    .ZN(_13697_));
 NOR2_X1 _19653_ (.A1(_12401_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .ZN(_13698_));
 AOI21_X1 _19654_ (.A(_13698_),
    .B1(_01004_),
    .B2(_12547_),
    .ZN(_13699_));
 AOI221_X2 _19655_ (.A(_12372_),
    .B1(_13697_),
    .B2(_12373_),
    .C1(_13699_),
    .C2(_12445_),
    .ZN(_13700_));
 NOR3_X2 _19656_ (.A1(_12423_),
    .A2(_13696_),
    .A3(_13700_),
    .ZN(_13701_));
 MUX2_X1 _19657_ (.A(_01013_),
    .B(_01015_),
    .S(_13278_),
    .Z(_13702_));
 MUX2_X1 _19658_ (.A(_01014_),
    .B(_01016_),
    .S(_13278_),
    .Z(_13703_));
 MUX2_X1 _19659_ (.A(_13702_),
    .B(_13703_),
    .S(_13281_),
    .Z(_13704_));
 MUX2_X1 _19660_ (.A(_01005_),
    .B(_01007_),
    .S(_13278_),
    .Z(_13705_));
 MUX2_X1 _19661_ (.A(_01006_),
    .B(_01008_),
    .S(_12563_),
    .Z(_13706_));
 MUX2_X1 _19662_ (.A(_13705_),
    .B(_13706_),
    .S(_13281_),
    .Z(_13707_));
 MUX2_X1 _19663_ (.A(_13704_),
    .B(_13707_),
    .S(_12357_),
    .Z(_13708_));
 NOR2_X1 _19664_ (.A1(_12807_),
    .A2(_13708_),
    .ZN(_13709_));
 NOR3_X4 _19665_ (.A1(_12354_),
    .A2(_13701_),
    .A3(_13709_),
    .ZN(_13710_));
 MUX2_X1 _19666_ (.A(_01025_),
    .B(_01027_),
    .S(_13289_),
    .Z(_13711_));
 MUX2_X1 _19667_ (.A(_01026_),
    .B(_01028_),
    .S(_13289_),
    .Z(_13712_));
 MUX2_X1 _19668_ (.A(_13711_),
    .B(_13712_),
    .S(_12360_),
    .Z(_13713_));
 MUX2_X1 _19669_ (.A(_01017_),
    .B(_01019_),
    .S(_13289_),
    .Z(_13714_));
 MUX2_X1 _19670_ (.A(_01018_),
    .B(_01020_),
    .S(_13291_),
    .Z(_13715_));
 MUX2_X1 _19671_ (.A(_13714_),
    .B(_13715_),
    .S(_12360_),
    .Z(_13716_));
 MUX2_X1 _19672_ (.A(_13713_),
    .B(_13716_),
    .S(_13297_),
    .Z(_03095_));
 MUX2_X1 _19673_ (.A(_01029_),
    .B(_01031_),
    .S(_13291_),
    .Z(_03096_));
 MUX2_X1 _19674_ (.A(_01030_),
    .B(_01032_),
    .S(_13291_),
    .Z(_03097_));
 MUX2_X1 _19675_ (.A(_03096_),
    .B(_03097_),
    .S(_12911_),
    .Z(_03098_));
 MUX2_X1 _19676_ (.A(_01021_),
    .B(_01023_),
    .S(_13291_),
    .Z(_03099_));
 MUX2_X1 _19677_ (.A(_01022_),
    .B(_01024_),
    .S(_12434_),
    .Z(_03100_));
 MUX2_X1 _19678_ (.A(_03099_),
    .B(_03100_),
    .S(_12911_),
    .Z(_03101_));
 MUX2_X1 _19679_ (.A(_03098_),
    .B(_03101_),
    .S(_13297_),
    .Z(_03102_));
 MUX2_X1 _19680_ (.A(_03095_),
    .B(_03102_),
    .S(_13115_),
    .Z(_03103_));
 AOI21_X4 _19681_ (.A(_13710_),
    .B1(_03103_),
    .B2(_13117_),
    .ZN(_03104_));
 OAI21_X1 _19682_ (.A(_13077_),
    .B1(_13078_),
    .B2(_03104_),
    .ZN(_03105_));
 OR2_X1 _19683_ (.A1(_13691_),
    .A2(_03105_),
    .ZN(_16458_));
 INV_X1 _19684_ (.A(_16458_),
    .ZN(_16454_));
 MUX2_X1 _19685_ (.A(_01009_),
    .B(_01011_),
    .S(_12666_),
    .Z(_03106_));
 NOR2_X1 _19686_ (.A1(_11027_),
    .A2(_03106_),
    .ZN(_03107_));
 MUX2_X1 _19687_ (.A(_01010_),
    .B(_01012_),
    .S(_11240_),
    .Z(_03108_));
 NOR2_X1 _19688_ (.A1(_11012_),
    .A2(_03108_),
    .ZN(_03109_));
 NOR3_X1 _19689_ (.A1(_12104_),
    .A2(_03107_),
    .A3(_03109_),
    .ZN(_03110_));
 NOR2_X1 _19690_ (.A1(_11207_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .ZN(_03111_));
 AOI21_X1 _19691_ (.A(_03111_),
    .B1(_01004_),
    .B2(_11006_),
    .ZN(_03112_));
 AOI221_X2 _19692_ (.A(_11021_),
    .B1(_13697_),
    .B2(_11030_),
    .C1(_03112_),
    .C2(_12098_),
    .ZN(_03113_));
 NOR3_X2 _19693_ (.A1(_11057_),
    .A2(_03110_),
    .A3(_03113_),
    .ZN(_03114_));
 MUX2_X1 _19694_ (.A(_01013_),
    .B(_01015_),
    .S(_11239_),
    .Z(_03115_));
 MUX2_X1 _19695_ (.A(_01014_),
    .B(_01016_),
    .S(_11239_),
    .Z(_03116_));
 MUX2_X1 _19696_ (.A(_03115_),
    .B(_03116_),
    .S(_11059_),
    .Z(_03117_));
 MUX2_X1 _19697_ (.A(_01005_),
    .B(_01007_),
    .S(_11239_),
    .Z(_03118_));
 MUX2_X1 _19698_ (.A(_01006_),
    .B(_01008_),
    .S(_11239_),
    .Z(_03119_));
 MUX2_X1 _19699_ (.A(_03118_),
    .B(_03119_),
    .S(_11059_),
    .Z(_03120_));
 MUX2_X1 _19700_ (.A(_03117_),
    .B(_03120_),
    .S(_10992_),
    .Z(_03121_));
 NOR2_X1 _19701_ (.A1(_11037_),
    .A2(_03121_),
    .ZN(_03122_));
 NOR3_X4 _19702_ (.A1(_11052_),
    .A2(_03114_),
    .A3(_03122_),
    .ZN(_03123_));
 MUX2_X1 _19703_ (.A(_01025_),
    .B(_01027_),
    .S(_12085_),
    .Z(_03124_));
 MUX2_X1 _19704_ (.A(_01026_),
    .B(_01028_),
    .S(_12085_),
    .Z(_03125_));
 MUX2_X1 _19705_ (.A(_03124_),
    .B(_03125_),
    .S(_11041_),
    .Z(_03126_));
 MUX2_X1 _19706_ (.A(_01017_),
    .B(_01019_),
    .S(_12085_),
    .Z(_03127_));
 MUX2_X1 _19707_ (.A(_01018_),
    .B(_01020_),
    .S(_12085_),
    .Z(_03128_));
 MUX2_X1 _19708_ (.A(_03127_),
    .B(_03128_),
    .S(_11041_),
    .Z(_03129_));
 MUX2_X1 _19709_ (.A(_03126_),
    .B(_03129_),
    .S(_12068_),
    .Z(_03130_));
 MUX2_X1 _19710_ (.A(_01029_),
    .B(_01031_),
    .S(_12085_),
    .Z(_03131_));
 MUX2_X1 _19711_ (.A(_01030_),
    .B(_01032_),
    .S(_12085_),
    .Z(_03132_));
 MUX2_X1 _19712_ (.A(_03131_),
    .B(_03132_),
    .S(_11026_),
    .Z(_03133_));
 MUX2_X1 _19713_ (.A(_01021_),
    .B(_01023_),
    .S(_12085_),
    .Z(_03134_));
 MUX2_X1 _19714_ (.A(_01022_),
    .B(_01024_),
    .S(_12061_),
    .Z(_03135_));
 MUX2_X1 _19715_ (.A(_03134_),
    .B(_03135_),
    .S(_11026_),
    .Z(_03136_));
 MUX2_X1 _19716_ (.A(_03133_),
    .B(_03136_),
    .S(_12068_),
    .Z(_03137_));
 MUX2_X2 _19717_ (.A(_03130_),
    .B(_03137_),
    .S(_10987_),
    .Z(_03138_));
 AOI21_X4 _19718_ (.A(_03123_),
    .B1(_03138_),
    .B2(_11053_),
    .ZN(_03139_));
 AND2_X1 _19719_ (.A1(_11973_),
    .A2(_03139_),
    .ZN(_03140_));
 NAND2_X1 _19720_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(_10819_),
    .ZN(_03141_));
 CLKBUF_X2 _19721_ (.A(\cs_registers_i.pc_id_i[27] ),
    .Z(_03142_));
 NAND2_X1 _19722_ (.A1(_03142_),
    .A2(_11111_),
    .ZN(_03143_));
 OAI21_X1 _19723_ (.A(_03141_),
    .B1(_03143_),
    .B2(_11114_),
    .ZN(_03144_));
 OR2_X4 _19724_ (.A1(_03140_),
    .A2(_03144_),
    .ZN(_16453_));
 INV_X2 _19725_ (.A(_16453_),
    .ZN(_16457_));
 INV_X1 _19726_ (.A(_15880_),
    .ZN(_03145_));
 BUF_X2 _19727_ (.A(_15876_),
    .Z(_03146_));
 AOI21_X2 _19728_ (.A(_15875_),
    .B1(_15871_),
    .B2(_03146_),
    .ZN(_03147_));
 NAND2_X2 _19729_ (.A1(_15872_),
    .A2(_03146_),
    .ZN(_03148_));
 OAI21_X4 _19730_ (.A(_03147_),
    .B1(_13603_),
    .B2(_03148_),
    .ZN(_03149_));
 XNOR2_X2 _19731_ (.A(_03149_),
    .B(_03145_),
    .ZN(\alu_adder_result_ex[27] ));
 INV_X1 _19732_ (.A(_03146_),
    .ZN(_03150_));
 INV_X1 _19733_ (.A(_15867_),
    .ZN(_03151_));
 AOI21_X2 _19734_ (.A(_13596_),
    .B1(_15864_),
    .B2(_13427_),
    .ZN(_03152_));
 OAI21_X4 _19735_ (.A(_03151_),
    .B1(_03152_),
    .B2(_13604_),
    .ZN(_03153_));
 AOI21_X4 _19736_ (.A(_15871_),
    .B1(_15872_),
    .B2(_03153_),
    .ZN(_03154_));
 NOR2_X4 _19737_ (.A1(_03150_),
    .A2(_03154_),
    .ZN(_03155_));
 AND3_X2 _19738_ (.A1(_15864_),
    .A2(_15868_),
    .A3(_15872_),
    .ZN(_03156_));
 NOR2_X1 _19739_ (.A1(_03146_),
    .A2(_03156_),
    .ZN(_03157_));
 AOI21_X2 _19740_ (.A(_03155_),
    .B1(_03157_),
    .B2(_03154_),
    .ZN(_03158_));
 AND2_X1 _19741_ (.A1(_03150_),
    .A2(_03154_),
    .ZN(_03159_));
 OAI211_X2 _19742_ (.A(_13438_),
    .B(_03159_),
    .C1(_13440_),
    .C2(_12342_),
    .ZN(_03160_));
 NAND2_X2 _19743_ (.A1(_03146_),
    .A2(_03156_),
    .ZN(_03161_));
 OAI211_X4 _19744_ (.A(_03158_),
    .B(_03160_),
    .C1(_13612_),
    .C2(_03161_),
    .ZN(_03162_));
 INV_X4 _19745_ (.A(net391),
    .ZN(\alu_adder_result_ex[26] ));
 AOI21_X1 _19746_ (.A(_13073_),
    .B1(_13075_),
    .B2(_10876_),
    .ZN(_03163_));
 MUX2_X1 _19747_ (.A(_01040_),
    .B(_01042_),
    .S(_12736_),
    .Z(_03164_));
 NOR2_X1 _19748_ (.A1(_12361_),
    .A2(_03164_),
    .ZN(_03165_));
 MUX2_X1 _19749_ (.A(_01041_),
    .B(_01043_),
    .S(_13079_),
    .Z(_03166_));
 NOR2_X1 _19750_ (.A1(_12367_),
    .A2(_03166_),
    .ZN(_03167_));
 NOR3_X1 _19751_ (.A1(_12409_),
    .A2(_03165_),
    .A3(_03167_),
    .ZN(_03168_));
 INV_X1 _19752_ (.A(_01034_),
    .ZN(_03169_));
 NOR2_X1 _19753_ (.A1(_12401_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .ZN(_03170_));
 AOI21_X1 _19754_ (.A(_03170_),
    .B1(_01035_),
    .B2(_12547_),
    .ZN(_03171_));
 AOI221_X2 _19755_ (.A(_12372_),
    .B1(_03169_),
    .B2(_12373_),
    .C1(_03171_),
    .C2(_12445_),
    .ZN(_03172_));
 NOR3_X2 _19756_ (.A1(_12423_),
    .A2(_03168_),
    .A3(_03172_),
    .ZN(_03173_));
 MUX2_X1 _19757_ (.A(_01044_),
    .B(_01046_),
    .S(_13170_),
    .Z(_03174_));
 MUX2_X1 _19758_ (.A(_01045_),
    .B(_01047_),
    .S(_12919_),
    .Z(_03175_));
 MUX2_X1 _19759_ (.A(_03174_),
    .B(_03175_),
    .S(_13092_),
    .Z(_03176_));
 MUX2_X1 _19760_ (.A(_01036_),
    .B(_01038_),
    .S(_12919_),
    .Z(_03177_));
 MUX2_X1 _19761_ (.A(_01037_),
    .B(_01039_),
    .S(_13278_),
    .Z(_03178_));
 MUX2_X1 _19762_ (.A(_03177_),
    .B(_03178_),
    .S(_13281_),
    .Z(_03179_));
 MUX2_X1 _19763_ (.A(_03176_),
    .B(_03179_),
    .S(_12408_),
    .Z(_03180_));
 NOR2_X1 _19764_ (.A1(_12807_),
    .A2(_03180_),
    .ZN(_03181_));
 NOR3_X4 _19765_ (.A1(_12354_),
    .A2(_03173_),
    .A3(_03181_),
    .ZN(_03182_));
 MUX2_X1 _19766_ (.A(_01056_),
    .B(_01058_),
    .S(net343),
    .Z(_03183_));
 MUX2_X1 _19767_ (.A(_01057_),
    .B(_01059_),
    .S(_13472_),
    .Z(_03184_));
 MUX2_X1 _19768_ (.A(_03183_),
    .B(_03184_),
    .S(_13194_),
    .Z(_03185_));
 MUX2_X1 _19769_ (.A(_01048_),
    .B(_01050_),
    .S(_13472_),
    .Z(_03186_));
 MUX2_X1 _19770_ (.A(_01049_),
    .B(_01051_),
    .S(_13192_),
    .Z(_03187_));
 MUX2_X1 _19771_ (.A(_03186_),
    .B(_03187_),
    .S(_13194_),
    .Z(_03188_));
 MUX2_X1 _19772_ (.A(_03185_),
    .B(_03188_),
    .S(_13297_),
    .Z(_03189_));
 MUX2_X1 _19773_ (.A(_01060_),
    .B(_01062_),
    .S(_13472_),
    .Z(_03190_));
 MUX2_X1 _19774_ (.A(_01061_),
    .B(_01063_),
    .S(_13192_),
    .Z(_03191_));
 MUX2_X1 _19775_ (.A(_03190_),
    .B(_03191_),
    .S(_12360_),
    .Z(_03192_));
 MUX2_X1 _19776_ (.A(_01052_),
    .B(_01054_),
    .S(_13192_),
    .Z(_03193_));
 MUX2_X1 _19777_ (.A(_01053_),
    .B(_01055_),
    .S(_13289_),
    .Z(_03194_));
 MUX2_X1 _19778_ (.A(_03193_),
    .B(_03194_),
    .S(_12360_),
    .Z(_03195_));
 MUX2_X1 _19779_ (.A(_03192_),
    .B(_03195_),
    .S(_13297_),
    .Z(_03196_));
 MUX2_X1 _19780_ (.A(_03189_),
    .B(_03196_),
    .S(_13115_),
    .Z(_03197_));
 AOI21_X4 _19781_ (.A(_03182_),
    .B1(_03197_),
    .B2(_13117_),
    .ZN(_03198_));
 OAI21_X1 _19782_ (.A(_13077_),
    .B1(_13078_),
    .B2(_03198_),
    .ZN(_03199_));
 OR2_X1 _19783_ (.A1(_03163_),
    .A2(_03199_),
    .ZN(_16466_));
 INV_X1 _19784_ (.A(_16466_),
    .ZN(_16462_));
 NAND2_X1 _19785_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(_10957_),
    .ZN(_03200_));
 NOR2_X2 _19786_ (.A1(_11021_),
    .A2(_11051_),
    .ZN(_03201_));
 MUX2_X1 _19787_ (.A(_01036_),
    .B(_01038_),
    .S(_11017_),
    .Z(_03202_));
 NOR2_X1 _19788_ (.A1(_11002_),
    .A2(_03202_),
    .ZN(_03203_));
 MUX2_X1 _19789_ (.A(_01037_),
    .B(_01039_),
    .S(_11254_),
    .Z(_03204_));
 NOR2_X1 _19790_ (.A1(_11013_),
    .A2(_03204_),
    .ZN(_03205_));
 NOR3_X1 _19791_ (.A1(_11038_),
    .A2(_03203_),
    .A3(_03205_),
    .ZN(_03206_));
 NOR2_X1 _19792_ (.A1(_11209_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .ZN(_03207_));
 AOI21_X1 _19793_ (.A(_03207_),
    .B1(_01035_),
    .B2(_11188_),
    .ZN(_03208_));
 AOI221_X1 _19794_ (.A(_11057_),
    .B1(_03169_),
    .B2(_11032_),
    .C1(_03208_),
    .C2(_11094_),
    .ZN(_03209_));
 OAI21_X1 _19795_ (.A(_03201_),
    .B1(_03206_),
    .B2(_03209_),
    .ZN(_03210_));
 MUX2_X1 _19796_ (.A(_01052_),
    .B(_01054_),
    .S(_11097_),
    .Z(_03211_));
 MUX2_X1 _19797_ (.A(_01053_),
    .B(_01055_),
    .S(_11097_),
    .Z(_03212_));
 MUX2_X1 _19798_ (.A(_03211_),
    .B(_03212_),
    .S(_11061_),
    .Z(_03213_));
 MUX2_X1 _19799_ (.A(_01048_),
    .B(_01050_),
    .S(_11097_),
    .Z(_03214_));
 MUX2_X1 _19800_ (.A(_01049_),
    .B(_01051_),
    .S(_11097_),
    .Z(_03215_));
 MUX2_X1 _19801_ (.A(_03214_),
    .B(_03215_),
    .S(_11061_),
    .Z(_03216_));
 MUX2_X1 _19802_ (.A(_03213_),
    .B(_03216_),
    .S(_11223_),
    .Z(_03217_));
 NAND2_X1 _19803_ (.A1(_11931_),
    .A2(_03217_),
    .ZN(_03218_));
 MUX2_X1 _19804_ (.A(_01044_),
    .B(_01046_),
    .S(_12503_),
    .Z(_03219_));
 MUX2_X1 _19805_ (.A(_01045_),
    .B(_01047_),
    .S(_12503_),
    .Z(_03220_));
 MUX2_X1 _19806_ (.A(_03219_),
    .B(_03220_),
    .S(_11093_),
    .Z(_03221_));
 MUX2_X1 _19807_ (.A(_01040_),
    .B(_01042_),
    .S(_12503_),
    .Z(_03222_));
 MUX2_X1 _19808_ (.A(_01041_),
    .B(_01043_),
    .S(_11246_),
    .Z(_03223_));
 MUX2_X1 _19809_ (.A(_03222_),
    .B(_03223_),
    .S(_11093_),
    .Z(_03224_));
 MUX2_X1 _19810_ (.A(_03221_),
    .B(_03224_),
    .S(_11073_),
    .Z(_03225_));
 OAI21_X1 _19811_ (.A(_11055_),
    .B1(_11053_),
    .B2(_03225_),
    .ZN(_03226_));
 NAND3_X2 _19812_ (.A1(_03210_),
    .A2(_03218_),
    .A3(_03226_),
    .ZN(_03227_));
 MUX2_X1 _19813_ (.A(_01060_),
    .B(_01062_),
    .S(_11017_),
    .Z(_03228_));
 MUX2_X1 _19814_ (.A(_01061_),
    .B(_01063_),
    .S(_11017_),
    .Z(_03229_));
 MUX2_X1 _19815_ (.A(_03228_),
    .B(_03229_),
    .S(_11088_),
    .Z(_03230_));
 NAND2_X1 _19816_ (.A1(_10989_),
    .A2(_03230_),
    .ZN(_03231_));
 MUX2_X1 _19817_ (.A(_01056_),
    .B(_01058_),
    .S(_11017_),
    .Z(_03232_));
 MUX2_X1 _19818_ (.A(_01057_),
    .B(_01059_),
    .S(_11017_),
    .Z(_03233_));
 MUX2_X1 _19819_ (.A(_03232_),
    .B(_03233_),
    .S(_11088_),
    .Z(_03234_));
 NAND2_X1 _19820_ (.A1(_11038_),
    .A2(_03234_),
    .ZN(_03235_));
 NAND4_X2 _19821_ (.A1(_11056_),
    .A2(_11931_),
    .A3(_03231_),
    .A4(_03235_),
    .ZN(_03236_));
 AND2_X2 _19822_ (.A1(_03227_),
    .A2(_03236_),
    .ZN(_03237_));
 CLKBUF_X2 _19823_ (.A(\cs_registers_i.pc_id_i[28] ),
    .Z(_03238_));
 NAND2_X1 _19824_ (.A1(_03238_),
    .A2(_11113_),
    .ZN(_03239_));
 OAI221_X2 _19825_ (.A(_03200_),
    .B1(_03237_),
    .B2(_11818_),
    .C1(_03239_),
    .C2(_11115_),
    .ZN(_03240_));
 BUF_X4 _19826_ (.A(_03240_),
    .Z(_16461_));
 INV_X2 _19827_ (.A(_16461_),
    .ZN(_16465_));
 AOI21_X1 _19828_ (.A(_13073_),
    .B1(_13075_),
    .B2(_10875_),
    .ZN(_03241_));
 MUX2_X1 _19829_ (.A(_01071_),
    .B(_01073_),
    .S(_12736_),
    .Z(_03242_));
 NOR2_X1 _19830_ (.A1(_12361_),
    .A2(_03242_),
    .ZN(_03243_));
 MUX2_X1 _19831_ (.A(_01072_),
    .B(_01074_),
    .S(_13079_),
    .Z(_03244_));
 NOR2_X1 _19832_ (.A1(_12367_),
    .A2(_03244_),
    .ZN(_03245_));
 NOR3_X1 _19833_ (.A1(_12409_),
    .A2(_03243_),
    .A3(_03245_),
    .ZN(_03246_));
 INV_X1 _19834_ (.A(_01065_),
    .ZN(_03247_));
 NOR2_X1 _19835_ (.A1(_12401_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .ZN(_03248_));
 AOI21_X1 _19836_ (.A(_03248_),
    .B1(_01066_),
    .B2(_12547_),
    .ZN(_03249_));
 AOI221_X2 _19837_ (.A(_12372_),
    .B1(_03247_),
    .B2(_12373_),
    .C1(_03249_),
    .C2(_12445_),
    .ZN(_03250_));
 NOR3_X2 _19838_ (.A1(_12423_),
    .A2(_03246_),
    .A3(_03250_),
    .ZN(_03251_));
 MUX2_X1 _19839_ (.A(_01075_),
    .B(_01077_),
    .S(_13170_),
    .Z(_03252_));
 MUX2_X1 _19840_ (.A(_01076_),
    .B(_01078_),
    .S(_12919_),
    .Z(_03253_));
 MUX2_X1 _19841_ (.A(_03252_),
    .B(_03253_),
    .S(_13092_),
    .Z(_03254_));
 MUX2_X1 _19842_ (.A(_01067_),
    .B(_01069_),
    .S(_12919_),
    .Z(_03255_));
 MUX2_X1 _19843_ (.A(_01068_),
    .B(_01070_),
    .S(_13278_),
    .Z(_03256_));
 MUX2_X1 _19844_ (.A(_03255_),
    .B(_03256_),
    .S(_13281_),
    .Z(_03257_));
 MUX2_X1 _19845_ (.A(_03254_),
    .B(_03257_),
    .S(_12408_),
    .Z(_03258_));
 NOR2_X1 _19846_ (.A1(_12807_),
    .A2(_03258_),
    .ZN(_03259_));
 NOR3_X4 _19847_ (.A1(_12354_),
    .A2(_03251_),
    .A3(_03259_),
    .ZN(_03260_));
 MUX2_X1 _19848_ (.A(_01087_),
    .B(_01089_),
    .S(net343),
    .Z(_03261_));
 MUX2_X1 _19849_ (.A(_01088_),
    .B(_01090_),
    .S(_13472_),
    .Z(_03262_));
 MUX2_X1 _19850_ (.A(_03261_),
    .B(_03262_),
    .S(_13194_),
    .Z(_03263_));
 MUX2_X1 _19851_ (.A(_01079_),
    .B(_01081_),
    .S(_13472_),
    .Z(_03264_));
 MUX2_X1 _19852_ (.A(_01080_),
    .B(_01082_),
    .S(_13192_),
    .Z(_03265_));
 MUX2_X1 _19853_ (.A(_03264_),
    .B(_03265_),
    .S(_13194_),
    .Z(_03266_));
 MUX2_X1 _19854_ (.A(_03263_),
    .B(_03266_),
    .S(_13297_),
    .Z(_03267_));
 MUX2_X1 _19855_ (.A(_01091_),
    .B(_01093_),
    .S(_13472_),
    .Z(_03268_));
 MUX2_X1 _19856_ (.A(_01092_),
    .B(_01094_),
    .S(_13192_),
    .Z(_03269_));
 MUX2_X1 _19857_ (.A(_03268_),
    .B(_03269_),
    .S(_12360_),
    .Z(_03270_));
 MUX2_X1 _19858_ (.A(_01083_),
    .B(_01085_),
    .S(_13192_),
    .Z(_03271_));
 MUX2_X1 _19859_ (.A(_01084_),
    .B(_01086_),
    .S(_13289_),
    .Z(_03272_));
 MUX2_X1 _19860_ (.A(_03271_),
    .B(_03272_),
    .S(_12360_),
    .Z(_03273_));
 MUX2_X1 _19861_ (.A(_03270_),
    .B(_03273_),
    .S(_13297_),
    .Z(_03274_));
 MUX2_X1 _19862_ (.A(_03267_),
    .B(_03274_),
    .S(_13115_),
    .Z(_03275_));
 AOI21_X4 _19863_ (.A(_03260_),
    .B1(_03275_),
    .B2(_13117_),
    .ZN(_03276_));
 OAI21_X1 _19864_ (.A(_13077_),
    .B1(_13078_),
    .B2(_03276_),
    .ZN(_03277_));
 OR2_X2 _19865_ (.A1(_03241_),
    .A2(_03277_),
    .ZN(_16474_));
 INV_X1 _19866_ (.A(_16474_),
    .ZN(_16470_));
 NAND2_X1 _19867_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(_10957_),
    .ZN(_03278_));
 MUX2_X1 _19868_ (.A(_01071_),
    .B(_01073_),
    .S(_11017_),
    .Z(_03279_));
 NOR2_X1 _19869_ (.A1(_11088_),
    .A2(_03279_),
    .ZN(_03280_));
 MUX2_X1 _19870_ (.A(_01072_),
    .B(_01074_),
    .S(_11254_),
    .Z(_03281_));
 NOR2_X1 _19871_ (.A1(_11013_),
    .A2(_03281_),
    .ZN(_03282_));
 NOR3_X1 _19872_ (.A1(_10994_),
    .A2(_03280_),
    .A3(_03282_),
    .ZN(_03283_));
 NOR2_X1 _19873_ (.A1(_11209_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .ZN(_03284_));
 AOI21_X1 _19874_ (.A(_03284_),
    .B1(_01066_),
    .B2(_11008_),
    .ZN(_03285_));
 AOI221_X1 _19875_ (.A(_11022_),
    .B1(_03247_),
    .B2(_11032_),
    .C1(_03285_),
    .C2(_11001_),
    .ZN(_03286_));
 OR3_X1 _19876_ (.A1(_10989_),
    .A2(_03283_),
    .A3(_03286_),
    .ZN(_03287_));
 MUX2_X1 _19877_ (.A(_01075_),
    .B(_01077_),
    .S(_11188_),
    .Z(_03288_));
 MUX2_X1 _19878_ (.A(_01076_),
    .B(_01078_),
    .S(_11188_),
    .Z(_03289_));
 MUX2_X1 _19879_ (.A(_03288_),
    .B(_03289_),
    .S(_11002_),
    .Z(_03290_));
 NAND2_X1 _19880_ (.A1(_11056_),
    .A2(_03290_),
    .ZN(_03291_));
 MUX2_X1 _19881_ (.A(_01067_),
    .B(_01069_),
    .S(_11188_),
    .Z(_03292_));
 MUX2_X1 _19882_ (.A(_01068_),
    .B(_01070_),
    .S(_11188_),
    .Z(_03293_));
 MUX2_X1 _19883_ (.A(_03292_),
    .B(_03293_),
    .S(_11088_),
    .Z(_03294_));
 NAND2_X1 _19884_ (.A1(_10995_),
    .A2(_03294_),
    .ZN(_03295_));
 NAND3_X1 _19885_ (.A1(_10989_),
    .A2(_03291_),
    .A3(_03295_),
    .ZN(_03296_));
 AOI21_X2 _19886_ (.A(_11054_),
    .B1(_03287_),
    .B2(_03296_),
    .ZN(_03297_));
 MUX2_X1 _19887_ (.A(_01083_),
    .B(_01085_),
    .S(_11209_),
    .Z(_03298_));
 MUX2_X1 _19888_ (.A(_01084_),
    .B(_01086_),
    .S(_11209_),
    .Z(_03299_));
 MUX2_X1 _19889_ (.A(_03298_),
    .B(_03299_),
    .S(_11094_),
    .Z(_03300_));
 MUX2_X1 _19890_ (.A(_01079_),
    .B(_01080_),
    .S(_11001_),
    .Z(_03301_));
 MUX2_X1 _19891_ (.A(_01081_),
    .B(_01082_),
    .S(_11028_),
    .Z(_03302_));
 AOI222_X2 _19892_ (.A1(_11085_),
    .A2(_03300_),
    .B1(_03301_),
    .B2(_11091_),
    .C1(_03302_),
    .C2(_11100_),
    .ZN(_03303_));
 NAND2_X1 _19893_ (.A1(_11931_),
    .A2(_03303_),
    .ZN(_03304_));
 MUX2_X1 _19894_ (.A(_01093_),
    .B(_01094_),
    .S(_11805_),
    .Z(_03305_));
 AOI21_X2 _19895_ (.A(_11073_),
    .B1(_03305_),
    .B2(_11069_),
    .ZN(_03306_));
 MUX2_X1 _19896_ (.A(_01089_),
    .B(_01090_),
    .S(_11027_),
    .Z(_03307_));
 AOI21_X2 _19897_ (.A(_11057_),
    .B1(_03307_),
    .B2(_11068_),
    .ZN(_03308_));
 OAI21_X1 _19898_ (.A(_11081_),
    .B1(_03306_),
    .B2(_03308_),
    .ZN(_03309_));
 MUX2_X1 _19899_ (.A(_01087_),
    .B(_01088_),
    .S(_11805_),
    .Z(_03310_));
 INV_X1 _19900_ (.A(_03310_),
    .ZN(_03311_));
 MUX2_X1 _19901_ (.A(_01091_),
    .B(_01092_),
    .S(_11028_),
    .Z(_03312_));
 INV_X1 _19902_ (.A(_03312_),
    .ZN(_03313_));
 AOI221_X2 _19903_ (.A(_10994_),
    .B1(_03308_),
    .B2(_03311_),
    .C1(_03313_),
    .C2(_03306_),
    .ZN(_03314_));
 AOI21_X2 _19904_ (.A(_03304_),
    .B1(_03309_),
    .B2(_03314_),
    .ZN(_03315_));
 NOR2_X2 _19905_ (.A1(_03297_),
    .A2(_03315_),
    .ZN(_03316_));
 NAND2_X1 _19906_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(_11113_),
    .ZN(_03317_));
 OAI221_X2 _19907_ (.A(_03278_),
    .B1(_03316_),
    .B2(_11818_),
    .C1(_03317_),
    .C2(_11115_),
    .ZN(_03318_));
 BUF_X4 _19908_ (.A(_03318_),
    .Z(_16469_));
 INV_X1 _19909_ (.A(_16469_),
    .ZN(_16473_));
 CLKBUF_X3 _19910_ (.A(_15888_),
    .Z(_03319_));
 INV_X1 _19911_ (.A(_15883_),
    .ZN(_03320_));
 BUF_X2 _19912_ (.A(_15884_),
    .Z(_03321_));
 OAI21_X1 _19913_ (.A(_03321_),
    .B1(_15879_),
    .B2(_15880_),
    .ZN(_03322_));
 AOI21_X1 _19914_ (.A(_03319_),
    .B1(_03320_),
    .B2(_03322_),
    .ZN(_03323_));
 INV_X1 _19915_ (.A(_15879_),
    .ZN(_03324_));
 OAI21_X1 _19916_ (.A(_03324_),
    .B1(_03147_),
    .B2(_03145_),
    .ZN(_03325_));
 AOI21_X1 _19917_ (.A(_15883_),
    .B1(_03325_),
    .B2(_03321_),
    .ZN(_03326_));
 AOI21_X2 _19918_ (.A(_03323_),
    .B1(_03326_),
    .B2(_03319_),
    .ZN(_03327_));
 AND3_X1 _19919_ (.A1(_15880_),
    .A2(_03321_),
    .A3(_03319_),
    .ZN(_03328_));
 OR3_X4 _19920_ (.A1(_03148_),
    .A2(_13603_),
    .A3(_03328_),
    .ZN(_03329_));
 AOI21_X1 _19921_ (.A(_15883_),
    .B1(_15879_),
    .B2(_03321_),
    .ZN(_03330_));
 NAND2_X1 _19922_ (.A1(_03147_),
    .A2(_03330_),
    .ZN(_03331_));
 OAI22_X4 _19923_ (.A1(_13603_),
    .A2(_03148_),
    .B1(_03331_),
    .B2(_03319_),
    .ZN(_03332_));
 AOI21_X4 _19924_ (.A(_03327_),
    .B1(_03332_),
    .B2(_03329_),
    .ZN(\alu_adder_result_ex[29] ));
 OAI21_X4 _19925_ (.A(_15880_),
    .B1(_15875_),
    .B2(_03155_),
    .ZN(_03333_));
 NAND2_X4 _19926_ (.A1(_03333_),
    .A2(_03324_),
    .ZN(_03334_));
 NOR2_X1 _19927_ (.A1(_03145_),
    .A2(_03161_),
    .ZN(_03335_));
 AOI21_X4 _19928_ (.A(_03334_),
    .B1(_03335_),
    .B2(_13441_),
    .ZN(_03336_));
 XNOR2_X2 _19929_ (.A(_03336_),
    .B(_03321_),
    .ZN(\alu_adder_result_ex[28] ));
 AOI21_X1 _19930_ (.A(_13072_),
    .B1(_13074_),
    .B2(_10884_),
    .ZN(_03337_));
 MUX2_X1 _19931_ (.A(_01102_),
    .B(_01104_),
    .S(_12736_),
    .Z(_03338_));
 NOR2_X1 _19932_ (.A1(_12361_),
    .A2(_03338_),
    .ZN(_03339_));
 MUX2_X1 _19933_ (.A(_01103_),
    .B(_01105_),
    .S(_13079_),
    .Z(_03340_));
 NOR2_X1 _19934_ (.A1(_12367_),
    .A2(_03340_),
    .ZN(_03341_));
 NOR3_X1 _19935_ (.A1(_12409_),
    .A2(_03339_),
    .A3(_03341_),
    .ZN(_03342_));
 INV_X1 _19936_ (.A(_01096_),
    .ZN(_03343_));
 NOR2_X1 _19937_ (.A1(_12398_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .ZN(_03344_));
 AOI21_X1 _19938_ (.A(_03344_),
    .B1(_01097_),
    .B2(_12547_),
    .ZN(_03345_));
 AOI221_X2 _19939_ (.A(_10758_),
    .B1(_03343_),
    .B2(_12373_),
    .C1(_03345_),
    .C2(_12555_),
    .ZN(_03346_));
 NOR3_X2 _19940_ (.A1(_12423_),
    .A2(_03342_),
    .A3(_03346_),
    .ZN(_03347_));
 MUX2_X1 _19941_ (.A(_01106_),
    .B(_01108_),
    .S(_12400_),
    .Z(_03348_));
 MUX2_X1 _19942_ (.A(_01107_),
    .B(_01109_),
    .S(_13170_),
    .Z(_03349_));
 MUX2_X1 _19943_ (.A(_03348_),
    .B(_03349_),
    .S(_13092_),
    .Z(_03350_));
 MUX2_X1 _19944_ (.A(_01098_),
    .B(_01100_),
    .S(_13170_),
    .Z(_03351_));
 MUX2_X1 _19945_ (.A(_01099_),
    .B(_01101_),
    .S(_12919_),
    .Z(_03352_));
 MUX2_X1 _19946_ (.A(_03351_),
    .B(_03352_),
    .S(_13092_),
    .Z(_03353_));
 MUX2_X1 _19947_ (.A(_03350_),
    .B(_03353_),
    .S(_12408_),
    .Z(_03354_));
 NOR2_X2 _19948_ (.A1(_12807_),
    .A2(_03354_),
    .ZN(_03355_));
 NOR3_X4 _19949_ (.A1(_12354_),
    .A2(_03347_),
    .A3(_03355_),
    .ZN(_03356_));
 MUX2_X1 _19950_ (.A(_01118_),
    .B(_01120_),
    .S(_12385_),
    .Z(_03357_));
 MUX2_X1 _19951_ (.A(_01119_),
    .B(_01121_),
    .S(net343),
    .Z(_03358_));
 MUX2_X1 _19952_ (.A(_03357_),
    .B(_03358_),
    .S(_12392_),
    .Z(_03359_));
 MUX2_X1 _19953_ (.A(_01110_),
    .B(_01112_),
    .S(net343),
    .Z(_03360_));
 MUX2_X1 _19954_ (.A(_01111_),
    .B(_01113_),
    .S(net344),
    .Z(_03361_));
 MUX2_X1 _19955_ (.A(_03360_),
    .B(_03361_),
    .S(_12392_),
    .Z(_03362_));
 MUX2_X1 _19956_ (.A(_03359_),
    .B(_03362_),
    .S(_12394_),
    .Z(_03363_));
 MUX2_X1 _19957_ (.A(_01122_),
    .B(_01124_),
    .S(net343),
    .Z(_03364_));
 MUX2_X1 _19958_ (.A(_01123_),
    .B(_01125_),
    .S(_13472_),
    .Z(_03365_));
 MUX2_X1 _19959_ (.A(_03364_),
    .B(_03365_),
    .S(_12392_),
    .Z(_03366_));
 MUX2_X1 _19960_ (.A(_01114_),
    .B(_01116_),
    .S(net344),
    .Z(_03367_));
 MUX2_X1 _19961_ (.A(_01115_),
    .B(_01117_),
    .S(_13192_),
    .Z(_03368_));
 MUX2_X1 _19962_ (.A(_03367_),
    .B(_03368_),
    .S(_13194_),
    .Z(_03369_));
 MUX2_X1 _19963_ (.A(_03366_),
    .B(_03369_),
    .S(_12394_),
    .Z(_03370_));
 MUX2_X1 _19964_ (.A(_03363_),
    .B(_03370_),
    .S(_13115_),
    .Z(_03371_));
 AOI21_X4 _19965_ (.A(_03356_),
    .B1(_03371_),
    .B2(_13117_),
    .ZN(_03372_));
 OAI21_X1 _19966_ (.A(_10838_),
    .B1(_11121_),
    .B2(_03372_),
    .ZN(_03373_));
 OR2_X1 _19967_ (.A1(_03337_),
    .A2(_03373_),
    .ZN(_16477_));
 INV_X1 _19968_ (.A(_16477_),
    .ZN(_16481_));
 NAND2_X1 _19969_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(_10957_),
    .ZN(_03374_));
 MUX2_X1 _19970_ (.A(_01102_),
    .B(_01104_),
    .S(_11254_),
    .Z(_03375_));
 NOR2_X1 _19971_ (.A1(_11088_),
    .A2(_03375_),
    .ZN(_03376_));
 MUX2_X1 _19972_ (.A(_01103_),
    .B(_01105_),
    .S(_11254_),
    .Z(_03377_));
 NOR2_X1 _19973_ (.A1(_11013_),
    .A2(_03377_),
    .ZN(_03378_));
 NOR3_X1 _19974_ (.A1(_10994_),
    .A2(_03376_),
    .A3(_03378_),
    .ZN(_03379_));
 NOR2_X1 _19975_ (.A1(_11209_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .ZN(_03380_));
 AOI21_X1 _19976_ (.A(_03380_),
    .B1(_01097_),
    .B2(_11008_),
    .ZN(_03381_));
 AOI221_X1 _19977_ (.A(_11022_),
    .B1(_03343_),
    .B2(_11032_),
    .C1(_03381_),
    .C2(_11001_),
    .ZN(_03382_));
 OR3_X2 _19978_ (.A1(_10989_),
    .A2(_03379_),
    .A3(_03382_),
    .ZN(_03383_));
 MUX2_X1 _19979_ (.A(_01106_),
    .B(_01108_),
    .S(_11008_),
    .Z(_03384_));
 MUX2_X1 _19980_ (.A(_01107_),
    .B(_01109_),
    .S(_11188_),
    .Z(_03385_));
 MUX2_X1 _19981_ (.A(_03384_),
    .B(_03385_),
    .S(_11088_),
    .Z(_03386_));
 NAND2_X1 _19982_ (.A1(_11055_),
    .A2(_03386_),
    .ZN(_03387_));
 MUX2_X1 _19983_ (.A(_01098_),
    .B(_01100_),
    .S(_11008_),
    .Z(_03388_));
 MUX2_X1 _19984_ (.A(_01099_),
    .B(_01101_),
    .S(_11008_),
    .Z(_03389_));
 MUX2_X1 _19985_ (.A(_03388_),
    .B(_03389_),
    .S(_11088_),
    .Z(_03390_));
 NAND2_X1 _19986_ (.A1(_10995_),
    .A2(_03390_),
    .ZN(_03391_));
 NAND3_X2 _19987_ (.A1(_10989_),
    .A2(_03387_),
    .A3(_03391_),
    .ZN(_03392_));
 AOI21_X4 _19988_ (.A(_11054_),
    .B1(_03383_),
    .B2(_03392_),
    .ZN(_03393_));
 MUX2_X1 _19989_ (.A(_01114_),
    .B(_01116_),
    .S(_11254_),
    .Z(_03394_));
 MUX2_X1 _19990_ (.A(_01115_),
    .B(_01117_),
    .S(_11254_),
    .Z(_03395_));
 MUX2_X1 _19991_ (.A(_03394_),
    .B(_03395_),
    .S(_11094_),
    .Z(_03396_));
 MUX2_X1 _19992_ (.A(_01110_),
    .B(_01111_),
    .S(_11094_),
    .Z(_03397_));
 MUX2_X1 _19993_ (.A(_01112_),
    .B(_01113_),
    .S(_11001_),
    .Z(_03398_));
 AOI222_X2 _19994_ (.A1(_11085_),
    .A2(_03396_),
    .B1(_03397_),
    .B2(_11091_),
    .C1(_03398_),
    .C2(_11100_),
    .ZN(_03399_));
 MUX2_X1 _19995_ (.A(_01120_),
    .B(_01121_),
    .S(_11075_),
    .Z(_03400_));
 AOI21_X1 _19996_ (.A(_11058_),
    .B1(_03400_),
    .B2(_11069_),
    .ZN(_03401_));
 MUX2_X1 _19997_ (.A(_01124_),
    .B(_01125_),
    .S(_11093_),
    .Z(_03402_));
 AOI21_X1 _19998_ (.A(_11073_),
    .B1(_03402_),
    .B2(_11069_),
    .ZN(_03403_));
 OAI21_X1 _19999_ (.A(_11081_),
    .B1(_03401_),
    .B2(_03403_),
    .ZN(_03404_));
 NAND2_X1 _20000_ (.A1(_11013_),
    .A2(_01122_),
    .ZN(_03405_));
 NAND2_X1 _20001_ (.A1(_11002_),
    .A2(_01123_),
    .ZN(_03406_));
 NAND3_X1 _20002_ (.A1(_03403_),
    .A2(_03405_),
    .A3(_03406_),
    .ZN(_03407_));
 NAND2_X1 _20003_ (.A1(_11013_),
    .A2(_01118_),
    .ZN(_03408_));
 NAND2_X1 _20004_ (.A1(_11002_),
    .A2(_01119_),
    .ZN(_03409_));
 NAND3_X1 _20005_ (.A1(_03401_),
    .A2(_03408_),
    .A3(_03409_),
    .ZN(_03410_));
 NAND4_X1 _20006_ (.A1(_11056_),
    .A2(_03404_),
    .A3(_03407_),
    .A4(_03410_),
    .ZN(_03411_));
 AND3_X2 _20007_ (.A1(_11054_),
    .A2(_03399_),
    .A3(_03411_),
    .ZN(_03412_));
 NOR3_X2 _20008_ (.A1(_11215_),
    .A2(_03393_),
    .A3(_03412_),
    .ZN(_03413_));
 OAI21_X2 _20009_ (.A(_11113_),
    .B1(_11115_),
    .B2(\cs_registers_i.pc_id_i[30] ),
    .ZN(_03414_));
 OAI21_X4 _20010_ (.A(_03374_),
    .B1(_03413_),
    .B2(_03414_),
    .ZN(_16482_));
 INV_X2 _20011_ (.A(_16482_),
    .ZN(_16478_));
 AOI21_X1 _20012_ (.A(_11167_),
    .B1(_12345_),
    .B2(_12346_),
    .ZN(_03415_));
 NOR2_X1 _20013_ (.A1(_11727_),
    .A2(_11167_),
    .ZN(_03416_));
 MUX2_X1 _20014_ (.A(_01153_),
    .B(_01155_),
    .S(_11614_),
    .Z(_03417_));
 MUX2_X1 _20015_ (.A(_01154_),
    .B(_01156_),
    .S(_11614_),
    .Z(_03418_));
 MUX2_X1 _20016_ (.A(_03417_),
    .B(_03418_),
    .S(_10710_),
    .Z(_03419_));
 MUX2_X1 _20017_ (.A(_01137_),
    .B(_01139_),
    .S(net377),
    .Z(_03420_));
 MUX2_X1 _20018_ (.A(_01138_),
    .B(_01140_),
    .S(net377),
    .Z(_03421_));
 MUX2_X1 _20019_ (.A(_03420_),
    .B(_03421_),
    .S(_11316_),
    .Z(_03422_));
 MUX2_X1 _20020_ (.A(_03419_),
    .B(_03422_),
    .S(_10763_),
    .Z(_03423_));
 NAND3_X1 _20021_ (.A1(_10731_),
    .A2(_10747_),
    .A3(_03423_),
    .ZN(_03424_));
 MUX2_X1 _20022_ (.A(_01149_),
    .B(_01151_),
    .S(_11501_),
    .Z(_03425_));
 MUX2_X1 _20023_ (.A(_01150_),
    .B(_01152_),
    .S(_11501_),
    .Z(_03426_));
 MUX2_X1 _20024_ (.A(_03425_),
    .B(_03426_),
    .S(_10710_),
    .Z(_03427_));
 MUX2_X1 _20025_ (.A(_01133_),
    .B(_01135_),
    .S(_11501_),
    .Z(_03428_));
 MUX2_X1 _20026_ (.A(_01134_),
    .B(_01136_),
    .S(_11614_),
    .Z(_03429_));
 MUX2_X1 _20027_ (.A(_03428_),
    .B(_03429_),
    .S(_10710_),
    .Z(_03430_));
 MUX2_X1 _20028_ (.A(_03427_),
    .B(_03430_),
    .S(_10763_),
    .Z(_03431_));
 NAND3_X1 _20029_ (.A1(_10736_),
    .A2(_10747_),
    .A3(_03431_),
    .ZN(_03432_));
 MUX2_X1 _20030_ (.A(_01145_),
    .B(_01147_),
    .S(_11614_),
    .Z(_03433_));
 MUX2_X1 _20031_ (.A(_01129_),
    .B(_01131_),
    .S(_11614_),
    .Z(_03434_));
 MUX2_X1 _20032_ (.A(_03433_),
    .B(_03434_),
    .S(_10763_),
    .Z(_03435_));
 MUX2_X1 _20033_ (.A(_01146_),
    .B(_01148_),
    .S(_11614_),
    .Z(_03436_));
 MUX2_X1 _20034_ (.A(_01130_),
    .B(_01132_),
    .S(_11614_),
    .Z(_03437_));
 MUX2_X1 _20035_ (.A(_03436_),
    .B(_03437_),
    .S(_10763_),
    .Z(_03438_));
 MUX2_X1 _20036_ (.A(_03435_),
    .B(_03438_),
    .S(_10711_),
    .Z(_03439_));
 NAND2_X1 _20037_ (.A1(_11344_),
    .A2(_03439_),
    .ZN(_03440_));
 INV_X1 _20038_ (.A(_01127_),
    .ZN(_03441_));
 NOR2_X1 _20039_ (.A1(_11502_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .ZN(_03442_));
 AOI21_X1 _20040_ (.A(_03442_),
    .B1(_01128_),
    .B2(net378),
    .ZN(_03443_));
 AOI221_X2 _20041_ (.A(_11134_),
    .B1(_03441_),
    .B2(_11137_),
    .C1(_03443_),
    .C2(_11316_),
    .ZN(_03444_));
 MUX2_X1 _20042_ (.A(_01141_),
    .B(_01143_),
    .S(_11502_),
    .Z(_03445_));
 NOR2_X1 _20043_ (.A1(_10711_),
    .A2(_03445_),
    .ZN(_03446_));
 MUX2_X1 _20044_ (.A(_01142_),
    .B(_01144_),
    .S(_11502_),
    .Z(_03447_));
 NOR2_X1 _20045_ (.A1(_11130_),
    .A2(_03447_),
    .ZN(_03448_));
 NOR3_X1 _20046_ (.A1(_10763_),
    .A2(_03446_),
    .A3(_03448_),
    .ZN(_03449_));
 OAI21_X1 _20047_ (.A(_11388_),
    .B1(_03444_),
    .B2(_03449_),
    .ZN(_03450_));
 AND4_X1 _20048_ (.A1(_03424_),
    .A2(_03432_),
    .A3(_03440_),
    .A4(_03450_),
    .ZN(_03451_));
 BUF_X4 _20049_ (.A(_03451_),
    .Z(_03452_));
 AOI221_X2 _20050_ (.A(_03415_),
    .B1(_03416_),
    .B2(_12351_),
    .C1(_11167_),
    .C2(_03452_),
    .ZN(_15893_));
 INV_X1 _20051_ (.A(_15893_),
    .ZN(_15897_));
 MUX2_X1 _20052_ (.A(_01143_),
    .B(_01147_),
    .S(_10985_),
    .Z(_03453_));
 NOR3_X1 _20053_ (.A1(_11029_),
    .A2(_10990_),
    .A3(_03453_),
    .ZN(_03454_));
 MUX2_X1 _20054_ (.A(_01141_),
    .B(_01145_),
    .S(_10984_),
    .Z(_03455_));
 NOR3_X1 _20055_ (.A1(_11244_),
    .A2(_10990_),
    .A3(_03455_),
    .ZN(_03456_));
 MUX2_X1 _20056_ (.A(_01149_),
    .B(_01153_),
    .S(_10984_),
    .Z(_03457_));
 NOR3_X1 _20057_ (.A1(_11244_),
    .A2(_10991_),
    .A3(_03457_),
    .ZN(_03458_));
 MUX2_X1 _20058_ (.A(_01151_),
    .B(_01155_),
    .S(_10984_),
    .Z(_03459_));
 NOR3_X1 _20059_ (.A1(_11029_),
    .A2(_10991_),
    .A3(_03459_),
    .ZN(_03460_));
 NOR4_X1 _20060_ (.A1(_03454_),
    .A2(_03456_),
    .A3(_03458_),
    .A4(_03460_),
    .ZN(_03461_));
 NAND3_X1 _20061_ (.A1(_11012_),
    .A2(_11051_),
    .A3(_03461_),
    .ZN(_03462_));
 NOR2_X1 _20062_ (.A1(_11063_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .ZN(_03463_));
 AOI21_X1 _20063_ (.A(_03463_),
    .B1(_01128_),
    .B2(_11004_),
    .ZN(_03464_));
 AOI221_X1 _20064_ (.A(_10985_),
    .B1(_03441_),
    .B2(_11030_),
    .C1(_03464_),
    .C2(_10997_),
    .ZN(_03465_));
 MUX2_X1 _20065_ (.A(_01129_),
    .B(_01131_),
    .S(_11063_),
    .Z(_03466_));
 NOR2_X1 _20066_ (.A1(_11025_),
    .A2(_03466_),
    .ZN(_03467_));
 MUX2_X1 _20067_ (.A(_01130_),
    .B(_01132_),
    .S(_11063_),
    .Z(_03468_));
 NOR2_X1 _20068_ (.A1(_11011_),
    .A2(_03468_),
    .ZN(_03469_));
 NOR3_X1 _20069_ (.A1(_11036_),
    .A2(_03467_),
    .A3(_03469_),
    .ZN(_03470_));
 OAI21_X1 _20070_ (.A(_03201_),
    .B1(_03465_),
    .B2(_03470_),
    .ZN(_03471_));
 MUX2_X1 _20071_ (.A(_01150_),
    .B(_01154_),
    .S(_10984_),
    .Z(_03472_));
 MUX2_X1 _20072_ (.A(_01152_),
    .B(_01156_),
    .S(_10984_),
    .Z(_03473_));
 MUX2_X1 _20073_ (.A(_03472_),
    .B(_03473_),
    .S(_11238_),
    .Z(_03474_));
 MUX2_X1 _20074_ (.A(_01142_),
    .B(_01146_),
    .S(_10984_),
    .Z(_03475_));
 MUX2_X1 _20075_ (.A(_01144_),
    .B(_01148_),
    .S(_10984_),
    .Z(_03476_));
 MUX2_X1 _20076_ (.A(_03475_),
    .B(_03476_),
    .S(_11238_),
    .Z(_03477_));
 MUX2_X1 _20077_ (.A(_03474_),
    .B(_03477_),
    .S(_10991_),
    .Z(_03478_));
 NAND3_X1 _20078_ (.A1(_11026_),
    .A2(_11051_),
    .A3(_03478_),
    .ZN(_03479_));
 MUX2_X1 _20079_ (.A(_01135_),
    .B(_01139_),
    .S(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .Z(_03480_));
 MUX2_X1 _20080_ (.A(_01136_),
    .B(_01140_),
    .S(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .Z(_03481_));
 MUX2_X1 _20081_ (.A(_03480_),
    .B(_03481_),
    .S(_10996_),
    .Z(_03482_));
 MUX2_X1 _20082_ (.A(_01133_),
    .B(_01137_),
    .S(_10984_),
    .Z(_03483_));
 MUX2_X1 _20083_ (.A(_01134_),
    .B(_01138_),
    .S(_10984_),
    .Z(_03484_));
 MUX2_X1 _20084_ (.A(_03483_),
    .B(_03484_),
    .S(_10997_),
    .Z(_03485_));
 MUX2_X1 _20085_ (.A(_03482_),
    .B(_03485_),
    .S(_11029_),
    .Z(_03486_));
 NAND3_X1 _20086_ (.A1(_11021_),
    .A2(_10979_),
    .A3(_03486_),
    .ZN(_03487_));
 AND4_X4 _20087_ (.A1(_03462_),
    .A2(_03471_),
    .A3(_03479_),
    .A4(_03487_),
    .ZN(_03488_));
 MUX2_X1 _20088_ (.A(\cs_registers_i.pc_id_i[31] ),
    .B(_03488_),
    .S(_10977_),
    .Z(_03489_));
 AOI22_X4 _20089_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(_10819_),
    .B1(_11111_),
    .B2(_03489_),
    .ZN(_15894_));
 BUF_X2 _20090_ (.A(_00179_),
    .Z(_03490_));
 BUF_X4 _20091_ (.A(_00178_),
    .Z(_03491_));
 CLKBUF_X3 _20092_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Z(_03492_));
 BUF_X4 _20093_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .Z(_03493_));
 NOR2_X4 _20094_ (.A1(_03492_),
    .A2(_03493_),
    .ZN(_03494_));
 AND3_X2 _20095_ (.A1(_03490_),
    .A2(_03491_),
    .A3(_03494_),
    .ZN(_03495_));
 NAND2_X1 _20096_ (.A1(_03452_),
    .A2(_03495_),
    .ZN(_03496_));
 NAND3_X4 _20097_ (.A1(_03490_),
    .A2(_03491_),
    .A3(_03494_),
    .ZN(_03497_));
 INV_X4 _20098_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .ZN(_03498_));
 BUF_X2 _20099_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .Z(_03499_));
 OAI221_X1 _20100_ (.A(_03497_),
    .B1(_03494_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .C1(_03498_),
    .C2(_03499_),
    .ZN(_03500_));
 NOR2_X1 _20101_ (.A1(_03491_),
    .A2(_03488_),
    .ZN(_03501_));
 OAI21_X1 _20102_ (.A(_03496_),
    .B1(_03500_),
    .B2(_03501_),
    .ZN(_03502_));
 CLKBUF_X3 _20103_ (.A(_01157_),
    .Z(_03503_));
 BUF_X4 _20104_ (.A(_03494_),
    .Z(_03504_));
 NOR2_X1 _20105_ (.A1(_03503_),
    .A2(_03504_),
    .ZN(_03505_));
 XNOR2_X1 _20106_ (.A(_03502_),
    .B(_03505_),
    .ZN(_03506_));
 NOR2_X1 _20107_ (.A1(_11865_),
    .A2(_03506_),
    .ZN(_03507_));
 NOR2_X4 _20108_ (.A1(_11929_),
    .A2(_11918_),
    .ZN(_03508_));
 XOR2_X2 _20109_ (.A(_15893_),
    .B(_15894_),
    .Z(_03509_));
 XNOR2_X1 _20110_ (.A(_03508_),
    .B(_03509_),
    .ZN(_03510_));
 AOI21_X1 _20111_ (.A(_03507_),
    .B1(_03510_),
    .B2(_11865_),
    .ZN(_03511_));
 INV_X1 _20112_ (.A(_15891_),
    .ZN(_03512_));
 INV_X1 _20113_ (.A(_03330_),
    .ZN(_03513_));
 AOI221_X2 _20114_ (.A(_15887_),
    .B1(_03149_),
    .B2(_03328_),
    .C1(_03513_),
    .C2(_03319_),
    .ZN(_03514_));
 INV_X1 _20115_ (.A(_15892_),
    .ZN(_03515_));
 OAI21_X2 _20116_ (.A(_03512_),
    .B1(_03514_),
    .B2(_03515_),
    .ZN(_03516_));
 XOR2_X2 _20117_ (.A(_03511_),
    .B(_03516_),
    .Z(_03517_));
 BUF_X1 rebuffer14 (.A(_03517_),
    .Z(net288));
 AOI21_X2 _20119_ (.A(_15883_),
    .B1(_03334_),
    .B2(_03321_),
    .ZN(_03518_));
 INV_X1 _20120_ (.A(_03518_),
    .ZN(_03519_));
 AOI21_X2 _20121_ (.A(_15887_),
    .B1(_03519_),
    .B2(_03319_),
    .ZN(_03520_));
 NAND3_X1 _20122_ (.A1(_03146_),
    .A2(_03156_),
    .A3(_03328_),
    .ZN(_03521_));
 OAI21_X2 _20123_ (.A(_03520_),
    .B1(_03521_),
    .B2(_13612_),
    .ZN(_03522_));
 XNOR2_X2 _20124_ (.A(_03522_),
    .B(_03515_),
    .ZN(\alu_adder_result_ex[30] ));
 INV_X1 _20125_ (.A(_15894_),
    .ZN(_15898_));
 INV_X4 _20126_ (.A(_10768_),
    .ZN(_03523_));
 CLKBUF_X3 _20127_ (.A(_10767_),
    .Z(_03524_));
 NOR2_X2 _20128_ (.A1(_10771_),
    .A2(_03524_),
    .ZN(_03525_));
 INV_X2 _20129_ (.A(_03525_),
    .ZN(_03526_));
 NOR2_X4 _20130_ (.A1(_03523_),
    .A2(_03526_),
    .ZN(_03527_));
 NAND2_X2 _20131_ (.A1(net59),
    .A2(_03527_),
    .ZN(_03528_));
 NOR2_X2 _20132_ (.A1(net33),
    .A2(\load_store_unit_i.lsu_err_q ),
    .ZN(_03529_));
 NOR3_X2 _20133_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_03528_),
    .A3(_03529_),
    .ZN(\id_stage_i.controller_i.load_err_d ));
 NOR3_X2 _20134_ (.A1(_01159_),
    .A2(_03528_),
    .A3(_03529_),
    .ZN(\id_stage_i.controller_i.store_err_d ));
 CLKBUF_X3 _20135_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Z(_03530_));
 BUF_X4 _20136_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .Z(_03531_));
 INV_X4 _20137_ (.A(_03531_),
    .ZN(_03532_));
 INV_X2 _20138_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .ZN(_03533_));
 BUF_X4 _20139_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_03534_));
 NAND2_X1 _20140_ (.A1(_03533_),
    .A2(_03534_),
    .ZN(_03535_));
 NOR3_X4 _20141_ (.A1(_03530_),
    .A2(_03532_),
    .A3(_03535_),
    .ZN(_03536_));
 NAND2_X4 _20142_ (.A1(_11294_),
    .A2(_11326_),
    .ZN(_03537_));
 INV_X1 _20143_ (.A(_15906_),
    .ZN(_03538_));
 AOI21_X1 _20144_ (.A(_15903_),
    .B1(_03538_),
    .B2(_15904_),
    .ZN(_03539_));
 AOI21_X1 _20145_ (.A(_03539_),
    .B1(_15907_),
    .B2(_15904_),
    .ZN(_03540_));
 INV_X1 _20146_ (.A(_03540_),
    .ZN(_03541_));
 NOR4_X4 _20147_ (.A1(_11630_),
    .A2(_11638_),
    .A3(_11646_),
    .A4(_11647_),
    .ZN(_03542_));
 NOR4_X4 _20148_ (.A1(_11705_),
    .A2(_11713_),
    .A3(_11721_),
    .A4(_11722_),
    .ZN(_03543_));
 NAND2_X1 _20149_ (.A1(_10884_),
    .A2(_10805_),
    .ZN(_03544_));
 OAI33_X1 _20150_ (.A1(_10805_),
    .A2(_03542_),
    .A3(_03543_),
    .B1(_03544_),
    .B2(_11650_),
    .B3(_11649_),
    .ZN(_03545_));
 NAND2_X2 _20151_ (.A1(_16309_),
    .A2(net14),
    .ZN(_03546_));
 NOR2_X1 _20152_ (.A1(_11478_),
    .A2(_03546_),
    .ZN(_03547_));
 INV_X1 _20153_ (.A(_11489_),
    .ZN(_03548_));
 CLKBUF_X2 _20154_ (.A(_15914_),
    .Z(_03549_));
 INV_X1 _20155_ (.A(_03549_),
    .ZN(_03550_));
 NAND2_X4 _20156_ (.A1(_03548_),
    .A2(_03550_),
    .ZN(_03551_));
 CLKBUF_X3 _20157_ (.A(_15917_),
    .Z(_03552_));
 INV_X1 _20158_ (.A(_03552_),
    .ZN(_03553_));
 BUF_X4 _20159_ (.A(_15922_),
    .Z(_03554_));
 INV_X2 _20160_ (.A(_03554_),
    .ZN(_03555_));
 NAND2_X2 _20161_ (.A1(_03553_),
    .A2(_03555_),
    .ZN(_03556_));
 NOR2_X4 _20162_ (.A1(_03551_),
    .A2(_03556_),
    .ZN(_03557_));
 AOI21_X2 _20163_ (.A(_11536_),
    .B1(_11537_),
    .B2(_11481_),
    .ZN(_03558_));
 OAI21_X2 _20164_ (.A(_11573_),
    .B1(_11610_),
    .B2(_11570_),
    .ZN(_03559_));
 NAND2_X4 _20165_ (.A1(_03558_),
    .A2(_03559_),
    .ZN(_03560_));
 BUF_X4 _20166_ (.A(_11533_),
    .Z(_16278_));
 NAND2_X4 _20167_ (.A1(_11328_),
    .A2(_16278_),
    .ZN(_03561_));
 NOR4_X4 _20168_ (.A1(_16326_),
    .A2(_03557_),
    .A3(_03560_),
    .A4(_03561_),
    .ZN(_03562_));
 NAND3_X2 _20169_ (.A1(_11492_),
    .A2(_03547_),
    .A3(_03562_),
    .ZN(_03563_));
 BUF_X4 _20170_ (.A(\cs_registers_i.debug_mode_i ),
    .Z(_03564_));
 OAI21_X4 _20171_ (.A(_03541_),
    .B1(_03563_),
    .B2(_03564_),
    .ZN(_03565_));
 OAI21_X4 _20172_ (.A(_16298_),
    .B1(net10),
    .B2(_10819_),
    .ZN(_03566_));
 NAND2_X1 _20173_ (.A1(_10888_),
    .A2(_10805_),
    .ZN(_03567_));
 OAI33_X1 _20174_ (.A1(_10805_),
    .A2(_03542_),
    .A3(_11724_),
    .B1(_03567_),
    .B2(_11650_),
    .B3(_11649_),
    .ZN(_03568_));
 NAND2_X4 _20175_ (.A1(_16309_),
    .A2(net13),
    .ZN(_03569_));
 NOR2_X2 _20176_ (.A1(_11285_),
    .A2(_11289_),
    .ZN(_03570_));
 AND3_X4 _20177_ (.A1(_11282_),
    .A2(_03570_),
    .A3(_11326_),
    .ZN(_03571_));
 NAND2_X2 _20178_ (.A1(_03571_),
    .A2(_11534_),
    .ZN(_03572_));
 NOR4_X4 _20179_ (.A1(_16330_),
    .A2(_03566_),
    .A3(_03569_),
    .A4(_03572_),
    .ZN(_03573_));
 NAND2_X1 _20180_ (.A1(_03549_),
    .A2(_03571_),
    .ZN(_03574_));
 AOI211_X2 _20181_ (.A(_11477_),
    .B(_03574_),
    .C1(_11379_),
    .C2(_11434_),
    .ZN(_03575_));
 BUF_X4 _20182_ (.A(_03548_),
    .Z(_03576_));
 NOR2_X2 _20183_ (.A1(_03552_),
    .A2(_03554_),
    .ZN(_03577_));
 NAND2_X2 _20184_ (.A1(_03576_),
    .A2(_03577_),
    .ZN(_03578_));
 NAND3_X2 _20185_ (.A1(_11282_),
    .A2(_03570_),
    .A3(_11326_),
    .ZN(_03579_));
 BUF_X4 _20186_ (.A(_03579_),
    .Z(_03580_));
 NOR2_X1 _20187_ (.A1(_03580_),
    .A2(_03557_),
    .ZN(_03581_));
 MUX2_X1 _20188_ (.A(_03578_),
    .B(_03581_),
    .S(_11477_),
    .Z(_03582_));
 OAI21_X4 _20189_ (.A(_03573_),
    .B1(_03575_),
    .B2(_03582_),
    .ZN(_03583_));
 NOR2_X4 _20190_ (.A1(_03560_),
    .A2(_03569_),
    .ZN(_03584_));
 NOR2_X2 _20191_ (.A1(_03580_),
    .A2(_16330_),
    .ZN(_03585_));
 NAND2_X2 _20192_ (.A1(_03584_),
    .A2(_03585_),
    .ZN(_03586_));
 NOR2_X1 _20193_ (.A1(_16278_),
    .A2(_03557_),
    .ZN(_03587_));
 OAI21_X4 _20194_ (.A(_11328_),
    .B1(_11477_),
    .B2(_16278_),
    .ZN(_03588_));
 BUF_X4 _20195_ (.A(_03550_),
    .Z(_03589_));
 NOR3_X1 _20196_ (.A1(_03589_),
    .A2(_11477_),
    .A3(_16278_),
    .ZN(_03590_));
 BUF_X8 _20197_ (.A(_11479_),
    .Z(_03591_));
 AOI21_X2 _20198_ (.A(_03591_),
    .B1(_11379_),
    .B2(_11434_),
    .ZN(_03592_));
 AOI222_X2 _20199_ (.A1(_15909_),
    .A2(_03587_),
    .B1(_03578_),
    .B2(_03588_),
    .C1(_03590_),
    .C2(_03592_),
    .ZN(_03593_));
 OAI21_X4 _20200_ (.A(_03583_),
    .B1(_03586_),
    .B2(_03593_),
    .ZN(_03594_));
 AOI21_X4 _20201_ (.A(_03580_),
    .B1(_11434_),
    .B2(_11378_),
    .ZN(_03595_));
 NOR2_X2 _20202_ (.A1(_11489_),
    .A2(_03549_),
    .ZN(_03596_));
 AND3_X1 _20203_ (.A1(_03571_),
    .A2(_16309_),
    .A3(net14),
    .ZN(_03597_));
 NOR4_X1 _20204_ (.A1(_11221_),
    .A2(_03580_),
    .A3(net10),
    .A4(_16298_),
    .ZN(_03598_));
 NAND4_X1 _20205_ (.A1(_11476_),
    .A2(_16282_),
    .A3(_03597_),
    .A4(_03598_),
    .ZN(_03599_));
 NOR4_X1 _20206_ (.A1(_03595_),
    .A2(_16326_),
    .A3(_03596_),
    .A4(_03599_),
    .ZN(_03600_));
 OR3_X2 _20207_ (.A1(_16330_),
    .A2(_03566_),
    .A3(_03572_),
    .ZN(_03601_));
 AOI21_X2 _20208_ (.A(_10814_),
    .B1(_11334_),
    .B2(_11333_),
    .ZN(_03602_));
 NOR3_X4 _20209_ (.A1(_11122_),
    .A2(_11331_),
    .A3(_03602_),
    .ZN(_03603_));
 OR4_X4 _20210_ (.A1(_03576_),
    .A2(_11435_),
    .A3(_03579_),
    .A4(_03603_),
    .ZN(_03604_));
 NAND2_X1 _20211_ (.A1(_16270_),
    .A2(_03597_),
    .ZN(_03605_));
 NAND2_X1 _20212_ (.A1(_03596_),
    .A2(_03577_),
    .ZN(_03606_));
 AND2_X2 _20213_ (.A1(_16309_),
    .A2(net13),
    .ZN(_03607_));
 NAND2_X1 _20214_ (.A1(_03606_),
    .A2(_03607_),
    .ZN(_03608_));
 NAND2_X2 _20215_ (.A1(_03571_),
    .A2(_16278_),
    .ZN(_03609_));
 OR3_X2 _20216_ (.A1(_11770_),
    .A2(_03560_),
    .A3(_03609_),
    .ZN(_03610_));
 AOI21_X1 _20217_ (.A(_11477_),
    .B1(_11434_),
    .B2(_11379_),
    .ZN(_03611_));
 OAI33_X1 _20218_ (.A1(_03601_),
    .A2(_03604_),
    .A3(_03605_),
    .B1(_03608_),
    .B2(_03610_),
    .B3(_03611_),
    .ZN(_03612_));
 OAI21_X1 _20219_ (.A(_10838_),
    .B1(_11121_),
    .B2(_11427_),
    .ZN(_03613_));
 INV_X1 _20220_ (.A(_00139_),
    .ZN(_03614_));
 MUX2_X1 _20221_ (.A(_10758_),
    .B(_03614_),
    .S(_10859_),
    .Z(_03615_));
 AOI21_X1 _20222_ (.A(_10804_),
    .B1(_11481_),
    .B2(_03615_),
    .ZN(_03616_));
 NAND3_X1 _20223_ (.A1(_11308_),
    .A2(_11486_),
    .A3(_11487_),
    .ZN(_03617_));
 AOI211_X2 _20224_ (.A(_11479_),
    .B(_03613_),
    .C1(_03616_),
    .C2(_03617_),
    .ZN(_03618_));
 OR2_X1 _20225_ (.A1(_03557_),
    .A2(_03618_),
    .ZN(_03619_));
 NOR3_X2 _20226_ (.A1(_11489_),
    .A2(_03591_),
    .A3(_11378_),
    .ZN(_03620_));
 NAND3_X4 _20227_ (.A1(_16286_),
    .A2(_16298_),
    .A3(_16330_),
    .ZN(_03621_));
 OR3_X4 _20228_ (.A1(_11477_),
    .A2(_03569_),
    .A3(_03572_),
    .ZN(_03622_));
 NOR4_X1 _20229_ (.A1(_03619_),
    .A2(_03620_),
    .A3(_03621_),
    .A4(_03622_),
    .ZN(_03623_));
 NAND4_X1 _20230_ (.A1(_11477_),
    .A2(_16309_),
    .A3(net14),
    .A4(_03606_),
    .ZN(_03624_));
 AOI21_X2 _20231_ (.A(_11534_),
    .B1(_11379_),
    .B2(_11328_),
    .ZN(_03625_));
 OR4_X4 _20232_ (.A1(_03580_),
    .A2(_11770_),
    .A3(_03566_),
    .A4(_03569_),
    .ZN(_03626_));
 OAI21_X1 _20233_ (.A(_03548_),
    .B1(_03589_),
    .B2(_16278_),
    .ZN(_03627_));
 OAI211_X2 _20234_ (.A(_11476_),
    .B(_03627_),
    .C1(_03580_),
    .C2(_11434_),
    .ZN(_03628_));
 OAI33_X1 _20235_ (.A1(_03595_),
    .A2(_03610_),
    .A3(_03624_),
    .B1(_03625_),
    .B2(_03626_),
    .B3(_03628_),
    .ZN(_03629_));
 OR4_X1 _20236_ (.A1(_03600_),
    .A2(_03612_),
    .A3(_03623_),
    .A4(_03629_),
    .ZN(_03630_));
 BUF_X4 _20237_ (.A(_03591_),
    .Z(_03631_));
 NOR2_X2 _20238_ (.A1(_16253_),
    .A2(_11434_),
    .ZN(_03632_));
 NAND2_X2 _20239_ (.A1(_03589_),
    .A2(_03555_),
    .ZN(_03633_));
 NOR2_X2 _20240_ (.A1(_11379_),
    .A2(_11435_),
    .ZN(_03634_));
 AOI22_X2 _20241_ (.A1(_11489_),
    .A2(_03632_),
    .B1(_03633_),
    .B2(_03634_),
    .ZN(_03635_));
 BUF_X4 _20242_ (.A(_03549_),
    .Z(_03636_));
 NOR2_X1 _20243_ (.A1(_03636_),
    .A2(_03554_),
    .ZN(_03637_));
 AOI22_X1 _20244_ (.A1(_16266_),
    .A2(_11478_),
    .B1(_03637_),
    .B2(_03618_),
    .ZN(_03638_));
 OAI22_X1 _20245_ (.A1(_11329_),
    .A2(_16270_),
    .B1(_03638_),
    .B2(_16253_),
    .ZN(_03639_));
 NAND3_X4 _20246_ (.A1(_11328_),
    .A2(_16253_),
    .A3(_11434_),
    .ZN(_03640_));
 AOI21_X1 _20247_ (.A(_11489_),
    .B1(_03633_),
    .B2(_03640_),
    .ZN(_03641_));
 OAI221_X2 _20248_ (.A(_03553_),
    .B1(_03631_),
    .B2(_03635_),
    .C1(_03639_),
    .C2(_03641_),
    .ZN(_03642_));
 NOR2_X1 _20249_ (.A1(_03609_),
    .A2(_03626_),
    .ZN(_03643_));
 AOI211_X2 _20250_ (.A(_03594_),
    .B(_03630_),
    .C1(_03642_),
    .C2(_03643_),
    .ZN(_03644_));
 INV_X1 _20251_ (.A(_16322_),
    .ZN(_16318_));
 NAND2_X2 _20252_ (.A1(_16318_),
    .A2(_16326_),
    .ZN(_03645_));
 CLKBUF_X2 _20253_ (.A(_15929_),
    .Z(_03646_));
 CLKBUF_X3 _20254_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .Z(_03647_));
 INV_X2 _20255_ (.A(_03647_),
    .ZN(_03648_));
 INV_X4 _20256_ (.A(_03534_),
    .ZN(_03649_));
 NOR3_X4 _20257_ (.A1(_03531_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A3(_03649_),
    .ZN(_03650_));
 AND2_X1 _20258_ (.A1(_03530_),
    .A2(_03650_),
    .ZN(_03651_));
 BUF_X4 _20259_ (.A(_03651_),
    .Z(_03652_));
 NAND3_X4 _20260_ (.A1(_10794_),
    .A2(_03648_),
    .A3(_03652_),
    .ZN(_03653_));
 OR3_X2 _20261_ (.A1(_03646_),
    .A2(_03580_),
    .A3(_03653_),
    .ZN(_03654_));
 NOR2_X1 _20262_ (.A1(_03645_),
    .A2(_03654_),
    .ZN(_03655_));
 NOR4_X1 _20263_ (.A1(_03537_),
    .A2(_03565_),
    .A3(_03644_),
    .A4(_03655_),
    .ZN(_03656_));
 INV_X1 _20264_ (.A(_01161_),
    .ZN(_03657_));
 OAI21_X1 _20265_ (.A(_03657_),
    .B1(_11282_),
    .B2(_03537_),
    .ZN(_03658_));
 NOR2_X1 _20266_ (.A1(_03656_),
    .A2(_03658_),
    .ZN(_03659_));
 BUF_X1 _20267_ (.A(\cs_registers_i.priv_lvl_q[0] ),
    .Z(_03660_));
 CLKBUF_X2 _20268_ (.A(\cs_registers_i.priv_lvl_q[1] ),
    .Z(_03661_));
 NAND2_X2 _20269_ (.A1(_03660_),
    .A2(_03661_),
    .ZN(_03662_));
 NOR2_X2 _20270_ (.A1(_11280_),
    .A2(_10972_),
    .ZN(_03663_));
 NAND3_X2 _20271_ (.A1(_11319_),
    .A2(_11320_),
    .A3(_03663_),
    .ZN(_03664_));
 NOR4_X4 _20272_ (.A1(_10875_),
    .A2(_01161_),
    .A3(_11317_),
    .A4(_03664_),
    .ZN(_03665_));
 NAND3_X1 _20273_ (.A1(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(_03662_),
    .A3(_03665_),
    .ZN(_03666_));
 AND3_X2 _20274_ (.A1(_10794_),
    .A2(_10917_),
    .A3(_10967_),
    .ZN(_03667_));
 NAND3_X4 _20275_ (.A1(_10971_),
    .A2(_11324_),
    .A3(_03667_),
    .ZN(_03668_));
 NAND2_X4 _20276_ (.A1(net300),
    .A2(_11303_),
    .ZN(_03669_));
 NOR2_X1 _20277_ (.A1(_03564_),
    .A2(_03669_),
    .ZN(_03670_));
 AOI21_X1 _20278_ (.A(_03670_),
    .B1(_03662_),
    .B2(_11319_),
    .ZN(_03671_));
 OAI21_X2 _20279_ (.A(_03666_),
    .B1(_03668_),
    .B2(_03671_),
    .ZN(_03672_));
 NOR2_X1 _20280_ (.A1(_03659_),
    .A2(_03672_),
    .ZN(_03673_));
 NOR2_X1 _20281_ (.A1(_03536_),
    .A2(_03673_),
    .ZN(\id_stage_i.controller_i.illegal_insn_d ));
 NAND2_X2 _20282_ (.A1(_11319_),
    .A2(_11320_),
    .ZN(_03674_));
 NAND3_X4 _20283_ (.A1(_10794_),
    .A2(_10917_),
    .A3(_10967_),
    .ZN(_03675_));
 NAND2_X2 _20284_ (.A1(_10736_),
    .A2(_10877_),
    .ZN(_03676_));
 NOR4_X2 _20285_ (.A1(_11280_),
    .A2(_03674_),
    .A3(_03675_),
    .A4(_03676_),
    .ZN(_03677_));
 NAND2_X2 _20286_ (.A1(_10711_),
    .A2(_03677_),
    .ZN(_03678_));
 NOR2_X1 _20287_ (.A1(_03664_),
    .A2(_03676_),
    .ZN(_03679_));
 AOI21_X1 _20288_ (.A(_03647_),
    .B1(_03679_),
    .B2(_12367_),
    .ZN(_03680_));
 OAI21_X2 _20289_ (.A(_03678_),
    .B1(_03680_),
    .B2(_10810_),
    .ZN(_03681_));
 NOR3_X1 _20290_ (.A1(_03659_),
    .A2(_03672_),
    .A3(_03681_),
    .ZN(_03682_));
 NOR2_X1 _20291_ (.A1(_03536_),
    .A2(_03682_),
    .ZN(\id_stage_i.controller_i.exc_req_d ));
 CLKBUF_X3 _20292_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .Z(_03683_));
 AND2_X1 _20293_ (.A1(net414),
    .A2(_11863_),
    .ZN(_03684_));
 NAND3_X4 _20294_ (.A1(_11878_),
    .A2(_10955_),
    .A3(_03684_),
    .ZN(_03685_));
 BUF_X4 _20295_ (.A(_03685_),
    .Z(_03686_));
 INV_X2 _20296_ (.A(_03653_),
    .ZN(_03687_));
 NAND3_X4 _20297_ (.A1(_11294_),
    .A2(_11326_),
    .A3(_03687_),
    .ZN(_03688_));
 NOR2_X4 _20298_ (.A1(_03686_),
    .A2(_03688_),
    .ZN(_03689_));
 NAND2_X1 _20299_ (.A1(_03683_),
    .A2(_03689_),
    .ZN(_03690_));
 CLKBUF_X3 _20300_ (.A(_03690_),
    .Z(_03691_));
 CLKBUF_X3 _20301_ (.A(_03691_),
    .Z(_03692_));
 BUF_X4 _20302_ (.A(_15948_),
    .Z(_03693_));
 BUF_X4 _20303_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .Z(_03694_));
 BUF_X4 _20304_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Z(_03695_));
 NOR2_X1 _20305_ (.A1(_03694_),
    .A2(_03695_),
    .ZN(_03696_));
 AND3_X1 _20306_ (.A1(_01162_),
    .A2(_03693_),
    .A3(_03696_),
    .ZN(_03697_));
 AND2_X1 _20307_ (.A1(_03689_),
    .A2(_03697_),
    .ZN(_03698_));
 INV_X1 _20308_ (.A(_03493_),
    .ZN(_03699_));
 BUF_X4 _20309_ (.A(_03699_),
    .Z(_03700_));
 OAI21_X1 _20310_ (.A(_03692_),
    .B1(_03698_),
    .B2(_03700_),
    .ZN(_00005_));
 CLKBUF_X3 _20311_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .Z(_03701_));
 CLKBUF_X3 _20312_ (.A(_03689_),
    .Z(_03702_));
 OR4_X2 _20313_ (.A1(\alu_adder_result_ex[27] ),
    .A2(\alu_adder_result_ex[29] ),
    .A3(\alu_adder_result_ex[28] ),
    .A4(\alu_adder_result_ex[30] ),
    .ZN(_03703_));
 CLKBUF_X3 _20314_ (.A(_16507_),
    .Z(_03704_));
 INV_X1 _20315_ (.A(_03704_),
    .ZN(_03705_));
 OAI21_X1 _20316_ (.A(_15788_),
    .B1(_15783_),
    .B2(_12154_),
    .ZN(_03706_));
 NAND2_X1 _20317_ (.A1(_12158_),
    .A2(_03706_),
    .ZN(_03707_));
 XOR2_X2 _20318_ (.A(_12142_),
    .B(_03707_),
    .Z(\alu_adder_result_ex[5] ));
 XOR2_X2 _20319_ (.A(_12148_),
    .B(_12153_),
    .Z(\alu_adder_result_ex[3] ));
 OR4_X2 _20320_ (.A1(_03705_),
    .A2(\alu_adder_result_ex[7] ),
    .A3(\alu_adder_result_ex[5] ),
    .A4(\alu_adder_result_ex[3] ),
    .ZN(_03708_));
 NOR3_X1 _20321_ (.A1(\alu_adder_result_ex[11] ),
    .A2(\alu_adder_result_ex[13] ),
    .A3(_03708_),
    .ZN(_03709_));
 NAND3_X1 _20322_ (.A1(_12271_),
    .A2(_12881_),
    .A3(_03709_),
    .ZN(_03710_));
 NOR2_X1 _20323_ (.A1(_12151_),
    .A2(_12166_),
    .ZN(_03711_));
 MUX2_X1 _20324_ (.A(_03711_),
    .B(_12151_),
    .S(_12181_),
    .Z(_03712_));
 NAND3_X1 _20325_ (.A1(_12152_),
    .A2(_12168_),
    .A3(_12167_),
    .ZN(_03713_));
 AOI21_X2 _20326_ (.A(_03713_),
    .B1(_12177_),
    .B2(_12176_),
    .ZN(_03714_));
 NOR4_X2 _20327_ (.A1(_12152_),
    .A2(net360),
    .A3(_11918_),
    .A4(_12171_),
    .ZN(_03715_));
 NOR3_X4 _20328_ (.A1(_03712_),
    .A2(_03714_),
    .A3(_03715_),
    .ZN(\alu_adder_result_ex[2] ));
 NOR4_X1 _20329_ (.A1(\alu_adder_result_ex[10] ),
    .A2(\alu_adder_result_ex[12] ),
    .A3(_03710_),
    .A4(\alu_adder_result_ex[2] ),
    .ZN(_03716_));
 OAI21_X1 _20330_ (.A(_12149_),
    .B1(_12168_),
    .B2(_12152_),
    .ZN(_03717_));
 AOI21_X2 _20331_ (.A(_15783_),
    .B1(_03717_),
    .B2(_12148_),
    .ZN(_03718_));
 NAND3_X1 _20332_ (.A1(_12151_),
    .A2(_12148_),
    .A3(_12166_),
    .ZN(_03719_));
 NAND3_X1 _20333_ (.A1(net348),
    .A2(_03718_),
    .A3(_03719_),
    .ZN(_03720_));
 OAI21_X1 _20334_ (.A(_03720_),
    .B1(_03718_),
    .B2(net348),
    .ZN(_03721_));
 NAND3_X1 _20335_ (.A1(net348),
    .A2(_11864_),
    .A3(_03718_),
    .ZN(_03722_));
 AOI21_X1 _20336_ (.A(_03722_),
    .B1(_12177_),
    .B2(_12176_),
    .ZN(_03723_));
 NOR2_X1 _20337_ (.A1(net348),
    .A2(_03719_),
    .ZN(_03724_));
 AOI211_X2 _20338_ (.A(_03721_),
    .B(_03723_),
    .C1(_14464_),
    .C2(_03724_),
    .ZN(_03725_));
 INV_X4 _20339_ (.A(_03725_),
    .ZN(\alu_adder_result_ex[4] ));
 NOR4_X2 _20340_ (.A1(net8),
    .A2(\alu_adder_result_ex[8] ),
    .A3(\alu_adder_result_ex[21] ),
    .A4(\alu_adder_result_ex[4] ),
    .ZN(_03726_));
 NOR4_X2 _20341_ (.A1(\alu_adder_result_ex[15] ),
    .A2(\alu_adder_result_ex[14] ),
    .A3(\alu_adder_result_ex[18] ),
    .A4(\alu_adder_result_ex[23] ),
    .ZN(_03727_));
 NAND3_X2 _20342_ (.A1(_03716_),
    .A2(_03726_),
    .A3(_03727_),
    .ZN(_03728_));
 NOR4_X2 _20343_ (.A1(\alu_adder_result_ex[16] ),
    .A2(\alu_adder_result_ex[19] ),
    .A3(\alu_adder_result_ex[22] ),
    .A4(\alu_adder_result_ex[25] ),
    .ZN(_03729_));
 NAND2_X2 _20344_ (.A1(net391),
    .A2(_03729_),
    .ZN(_03730_));
 OR3_X2 _20345_ (.A1(\alu_adder_result_ex[20] ),
    .A2(\alu_adder_result_ex[24] ),
    .A3(_03517_),
    .ZN(_03731_));
 OR4_X4 _20346_ (.A1(_03703_),
    .A2(_03728_),
    .A3(_03730_),
    .A4(_03731_),
    .ZN(_03732_));
 NAND3_X1 _20347_ (.A1(_03701_),
    .A2(_03702_),
    .A3(_03732_),
    .ZN(_03733_));
 CLKBUF_X2 _20348_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Z(_03734_));
 INV_X1 _20349_ (.A(_03734_),
    .ZN(_03735_));
 OAI21_X1 _20350_ (.A(_03733_),
    .B1(_03702_),
    .B2(_03735_),
    .ZN(_00004_));
 NAND2_X2 _20351_ (.A1(net414),
    .A2(_11863_),
    .ZN(_03736_));
 NOR3_X4 _20352_ (.A1(_10869_),
    .A2(_10872_),
    .A3(_03736_),
    .ZN(_03737_));
 BUF_X4 _20353_ (.A(_03737_),
    .Z(_03738_));
 NOR2_X4 _20354_ (.A1(_03537_),
    .A2(_03653_),
    .ZN(_03739_));
 NAND2_X4 _20355_ (.A1(_03738_),
    .A2(_03739_),
    .ZN(_03740_));
 NAND2_X1 _20356_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .A2(_03740_),
    .ZN(_03741_));
 BUF_X4 _20357_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Z(_03742_));
 BUF_X4 _20358_ (.A(_03742_),
    .Z(_03743_));
 BUF_X4 _20359_ (.A(_03743_),
    .Z(_03744_));
 NOR4_X4 _20360_ (.A1(_03703_),
    .A2(_03728_),
    .A3(_03730_),
    .A4(_03731_),
    .ZN(_03745_));
 AOI21_X1 _20361_ (.A(_03744_),
    .B1(_03701_),
    .B2(_03745_),
    .ZN(_03746_));
 OAI21_X1 _20362_ (.A(_03741_),
    .B1(_03746_),
    .B2(_03740_),
    .ZN(_00003_));
 AND2_X2 _20363_ (.A1(_10828_),
    .A2(_10869_),
    .ZN(_03747_));
 OAI21_X2 _20364_ (.A(_10826_),
    .B1(_10885_),
    .B2(_03747_),
    .ZN(_03748_));
 AND2_X1 _20365_ (.A1(_12276_),
    .A2(_03748_),
    .ZN(_03749_));
 CLKBUF_X3 _20366_ (.A(_03749_),
    .Z(_03750_));
 CLKBUF_X2 _20367_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Z(_03751_));
 BUF_X4 _20368_ (.A(_03751_),
    .Z(_03752_));
 INV_X1 _20369_ (.A(_03752_),
    .ZN(_03753_));
 OAI21_X1 _20370_ (.A(_01163_),
    .B1(_03750_),
    .B2(_03753_),
    .ZN(_03754_));
 BUF_X4 _20371_ (.A(_12276_),
    .Z(_03755_));
 XNOR2_X2 _20372_ (.A(_10828_),
    .B(_10951_),
    .ZN(_03756_));
 NAND3_X4 _20373_ (.A1(_11878_),
    .A2(_12276_),
    .A3(_03756_),
    .ZN(_03757_));
 INV_X1 _20374_ (.A(_03757_),
    .ZN(_03758_));
 AND2_X1 _20375_ (.A1(_03488_),
    .A2(_03758_),
    .ZN(_03759_));
 BUF_X4 _20376_ (.A(_03759_),
    .Z(_03760_));
 NAND2_X4 _20377_ (.A1(_10826_),
    .A2(_03737_),
    .ZN(_03761_));
 AOI21_X1 _20378_ (.A(_03498_),
    .B1(_03760_),
    .B2(_03761_),
    .ZN(_03762_));
 NOR2_X1 _20379_ (.A1(_10921_),
    .A2(_10869_),
    .ZN(_03763_));
 AOI22_X4 _20380_ (.A1(_10921_),
    .A2(_10849_),
    .B1(_11866_),
    .B2(_03763_),
    .ZN(_03764_));
 NOR2_X4 _20381_ (.A1(_11865_),
    .A2(_03764_),
    .ZN(_03765_));
 NAND2_X4 _20382_ (.A1(_03452_),
    .A2(_03765_),
    .ZN(_03766_));
 NOR3_X1 _20383_ (.A1(_03760_),
    .A2(_03761_),
    .A3(_03766_),
    .ZN(_03767_));
 AOI21_X1 _20384_ (.A(_03767_),
    .B1(_03766_),
    .B2(_03760_),
    .ZN(_03768_));
 OAI21_X1 _20385_ (.A(_03762_),
    .B1(_03768_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .ZN(_03769_));
 INV_X1 _20386_ (.A(_03683_),
    .ZN(_03770_));
 NAND3_X4 _20387_ (.A1(_03498_),
    .A2(_03770_),
    .A3(_03504_),
    .ZN(_03771_));
 OAI21_X1 _20388_ (.A(_03769_),
    .B1(_03771_),
    .B2(_03701_),
    .ZN(_03772_));
 NAND2_X1 _20389_ (.A1(net307),
    .A2(_03772_),
    .ZN(_03773_));
 NAND3_X4 _20390_ (.A1(_03755_),
    .A2(_03739_),
    .A3(_03773_),
    .ZN(_03774_));
 NOR2_X4 _20391_ (.A1(_03738_),
    .A2(_03774_),
    .ZN(_03775_));
 MUX2_X1 _20392_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .B(_03754_),
    .S(_03775_),
    .Z(_00000_));
 BUF_X4 _20393_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Z(_03776_));
 NAND4_X4 _20394_ (.A1(net298),
    .A2(_10871_),
    .A3(_11863_),
    .A4(_03748_),
    .ZN(_03777_));
 BUF_X2 _20395_ (.A(_03777_),
    .Z(_03778_));
 NOR2_X2 _20396_ (.A1(_03753_),
    .A2(_03778_),
    .ZN(_03779_));
 MUX2_X1 _20397_ (.A(_03776_),
    .B(_03779_),
    .S(_03775_),
    .Z(_00001_));
 BUF_X4 _20398_ (.A(_03492_),
    .Z(_03780_));
 CLKBUF_X3 _20399_ (.A(_03780_),
    .Z(_03781_));
 NAND2_X1 _20400_ (.A1(_03781_),
    .A2(_03740_),
    .ZN(_03782_));
 BUF_X4 _20401_ (.A(_03493_),
    .Z(_03783_));
 BUF_X4 _20402_ (.A(_03783_),
    .Z(_03784_));
 NAND2_X1 _20403_ (.A1(_03784_),
    .A2(_03697_),
    .ZN(_03785_));
 OAI21_X1 _20404_ (.A(_03782_),
    .B1(_03785_),
    .B2(_03740_),
    .ZN(_00002_));
 BUF_X4 _20405_ (.A(\alu_adder_result_ex[0] ),
    .Z(_03786_));
 INV_X2 _20406_ (.A(_03786_),
    .ZN(_16502_));
 OR2_X1 _20407_ (.A1(_03776_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .ZN(_03787_));
 CLKBUF_X3 _20408_ (.A(_03787_),
    .Z(_03788_));
 BUF_X4 _20409_ (.A(_03788_),
    .Z(_03789_));
 MUX2_X2 _20410_ (.A(net276),
    .B(_12752_),
    .S(_03789_),
    .Z(_03790_));
 INV_X1 _20411_ (.A(_03790_),
    .ZN(_03791_));
 OR2_X1 _20412_ (.A1(_03752_),
    .A2(_03776_),
    .ZN(_03792_));
 BUF_X2 _20413_ (.A(_03792_),
    .Z(_03793_));
 BUF_X4 _20414_ (.A(_03793_),
    .Z(_03794_));
 NAND2_X1 _20415_ (.A1(_12790_),
    .A2(_03794_),
    .ZN(_03795_));
 OAI21_X4 _20416_ (.A(_11195_),
    .B1(_11213_),
    .B2(_11054_),
    .ZN(_03796_));
 OAI21_X4 _20417_ (.A(_03795_),
    .B1(_03794_),
    .B2(_03796_),
    .ZN(_03797_));
 NOR2_X1 _20418_ (.A1(_03791_),
    .A2(_03797_),
    .ZN(_15952_));
 BUF_X4 _20419_ (.A(_03788_),
    .Z(_03798_));
 OR2_X1 _20420_ (.A1(_00217_),
    .A2(_03777_),
    .ZN(_03799_));
 CLKBUF_X3 _20421_ (.A(_00692_),
    .Z(_03800_));
 OAI21_X1 _20422_ (.A(_03799_),
    .B1(_03750_),
    .B2(_03800_),
    .ZN(_03801_));
 AOI22_X1 _20423_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .A2(_03798_),
    .B1(_03801_),
    .B2(_03752_),
    .ZN(_03802_));
 INV_X1 _20424_ (.A(_03802_),
    .ZN(_15953_));
 INV_X1 _20425_ (.A(_03797_),
    .ZN(_03803_));
 OR2_X1 _20426_ (.A1(net301),
    .A2(_03789_),
    .ZN(_03804_));
 NOR2_X4 _20427_ (.A1(_03776_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .ZN(_03805_));
 OAI21_X4 _20428_ (.A(_03804_),
    .B1(_12825_),
    .B2(_03805_),
    .ZN(_03806_));
 NAND2_X1 _20429_ (.A1(_03803_),
    .A2(_03806_),
    .ZN(_14470_));
 CLKBUF_X3 _20430_ (.A(_03797_),
    .Z(_03807_));
 AND2_X1 _20431_ (.A1(net364),
    .A2(_03805_),
    .ZN(_03808_));
 AOI21_X4 _20432_ (.A(_03808_),
    .B1(_03798_),
    .B2(net286),
    .ZN(_03809_));
 NOR2_X1 _20433_ (.A1(_03807_),
    .A2(_03809_),
    .ZN(_15965_));
 BUF_X4 _20434_ (.A(_03806_),
    .Z(_03810_));
 NAND2_X4 _20435_ (.A1(_11050_),
    .A2(_11103_),
    .ZN(_03811_));
 OR2_X2 _20436_ (.A1(_12848_),
    .A2(_12866_),
    .ZN(_03812_));
 MUX2_X1 _20437_ (.A(_03811_),
    .B(_03812_),
    .S(_03793_),
    .Z(_03813_));
 CLKBUF_X3 _20438_ (.A(_03813_),
    .Z(_03814_));
 NAND2_X1 _20439_ (.A1(_03810_),
    .A2(_03814_),
    .ZN(_14474_));
 NOR4_X4 _20440_ (.A1(_11407_),
    .A2(_11416_),
    .A3(_11425_),
    .A4(_11426_),
    .ZN(_03815_));
 NOR2_X1 _20441_ (.A1(_03815_),
    .A2(_03789_),
    .ZN(_03816_));
 AOI21_X4 _20442_ (.A(_03816_),
    .B1(_03789_),
    .B2(_13012_),
    .ZN(_03817_));
 NOR2_X1 _20443_ (.A1(_03807_),
    .A2(_03817_),
    .ZN(_15969_));
 BUF_X4 _20444_ (.A(_03809_),
    .Z(_03818_));
 INV_X2 _20445_ (.A(_03814_),
    .ZN(_03819_));
 NOR2_X1 _20446_ (.A1(_03818_),
    .A2(_03819_),
    .ZN(_15968_));
 AND2_X2 _20447_ (.A1(_11837_),
    .A2(_11859_),
    .ZN(_03820_));
 AOI21_X2 _20448_ (.A(_10983_),
    .B1(_12964_),
    .B2(_12970_),
    .ZN(_03821_));
 AOI21_X4 _20449_ (.A(_03821_),
    .B1(_12953_),
    .B2(_10983_),
    .ZN(_03822_));
 MUX2_X1 _20450_ (.A(_03820_),
    .B(_03822_),
    .S(_03794_),
    .Z(_03823_));
 CLKBUF_X3 _20451_ (.A(_03823_),
    .Z(_03824_));
 NAND2_X1 _20452_ (.A1(_03810_),
    .A2(_03824_),
    .ZN(_14478_));
 AND2_X1 _20453_ (.A1(net330),
    .A2(_03805_),
    .ZN(_03825_));
 AOI21_X4 _20454_ (.A(_03825_),
    .B1(_03798_),
    .B2(net312),
    .ZN(_03826_));
 NOR2_X1 _20455_ (.A1(_03807_),
    .A2(_03826_),
    .ZN(_14484_));
 NOR2_X1 _20456_ (.A1(_03819_),
    .A2(_03817_),
    .ZN(_14483_));
 INV_X2 _20457_ (.A(_03823_),
    .ZN(_03827_));
 NOR2_X1 _20458_ (.A1(_03818_),
    .A2(_03827_),
    .ZN(_14485_));
 NOR2_X2 _20459_ (.A1(_13030_),
    .A2(_13048_),
    .ZN(_03828_));
 MUX2_X1 _20460_ (.A(_11967_),
    .B(_03828_),
    .S(_03794_),
    .Z(_03829_));
 CLKBUF_X3 _20461_ (.A(_03829_),
    .Z(_03830_));
 NAND2_X1 _20462_ (.A1(_03810_),
    .A2(_03830_),
    .ZN(_14489_));
 OR2_X4 _20463_ (.A1(_11510_),
    .A2(_11528_),
    .ZN(_03831_));
 MUX2_X2 _20464_ (.A(_03831_),
    .B(_13198_),
    .S(_03789_),
    .Z(_03832_));
 INV_X1 _20465_ (.A(_03832_),
    .ZN(_03833_));
 NOR2_X1 _20466_ (.A1(_03807_),
    .A2(_03833_),
    .ZN(_15991_));
 NOR2_X1 _20467_ (.A1(_03819_),
    .A2(_03826_),
    .ZN(_14504_));
 BUF_X4 _20468_ (.A(_03817_),
    .Z(_03834_));
 NOR2_X1 _20469_ (.A1(_03834_),
    .A2(_03827_),
    .ZN(_14503_));
 INV_X2 _20470_ (.A(_03829_),
    .ZN(_03835_));
 NOR2_X1 _20471_ (.A1(_03818_),
    .A2(_03835_),
    .ZN(_14505_));
 NOR2_X4 _20472_ (.A1(_13137_),
    .A2(_13155_),
    .ZN(_03836_));
 BUF_X4 _20473_ (.A(_03793_),
    .Z(_03837_));
 MUX2_X1 _20474_ (.A(_12008_),
    .B(_03836_),
    .S(_03837_),
    .Z(_03838_));
 CLKBUF_X3 _20475_ (.A(_03838_),
    .Z(_03839_));
 NAND2_X1 _20476_ (.A1(_03810_),
    .A2(_03839_),
    .ZN(_14508_));
 MUX2_X2 _20477_ (.A(net361),
    .B(_13307_),
    .S(_03788_),
    .Z(_03840_));
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 INV_X1 _20479_ (.A(net322),
    .ZN(_03842_));
 NOR2_X1 _20480_ (.A1(_03807_),
    .A2(_03842_),
    .ZN(_16003_));
 NOR2_X1 _20481_ (.A1(_03819_),
    .A2(_03833_),
    .ZN(_16004_));
 NOR2_X1 _20482_ (.A1(_03827_),
    .A2(_03826_),
    .ZN(_14527_));
 NOR2_X1 _20483_ (.A1(_03834_),
    .A2(_03835_),
    .ZN(_14526_));
 NOR2_X4 _20484_ (.A1(_03751_),
    .A2(_03776_),
    .ZN(_03843_));
 NOR2_X1 _20485_ (.A1(_13156_),
    .A2(_03843_),
    .ZN(_03844_));
 AOI21_X4 _20486_ (.A(_03844_),
    .B1(_03843_),
    .B2(_12008_),
    .ZN(_03845_));
 NOR2_X1 _20487_ (.A1(_03818_),
    .A2(_03845_),
    .ZN(_14528_));
 NOR2_X2 _20488_ (.A1(_13217_),
    .A2(_13235_),
    .ZN(_03846_));
 MUX2_X1 _20489_ (.A(_12051_),
    .B(_03846_),
    .S(_03794_),
    .Z(_03847_));
 CLKBUF_X3 _20490_ (.A(_03847_),
    .Z(_03848_));
 NAND2_X1 _20491_ (.A1(_03810_),
    .A2(_03848_),
    .ZN(_14533_));
 OR2_X4 _20492_ (.A1(_11598_),
    .A2(_11609_),
    .ZN(_03849_));
 MUX2_X2 _20493_ (.A(_03849_),
    .B(_13384_),
    .S(_03789_),
    .Z(_03850_));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 NAND2_X1 _20495_ (.A1(_03803_),
    .A2(net317),
    .ZN(_14544_));
 BUF_X4 _20496_ (.A(_03826_),
    .Z(_03852_));
 NOR2_X1 _20497_ (.A1(_03852_),
    .A2(_03835_),
    .ZN(_14550_));
 NOR2_X1 _20498_ (.A1(_03834_),
    .A2(_03845_),
    .ZN(_14549_));
 INV_X2 _20499_ (.A(_03847_),
    .ZN(_03853_));
 NOR2_X1 _20500_ (.A1(_03818_),
    .A2(_03853_),
    .ZN(_14551_));
 NOR2_X2 _20501_ (.A1(_12071_),
    .A2(_12091_),
    .ZN(_03854_));
 NOR2_X2 _20502_ (.A1(_13327_),
    .A2(_13345_),
    .ZN(_03855_));
 MUX2_X1 _20503_ (.A(_03854_),
    .B(_03855_),
    .S(_03837_),
    .Z(_03856_));
 CLKBUF_X3 _20504_ (.A(_03856_),
    .Z(_03857_));
 NAND2_X1 _20505_ (.A1(_03810_),
    .A2(_03857_),
    .ZN(_14559_));
 MUX2_X2 _20506_ (.A(_11648_),
    .B(_13480_),
    .S(_03789_),
    .Z(_03858_));
 INV_X1 _20507_ (.A(_03858_),
    .ZN(_03859_));
 NOR2_X1 _20508_ (.A1(_03807_),
    .A2(_03859_),
    .ZN(_16037_));
 NAND2_X1 _20509_ (.A1(_03814_),
    .A2(net317),
    .ZN(_14577_));
 NOR2_X1 _20510_ (.A1(_03852_),
    .A2(_03845_),
    .ZN(_14581_));
 NOR2_X1 _20511_ (.A1(_03834_),
    .A2(_03853_),
    .ZN(_14583_));
 MUX2_X2 _20512_ (.A(_12092_),
    .B(_13346_),
    .S(_03837_),
    .Z(_03860_));
 NOR2_X1 _20513_ (.A1(_03818_),
    .A2(_03860_),
    .ZN(_14582_));
 NOR2_X4 _20514_ (.A1(_12116_),
    .A2(_12135_),
    .ZN(_03861_));
 NOR2_X2 _20515_ (.A1(_13403_),
    .A2(_13421_),
    .ZN(_03862_));
 MUX2_X1 _20516_ (.A(_03861_),
    .B(_03862_),
    .S(_03837_),
    .Z(_03863_));
 BUF_X4 _20517_ (.A(_03863_),
    .Z(_03864_));
 NAND2_X1 _20518_ (.A1(_03810_),
    .A2(_03864_),
    .ZN(_14589_));
 NAND2_X1 _20519_ (.A1(_12425_),
    .A2(_11685_),
    .ZN(_03865_));
 AOI21_X2 _20520_ (.A(_11659_),
    .B1(_11667_),
    .B2(_11677_),
    .ZN(_03866_));
 NAND2_X4 _20521_ (.A1(_03865_),
    .A2(_03866_),
    .ZN(_03867_));
 MUX2_X1 _20522_ (.A(_03867_),
    .B(_13555_),
    .S(_03788_),
    .Z(_03868_));
 CLKBUF_X3 _20523_ (.A(_03868_),
    .Z(_03869_));
 INV_X1 _20524_ (.A(_03869_),
    .ZN(_03870_));
 NOR2_X1 _20525_ (.A1(_03807_),
    .A2(_03870_),
    .ZN(_16048_));
 NOR2_X1 _20526_ (.A1(_03819_),
    .A2(_03859_),
    .ZN(_16047_));
 NAND2_X1 _20527_ (.A1(_03824_),
    .A2(net317),
    .ZN(_14609_));
 NOR2_X1 _20528_ (.A1(_03852_),
    .A2(_03853_),
    .ZN(_14613_));
 NOR2_X1 _20529_ (.A1(_03834_),
    .A2(_03860_),
    .ZN(_14612_));
 MUX2_X2 _20530_ (.A(_12136_),
    .B(_13422_),
    .S(_03837_),
    .Z(_03871_));
 NOR2_X1 _20531_ (.A1(_03818_),
    .A2(_03871_),
    .ZN(_14614_));
 INV_X2 _20532_ (.A(_12217_),
    .ZN(_03872_));
 NOR2_X4 _20533_ (.A1(_13499_),
    .A2(_13517_),
    .ZN(_03873_));
 MUX2_X1 _20534_ (.A(_03872_),
    .B(_03873_),
    .S(_03837_),
    .Z(_03874_));
 BUF_X4 _20535_ (.A(_03874_),
    .Z(_03875_));
 NAND2_X1 _20536_ (.A1(_03810_),
    .A2(_03875_),
    .ZN(_14622_));
 MUX2_X1 _20537_ (.A(_11724_),
    .B(_13648_),
    .S(_03788_),
    .Z(_03876_));
 CLKBUF_X3 _20538_ (.A(_03876_),
    .Z(_03877_));
 BUF_X4 _20539_ (.A(_03877_),
    .Z(_03878_));
 NAND2_X1 _20540_ (.A1(_03803_),
    .A2(_03878_),
    .ZN(_14644_));
 NAND2_X1 _20541_ (.A1(_03830_),
    .A2(_03850_),
    .ZN(_14649_));
 NOR2_X1 _20542_ (.A1(_03852_),
    .A2(_03860_),
    .ZN(_14653_));
 NOR2_X1 _20543_ (.A1(_03834_),
    .A2(_03871_),
    .ZN(_14652_));
 MUX2_X2 _20544_ (.A(_12217_),
    .B(_13518_),
    .S(_03837_),
    .Z(_03879_));
 NOR2_X1 _20545_ (.A1(_03818_),
    .A2(_03879_),
    .ZN(_14654_));
 NOR2_X4 _20546_ (.A1(_12241_),
    .A2(_12259_),
    .ZN(_03880_));
 NOR2_X4 _20547_ (.A1(_13574_),
    .A2(_13592_),
    .ZN(_03881_));
 MUX2_X1 _20548_ (.A(_03880_),
    .B(_03881_),
    .S(_03794_),
    .Z(_03882_));
 BUF_X4 _20549_ (.A(_03882_),
    .Z(_03883_));
 NAND2_X1 _20550_ (.A1(_03810_),
    .A2(_03883_),
    .ZN(_14662_));
 NOR3_X2 _20551_ (.A1(_11749_),
    .A2(_11768_),
    .A3(_03788_),
    .ZN(_03884_));
 AOI21_X2 _20552_ (.A(_03884_),
    .B1(_03789_),
    .B2(_03104_),
    .ZN(_03885_));
 CLKBUF_X3 _20553_ (.A(_03885_),
    .Z(_03886_));
 NOR2_X1 _20554_ (.A1(_03807_),
    .A2(_03886_),
    .ZN(_16079_));
 NAND2_X1 _20555_ (.A1(_03814_),
    .A2(_03878_),
    .ZN(_14684_));
 NAND2_X1 _20556_ (.A1(_03839_),
    .A2(_03850_),
    .ZN(_14689_));
 NOR2_X1 _20557_ (.A1(_03852_),
    .A2(_03871_),
    .ZN(_14693_));
 NOR2_X1 _20558_ (.A1(_03834_),
    .A2(_03879_),
    .ZN(_14692_));
 MUX2_X2 _20559_ (.A(_12260_),
    .B(_13593_),
    .S(_03837_),
    .Z(_03887_));
 NOR2_X1 _20560_ (.A1(_03818_),
    .A2(_03887_),
    .ZN(_14694_));
 AOI21_X2 _20561_ (.A(_10983_),
    .B1(_12315_),
    .B2(_12321_),
    .ZN(_03888_));
 AOI21_X4 _20562_ (.A(_03888_),
    .B1(_12304_),
    .B2(_10983_),
    .ZN(_03889_));
 MUX2_X2 _20563_ (.A(_03889_),
    .B(_13686_),
    .S(_03794_),
    .Z(_03890_));
 CLKBUF_X3 _20564_ (.A(_03890_),
    .Z(_03891_));
 NAND2_X1 _20565_ (.A1(_03810_),
    .A2(_03891_),
    .ZN(_14705_));
 AND2_X1 _20566_ (.A1(_12420_),
    .A2(_03805_),
    .ZN(_03892_));
 AOI21_X2 _20567_ (.A(_03892_),
    .B1(_03789_),
    .B2(_03198_),
    .ZN(_03893_));
 BUF_X4 _20568_ (.A(_03893_),
    .Z(_03894_));
 NOR2_X1 _20569_ (.A1(_03807_),
    .A2(_03894_),
    .ZN(_16090_));
 NOR2_X1 _20570_ (.A1(_03819_),
    .A2(_03886_),
    .ZN(_16089_));
 NAND2_X1 _20571_ (.A1(_03824_),
    .A2(_03878_),
    .ZN(_14726_));
 NAND2_X1 _20572_ (.A1(_03848_),
    .A2(_03850_),
    .ZN(_14732_));
 NOR2_X2 _20573_ (.A1(_03852_),
    .A2(_03879_),
    .ZN(_14736_));
 NOR2_X2 _20574_ (.A1(_03834_),
    .A2(_03887_),
    .ZN(_14735_));
 INV_X2 _20575_ (.A(_03890_),
    .ZN(_03895_));
 NOR2_X1 _20576_ (.A1(_03818_),
    .A2(_03895_),
    .ZN(_14737_));
 NOR2_X4 _20577_ (.A1(_11792_),
    .A2(_11816_),
    .ZN(_03896_));
 MUX2_X2 _20578_ (.A(_03896_),
    .B(_03139_),
    .S(_03794_),
    .Z(_03897_));
 CLKBUF_X3 _20579_ (.A(_03897_),
    .Z(_03898_));
 NAND2_X1 _20580_ (.A1(_03806_),
    .A2(_03898_),
    .ZN(_14751_));
 AND2_X1 _20581_ (.A1(_12473_),
    .A2(_03805_),
    .ZN(_03899_));
 AOI21_X2 _20582_ (.A(_03899_),
    .B1(_03798_),
    .B2(_03276_),
    .ZN(_03900_));
 BUF_X4 _20583_ (.A(_03900_),
    .Z(_03901_));
 NOR2_X1 _20584_ (.A1(_03797_),
    .A2(_03901_),
    .ZN(_14772_));
 NOR2_X1 _20585_ (.A1(_03819_),
    .A2(_03894_),
    .ZN(_14771_));
 NOR2_X1 _20586_ (.A1(_03827_),
    .A2(_03886_),
    .ZN(_14773_));
 NAND2_X1 _20587_ (.A1(_03830_),
    .A2(_03877_),
    .ZN(_14778_));
 BUF_X8 _20588_ (.A(_03850_),
    .Z(_03902_));
 NAND2_X2 _20589_ (.A1(_03902_),
    .A2(_03857_),
    .ZN(_14784_));
 NOR2_X1 _20590_ (.A1(_03852_),
    .A2(_03887_),
    .ZN(_14791_));
 NOR2_X2 _20591_ (.A1(_03834_),
    .A2(_03895_),
    .ZN(_14790_));
 INV_X1 _20592_ (.A(_03897_),
    .ZN(_03903_));
 NOR2_X1 _20593_ (.A1(_03809_),
    .A2(_03903_),
    .ZN(_14789_));
 AOI21_X2 _20594_ (.A(_10983_),
    .B1(_11266_),
    .B2(_11274_),
    .ZN(_03904_));
 AOI21_X4 _20595_ (.A(_03904_),
    .B1(_11251_),
    .B2(_10983_),
    .ZN(_03905_));
 NAND2_X2 _20596_ (.A1(_03227_),
    .A2(_03236_),
    .ZN(_03906_));
 MUX2_X2 _20597_ (.A(_03905_),
    .B(_03906_),
    .S(_03794_),
    .Z(_03907_));
 CLKBUF_X3 _20598_ (.A(_03907_),
    .Z(_03908_));
 NAND2_X1 _20599_ (.A1(_03806_),
    .A2(_03908_),
    .ZN(_14805_));
 MUX2_X2 _20600_ (.A(_12580_),
    .B(_03372_),
    .S(_03789_),
    .Z(_03909_));
 INV_X1 _20601_ (.A(_03909_),
    .ZN(_03910_));
 NOR2_X1 _20602_ (.A1(_03797_),
    .A2(_03910_),
    .ZN(_16111_));
 INV_X2 _20603_ (.A(_03900_),
    .ZN(_03911_));
 NAND2_X1 _20604_ (.A1(_03814_),
    .A2(_03911_),
    .ZN(_14828_));
 NAND2_X1 _20605_ (.A1(_03839_),
    .A2(_03877_),
    .ZN(_14832_));
 NAND2_X1 _20606_ (.A1(_03902_),
    .A2(_03864_),
    .ZN(_14840_));
 NOR2_X1 _20607_ (.A1(_03852_),
    .A2(_03895_),
    .ZN(_14847_));
 NOR2_X1 _20608_ (.A1(_03834_),
    .A2(_03903_),
    .ZN(_14846_));
 INV_X1 _20609_ (.A(_03907_),
    .ZN(_03912_));
 NOR2_X1 _20610_ (.A1(_03809_),
    .A2(_03912_),
    .ZN(_14845_));
 AOI21_X2 _20611_ (.A(_10983_),
    .B1(_12501_),
    .B2(_12509_),
    .ZN(_03913_));
 AOI21_X4 _20612_ (.A(_03913_),
    .B1(_12490_),
    .B2(_10983_),
    .ZN(_03914_));
 OR2_X2 _20613_ (.A1(_03297_),
    .A2(_03315_),
    .ZN(_03915_));
 MUX2_X2 _20614_ (.A(_03914_),
    .B(_03915_),
    .S(_03794_),
    .Z(_03916_));
 CLKBUF_X3 _20615_ (.A(_03916_),
    .Z(_03917_));
 NAND2_X1 _20616_ (.A1(_03806_),
    .A2(_03917_),
    .ZN(_14860_));
 MUX2_X1 _20617_ (.A(_12656_),
    .B(_03452_),
    .S(_03788_),
    .Z(_03918_));
 BUF_X4 _20618_ (.A(_03918_),
    .Z(_03919_));
 AND2_X1 _20619_ (.A1(_03803_),
    .A2(_03919_),
    .ZN(_16121_));
 NOR2_X1 _20620_ (.A1(_03819_),
    .A2(_03910_),
    .ZN(_16120_));
 NOR2_X1 _20621_ (.A1(_03827_),
    .A2(_03901_),
    .ZN(_14882_));
 NOR2_X1 _20622_ (.A1(_03835_),
    .A2(_03894_),
    .ZN(_14881_));
 NOR2_X1 _20623_ (.A1(_03845_),
    .A2(_03886_),
    .ZN(_14883_));
 NAND2_X1 _20624_ (.A1(_03848_),
    .A2(_03877_),
    .ZN(_14887_));
 NAND2_X1 _20625_ (.A1(_03902_),
    .A2(_03875_),
    .ZN(_14899_));
 NOR2_X1 _20626_ (.A1(_03852_),
    .A2(_03903_),
    .ZN(_14903_));
 NOR2_X1 _20627_ (.A1(_03817_),
    .A2(_03912_),
    .ZN(_14905_));
 INV_X1 _20628_ (.A(_03916_),
    .ZN(_03920_));
 NOR2_X1 _20629_ (.A1(_03809_),
    .A2(_03920_),
    .ZN(_14904_));
 NOR2_X4 _20630_ (.A1(_12598_),
    .A2(_12616_),
    .ZN(_03921_));
 OR2_X2 _20631_ (.A1(_03393_),
    .A2(_03412_),
    .ZN(_03922_));
 MUX2_X2 _20632_ (.A(_03921_),
    .B(_03922_),
    .S(_03793_),
    .Z(_03923_));
 CLKBUF_X3 _20633_ (.A(_03923_),
    .Z(_03924_));
 NAND2_X1 _20634_ (.A1(_03806_),
    .A2(_03924_),
    .ZN(_14917_));
 BUF_X4 _20635_ (.A(_03766_),
    .Z(_03925_));
 NOR2_X4 _20636_ (.A1(_03925_),
    .A2(_03805_),
    .ZN(_03926_));
 CLKBUF_X3 _20637_ (.A(_03926_),
    .Z(_14992_));
 NAND2_X1 _20638_ (.A1(_03807_),
    .A2(_14992_),
    .ZN(_14940_));
 NOR2_X1 _20639_ (.A1(_03835_),
    .A2(_03901_),
    .ZN(_14943_));
 NOR2_X1 _20640_ (.A1(_03845_),
    .A2(_03894_),
    .ZN(_14945_));
 NOR2_X1 _20641_ (.A1(_03853_),
    .A2(_03886_),
    .ZN(_14944_));
 NAND2_X1 _20642_ (.A1(_03857_),
    .A2(_03877_),
    .ZN(_14953_));
 NAND2_X1 _20643_ (.A1(net316),
    .A2(_03883_),
    .ZN(_14966_));
 NOR2_X1 _20644_ (.A1(_03852_),
    .A2(_03912_),
    .ZN(_14970_));
 NOR2_X1 _20645_ (.A1(_03817_),
    .A2(_03920_),
    .ZN(_14969_));
 INV_X1 _20646_ (.A(_03923_),
    .ZN(_03927_));
 NOR2_X1 _20647_ (.A1(_03809_),
    .A2(_03927_),
    .ZN(_14971_));
 NOR2_X4 _20648_ (.A1(_12675_),
    .A2(_12694_),
    .ZN(_03928_));
 MUX2_X2 _20649_ (.A(_03928_),
    .B(_03488_),
    .S(_03793_),
    .Z(_03929_));
 AND2_X1 _20650_ (.A1(_03806_),
    .A2(_03929_),
    .ZN(_14984_));
 BUF_X4 _20651_ (.A(_03760_),
    .Z(_03930_));
 NAND2_X4 _20652_ (.A1(_03930_),
    .A2(_03837_),
    .ZN(_03931_));
 NOR2_X4 _20653_ (.A1(_03931_),
    .A2(_03791_),
    .ZN(_14983_));
 NAND2_X1 _20654_ (.A1(_03776_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .ZN(_03932_));
 NAND2_X1 _20655_ (.A1(_03751_),
    .A2(_03750_),
    .ZN(_03933_));
 CLKBUF_X3 _20656_ (.A(_03933_),
    .Z(_03934_));
 OAI21_X1 _20657_ (.A(_03932_),
    .B1(_03934_),
    .B2(_03800_),
    .ZN(_14985_));
 NAND2_X1 _20658_ (.A1(_03819_),
    .A2(_14992_),
    .ZN(_15008_));
 NOR2_X1 _20659_ (.A1(_03845_),
    .A2(_03901_),
    .ZN(_15015_));
 NOR2_X1 _20660_ (.A1(_03853_),
    .A2(_03894_),
    .ZN(_15014_));
 NOR2_X1 _20661_ (.A1(_03860_),
    .A2(_03886_),
    .ZN(_15013_));
 NAND2_X1 _20662_ (.A1(_03864_),
    .A2(_03877_),
    .ZN(_15022_));
 NAND2_X1 _20663_ (.A1(net316),
    .A2(_03891_),
    .ZN(_15032_));
 NOR2_X1 _20664_ (.A1(_03826_),
    .A2(_03920_),
    .ZN(_15039_));
 NOR2_X1 _20665_ (.A1(_03817_),
    .A2(_03927_),
    .ZN(_15038_));
 INV_X1 _20666_ (.A(_03929_),
    .ZN(_03935_));
 NOR2_X1 _20667_ (.A1(_03809_),
    .A2(_03935_),
    .ZN(_15037_));
 INV_X1 _20668_ (.A(_03760_),
    .ZN(_03936_));
 NOR2_X2 _20669_ (.A1(_03936_),
    .A2(_03843_),
    .ZN(_03937_));
 BUF_X4 _20670_ (.A(_03937_),
    .Z(_03938_));
 AND2_X4 _20671_ (.A1(_03806_),
    .A2(_03938_),
    .ZN(_15050_));
 NAND2_X1 _20672_ (.A1(_03776_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .ZN(_03939_));
 CLKBUF_X3 _20673_ (.A(_00723_),
    .Z(_03940_));
 OAI21_X2 _20674_ (.A(_03939_),
    .B1(_03934_),
    .B2(_03940_),
    .ZN(_15051_));
 NAND2_X1 _20675_ (.A1(_03827_),
    .A2(_14992_),
    .ZN(_15069_));
 NOR2_X1 _20676_ (.A1(_03853_),
    .A2(_03901_),
    .ZN(_15074_));
 NOR2_X1 _20677_ (.A1(_03860_),
    .A2(_03894_),
    .ZN(_15073_));
 NOR2_X1 _20678_ (.A1(_03871_),
    .A2(_03886_),
    .ZN(_15075_));
 NAND2_X1 _20679_ (.A1(_03875_),
    .A2(_03877_),
    .ZN(_15081_));
 NAND2_X1 _20680_ (.A1(_03902_),
    .A2(_03898_),
    .ZN(_15092_));
 NOR2_X1 _20681_ (.A1(_03826_),
    .A2(_03927_),
    .ZN(_15097_));
 NOR2_X1 _20682_ (.A1(_03817_),
    .A2(_03935_),
    .ZN(_15096_));
 OR2_X1 _20683_ (.A1(_03809_),
    .A2(_03931_),
    .ZN(_15156_));
 INV_X1 _20684_ (.A(_15156_),
    .ZN(_15098_));
 CLKBUF_X2 _20685_ (.A(_03837_),
    .Z(_03941_));
 OR3_X2 _20686_ (.A1(_01163_),
    .A2(_00132_),
    .A3(_03757_),
    .ZN(_03942_));
 CLKBUF_X3 _20687_ (.A(_03942_),
    .Z(_03943_));
 CLKBUF_X3 _20688_ (.A(_00754_),
    .Z(_03944_));
 OAI21_X1 _20689_ (.A(_03943_),
    .B1(_03934_),
    .B2(_03944_),
    .ZN(_03945_));
 AND2_X1 _20690_ (.A1(_03941_),
    .A2(_03945_),
    .ZN(_15108_));
 NAND2_X1 _20691_ (.A1(_03835_),
    .A2(_14992_),
    .ZN(_15127_));
 NOR2_X1 _20692_ (.A1(_03860_),
    .A2(_03901_),
    .ZN(_15132_));
 NOR2_X1 _20693_ (.A1(_03871_),
    .A2(_03894_),
    .ZN(_15131_));
 NOR2_X1 _20694_ (.A1(_03879_),
    .A2(_03886_),
    .ZN(_15133_));
 NAND2_X1 _20695_ (.A1(_03878_),
    .A2(_03883_),
    .ZN(_15139_));
 NAND2_X1 _20696_ (.A1(net316),
    .A2(_03908_),
    .ZN(_15150_));
 OR2_X1 _20697_ (.A1(_03826_),
    .A2(_03935_),
    .ZN(_15155_));
 OR2_X1 _20698_ (.A1(_03817_),
    .A2(_03931_),
    .ZN(_15154_));
 INV_X1 _20699_ (.A(_15154_),
    .ZN(_15212_));
 BUF_X2 _20700_ (.A(_00785_),
    .Z(_03946_));
 OAI21_X1 _20701_ (.A(_03943_),
    .B1(_03934_),
    .B2(_03946_),
    .ZN(_03947_));
 AND2_X1 _20702_ (.A1(_03941_),
    .A2(_03947_),
    .ZN(_15165_));
 NAND2_X1 _20703_ (.A1(_03845_),
    .A2(_14992_),
    .ZN(_15184_));
 NOR2_X1 _20704_ (.A1(_03871_),
    .A2(_03901_),
    .ZN(_15191_));
 NOR2_X1 _20705_ (.A1(_03879_),
    .A2(_03894_),
    .ZN(_15190_));
 NOR2_X1 _20706_ (.A1(_03887_),
    .A2(_03885_),
    .ZN(_15189_));
 NAND2_X1 _20707_ (.A1(_03878_),
    .A2(_03891_),
    .ZN(_15198_));
 NAND2_X1 _20708_ (.A1(net316),
    .A2(_03917_),
    .ZN(_15207_));
 NOR2_X1 _20709_ (.A1(_03826_),
    .A2(_03931_),
    .ZN(_15213_));
 CLKBUF_X3 _20710_ (.A(_00816_),
    .Z(_03948_));
 OAI21_X1 _20711_ (.A(_03943_),
    .B1(_03934_),
    .B2(_03948_),
    .ZN(_03949_));
 AND2_X1 _20712_ (.A1(_03941_),
    .A2(_03949_),
    .ZN(_15223_));
 NAND2_X1 _20713_ (.A1(_03853_),
    .A2(_14992_),
    .ZN(_15243_));
 NOR2_X1 _20714_ (.A1(_03879_),
    .A2(_03901_),
    .ZN(_15247_));
 NOR2_X1 _20715_ (.A1(_03887_),
    .A2(_03894_),
    .ZN(_15246_));
 NOR2_X1 _20716_ (.A1(_03886_),
    .A2(_03895_),
    .ZN(_15248_));
 NAND2_X1 _20717_ (.A1(_03878_),
    .A2(_03898_),
    .ZN(_15255_));
 NAND2_X1 _20718_ (.A1(net316),
    .A2(_03924_),
    .ZN(_15266_));
 NAND2_X2 _20719_ (.A1(_03832_),
    .A2(_03938_),
    .ZN(_15264_));
 INV_X1 _20720_ (.A(_15264_),
    .ZN(_15370_));
 CLKBUF_X3 _20721_ (.A(_00847_),
    .Z(_03950_));
 OAI21_X1 _20722_ (.A(_03943_),
    .B1(_03934_),
    .B2(_03950_),
    .ZN(_03951_));
 AND2_X1 _20723_ (.A1(_03941_),
    .A2(_03951_),
    .ZN(_15275_));
 NAND2_X1 _20724_ (.A1(_03860_),
    .A2(_14992_),
    .ZN(_15295_));
 NOR2_X1 _20725_ (.A1(_03887_),
    .A2(_03901_),
    .ZN(_15300_));
 NOR2_X1 _20726_ (.A1(_03895_),
    .A2(_03894_),
    .ZN(_15299_));
 NOR2_X1 _20727_ (.A1(_03886_),
    .A2(_03903_),
    .ZN(_15301_));
 NAND2_X1 _20728_ (.A1(_03878_),
    .A2(_03908_),
    .ZN(_15307_));
 CLKBUF_X3 _20729_ (.A(_03929_),
    .Z(_03952_));
 NAND2_X1 _20730_ (.A1(_03902_),
    .A2(_03952_),
    .ZN(_15318_));
 NAND2_X1 _20731_ (.A1(_03840_),
    .A2(_03938_),
    .ZN(_15317_));
 INV_X1 _20732_ (.A(_15317_),
    .ZN(_15371_));
 INV_X2 _20733_ (.A(_00878_),
    .ZN(_03953_));
 NAND2_X1 _20734_ (.A1(_03953_),
    .A2(_03779_),
    .ZN(_03954_));
 AOI21_X1 _20735_ (.A(_03843_),
    .B1(_03943_),
    .B2(_03954_),
    .ZN(_15330_));
 NAND2_X1 _20736_ (.A1(_03871_),
    .A2(_03926_),
    .ZN(_15348_));
 NAND2_X1 _20737_ (.A1(_03891_),
    .A2(_03911_),
    .ZN(_15355_));
 NAND2_X1 _20738_ (.A1(_03878_),
    .A2(_03917_),
    .ZN(_15361_));
 AND2_X1 _20739_ (.A1(net317),
    .A2(_03938_),
    .ZN(_15372_));
 CLKBUF_X3 _20740_ (.A(_00909_),
    .Z(_03955_));
 OAI21_X1 _20741_ (.A(_03943_),
    .B1(_03934_),
    .B2(_03955_),
    .ZN(_03956_));
 AND2_X1 _20742_ (.A1(_03941_),
    .A2(_03956_),
    .ZN(_15383_));
 NAND2_X1 _20743_ (.A1(_03879_),
    .A2(_03926_),
    .ZN(_15403_));
 NAND2_X1 _20744_ (.A1(_03898_),
    .A2(_03911_),
    .ZN(_15407_));
 NAND2_X1 _20745_ (.A1(_03878_),
    .A2(_03924_),
    .ZN(_15414_));
 NAND2_X2 _20746_ (.A1(_03858_),
    .A2(_03938_),
    .ZN(_15415_));
 INV_X1 _20747_ (.A(_15415_),
    .ZN(_15503_));
 CLKBUF_X3 _20748_ (.A(_00940_),
    .Z(_03957_));
 OAI21_X1 _20749_ (.A(_03942_),
    .B1(_03934_),
    .B2(_03957_),
    .ZN(_03958_));
 AND2_X1 _20750_ (.A1(_03941_),
    .A2(_03958_),
    .ZN(_15429_));
 NAND2_X1 _20751_ (.A1(_03887_),
    .A2(_03926_),
    .ZN(_15448_));
 NAND2_X1 _20752_ (.A1(_03911_),
    .A2(_03908_),
    .ZN(_15453_));
 NAND2_X1 _20753_ (.A1(_03878_),
    .A2(_03952_),
    .ZN(_15459_));
 NAND2_X1 _20754_ (.A1(_03869_),
    .A2(_03938_),
    .ZN(_15460_));
 INV_X1 _20755_ (.A(_15460_),
    .ZN(_15504_));
 CLKBUF_X3 _20756_ (.A(_00971_),
    .Z(_03959_));
 OAI21_X1 _20757_ (.A(_03942_),
    .B1(_03934_),
    .B2(_03959_),
    .ZN(_03960_));
 AND2_X1 _20758_ (.A1(_03941_),
    .A2(_03960_),
    .ZN(_15472_));
 NAND2_X1 _20759_ (.A1(_03895_),
    .A2(_03926_),
    .ZN(_15492_));
 NAND2_X1 _20760_ (.A1(_03911_),
    .A2(_03917_),
    .ZN(_15497_));
 AND2_X1 _20761_ (.A1(_03877_),
    .A2(_03938_),
    .ZN(_15502_));
 INV_X2 _20762_ (.A(_01002_),
    .ZN(_03961_));
 NAND2_X1 _20763_ (.A1(_03961_),
    .A2(_03779_),
    .ZN(_03962_));
 AOI21_X1 _20764_ (.A(_03843_),
    .B1(_03943_),
    .B2(_03962_),
    .ZN(_15516_));
 NAND2_X1 _20765_ (.A1(_03903_),
    .A2(_03926_),
    .ZN(_15535_));
 NAND2_X1 _20766_ (.A1(_03911_),
    .A2(_03924_),
    .ZN(_15540_));
 INV_X2 _20767_ (.A(_03885_),
    .ZN(_03963_));
 NAND2_X1 _20768_ (.A1(_03963_),
    .A2(_03938_),
    .ZN(_15541_));
 INV_X1 _20769_ (.A(_15541_),
    .ZN(_15617_));
 INV_X1 _20770_ (.A(_01033_),
    .ZN(_03964_));
 NAND2_X1 _20771_ (.A1(_03964_),
    .A2(_03779_),
    .ZN(_03965_));
 AOI21_X2 _20772_ (.A(_03843_),
    .B1(_03943_),
    .B2(_03965_),
    .ZN(_15555_));
 NAND2_X1 _20773_ (.A1(_03912_),
    .A2(_03926_),
    .ZN(_15574_));
 NAND2_X1 _20774_ (.A1(_03911_),
    .A2(_03952_),
    .ZN(_15579_));
 INV_X2 _20775_ (.A(_03893_),
    .ZN(_03966_));
 NAND2_X1 _20776_ (.A1(_03966_),
    .A2(_03937_),
    .ZN(_15578_));
 INV_X1 _20777_ (.A(_15578_),
    .ZN(_15615_));
 CLKBUF_X3 _20778_ (.A(_01064_),
    .Z(_03967_));
 OAI21_X1 _20779_ (.A(_03942_),
    .B1(_03934_),
    .B2(_03967_),
    .ZN(_03968_));
 AND2_X1 _20780_ (.A1(_03941_),
    .A2(_03968_),
    .ZN(_15592_));
 NAND2_X1 _20781_ (.A1(_03920_),
    .A2(_03926_),
    .ZN(_15610_));
 NOR2_X1 _20782_ (.A1(_03901_),
    .A2(_03931_),
    .ZN(_15616_));
 INV_X1 _20783_ (.A(_01095_),
    .ZN(_03969_));
 NAND2_X1 _20784_ (.A1(_03969_),
    .A2(_03779_),
    .ZN(_03970_));
 AOI21_X2 _20785_ (.A(_03843_),
    .B1(_03943_),
    .B2(_03970_),
    .ZN(_15631_));
 NAND2_X1 _20786_ (.A1(_03927_),
    .A2(_03926_),
    .ZN(_15650_));
 CLKBUF_X3 _20787_ (.A(_01126_),
    .Z(_03971_));
 OAI21_X1 _20788_ (.A(_03942_),
    .B1(_03933_),
    .B2(_03971_),
    .ZN(_03972_));
 AND2_X1 _20789_ (.A1(_03941_),
    .A2(_03972_),
    .ZN(_15670_));
 NAND2_X1 _20790_ (.A1(_14992_),
    .A2(_03935_),
    .ZN(_15689_));
 OAI21_X1 _20791_ (.A(_03942_),
    .B1(_03933_),
    .B2(_03503_),
    .ZN(_03973_));
 AND2_X1 _20792_ (.A1(_03941_),
    .A2(_03973_),
    .ZN(_15706_));
 NAND2_X1 _20793_ (.A1(_14992_),
    .A2(_03931_),
    .ZN(_15723_));
 NAND2_X1 _20794_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(_03779_),
    .ZN(_03974_));
 AOI21_X2 _20795_ (.A(_03843_),
    .B1(_03943_),
    .B2(_03974_),
    .ZN(_15738_));
 INV_X1 _20796_ (.A(_15725_),
    .ZN(_15726_));
 INV_X1 _20797_ (.A(_15619_),
    .ZN(_15620_));
 INV_X4 _20798_ (.A(_15214_),
    .ZN(_15279_));
 INV_X1 _20799_ (.A(_03564_),
    .ZN(_03975_));
 NAND2_X1 _20800_ (.A1(_03530_),
    .A2(_03975_),
    .ZN(_03976_));
 INV_X2 _20801_ (.A(\cs_registers_i.nmi_mode_i ),
    .ZN(_03977_));
 OAI21_X2 _20802_ (.A(_03977_),
    .B1(net141),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .ZN(_03978_));
 NAND2_X2 _20803_ (.A1(_03531_),
    .A2(_03533_),
    .ZN(_03979_));
 OR4_X2 _20804_ (.A1(_03649_),
    .A2(_03976_),
    .A3(_03978_),
    .A4(_03979_),
    .ZN(_03980_));
 AOI22_X4 _20805_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net137),
    .B1(\cs_registers_i.mie_q[7] ),
    .B2(net138),
    .ZN(_03981_));
 AOI22_X4 _20806_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net135),
    .B1(\cs_registers_i.mie_q[5] ),
    .B2(net136),
    .ZN(_03982_));
 AOI22_X2 _20807_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net133),
    .B1(\cs_registers_i.mie_q[3] ),
    .B2(net134),
    .ZN(_03983_));
 AOI22_X2 _20808_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(net126),
    .B1(\cs_registers_i.mie_q[1] ),
    .B2(net132),
    .ZN(_03984_));
 NAND4_X2 _20809_ (.A1(_03981_),
    .A2(_03982_),
    .A3(_03983_),
    .A4(_03984_),
    .ZN(_03985_));
 AOI22_X4 _20810_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net127),
    .B1(\cs_registers_i.mie_q[11] ),
    .B2(net128),
    .ZN(_03986_));
 AOI22_X4 _20811_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net139),
    .B1(\cs_registers_i.mie_q[9] ),
    .B2(net140),
    .ZN(_03987_));
 AOI22_X4 _20812_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(net129),
    .B1(\cs_registers_i.mie_q[13] ),
    .B2(net130),
    .ZN(_03988_));
 NAND2_X2 _20813_ (.A1(\cs_registers_i.mie_q[14] ),
    .A2(net131),
    .ZN(_03989_));
 NAND4_X2 _20814_ (.A1(_03986_),
    .A2(_03987_),
    .A3(_03988_),
    .A4(_03989_),
    .ZN(_03990_));
 NOR2_X2 _20815_ (.A1(_03985_),
    .A2(_03990_),
    .ZN(_03991_));
 AOI21_X1 _20816_ (.A(net141),
    .B1(\cs_registers_i.mie_q[16] ),
    .B2(net143),
    .ZN(_03992_));
 AOI22_X2 _20817_ (.A1(net125),
    .A2(\cs_registers_i.mie_q[15] ),
    .B1(\cs_registers_i.mie_q[17] ),
    .B2(net142),
    .ZN(_03993_));
 AND3_X4 _20818_ (.A1(_03991_),
    .A2(_03992_),
    .A3(_03993_),
    .ZN(_03994_));
 NOR2_X2 _20819_ (.A1(_03980_),
    .A2(_03994_),
    .ZN(_03995_));
 NAND2_X4 _20820_ (.A1(_03532_),
    .A2(_03649_),
    .ZN(_03996_));
 BUF_X2 _20821_ (.A(\cs_registers_i.dcsr_q[2] ),
    .Z(_03997_));
 CLKBUF_X3 _20822_ (.A(debug_req_i),
    .Z(_03998_));
 NOR3_X2 _20823_ (.A1(_03530_),
    .A2(_03997_),
    .A3(_03998_),
    .ZN(_03999_));
 BUF_X4 _20824_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .Z(_04000_));
 AOI21_X1 _20825_ (.A(_03996_),
    .B1(_03999_),
    .B2(_04000_),
    .ZN(_04001_));
 OR2_X1 _20826_ (.A1(_03995_),
    .A2(_04001_),
    .ZN(_04002_));
 INV_X1 _20827_ (.A(\id_stage_i.branch_set ),
    .ZN(_04003_));
 OAI21_X1 _20828_ (.A(_10823_),
    .B1(_10830_),
    .B2(_10831_),
    .ZN(_04004_));
 NAND2_X1 _20829_ (.A1(_10834_),
    .A2(_04004_),
    .ZN(_04005_));
 NOR2_X4 _20830_ (.A1(_10780_),
    .A2(net306),
    .ZN(_04006_));
 OR4_X1 _20831_ (.A1(_10795_),
    .A2(_03653_),
    .A3(_04005_),
    .A4(_04006_),
    .ZN(_04007_));
 OAI21_X2 _20832_ (.A(_04003_),
    .B1(_03537_),
    .B2(_04007_),
    .ZN(_04008_));
 BUF_X4 _20833_ (.A(_03530_),
    .Z(_04009_));
 NAND2_X4 _20834_ (.A1(_04009_),
    .A2(_03650_),
    .ZN(_04010_));
 NOR2_X4 _20835_ (.A1(_10810_),
    .A2(_03648_),
    .ZN(_04011_));
 NOR2_X1 _20836_ (.A1(_04010_),
    .A2(_04011_),
    .ZN(_04012_));
 INV_X1 _20837_ (.A(_03530_),
    .ZN(_04013_));
 NAND4_X4 _20838_ (.A1(_04013_),
    .A2(_03531_),
    .A3(_03533_),
    .A4(_03534_),
    .ZN(_04014_));
 OR3_X2 _20839_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.exc_req_q ),
    .A3(\id_stage_i.controller_i.load_err_q ),
    .ZN(_04015_));
 BUF_X1 _20840_ (.A(_00557_),
    .Z(_04016_));
 OR3_X1 _20841_ (.A1(_00549_),
    .A2(_03660_),
    .A3(_03661_),
    .ZN(_04017_));
 OAI21_X4 _20842_ (.A(_04017_),
    .B1(_03662_),
    .B2(_00556_),
    .ZN(_04018_));
 OR2_X1 _20843_ (.A1(_03564_),
    .A2(_04018_),
    .ZN(_04019_));
 NAND2_X4 _20844_ (.A1(_10794_),
    .A2(_03647_),
    .ZN(_04020_));
 AND3_X1 _20845_ (.A1(_04016_),
    .A2(_04019_),
    .A3(_04020_),
    .ZN(_04021_));
 NAND2_X1 _20846_ (.A1(_04015_),
    .A2(_04021_),
    .ZN(_04022_));
 NOR4_X2 _20847_ (.A1(_11280_),
    .A2(_03674_),
    .A3(_03675_),
    .A4(_03676_),
    .ZN(_04023_));
 NOR2_X1 _20848_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_04011_),
    .ZN(_04024_));
 NAND3_X1 _20849_ (.A1(_10711_),
    .A2(_04023_),
    .A3(_04024_),
    .ZN(_04025_));
 NOR2_X2 _20850_ (.A1(_04022_),
    .A2(_04025_),
    .ZN(_04026_));
 NOR2_X2 _20851_ (.A1(_04014_),
    .A2(_04026_),
    .ZN(_04027_));
 OR4_X2 _20852_ (.A1(_10711_),
    .A2(_11136_),
    .A3(_11322_),
    .A4(_11323_),
    .ZN(_04028_));
 NOR4_X4 _20853_ (.A1(_11280_),
    .A2(_04028_),
    .A3(_11304_),
    .A4(_03675_),
    .ZN(_04029_));
 OR2_X2 _20854_ (.A1(_04015_),
    .A2(_04029_),
    .ZN(_04030_));
 AOI221_X2 _20855_ (.A(_04002_),
    .B1(_04008_),
    .B2(_04012_),
    .C1(_04027_),
    .C2(_04030_),
    .ZN(_04031_));
 BUF_X4 _20856_ (.A(_04031_),
    .Z(_04032_));
 NOR2_X2 _20857_ (.A1(_04014_),
    .A2(_04015_),
    .ZN(_04033_));
 AOI21_X4 _20858_ (.A(_03652_),
    .B1(_04029_),
    .B2(_04033_),
    .ZN(_04034_));
 NOR2_X4 _20859_ (.A1(_03533_),
    .A2(_03996_),
    .ZN(_04035_));
 NOR2_X1 _20860_ (.A1(_03530_),
    .A2(_04015_),
    .ZN(_04036_));
 INV_X2 _20861_ (.A(_11319_),
    .ZN(_04037_));
 OAI21_X2 _20862_ (.A(_04036_),
    .B1(_03668_),
    .B2(_04037_),
    .ZN(_04038_));
 NOR2_X2 _20863_ (.A1(_03649_),
    .A2(_03979_),
    .ZN(_04039_));
 AOI21_X4 _20864_ (.A(_04035_),
    .B1(_04038_),
    .B2(_04039_),
    .ZN(_04040_));
 AND2_X1 _20865_ (.A1(_04034_),
    .A2(_04040_),
    .ZN(_04041_));
 BUF_X4 _20866_ (.A(_04041_),
    .Z(_04042_));
 NOR2_X4 _20867_ (.A1(_04032_),
    .A2(_04042_),
    .ZN(_04043_));
 OR2_X1 _20868_ (.A1(_03980_),
    .A2(_03994_),
    .ZN(_04044_));
 NAND2_X1 _20869_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net137),
    .ZN(_04045_));
 NAND2_X1 _20870_ (.A1(\cs_registers_i.mie_q[5] ),
    .A2(net136),
    .ZN(_04046_));
 AND2_X1 _20871_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net135),
    .ZN(_04047_));
 NAND2_X1 _20872_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(net132),
    .ZN(_04048_));
 AOI21_X1 _20873_ (.A(_04048_),
    .B1(net133),
    .B2(\cs_registers_i.mie_q[2] ),
    .ZN(_04049_));
 AOI21_X1 _20874_ (.A(_04049_),
    .B1(net134),
    .B2(\cs_registers_i.mie_q[3] ),
    .ZN(_04050_));
 OAI21_X1 _20875_ (.A(_04046_),
    .B1(_04047_),
    .B2(_04050_),
    .ZN(_04051_));
 AOI22_X2 _20876_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(net138),
    .B1(_04045_),
    .B2(_04051_),
    .ZN(_04052_));
 AOI21_X1 _20877_ (.A(_04052_),
    .B1(net139),
    .B2(\cs_registers_i.mie_q[8] ),
    .ZN(_04053_));
 AOI21_X1 _20878_ (.A(_04053_),
    .B1(net140),
    .B2(\cs_registers_i.mie_q[9] ),
    .ZN(_04054_));
 AOI21_X1 _20879_ (.A(_04054_),
    .B1(net127),
    .B2(\cs_registers_i.mie_q[10] ),
    .ZN(_04055_));
 AOI21_X1 _20880_ (.A(_04055_),
    .B1(net128),
    .B2(\cs_registers_i.mie_q[11] ),
    .ZN(_04056_));
 AOI21_X1 _20881_ (.A(_04056_),
    .B1(net129),
    .B2(\cs_registers_i.mie_q[12] ),
    .ZN(_04057_));
 AND2_X1 _20882_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(net130),
    .ZN(_04058_));
 OAI21_X1 _20883_ (.A(_03989_),
    .B1(_04057_),
    .B2(_04058_),
    .ZN(_04059_));
 INV_X1 _20884_ (.A(net141),
    .ZN(_04060_));
 NOR2_X2 _20885_ (.A1(\cs_registers_i.nmi_mode_i ),
    .A2(_04060_),
    .ZN(_04061_));
 NOR2_X1 _20886_ (.A1(_03991_),
    .A2(_04061_),
    .ZN(_04062_));
 AOI21_X2 _20887_ (.A(_04044_),
    .B1(_04059_),
    .B2(_04062_),
    .ZN(_04063_));
 NOR3_X4 _20888_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.exc_req_q ),
    .A3(\id_stage_i.controller_i.load_err_q ),
    .ZN(_04064_));
 NAND2_X2 _20889_ (.A1(_03536_),
    .A2(_04064_),
    .ZN(_04065_));
 NOR3_X4 _20890_ (.A1(_03669_),
    .A2(_03668_),
    .A3(_04065_),
    .ZN(_04066_));
 BUF_X4 _20891_ (.A(_04066_),
    .Z(_04067_));
 NOR3_X4 _20892_ (.A1(_04037_),
    .A2(_03668_),
    .A3(_04065_),
    .ZN(_04068_));
 BUF_X4 _20893_ (.A(_04068_),
    .Z(_04069_));
 BUF_X4 _20894_ (.A(_04069_),
    .Z(_04070_));
 AOI221_X2 _20895_ (.A(_04063_),
    .B1(_04067_),
    .B2(\cs_registers_i.csr_depc_o[2] ),
    .C1(_04070_),
    .C2(\cs_registers_i.csr_mepc_o[2] ),
    .ZN(_04071_));
 INV_X1 _20896_ (.A(\alu_adder_result_ex[2] ),
    .ZN(_04072_));
 BUF_X4 _20897_ (.A(_04010_),
    .Z(_04073_));
 OAI21_X1 _20898_ (.A(_04071_),
    .B1(_04072_),
    .B2(_04073_),
    .ZN(_04074_));
 NAND2_X1 _20899_ (.A1(_04043_),
    .A2(_04074_),
    .ZN(_04075_));
 AOI21_X2 _20900_ (.A(_04002_),
    .B1(_04027_),
    .B2(_04030_),
    .ZN(_04076_));
 NAND2_X1 _20901_ (.A1(_04008_),
    .A2(_04012_),
    .ZN(_04077_));
 NAND2_X4 _20902_ (.A1(_04076_),
    .A2(_04077_),
    .ZN(_04078_));
 BUF_X4 _20903_ (.A(_04078_),
    .Z(_04079_));
 BUF_X4 _20904_ (.A(_04079_),
    .Z(_04080_));
 BUF_X4 _20905_ (.A(_04080_),
    .Z(_04081_));
 INV_X1 _20906_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .ZN(_04082_));
 OAI21_X1 _20907_ (.A(_04075_),
    .B1(_04081_),
    .B2(_04082_),
    .ZN(_16510_));
 CLKBUF_X3 _20908_ (.A(_03652_),
    .Z(_04083_));
 NOR2_X4 _20909_ (.A1(_04014_),
    .A2(_04064_),
    .ZN(_04084_));
 BUF_X2 _20910_ (.A(_01160_),
    .Z(_04085_));
 INV_X2 _20911_ (.A(_04085_),
    .ZN(_04086_));
 AOI22_X1 _20912_ (.A1(_04083_),
    .A2(\alu_adder_result_ex[3] ),
    .B1(_04084_),
    .B2(_04086_),
    .ZN(_04087_));
 INV_X1 _20913_ (.A(_03991_),
    .ZN(_04088_));
 NAND2_X1 _20914_ (.A1(_03977_),
    .A2(net141),
    .ZN(_04089_));
 INV_X1 _20915_ (.A(_03982_),
    .ZN(_04090_));
 OAI21_X1 _20916_ (.A(_03981_),
    .B1(_04090_),
    .B2(_03983_),
    .ZN(_04091_));
 NAND2_X1 _20917_ (.A1(_03987_),
    .A2(_04091_),
    .ZN(_04092_));
 NAND2_X1 _20918_ (.A1(_03986_),
    .A2(_04092_),
    .ZN(_04093_));
 NAND2_X1 _20919_ (.A1(_03988_),
    .A2(_04093_),
    .ZN(_04094_));
 NAND4_X1 _20920_ (.A1(_03989_),
    .A2(_04088_),
    .A3(_04089_),
    .A4(_04094_),
    .ZN(_04095_));
 NAND2_X1 _20921_ (.A1(_03995_),
    .A2(_04095_),
    .ZN(_04096_));
 INV_X1 _20922_ (.A(_01165_),
    .ZN(_04097_));
 AOI22_X2 _20923_ (.A1(_04097_),
    .A2(_04067_),
    .B1(_04069_),
    .B2(\cs_registers_i.csr_mepc_o[3] ),
    .ZN(_04098_));
 AND4_X1 _20924_ (.A1(_04078_),
    .A2(_04087_),
    .A3(_04096_),
    .A4(_04098_),
    .ZN(_04099_));
 BUF_X4 _20925_ (.A(_04032_),
    .Z(_04100_));
 INV_X1 _20926_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .ZN(_04101_));
 AOI21_X2 _20927_ (.A(_04099_),
    .B1(_04100_),
    .B2(_04101_),
    .ZN(_16512_));
 OAI21_X1 _20928_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_04081_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .ZN(_04102_));
 INV_X1 _20929_ (.A(_04102_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 BUF_X4 _20930_ (.A(\cs_registers_i.pc_if_i[1] ),
    .Z(_04103_));
 BUF_X4 _20931_ (.A(_04103_),
    .Z(_04104_));
 BUF_X4 _20932_ (.A(_04104_),
    .Z(_04105_));
 BUF_X4 _20933_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_04106_));
 INV_X8 _20934_ (.A(_04106_),
    .ZN(_04107_));
 BUF_X2 _20935_ (.A(instr_err_i),
    .Z(_04108_));
 CLKBUF_X2 _20936_ (.A(instr_rdata_i[17]),
    .Z(_04109_));
 CLKBUF_X2 _20937_ (.A(instr_rdata_i[16]),
    .Z(_04110_));
 AOI21_X1 _20938_ (.A(_04108_),
    .B1(_04109_),
    .B2(_04110_),
    .ZN(_04111_));
 AND2_X1 _20939_ (.A1(_04107_),
    .A2(_04111_),
    .ZN(_04112_));
 BUF_X2 _20940_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .Z(_04113_));
 AOI21_X2 _20941_ (.A(_04113_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .ZN(_04114_));
 AOI21_X4 _20942_ (.A(_04112_),
    .B1(_04114_),
    .B2(_04106_),
    .ZN(_04115_));
 NAND2_X1 _20943_ (.A1(_04105_),
    .A2(_04115_),
    .ZN(_04116_));
 AOI21_X1 _20944_ (.A(_04108_),
    .B1(net103),
    .B2(net94),
    .ZN(_04117_));
 AOI21_X1 _20945_ (.A(_04113_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .ZN(_04118_));
 CLKBUF_X3 _20946_ (.A(_04106_),
    .Z(_04119_));
 CLKBUF_X3 _20947_ (.A(_04119_),
    .Z(_04120_));
 BUF_X4 _20948_ (.A(_04120_),
    .Z(_04121_));
 MUX2_X2 _20949_ (.A(_04117_),
    .B(_04118_),
    .S(_04121_),
    .Z(_04122_));
 BUF_X4 _20950_ (.A(_04105_),
    .Z(_04123_));
 OAI21_X4 _20951_ (.A(_04116_),
    .B1(_04122_),
    .B2(_04123_),
    .ZN(_16232_));
 INV_X1 _20952_ (.A(_16232_),
    .ZN(_15755_));
 NOR2_X1 _20953_ (.A1(_03998_),
    .A2(core_busy_q),
    .ZN(_04124_));
 NAND2_X2 _20954_ (.A1(_03994_),
    .A2(_04124_),
    .ZN(_04125_));
 AOI21_X1 _20955_ (.A(net145),
    .B1(_04125_),
    .B2(fetch_enable_q),
    .ZN(_04126_));
 INV_X1 _20956_ (.A(_04126_),
    .ZN(_00006_));
 BUF_X8 _20957_ (.A(_03790_),
    .Z(_04127_));
 NAND2_X1 _20958_ (.A1(_04127_),
    .A2(_03814_),
    .ZN(_14468_));
 BUF_X4 _20959_ (.A(_03798_),
    .Z(_04128_));
 BUF_X2 _20960_ (.A(_03777_),
    .Z(_04129_));
 OR2_X1 _20961_ (.A1(_00558_),
    .A2(_04129_),
    .ZN(_04130_));
 CLKBUF_X3 _20962_ (.A(_03750_),
    .Z(_04131_));
 OAI21_X1 _20963_ (.A(_04130_),
    .B1(_04131_),
    .B2(_03944_),
    .ZN(_04132_));
 BUF_X4 _20964_ (.A(_03752_),
    .Z(_04133_));
 AOI22_X2 _20965_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A2(_04128_),
    .B1(_04132_),
    .B2(_04133_),
    .ZN(_14473_));
 OR2_X1 _20966_ (.A1(_00560_),
    .A2(_04129_),
    .ZN(_04134_));
 OAI21_X1 _20967_ (.A(_04134_),
    .B1(_04131_),
    .B2(_03948_),
    .ZN(_04135_));
 AOI22_X2 _20968_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_04128_),
    .B1(_04135_),
    .B2(_04133_),
    .ZN(_14488_));
 INV_X1 _20969_ (.A(_15979_),
    .ZN(_14498_));
 NAND2_X1 _20970_ (.A1(_04127_),
    .A2(_03857_),
    .ZN(_14531_));
 INV_X1 _20971_ (.A(_15999_),
    .ZN(_14539_));
 OR2_X1 _20972_ (.A1(_00563_),
    .A2(_03778_),
    .ZN(_04136_));
 OAI21_X1 _20973_ (.A(_04136_),
    .B1(_04131_),
    .B2(_03955_),
    .ZN(_04137_));
 AOI22_X2 _20974_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(_04128_),
    .B1(_04137_),
    .B2(_04133_),
    .ZN(_14558_));
 NAND2_X1 _20975_ (.A1(_03824_),
    .A2(net322),
    .ZN(_14576_));
 INV_X1 _20976_ (.A(_16022_),
    .ZN(_14597_));
 BUF_X8 _20977_ (.A(_03832_),
    .Z(_04138_));
 NAND2_X1 _20978_ (.A1(net373),
    .A2(_03839_),
    .ZN(_14607_));
 NAND2_X1 _20979_ (.A1(_04127_),
    .A2(_03883_),
    .ZN(_14620_));
 INV_X1 _20980_ (.A(_16041_),
    .ZN(_14628_));
 CLKBUF_X3 _20981_ (.A(_03858_),
    .Z(_04139_));
 NAND2_X1 _20982_ (.A1(_03824_),
    .A2(_04139_),
    .ZN(_14642_));
 NAND2_X1 _20983_ (.A1(net373),
    .A2(_03848_),
    .ZN(_14647_));
 NAND2_X1 _20984_ (.A1(_04127_),
    .A2(_03891_),
    .ZN(_14660_));
 INV_X1 _20985_ (.A(_16057_),
    .ZN(_14668_));
 NAND2_X1 _20986_ (.A1(_03830_),
    .A2(_03858_),
    .ZN(_14682_));
 NAND2_X1 _20987_ (.A1(_04138_),
    .A2(_03857_),
    .ZN(_14687_));
 NAND2_X1 _20988_ (.A1(_04127_),
    .A2(_03898_),
    .ZN(_14703_));
 INV_X1 _20989_ (.A(_16070_),
    .ZN(_14711_));
 CLKBUF_X3 _20990_ (.A(_03869_),
    .Z(_04140_));
 NAND2_X1 _20991_ (.A1(_03830_),
    .A2(_04140_),
    .ZN(_14725_));
 NAND2_X4 _20992_ (.A1(_04138_),
    .A2(_03864_),
    .ZN(_14730_));
 NAND2_X1 _20993_ (.A1(_03848_),
    .A2(_03858_),
    .ZN(_14776_));
 NAND2_X1 _20994_ (.A1(_03824_),
    .A2(_03966_),
    .ZN(_14827_));
 NAND2_X1 _20995_ (.A1(_03857_),
    .A2(_04140_),
    .ZN(_14886_));
 BUF_X8 _20996_ (.A(_03840_),
    .Z(_04141_));
 NAND2_X1 _20997_ (.A1(_04141_),
    .A2(_03883_),
    .ZN(_14898_));
 BUF_X4 _20998_ (.A(_03909_),
    .Z(_04142_));
 NAND2_X1 _20999_ (.A1(_03824_),
    .A2(_04142_),
    .ZN(_14938_));
 NAND2_X1 _21000_ (.A1(_03864_),
    .A2(_03869_),
    .ZN(_14952_));
 NAND2_X1 _21001_ (.A1(net373),
    .A2(_03898_),
    .ZN(_14964_));
 NAND2_X1 _21002_ (.A1(_04140_),
    .A2(_03875_),
    .ZN(_15021_));
 BUF_X4 _21003_ (.A(_03919_),
    .Z(_04143_));
 NAND2_X1 _21004_ (.A1(_03830_),
    .A2(_04143_),
    .ZN(_15068_));
 NAND2_X1 _21005_ (.A1(net321),
    .A2(_03908_),
    .ZN(_15091_));
 NAND2_X1 _21006_ (.A1(_03839_),
    .A2(_04143_),
    .ZN(_15126_));
 NAND2_X1 _21007_ (.A1(net321),
    .A2(_03917_),
    .ZN(_15149_));
 NAND2_X1 _21008_ (.A1(_04140_),
    .A2(_03898_),
    .ZN(_15197_));
 NAND2_X1 _21009_ (.A1(_03864_),
    .A2(_04142_),
    .ZN(_15241_));
 NAND2_X1 _21010_ (.A1(_04140_),
    .A2(_03908_),
    .ZN(_15254_));
 NAND2_X1 _21011_ (.A1(_03864_),
    .A2(_04143_),
    .ZN(_15294_));
 NAND2_X1 _21012_ (.A1(_03963_),
    .A2(_03908_),
    .ZN(_15353_));
 NAND2_X1 _21013_ (.A1(_04140_),
    .A2(_03924_),
    .ZN(_15360_));
 NAND2_X1 _21014_ (.A1(_03891_),
    .A2(_04142_),
    .ZN(_15401_));
 NAND2_X1 _21015_ (.A1(_03966_),
    .A2(_03908_),
    .ZN(_15406_));
 NAND2_X1 _21016_ (.A1(_04140_),
    .A2(_03952_),
    .ZN(_15413_));
 INV_X1 _21017_ (.A(_15374_),
    .ZN(_15375_));
 NAND2_X1 _21018_ (.A1(_03891_),
    .A2(_04143_),
    .ZN(_15447_));
 NAND2_X1 _21019_ (.A1(_03966_),
    .A2(_03917_),
    .ZN(_15452_));
 NAND2_X1 _21020_ (.A1(_03908_),
    .A2(_04142_),
    .ZN(_15490_));
 NAND2_X1 _21021_ (.A1(_03963_),
    .A2(_03952_),
    .ZN(_15495_));
 NAND2_X1 _21022_ (.A1(_03908_),
    .A2(_04143_),
    .ZN(_15534_));
 NAND2_X1 _21023_ (.A1(_03966_),
    .A2(_03952_),
    .ZN(_15539_));
 NAND2_X1 _21024_ (.A1(_03917_),
    .A2(_04143_),
    .ZN(_15573_));
 NAND2_X1 _21025_ (.A1(_04143_),
    .A2(_03952_),
    .ZN(_15649_));
 INV_X2 _21026_ (.A(_15423_),
    .ZN(_15424_));
 NAND2_X1 _21027_ (.A1(_04143_),
    .A2(_03938_),
    .ZN(_15688_));
 OR2_X1 _21028_ (.A1(_00185_),
    .A2(_03778_),
    .ZN(_04144_));
 OAI21_X1 _21029_ (.A(_04144_),
    .B1(_04131_),
    .B2(_03940_),
    .ZN(_04145_));
 AOI22_X2 _21030_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A2(_04128_),
    .B1(_04145_),
    .B2(_04133_),
    .ZN(_14469_));
 NAND2_X1 _21031_ (.A1(_04127_),
    .A2(_03829_),
    .ZN(_14479_));
 NAND2_X1 _21032_ (.A1(_04127_),
    .A2(_03848_),
    .ZN(_14509_));
 INV_X1 _21033_ (.A(_15985_),
    .ZN(_14517_));
 NAND2_X1 _21034_ (.A1(_03953_),
    .A2(_04129_),
    .ZN(_04146_));
 OAI21_X1 _21035_ (.A(_04146_),
    .B1(_04129_),
    .B2(_00562_),
    .ZN(_04147_));
 AOI22_X2 _21036_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_04128_),
    .B1(_04147_),
    .B2(_04133_),
    .ZN(_14532_));
 NAND2_X1 _21037_ (.A1(_03824_),
    .A2(_03832_),
    .ZN(_14545_));
 INV_X1 _21038_ (.A(_16008_),
    .ZN(_14567_));
 INV_X1 _21039_ (.A(_16014_),
    .ZN(_14572_));
 NAND2_X1 _21040_ (.A1(_04127_),
    .A2(_03875_),
    .ZN(_14590_));
 INV_X1 _21041_ (.A(_16026_),
    .ZN(_14598_));
 NAND2_X1 _21042_ (.A1(_03830_),
    .A2(_03840_),
    .ZN(_14608_));
 OR2_X1 _21043_ (.A1(_00565_),
    .A2(_03778_),
    .ZN(_04148_));
 OAI21_X1 _21044_ (.A(_04148_),
    .B1(_04131_),
    .B2(_03959_),
    .ZN(_04149_));
 AOI22_X2 _21045_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(_04128_),
    .B1(_04149_),
    .B2(_04133_),
    .ZN(_14621_));
 NAND2_X1 _21046_ (.A1(_03814_),
    .A2(_03869_),
    .ZN(_14643_));
 NAND2_X1 _21047_ (.A1(_03839_),
    .A2(_03840_),
    .ZN(_14648_));
 NAND2_X1 _21048_ (.A1(_03961_),
    .A2(_04129_),
    .ZN(_04150_));
 OAI21_X1 _21049_ (.A(_04150_),
    .B1(_04129_),
    .B2(_00566_),
    .ZN(_04151_));
 AOI22_X2 _21050_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A2(_04128_),
    .B1(_04151_),
    .B2(_04133_),
    .ZN(_14661_));
 NAND2_X1 _21051_ (.A1(_03824_),
    .A2(_03869_),
    .ZN(_14683_));
 NAND2_X1 _21052_ (.A1(_04141_),
    .A2(_03848_),
    .ZN(_14688_));
 NAND2_X1 _21053_ (.A1(_03964_),
    .A2(_04129_),
    .ZN(_04152_));
 OAI21_X1 _21054_ (.A(_04152_),
    .B1(_04129_),
    .B2(_00567_),
    .ZN(_04153_));
 AOI22_X2 _21055_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A2(_04128_),
    .B1(_04153_),
    .B2(_04133_),
    .ZN(_14704_));
 NAND2_X1 _21056_ (.A1(_04141_),
    .A2(_03857_),
    .ZN(_14731_));
 NAND2_X1 _21057_ (.A1(_04127_),
    .A2(_03907_),
    .ZN(_14752_));
 NAND2_X1 _21058_ (.A1(_03839_),
    .A2(_03869_),
    .ZN(_14777_));
 NAND2_X4 _21059_ (.A1(_04138_),
    .A2(_03875_),
    .ZN(_14785_));
 NAND2_X1 _21060_ (.A1(_04127_),
    .A2(_03917_),
    .ZN(_14806_));
 NAND2_X1 _21061_ (.A1(_03857_),
    .A2(_03858_),
    .ZN(_14833_));
 NAND2_X4 _21062_ (.A1(_04138_),
    .A2(_03883_),
    .ZN(_14841_));
 NAND2_X1 _21063_ (.A1(_03790_),
    .A2(_03924_),
    .ZN(_14861_));
 NAND2_X1 _21064_ (.A1(_03790_),
    .A2(_03952_),
    .ZN(_14918_));
 NAND2_X1 _21065_ (.A1(_03814_),
    .A2(_04143_),
    .ZN(_14939_));
 NAND2_X1 _21066_ (.A1(net321),
    .A2(_03891_),
    .ZN(_14965_));
 NAND2_X1 _21067_ (.A1(_03830_),
    .A2(_04142_),
    .ZN(_15009_));
 NAND2_X1 _21068_ (.A1(net373),
    .A2(_03907_),
    .ZN(_15033_));
 NAND2_X1 _21069_ (.A1(_04139_),
    .A2(_03891_),
    .ZN(_15082_));
 NAND2_X1 _21070_ (.A1(_04139_),
    .A2(_03898_),
    .ZN(_15140_));
 NAND2_X1 _21071_ (.A1(_03857_),
    .A2(_04142_),
    .ZN(_15185_));
 NAND2_X1 _21072_ (.A1(net373),
    .A2(_03952_),
    .ZN(_15208_));
 NAND2_X1 _21073_ (.A1(_03857_),
    .A2(_03919_),
    .ZN(_15242_));
 NAND2_X1 _21074_ (.A1(net321),
    .A2(_03952_),
    .ZN(_15265_));
 NAND2_X1 _21075_ (.A1(_04139_),
    .A2(_03924_),
    .ZN(_15308_));
 NAND2_X1 _21076_ (.A1(_03883_),
    .A2(_03909_),
    .ZN(_15349_));
 NAND2_X1 _21077_ (.A1(_03966_),
    .A2(_03897_),
    .ZN(_15354_));
 NAND2_X1 _21078_ (.A1(_03883_),
    .A2(_03919_),
    .ZN(_15402_));
 NAND2_X1 _21079_ (.A1(_03898_),
    .A2(_03919_),
    .ZN(_15491_));
 NAND2_X1 _21080_ (.A1(_03966_),
    .A2(_03924_),
    .ZN(_15496_));
 NAND2_X1 _21081_ (.A1(_04142_),
    .A2(_03929_),
    .ZN(_15611_));
 NAND2_X1 _21082_ (.A1(_03790_),
    .A2(_03823_),
    .ZN(_14475_));
 OR2_X1 _21083_ (.A1(_00559_),
    .A2(_03778_),
    .ZN(_04154_));
 OAI21_X1 _21084_ (.A(_04154_),
    .B1(_04131_),
    .B2(_03946_),
    .ZN(_04155_));
 AOI22_X2 _21085_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A2(_04128_),
    .B1(_04155_),
    .B2(_04133_),
    .ZN(_14480_));
 NAND2_X1 _21086_ (.A1(_03790_),
    .A2(_03839_),
    .ZN(_14490_));
 INV_X1 _21087_ (.A(_15977_),
    .ZN(_14500_));
 OR2_X1 _21088_ (.A1(_00561_),
    .A2(_03778_),
    .ZN(_04156_));
 OAI21_X1 _21089_ (.A(_04156_),
    .B1(_04131_),
    .B2(_03950_),
    .ZN(_04157_));
 AOI22_X2 _21090_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A2(_04128_),
    .B1(_04157_),
    .B2(_04133_),
    .ZN(_14510_));
 INV_X1 _21091_ (.A(_15987_),
    .ZN(_14518_));
 INV_X1 _21092_ (.A(_15997_),
    .ZN(_14541_));
 NAND2_X1 _21093_ (.A1(_03814_),
    .A2(net322),
    .ZN(_14546_));
 NAND2_X1 _21094_ (.A1(_03790_),
    .A2(_03864_),
    .ZN(_14560_));
 INV_X1 _21095_ (.A(_16012_),
    .ZN(_14568_));
 INV_X1 _21096_ (.A(_16016_),
    .ZN(_14573_));
 NAND2_X1 _21097_ (.A1(_03830_),
    .A2(_03832_),
    .ZN(_14578_));
 OR2_X1 _21098_ (.A1(_00564_),
    .A2(_03778_),
    .ZN(_04158_));
 OAI21_X1 _21099_ (.A(_04158_),
    .B1(_04131_),
    .B2(_03957_),
    .ZN(_04159_));
 AOI22_X2 _21100_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A2(_03798_),
    .B1(_04159_),
    .B2(_03752_),
    .ZN(_14591_));
 INV_X1 _21101_ (.A(_16035_),
    .ZN(_14630_));
 INV_X1 _21102_ (.A(_16053_),
    .ZN(_14670_));
 INV_X1 _21103_ (.A(_16066_),
    .ZN(_14713_));
 NAND2_X1 _21104_ (.A1(_03839_),
    .A2(_03858_),
    .ZN(_14727_));
 OR2_X1 _21105_ (.A1(_00568_),
    .A2(_03778_),
    .ZN(_04160_));
 OAI21_X1 _21106_ (.A(_04160_),
    .B1(_04131_),
    .B2(_03967_),
    .ZN(_04161_));
 AOI22_X2 _21107_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A2(_03798_),
    .B1(_04161_),
    .B2(_03752_),
    .ZN(_14753_));
 NAND2_X1 _21108_ (.A1(_04141_),
    .A2(_03864_),
    .ZN(_14786_));
 NAND2_X1 _21109_ (.A1(_03969_),
    .A2(_04129_),
    .ZN(_04162_));
 BUF_X2 _21110_ (.A(_00599_),
    .Z(_04163_));
 OAI21_X1 _21111_ (.A(_04162_),
    .B1(_04129_),
    .B2(_04163_),
    .ZN(_04164_));
 AOI22_X2 _21112_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(_03798_),
    .B1(_04164_),
    .B2(_03752_),
    .ZN(_14807_));
 NAND2_X1 _21113_ (.A1(_03830_),
    .A2(_03963_),
    .ZN(_14829_));
 NAND2_X1 _21114_ (.A1(_03848_),
    .A2(_03869_),
    .ZN(_14834_));
 NAND2_X1 _21115_ (.A1(_04141_),
    .A2(_03875_),
    .ZN(_14842_));
 OR2_X1 _21116_ (.A1(_00630_),
    .A2(_03778_),
    .ZN(_04165_));
 OAI21_X1 _21117_ (.A(_04165_),
    .B1(_04131_),
    .B2(_03971_),
    .ZN(_04166_));
 AOI22_X2 _21118_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(_03798_),
    .B1(_04166_),
    .B2(_03752_),
    .ZN(_14862_));
 NAND2_X1 _21119_ (.A1(_04139_),
    .A2(_03864_),
    .ZN(_14888_));
 NAND2_X1 _21120_ (.A1(_04138_),
    .A2(_03891_),
    .ZN(_14900_));
 OR2_X1 _21121_ (.A1(_00661_),
    .A2(_03778_),
    .ZN(_04167_));
 OAI21_X1 _21122_ (.A(_04167_),
    .B1(_03750_),
    .B2(_03503_),
    .ZN(_04168_));
 AOI22_X2 _21123_ (.A1(_03499_),
    .A2(_03798_),
    .B1(_04168_),
    .B2(_03752_),
    .ZN(_14919_));
 NAND2_X1 _21124_ (.A1(_04139_),
    .A2(_03875_),
    .ZN(_14954_));
 NAND2_X1 _21125_ (.A1(_03824_),
    .A2(_03919_),
    .ZN(_15010_));
 NAND2_X1 _21126_ (.A1(_04139_),
    .A2(_03883_),
    .ZN(_15023_));
 NAND2_X1 _21127_ (.A1(net321),
    .A2(_03897_),
    .ZN(_15034_));
 NAND2_X1 _21128_ (.A1(_03839_),
    .A2(_03909_),
    .ZN(_15070_));
 NAND2_X1 _21129_ (.A1(_04140_),
    .A2(_03883_),
    .ZN(_15083_));
 NAND2_X1 _21130_ (.A1(_03832_),
    .A2(_03917_),
    .ZN(_15093_));
 NAND2_X1 _21131_ (.A1(_03848_),
    .A2(_03909_),
    .ZN(_15128_));
 NAND2_X1 _21132_ (.A1(_04140_),
    .A2(_03890_),
    .ZN(_15141_));
 NAND2_X1 _21133_ (.A1(_03832_),
    .A2(_03924_),
    .ZN(_15151_));
 NAND2_X1 _21134_ (.A1(_03848_),
    .A2(_03919_),
    .ZN(_15186_));
 NAND2_X1 _21135_ (.A1(_04139_),
    .A2(_03907_),
    .ZN(_15199_));
 NAND2_X1 _21136_ (.A1(net322),
    .A2(_03924_),
    .ZN(_15209_));
 NAND2_X1 _21137_ (.A1(_04139_),
    .A2(_03917_),
    .ZN(_15256_));
 NAND2_X1 _21138_ (.A1(_03875_),
    .A2(_03909_),
    .ZN(_15296_));
 NAND2_X1 _21139_ (.A1(_04140_),
    .A2(_03916_),
    .ZN(_15309_));
 NAND2_X1 _21140_ (.A1(_03875_),
    .A2(_03919_),
    .ZN(_15350_));
 NAND2_X1 _21141_ (.A1(_04139_),
    .A2(_03929_),
    .ZN(_15362_));
 NAND2_X1 _21142_ (.A1(_03963_),
    .A2(_03916_),
    .ZN(_15408_));
 INV_X1 _21143_ (.A(_15215_),
    .ZN(_15216_));
 NAND2_X1 _21144_ (.A1(_03898_),
    .A2(_03909_),
    .ZN(_15449_));
 NAND2_X1 _21145_ (.A1(_03963_),
    .A2(_03923_),
    .ZN(_15454_));
 NAND2_X1 _21146_ (.A1(_04142_),
    .A2(_03916_),
    .ZN(_15536_));
 NAND2_X1 _21147_ (.A1(_04142_),
    .A2(_03923_),
    .ZN(_15575_));
 NAND2_X1 _21148_ (.A1(_04143_),
    .A2(_03923_),
    .ZN(_15612_));
 INV_X2 _21149_ (.A(_15422_),
    .ZN(_15467_));
 NAND2_X2 _21150_ (.A1(_04142_),
    .A2(_03938_),
    .ZN(_15651_));
 NOR2_X2 _21151_ (.A1(_00137_),
    .A2(_04115_),
    .ZN(_04169_));
 INV_X1 _21152_ (.A(_04169_),
    .ZN(_15756_));
 INV_X1 _21153_ (.A(_14585_),
    .ZN(_14586_));
 INV_X1 _21154_ (.A(_14616_),
    .ZN(_14617_));
 INV_X1 _21155_ (.A(_14656_),
    .ZN(_14657_));
 INV_X1 _21156_ (.A(_14677_),
    .ZN(_14678_));
 INV_X1 _21157_ (.A(_14696_),
    .ZN(_14697_));
 INV_X1 _21158_ (.A(_14720_),
    .ZN(_14721_));
 INV_X1 _21159_ (.A(_14739_),
    .ZN(_14740_));
 INV_X2 _21160_ (.A(_14766_),
    .ZN(_14767_));
 INV_X1 _21161_ (.A(_14793_),
    .ZN(_14794_));
 INV_X2 _21162_ (.A(_14804_),
    .ZN(_14818_));
 INV_X1 _21163_ (.A(_14817_),
    .ZN(_14819_));
 INV_X1 _21164_ (.A(_14849_),
    .ZN(_14850_));
 INV_X2 _21165_ (.A(_14859_),
    .ZN(_14873_));
 INV_X1 _21166_ (.A(_14872_),
    .ZN(_14874_));
 INV_X1 _21167_ (.A(_14907_),
    .ZN(_14908_));
 INV_X1 _21168_ (.A(_14916_),
    .ZN(_14930_));
 INV_X1 _21169_ (.A(_14929_),
    .ZN(_14931_));
 INV_X1 _21170_ (.A(_14963_),
    .ZN(_14980_));
 INV_X1 _21171_ (.A(_14973_),
    .ZN(_14974_));
 INV_X1 _21172_ (.A(_14987_),
    .ZN(_14989_));
 INV_X1 _21173_ (.A(_15000_),
    .ZN(_15002_));
 INV_X1 _21174_ (.A(_15017_),
    .ZN(_15018_));
 INV_X1 _21175_ (.A(_15041_),
    .ZN(_15042_));
 INV_X1 _21176_ (.A(_15053_),
    .ZN(_15055_));
 INV_X1 _21177_ (.A(_15077_),
    .ZN(_15078_));
 INV_X1 _21178_ (.A(_15100_),
    .ZN(_15101_));
 INV_X1 _21179_ (.A(_15110_),
    .ZN(_15112_));
 INV_X1 _21180_ (.A(_15120_),
    .ZN(_15121_));
 INV_X1 _21181_ (.A(_15135_),
    .ZN(_15136_));
 INV_X1 _21182_ (.A(_15167_),
    .ZN(_15168_));
 INV_X1 _21183_ (.A(_15177_),
    .ZN(_15178_));
 INV_X1 _21184_ (.A(_15193_),
    .ZN(_15194_));
 INV_X1 _21185_ (.A(_15225_),
    .ZN(_15227_));
 INV_X1 _21186_ (.A(_15234_),
    .ZN(_15235_));
 INV_X1 _21187_ (.A(_15250_),
    .ZN(_15251_));
 INV_X1 _21188_ (.A(_15277_),
    .ZN(_15278_));
 INV_X1 _21189_ (.A(_15287_),
    .ZN(_15288_));
 INV_X1 _21190_ (.A(_15303_),
    .ZN(_15304_));
 INV_X1 _21191_ (.A(_15324_),
    .ZN(_15325_));
 INV_X1 _21192_ (.A(_15332_),
    .ZN(_15334_));
 INV_X1 _21193_ (.A(_15341_),
    .ZN(_15342_));
 INV_X1 _21194_ (.A(_15385_),
    .ZN(_15386_));
 INV_X1 _21195_ (.A(_15394_),
    .ZN(_15395_));
 INV_X1 _21196_ (.A(_15431_),
    .ZN(_15432_));
 INV_X1 _21197_ (.A(_15440_),
    .ZN(_15441_));
 INV_X1 _21198_ (.A(_15474_),
    .ZN(_15476_));
 INV_X1 _21199_ (.A(_15483_),
    .ZN(_15484_));
 INV_X2 _21200_ (.A(_15506_),
    .ZN(_15507_));
 INV_X1 _21201_ (.A(_15518_),
    .ZN(_15519_));
 INV_X1 _21202_ (.A(_15527_),
    .ZN(_15528_));
 INV_X1 _21203_ (.A(_15557_),
    .ZN(_15558_));
 INV_X1 _21204_ (.A(_15566_),
    .ZN(_15567_));
 INV_X1 _21205_ (.A(_15594_),
    .ZN(_15596_));
 INV_X1 _21206_ (.A(_15603_),
    .ZN(_15604_));
 INV_X1 _21207_ (.A(_15633_),
    .ZN(_15634_));
 INV_X1 _21208_ (.A(_15642_),
    .ZN(_15643_));
 INV_X1 _21209_ (.A(_15657_),
    .ZN(_15661_));
 INV_X1 _21210_ (.A(_15666_),
    .ZN(_15667_));
 INV_X1 _21211_ (.A(_15672_),
    .ZN(_15673_));
 INV_X1 _21212_ (.A(_15681_),
    .ZN(_15682_));
 INV_X1 _21213_ (.A(_15695_),
    .ZN(_15696_));
 INV_X1 _21214_ (.A(_15702_),
    .ZN(_15703_));
 INV_X1 _21215_ (.A(_15708_),
    .ZN(_15709_));
 INV_X1 _21216_ (.A(_15716_),
    .ZN(_15717_));
 INV_X1 _21217_ (.A(_15729_),
    .ZN(_15730_));
 INV_X1 _21218_ (.A(_15737_),
    .ZN(_15747_));
 INV_X1 _21219_ (.A(_15746_),
    .ZN(_15748_));
 INV_X1 _21220_ (.A(_14486_),
    .ZN(_14513_));
 INV_X1 _21221_ (.A(_14506_),
    .ZN(_14536_));
 INV_X1 _21222_ (.A(_14529_),
    .ZN(_14563_));
 INV_X1 _21223_ (.A(_14552_),
    .ZN(_14594_));
 INV_X1 _21224_ (.A(_14584_),
    .ZN(_14625_));
 INV_X1 _21225_ (.A(_14615_),
    .ZN(_14665_));
 INV_X1 _21226_ (.A(_14636_),
    .ZN(_14679_));
 INV_X1 _21227_ (.A(_14655_),
    .ZN(_14708_));
 INV_X1 _21228_ (.A(_14676_),
    .ZN(_14722_));
 INV_X1 _21229_ (.A(_14695_),
    .ZN(_14756_));
 INV_X1 _21230_ (.A(_14719_),
    .ZN(_14768_));
 INV_X1 _21231_ (.A(_14738_),
    .ZN(_14810_));
 INV_X1 _21232_ (.A(_14749_),
    .ZN(_14820_));
 INV_X1 _21233_ (.A(_14762_),
    .ZN(_14824_));
 INV_X1 _21234_ (.A(_14765_),
    .ZN(_14823_));
 INV_X1 _21235_ (.A(_14774_),
    .ZN(_14837_));
 INV_X1 _21236_ (.A(_14792_),
    .ZN(_14865_));
 INV_X1 _21237_ (.A(_14803_),
    .ZN(_14875_));
 INV_X1 _21238_ (.A(_14816_),
    .ZN(_14878_));
 INV_X1 _21239_ (.A(_14848_),
    .ZN(_14922_));
 INV_X1 _21240_ (.A(_14858_),
    .ZN(_14932_));
 INV_X1 _21241_ (.A(_14871_),
    .ZN(_14935_));
 INV_X1 _21242_ (.A(_14884_),
    .ZN(_14957_));
 INV_X1 _21243_ (.A(_14896_),
    .ZN(_14979_));
 INV_X1 _21244_ (.A(_14906_),
    .ZN(_14988_));
 INV_X1 _21245_ (.A(_14915_),
    .ZN(_15001_));
 INV_X1 _21246_ (.A(_14928_),
    .ZN(_15005_));
 INV_X1 _21247_ (.A(_14946_),
    .ZN(_15026_));
 INV_X1 _21248_ (.A(_14950_),
    .ZN(_15029_));
 INV_X1 _21249_ (.A(_14962_),
    .ZN(_15047_));
 INV_X1 _21250_ (.A(_14972_),
    .ZN(_15054_));
 INV_X1 _21251_ (.A(_14986_),
    .ZN(_15056_));
 INV_X1 _21252_ (.A(_14995_),
    .ZN(_15060_));
 INV_X1 _21253_ (.A(_14999_),
    .ZN(_15065_));
 INV_X1 _21254_ (.A(_15016_),
    .ZN(_15086_));
 INV_X1 _21255_ (.A(_15040_),
    .ZN(_15111_));
 INV_X1 _21256_ (.A(_15052_),
    .ZN(_15113_));
 INV_X1 _21257_ (.A(_15076_),
    .ZN(_15144_));
 INV_X1 _21258_ (.A(_15099_),
    .ZN(_15169_));
 INV_X1 _21259_ (.A(_15109_),
    .ZN(_15170_));
 INV_X1 _21260_ (.A(_15119_),
    .ZN(_15181_));
 INV_X1 _21261_ (.A(_15134_),
    .ZN(_15202_));
 INV_X1 _21262_ (.A(_15166_),
    .ZN(_15226_));
 INV_X1 _21263_ (.A(_15176_),
    .ZN(_15238_));
 INV_X1 _21264_ (.A(_15192_),
    .ZN(_15259_));
 INV_X1 _21265_ (.A(_15224_),
    .ZN(_15280_));
 INV_X1 _21266_ (.A(_15233_),
    .ZN(_15291_));
 INV_X1 _21267_ (.A(_15249_),
    .ZN(_15312_));
 INV_X1 _21268_ (.A(_15276_),
    .ZN(_15333_));
 INV_X1 _21269_ (.A(_15286_),
    .ZN(_15345_));
 INV_X1 _21270_ (.A(_15302_),
    .ZN(_15365_));
 INV_X1 _21271_ (.A(_15323_),
    .ZN(_15378_));
 INV_X1 _21272_ (.A(_15331_),
    .ZN(_15387_));
 INV_X1 _21273_ (.A(_15340_),
    .ZN(_15398_));
 INV_X1 _21274_ (.A(_15384_),
    .ZN(_15433_));
 INV_X1 _21275_ (.A(_15393_),
    .ZN(_15444_));
 INV_X1 _21276_ (.A(_15430_),
    .ZN(_15475_));
 INV_X1 _21277_ (.A(_15439_),
    .ZN(_15487_));
 INV_X1 _21278_ (.A(_15473_),
    .ZN(_15520_));
 INV_X1 _21279_ (.A(_15482_),
    .ZN(_15531_));
 INV_X2 _21280_ (.A(_15505_),
    .ZN(_15546_));
 INV_X1 _21281_ (.A(_15517_),
    .ZN(_15559_));
 INV_X1 _21282_ (.A(_15526_),
    .ZN(_15570_));
 INV_X1 _21283_ (.A(_15556_),
    .ZN(_15595_));
 INV_X1 _21284_ (.A(_15565_),
    .ZN(_15607_));
 INV_X1 _21285_ (.A(_15593_),
    .ZN(_15635_));
 INV_X1 _21286_ (.A(_15602_),
    .ZN(_15646_));
 INV_X1 _21287_ (.A(_15618_),
    .ZN(_15658_));
 INV_X1 _21288_ (.A(_15632_),
    .ZN(_15674_));
 INV_X1 _21289_ (.A(_15641_),
    .ZN(_15685_));
 INV_X1 _21290_ (.A(_15656_),
    .ZN(_15697_));
 INV_X1 _21291_ (.A(_15671_),
    .ZN(_15710_));
 INV_X1 _21292_ (.A(_15680_),
    .ZN(_15720_));
 INV_X1 _21293_ (.A(_15694_),
    .ZN(_15731_));
 INV_X1 _21294_ (.A(_15715_),
    .ZN(_15751_));
 BUF_X4 _21295_ (.A(_11865_),
    .Z(_04170_));
 CLKBUF_X3 _21296_ (.A(_04170_),
    .Z(_04171_));
 BUF_X2 _21297_ (.A(_04171_),
    .Z(_04172_));
 CLKBUF_X3 _21298_ (.A(_03504_),
    .Z(_04173_));
 CLKBUF_X2 _21299_ (.A(_04173_),
    .Z(_04174_));
 OR3_X1 _21300_ (.A1(_00185_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04175_));
 BUF_X4 _21301_ (.A(_03755_),
    .Z(_04176_));
 CLKBUF_X3 _21302_ (.A(_04176_),
    .Z(_04177_));
 CLKBUF_X3 _21303_ (.A(_04177_),
    .Z(_04178_));
 OAI21_X1 _21304_ (.A(_04175_),
    .B1(_04178_),
    .B2(_16250_),
    .ZN(_15771_));
 CLKBUF_X3 _21305_ (.A(_04176_),
    .Z(_04179_));
 BUF_X8 _21306_ (.A(_03508_),
    .Z(_04180_));
 XNOR2_X1 _21307_ (.A(_11173_),
    .B(_04180_),
    .ZN(_04181_));
 NOR2_X2 _21308_ (.A1(_04181_),
    .A2(_04179_),
    .ZN(_04182_));
 NAND2_X1 _21309_ (.A1(net278),
    .A2(_03495_),
    .ZN(_04183_));
 BUF_X4 _21310_ (.A(_03498_),
    .Z(_04184_));
 BUF_X4 _21311_ (.A(_03491_),
    .Z(_04185_));
 OAI222_X2 _21312_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .B2(_04173_),
    .C1(_03796_),
    .C2(_04185_),
    .ZN(_04186_));
 OAI21_X2 _21313_ (.A(_04183_),
    .B1(_04186_),
    .B2(_03495_),
    .ZN(_04187_));
 AOI21_X2 _21314_ (.A(_04182_),
    .B1(_04187_),
    .B2(_04178_),
    .ZN(_14465_));
 XNOR2_X1 _21315_ (.A(_11379_),
    .B(_04180_),
    .ZN(_04188_));
 NOR2_X1 _21316_ (.A1(_04179_),
    .A2(_04188_),
    .ZN(_04189_));
 BUF_X2 _21317_ (.A(_03497_),
    .Z(_04190_));
 OAI22_X1 _21318_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .A2(_04173_),
    .B1(_04190_),
    .B2(net364),
    .ZN(_04191_));
 OAI22_X1 _21319_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .B1(_03820_),
    .B2(_04185_),
    .ZN(_04192_));
 CLKBUF_X3 _21320_ (.A(_03497_),
    .Z(_04193_));
 CLKBUF_X3 _21321_ (.A(_04193_),
    .Z(_04194_));
 AOI21_X1 _21322_ (.A(_04191_),
    .B1(_04192_),
    .B2(_04194_),
    .ZN(_04195_));
 AOI21_X1 _21323_ (.A(_04189_),
    .B1(_04195_),
    .B2(_04178_),
    .ZN(_15777_));
 BUF_X4 _21324_ (.A(_03508_),
    .Z(_04196_));
 XNOR2_X1 _21325_ (.A(_16266_),
    .B(_04196_),
    .ZN(_04197_));
 BUF_X4 _21326_ (.A(_03498_),
    .Z(_04198_));
 BUF_X4 _21327_ (.A(_03504_),
    .Z(_04199_));
 BUF_X4 _21328_ (.A(_03491_),
    .Z(_04200_));
 OAI222_X2 _21329_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .B2(_04199_),
    .C1(_11967_),
    .C2(_04200_),
    .ZN(_04201_));
 MUX2_X1 _21330_ (.A(_03815_),
    .B(_04201_),
    .S(_04193_),
    .Z(_04202_));
 CLKBUF_X3 _21331_ (.A(_04176_),
    .Z(_04203_));
 MUX2_X1 _21332_ (.A(_04197_),
    .B(_04202_),
    .S(_04203_),
    .Z(_15781_));
 XNOR2_X1 _21333_ (.A(_16274_),
    .B(net290),
    .ZN(_04204_));
 OAI222_X2 _21334_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .B2(_04173_),
    .C1(_12008_),
    .C2(_04185_),
    .ZN(_04205_));
 NAND2_X1 _21335_ (.A1(_04190_),
    .A2(_04205_),
    .ZN(_04206_));
 OAI21_X1 _21336_ (.A(_04206_),
    .B1(_04194_),
    .B2(net330),
    .ZN(_04207_));
 MUX2_X1 _21337_ (.A(_04204_),
    .B(_04207_),
    .S(_04203_),
    .Z(_15785_));
 XNOR2_X1 _21338_ (.A(_16282_),
    .B(net290),
    .ZN(_04208_));
 NOR2_X1 _21339_ (.A1(_04203_),
    .A2(_04208_),
    .ZN(_04209_));
 OAI22_X1 _21340_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .A2(_04173_),
    .B1(_04190_),
    .B2(_03831_),
    .ZN(_04210_));
 OAI22_X1 _21341_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .B1(_12051_),
    .B2(_04185_),
    .ZN(_04211_));
 AOI21_X1 _21342_ (.A(_04210_),
    .B1(_04211_),
    .B2(_04194_),
    .ZN(_04212_));
 AOI21_X2 _21343_ (.A(_04209_),
    .B1(_04212_),
    .B2(_04178_),
    .ZN(_15789_));
 XNOR2_X1 _21344_ (.A(_16290_),
    .B(_04180_),
    .ZN(_04213_));
 OAI222_X2 _21345_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .B2(_04173_),
    .C1(_03854_),
    .C2(_04185_),
    .ZN(_04214_));
 NAND2_X1 _21346_ (.A1(_04190_),
    .A2(_04214_),
    .ZN(_04215_));
 OAI21_X1 _21347_ (.A(_04215_),
    .B1(_04194_),
    .B2(net361),
    .ZN(_04216_));
 MUX2_X1 _21348_ (.A(_04213_),
    .B(_04216_),
    .S(_04203_),
    .Z(_15793_));
 XNOR2_X1 _21349_ (.A(_16298_),
    .B(_04180_),
    .ZN(_04217_));
 OAI222_X2 _21350_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .B2(_03504_),
    .C1(_03861_),
    .C2(_03491_),
    .ZN(_04218_));
 NOR2_X1 _21351_ (.A1(_03495_),
    .A2(_04218_),
    .ZN(_04219_));
 AOI21_X1 _21352_ (.A(_04219_),
    .B1(_03495_),
    .B2(_03849_),
    .ZN(_04220_));
 MUX2_X1 _21353_ (.A(_04217_),
    .B(_04220_),
    .S(_04203_),
    .Z(_15797_));
 OR3_X1 _21354_ (.A1(_00564_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04221_));
 OAI21_X1 _21355_ (.A(_04221_),
    .B1(_16306_),
    .B2(_04178_),
    .ZN(_15801_));
 XNOR2_X1 _21356_ (.A(_16313_),
    .B(_03508_),
    .ZN(_04222_));
 NOR2_X1 _21357_ (.A1(_04203_),
    .A2(_04222_),
    .ZN(_04223_));
 OAI22_X1 _21358_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .A2(_04173_),
    .B1(_04190_),
    .B2(_03867_),
    .ZN(_04224_));
 OAI22_X1 _21359_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B1(_03880_),
    .B2(_04185_),
    .ZN(_04225_));
 AOI21_X1 _21360_ (.A(_04224_),
    .B1(_04225_),
    .B2(_04194_),
    .ZN(_04226_));
 AOI21_X1 _21361_ (.A(_04223_),
    .B1(_04226_),
    .B2(_04178_),
    .ZN(_15805_));
 XNOR2_X1 _21362_ (.A(_16322_),
    .B(net290),
    .ZN(_04227_));
 OAI222_X2 _21363_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .B2(_04199_),
    .C1(_03889_),
    .C2(_04200_),
    .ZN(_04228_));
 MUX2_X1 _21364_ (.A(_03543_),
    .B(_04228_),
    .S(_04193_),
    .Z(_04229_));
 MUX2_X1 _21365_ (.A(_04227_),
    .B(_04229_),
    .S(_04203_),
    .Z(_15809_));
 OR3_X1 _21366_ (.A1(_00567_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04230_));
 OAI21_X1 _21367_ (.A(_04230_),
    .B1(_04178_),
    .B2(_16329_),
    .ZN(_15813_));
 OR3_X1 _21368_ (.A1(_00568_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04231_));
 OAI21_X1 _21369_ (.A(_04231_),
    .B1(_04178_),
    .B2(_16337_),
    .ZN(_15817_));
 BUF_X4 _21370_ (.A(_03508_),
    .Z(_04232_));
 XNOR2_X1 _21371_ (.A(_04232_),
    .B(_16341_),
    .ZN(_04233_));
 BUF_X4 _21372_ (.A(_03504_),
    .Z(_04234_));
 OAI222_X2 _21373_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .B2(_04234_),
    .C1(_03914_),
    .C2(_04185_),
    .ZN(_04235_));
 NAND2_X1 _21374_ (.A1(_04190_),
    .A2(_04235_),
    .ZN(_04236_));
 OAI21_X1 _21375_ (.A(_04236_),
    .B1(_04194_),
    .B2(_12473_),
    .ZN(_04237_));
 MUX2_X1 _21376_ (.A(_04233_),
    .B(_04237_),
    .S(_04203_),
    .Z(_15821_));
 XNOR2_X1 _21377_ (.A(_04232_),
    .B(_16349_),
    .ZN(_04238_));
 OAI222_X2 _21378_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .B2(_04234_),
    .C1(_03921_),
    .C2(_04185_),
    .ZN(_04239_));
 NAND2_X1 _21379_ (.A1(_04190_),
    .A2(_04239_),
    .ZN(_04240_));
 OAI21_X1 _21380_ (.A(_04240_),
    .B1(_04194_),
    .B2(_12580_),
    .ZN(_04241_));
 MUX2_X1 _21381_ (.A(_04238_),
    .B(_04241_),
    .S(_04203_),
    .Z(_15825_));
 XNOR2_X1 _21382_ (.A(_04232_),
    .B(_16357_),
    .ZN(_04242_));
 BUF_X2 _21383_ (.A(_03497_),
    .Z(_04243_));
 OAI222_X2 _21384_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .B2(_04234_),
    .C1(_03928_),
    .C2(_04185_),
    .ZN(_04244_));
 NAND2_X1 _21385_ (.A1(_04243_),
    .A2(_04244_),
    .ZN(_04245_));
 OAI21_X1 _21386_ (.A(_04245_),
    .B1(_04194_),
    .B2(_12656_),
    .ZN(_04246_));
 MUX2_X1 _21387_ (.A(_04242_),
    .B(_04246_),
    .S(_04203_),
    .Z(_15829_));
 OR3_X1 _21388_ (.A1(_03800_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04247_));
 BUF_X2 _21389_ (.A(_04176_),
    .Z(_04248_));
 OAI21_X1 _21390_ (.A(_04247_),
    .B1(_16369_),
    .B2(_04248_),
    .ZN(_15833_));
 XNOR2_X1 _21391_ (.A(_04232_),
    .B(_16378_),
    .ZN(_04249_));
 OAI222_X2 _21392_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .B2(_03504_),
    .C1(_03812_),
    .C2(_04200_),
    .ZN(_04250_));
 MUX2_X1 _21393_ (.A(_12825_),
    .B(_04250_),
    .S(_03497_),
    .Z(_04251_));
 CLKBUF_X3 _21394_ (.A(_04176_),
    .Z(_04252_));
 MUX2_X1 _21395_ (.A(_04249_),
    .B(_04251_),
    .S(_04252_),
    .Z(_15837_));
 XNOR2_X1 _21396_ (.A(_04232_),
    .B(_16386_),
    .ZN(_04253_));
 BUF_X4 _21397_ (.A(_03491_),
    .Z(_04254_));
 OAI222_X2 _21398_ (.A1(_04184_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .B2(_04234_),
    .C1(_03822_),
    .C2(_04254_),
    .ZN(_04255_));
 NAND2_X1 _21399_ (.A1(_04243_),
    .A2(_04255_),
    .ZN(_04256_));
 OAI21_X1 _21400_ (.A(_04256_),
    .B1(_04194_),
    .B2(net286),
    .ZN(_04257_));
 MUX2_X1 _21401_ (.A(_04253_),
    .B(_04257_),
    .S(_04252_),
    .Z(_15841_));
 XNOR2_X1 _21402_ (.A(_04232_),
    .B(_16394_),
    .ZN(_04258_));
 BUF_X4 _21403_ (.A(_03498_),
    .Z(_04259_));
 OAI222_X2 _21404_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .B2(_04234_),
    .C1(_03828_),
    .C2(_04254_),
    .ZN(_04260_));
 NAND2_X1 _21405_ (.A1(_04243_),
    .A2(_04260_),
    .ZN(_04261_));
 OAI21_X1 _21406_ (.A(_04261_),
    .B1(_04194_),
    .B2(net285),
    .ZN(_04262_));
 MUX2_X1 _21407_ (.A(_04258_),
    .B(_04262_),
    .S(_04252_),
    .Z(_15845_));
 OR3_X1 _21408_ (.A1(_03948_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04263_));
 OAI21_X1 _21409_ (.A(_04263_),
    .B1(_16398_),
    .B2(_04248_),
    .ZN(_15849_));
 XNOR2_X1 _21410_ (.A(_04232_),
    .B(_16405_),
    .ZN(_04264_));
 OAI222_X2 _21411_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .B2(_04234_),
    .C1(_03846_),
    .C2(_04254_),
    .ZN(_04265_));
 NAND2_X1 _21412_ (.A1(_04243_),
    .A2(_04265_),
    .ZN(_04266_));
 CLKBUF_X3 _21413_ (.A(_04193_),
    .Z(_04267_));
 OAI21_X1 _21414_ (.A(_04266_),
    .B1(_04267_),
    .B2(_13198_),
    .ZN(_04268_));
 MUX2_X1 _21415_ (.A(_04264_),
    .B(_04268_),
    .S(_04252_),
    .Z(_15853_));
 XNOR2_X1 _21416_ (.A(_04232_),
    .B(_16413_),
    .ZN(_04269_));
 OAI222_X2 _21417_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .B2(_04234_),
    .C1(_03855_),
    .C2(_04254_),
    .ZN(_04270_));
 NAND2_X1 _21418_ (.A1(_04243_),
    .A2(_04270_),
    .ZN(_04271_));
 OAI21_X1 _21419_ (.A(_04271_),
    .B1(_04267_),
    .B2(_13307_),
    .ZN(_04272_));
 MUX2_X1 _21420_ (.A(_04269_),
    .B(_04272_),
    .S(_04252_),
    .Z(_15857_));
 XNOR2_X1 _21421_ (.A(_04232_),
    .B(_16426_),
    .ZN(_04273_));
 OAI222_X2 _21422_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .B2(_04234_),
    .C1(_03862_),
    .C2(_04254_),
    .ZN(_04274_));
 NAND2_X1 _21423_ (.A1(_04243_),
    .A2(_04274_),
    .ZN(_04275_));
 OAI21_X1 _21424_ (.A(_04275_),
    .B1(_04267_),
    .B2(net350),
    .ZN(_04276_));
 MUX2_X1 _21425_ (.A(_04273_),
    .B(_04276_),
    .S(_04252_),
    .Z(_15861_));
 XNOR2_X1 _21426_ (.A(_04232_),
    .B(_16434_),
    .ZN(_04277_));
 OAI222_X2 _21427_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .B2(_04234_),
    .C1(_03873_),
    .C2(_04254_),
    .ZN(_04278_));
 NAND2_X1 _21428_ (.A1(_04243_),
    .A2(_04278_),
    .ZN(_04279_));
 OAI21_X1 _21429_ (.A(_04279_),
    .B1(_04267_),
    .B2(_13480_),
    .ZN(_04280_));
 MUX2_X1 _21430_ (.A(_04277_),
    .B(_04280_),
    .S(_04252_),
    .Z(_15865_));
 XNOR2_X1 _21431_ (.A(_04196_),
    .B(_16442_),
    .ZN(_04281_));
 OAI222_X2 _21432_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .B2(_04234_),
    .C1(_03881_),
    .C2(_04254_),
    .ZN(_04282_));
 NAND2_X1 _21433_ (.A1(_04243_),
    .A2(_04282_),
    .ZN(_04283_));
 OAI21_X1 _21434_ (.A(_04283_),
    .B1(_04267_),
    .B2(_13555_),
    .ZN(_04284_));
 MUX2_X1 _21435_ (.A(_04281_),
    .B(_04284_),
    .S(_04252_),
    .Z(_15869_));
 XNOR2_X1 _21436_ (.A(_04196_),
    .B(_16450_),
    .ZN(_04285_));
 OAI222_X2 _21437_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .B2(_04199_),
    .C1(_13686_),
    .C2(_04254_),
    .ZN(_04286_));
 NAND2_X1 _21438_ (.A1(_04243_),
    .A2(_04286_),
    .ZN(_04287_));
 OAI21_X1 _21439_ (.A(_04287_),
    .B1(_04267_),
    .B2(_13648_),
    .ZN(_04288_));
 MUX2_X1 _21440_ (.A(_04285_),
    .B(_04288_),
    .S(_04252_),
    .Z(_15873_));
 XNOR2_X1 _21441_ (.A(_04196_),
    .B(_16458_),
    .ZN(_04289_));
 OAI222_X2 _21442_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .B2(_04199_),
    .C1(_03139_),
    .C2(_04254_),
    .ZN(_04290_));
 NAND2_X1 _21443_ (.A1(_04243_),
    .A2(_04290_),
    .ZN(_04291_));
 OAI21_X1 _21444_ (.A(_04291_),
    .B1(_04267_),
    .B2(_03104_),
    .ZN(_04292_));
 MUX2_X1 _21445_ (.A(_04289_),
    .B(_04292_),
    .S(_04252_),
    .Z(_15877_));
 XNOR2_X1 _21446_ (.A(_04196_),
    .B(_16466_),
    .ZN(_04293_));
 OAI222_X2 _21447_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .B2(_04199_),
    .C1(_03906_),
    .C2(_04254_),
    .ZN(_04294_));
 NAND2_X1 _21448_ (.A1(_04193_),
    .A2(_04294_),
    .ZN(_04295_));
 OAI21_X1 _21449_ (.A(_04295_),
    .B1(_04267_),
    .B2(_03198_),
    .ZN(_04296_));
 MUX2_X1 _21450_ (.A(_04293_),
    .B(_04296_),
    .S(_04177_),
    .Z(_15881_));
 XNOR2_X1 _21451_ (.A(_04196_),
    .B(_16474_),
    .ZN(_04297_));
 OAI222_X2 _21452_ (.A1(_04259_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .B2(_04199_),
    .C1(_03915_),
    .C2(_04200_),
    .ZN(_04298_));
 NAND2_X1 _21453_ (.A1(_04193_),
    .A2(_04298_),
    .ZN(_04299_));
 OAI21_X1 _21454_ (.A(_04299_),
    .B1(_04267_),
    .B2(_03276_),
    .ZN(_04300_));
 MUX2_X1 _21455_ (.A(_04297_),
    .B(_04300_),
    .S(_04177_),
    .Z(_15885_));
 OR3_X1 _21456_ (.A1(_03971_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04301_));
 OAI21_X1 _21457_ (.A(_04301_),
    .B1(_16478_),
    .B2(_04248_),
    .ZN(_15889_));
 NOR2_X1 _21458_ (.A1(_03631_),
    .A2(_16313_),
    .ZN(_15901_));
 NAND2_X1 _21459_ (.A1(_11329_),
    .A2(_16301_),
    .ZN(_15905_));
 INV_X1 _21460_ (.A(_15919_),
    .ZN(_15912_));
 INV_X1 _21461_ (.A(_14472_),
    .ZN(_15956_));
 INV_X1 _21462_ (.A(_14502_),
    .ZN(_15989_));
 INV_X1 _21463_ (.A(_14520_),
    .ZN(_14522_));
 INV_X1 _21464_ (.A(_14543_),
    .ZN(_16018_));
 INV_X1 _21465_ (.A(_14565_),
    .ZN(_16024_));
 INV_X1 _21466_ (.A(_14575_),
    .ZN(_16030_));
 INV_X1 _21467_ (.A(_14596_),
    .ZN(_16039_));
 INV_X1 _21468_ (.A(_14564_),
    .ZN(_16040_));
 INV_X1 _21469_ (.A(_14601_),
    .ZN(_16043_));
 INV_X1 _21470_ (.A(_14619_),
    .ZN(_16051_));
 INV_X1 _21471_ (.A(_14627_),
    .ZN(_16055_));
 INV_X1 _21472_ (.A(_14659_),
    .ZN(_16064_));
 INV_X1 _21473_ (.A(_14667_),
    .ZN(_16068_));
 INV_X1 _21474_ (.A(_14681_),
    .ZN(_16072_));
 INV_X1 _21475_ (.A(_14645_),
    .ZN(_16075_));
 INV_X1 _21476_ (.A(_14702_),
    .ZN(_16081_));
 INV_X1 _21477_ (.A(_14710_),
    .ZN(_16082_));
 INV_X1 _21478_ (.A(_14724_),
    .ZN(_16085_));
 INV_X1 _21479_ (.A(_14729_),
    .ZN(_16093_));
 INV_X2 _21480_ (.A(_14745_),
    .ZN(_14747_));
 INV_X1 _21481_ (.A(_14758_),
    .ZN(_16097_));
 INV_X2 _21482_ (.A(_14770_),
    .ZN(_16099_));
 INV_X2 _21483_ (.A(_14799_),
    .ZN(_14802_));
 INV_X1 _21484_ (.A(_14812_),
    .ZN(_16104_));
 INV_X1 _21485_ (.A(_14757_),
    .ZN(_16105_));
 INV_X1 _21486_ (.A(_14744_),
    .ZN(_14813_));
 INV_X1 _21487_ (.A(_14769_),
    .ZN(_16106_));
 INV_X1 _21488_ (.A(_14831_),
    .ZN(_16110_));
 INV_X1 _21489_ (.A(_14867_),
    .ZN(_16114_));
 INV_X1 _21490_ (.A(_14811_),
    .ZN(_16115_));
 INV_X1 _21491_ (.A(_14798_),
    .ZN(_14868_));
 INV_X1 _21492_ (.A(_14825_),
    .ZN(_16116_));
 INV_X1 _21493_ (.A(_14892_),
    .ZN(_14895_));
 INV_X1 _21494_ (.A(_14924_),
    .ZN(_16123_));
 INV_X1 _21495_ (.A(_14937_),
    .ZN(_16125_));
 INV_X1 _21496_ (.A(_14959_),
    .ZN(_14960_));
 INV_X1 _21497_ (.A(_14991_),
    .ZN(_14993_));
 INV_X1 _21498_ (.A(_14911_),
    .ZN(_14998_));
 INV_X1 _21499_ (.A(_14936_),
    .ZN(_16129_));
 INV_X1 _21500_ (.A(_15058_),
    .ZN(_16135_));
 INV_X1 _21501_ (.A(_14990_),
    .ZN(_16136_));
 INV_X1 _21502_ (.A(_15067_),
    .ZN(_16138_));
 INV_X1 _21503_ (.A(_15115_),
    .ZN(_16142_));
 INV_X1 _21504_ (.A(_15125_),
    .ZN(_16144_));
 INV_X1 _21505_ (.A(_15172_),
    .ZN(_16148_));
 INV_X1 _21506_ (.A(_15114_),
    .ZN(_16149_));
 INV_X1 _21507_ (.A(_15104_),
    .ZN(_15173_));
 INV_X1 _21508_ (.A(_15124_),
    .ZN(_16150_));
 INV_X1 _21509_ (.A(_15229_),
    .ZN(_16154_));
 INV_X1 _21510_ (.A(_15240_),
    .ZN(_16156_));
 INV_X1 _21511_ (.A(_15282_),
    .ZN(_16160_));
 INV_X1 _21512_ (.A(_15293_),
    .ZN(_16162_));
 INV_X1 _21513_ (.A(_15320_),
    .ZN(_15321_));
 INV_X1 _21514_ (.A(_15336_),
    .ZN(_16166_));
 INV_X1 _21515_ (.A(_15271_),
    .ZN(_15337_));
 INV_X1 _21516_ (.A(_15347_),
    .ZN(_16168_));
 INV_X1 _21517_ (.A(_15389_),
    .ZN(_16172_));
 INV_X1 _21518_ (.A(_15400_),
    .ZN(_16174_));
 INV_X1 _21519_ (.A(_15435_),
    .ZN(_16178_));
 INV_X1 _21520_ (.A(_15446_),
    .ZN(_16180_));
 INV_X1 _21521_ (.A(_15434_),
    .ZN(_16184_));
 INV_X1 _21522_ (.A(_15425_),
    .ZN(_15480_));
 INV_X1 _21523_ (.A(_15489_),
    .ZN(_16186_));
 INV_X1 _21524_ (.A(_15522_),
    .ZN(_16190_));
 INV_X1 _21525_ (.A(_15468_),
    .ZN(_15524_));
 INV_X1 _21526_ (.A(_15533_),
    .ZN(_16192_));
 INV_X1 _21527_ (.A(_15561_),
    .ZN(_16196_));
 INV_X1 _21528_ (.A(_15512_),
    .ZN(_15563_));
 INV_X1 _21529_ (.A(_15572_),
    .ZN(_16198_));
 INV_X1 _21530_ (.A(_15598_),
    .ZN(_16202_));
 INV_X1 _21531_ (.A(_15551_),
    .ZN(_15599_));
 INV_X1 _21532_ (.A(_15609_),
    .ZN(_16204_));
 INV_X1 _21533_ (.A(_15637_),
    .ZN(_16208_));
 INV_X1 _21534_ (.A(_15648_),
    .ZN(_16210_));
 INV_X1 _21535_ (.A(_15653_),
    .ZN(_15654_));
 INV_X1 _21536_ (.A(_15623_),
    .ZN(_15664_));
 INV_X1 _21537_ (.A(_15676_),
    .ZN(_16214_));
 INV_X1 _21538_ (.A(_15687_),
    .ZN(_16216_));
 INV_X1 _21539_ (.A(_15691_),
    .ZN(_15692_));
 INV_X1 _21540_ (.A(_15659_),
    .ZN(_15700_));
 INV_X1 _21541_ (.A(_15722_),
    .ZN(_16222_));
 INV_X1 _21542_ (.A(_15733_),
    .ZN(_15734_));
 INV_X1 _21543_ (.A(_15753_),
    .ZN(_16228_));
 INV_X2 _21544_ (.A(_16281_),
    .ZN(_16277_));
 BUF_X4 _21545_ (.A(_03705_),
    .Z(_04302_));
 BUF_X4 _21546_ (.A(_04302_),
    .Z(_16485_));
 BUF_X4 _21547_ (.A(_04100_),
    .Z(_04303_));
 BUF_X4 _21548_ (.A(_04303_),
    .Z(_04304_));
 BUF_X2 _21549_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .Z(_04305_));
 BUF_X4 _21550_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_04306_));
 BUF_X4 _21551_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_04307_));
 BUF_X4 _21552_ (.A(_04307_),
    .Z(_04308_));
 OAI221_X1 _21553_ (.A(_04304_),
    .B1(_04305_),
    .B2(_04306_),
    .C1(_04308_),
    .C2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_04309_));
 NOR2_X1 _21554_ (.A1(_04009_),
    .A2(_04000_),
    .ZN(_04310_));
 OAI21_X1 _21555_ (.A(_03535_),
    .B1(_03996_),
    .B2(_04310_),
    .ZN(_04311_));
 AND3_X1 _21556_ (.A1(_00134_),
    .A2(_04309_),
    .A3(_04311_),
    .ZN(_04312_));
 NAND2_X4 _21557_ (.A1(_00133_),
    .A2(_04312_),
    .ZN(_04313_));
 INV_X2 _21558_ (.A(_04313_),
    .ZN(_16509_));
 XNOR2_X1 _21559_ (.A(_16236_),
    .B(_04180_),
    .ZN(_04314_));
 OAI222_X2 _21560_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .A2(_04198_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .B2(_03504_),
    .C1(_03811_),
    .C2(_04200_),
    .ZN(_04315_));
 MUX2_X1 _21561_ (.A(net301),
    .B(_04315_),
    .S(_03497_),
    .Z(_04316_));
 MUX2_X1 _21562_ (.A(_04314_),
    .B(_04316_),
    .S(_04177_),
    .Z(_15772_));
 OR3_X1 _21563_ (.A1(_00217_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04317_));
 OAI21_X2 _21564_ (.A(_04317_),
    .B1(_04178_),
    .B2(_16239_),
    .ZN(_14466_));
 OR3_X1 _21565_ (.A1(_00558_),
    .A2(_04172_),
    .A3(_04174_),
    .ZN(_04318_));
 OAI21_X1 _21566_ (.A(_04318_),
    .B1(_04178_),
    .B2(_16258_),
    .ZN(_15778_));
 CLKBUF_X2 _21567_ (.A(_04171_),
    .Z(_04319_));
 OR3_X1 _21568_ (.A1(_00559_),
    .A2(_04319_),
    .A3(_04174_),
    .ZN(_04320_));
 OAI21_X1 _21569_ (.A(_04320_),
    .B1(_16265_),
    .B2(_04248_),
    .ZN(_15782_));
 CLKBUF_X2 _21570_ (.A(_04173_),
    .Z(_04321_));
 OR3_X1 _21571_ (.A1(_00560_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04322_));
 OAI21_X1 _21572_ (.A(_04322_),
    .B1(_16273_),
    .B2(_04248_),
    .ZN(_15786_));
 OR3_X1 _21573_ (.A1(_00561_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04323_));
 OAI21_X1 _21574_ (.A(_04323_),
    .B1(_16281_),
    .B2(_04248_),
    .ZN(_15790_));
 OR3_X1 _21575_ (.A1(_00562_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04324_));
 OAI21_X1 _21576_ (.A(_04324_),
    .B1(_16289_),
    .B2(_04248_),
    .ZN(_15794_));
 OR3_X1 _21577_ (.A1(_00563_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04325_));
 OAI21_X1 _21578_ (.A(_04325_),
    .B1(_16297_),
    .B2(_04248_),
    .ZN(_15798_));
 XNOR2_X1 _21579_ (.A(_16305_),
    .B(net290),
    .ZN(_04326_));
 OAI222_X2 _21580_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .B2(_03504_),
    .C1(_03872_),
    .C2(_04200_),
    .ZN(_04327_));
 MUX2_X1 _21581_ (.A(_03542_),
    .B(_04327_),
    .S(_03497_),
    .Z(_04328_));
 MUX2_X1 _21582_ (.A(_04326_),
    .B(_04328_),
    .S(_04177_),
    .Z(_15802_));
 OR3_X1 _21583_ (.A1(_00565_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04329_));
 OAI21_X1 _21584_ (.A(_04329_),
    .B1(_16314_),
    .B2(_04248_),
    .ZN(_15806_));
 OR3_X1 _21585_ (.A1(_00566_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04330_));
 OAI21_X1 _21586_ (.A(_04330_),
    .B1(_16321_),
    .B2(_04248_),
    .ZN(_15810_));
 XNOR2_X1 _21587_ (.A(_16330_),
    .B(net290),
    .ZN(_04331_));
 OAI222_X2 _21588_ (.A1(_03498_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .B2(_03504_),
    .C1(_03896_),
    .C2(_03491_),
    .ZN(_04332_));
 NOR2_X1 _21589_ (.A1(_03495_),
    .A2(_04332_),
    .ZN(_04333_));
 AOI21_X1 _21590_ (.A(_04333_),
    .B1(_03495_),
    .B2(_11769_),
    .ZN(_04334_));
 MUX2_X1 _21591_ (.A(_04331_),
    .B(_04334_),
    .S(_04177_),
    .Z(_15814_));
 XNOR2_X1 _21592_ (.A(_04196_),
    .B(_16338_),
    .ZN(_04335_));
 OAI222_X2 _21593_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .B2(_04199_),
    .C1(_03905_),
    .C2(_04200_),
    .ZN(_04336_));
 NAND2_X1 _21594_ (.A1(_04193_),
    .A2(_04336_),
    .ZN(_04337_));
 OAI21_X1 _21595_ (.A(_04337_),
    .B1(_04267_),
    .B2(_12420_),
    .ZN(_04338_));
 MUX2_X1 _21596_ (.A(_04335_),
    .B(_04338_),
    .S(_04177_),
    .Z(_15818_));
 OR3_X1 _21597_ (.A1(_04163_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04339_));
 BUF_X2 _21598_ (.A(_04176_),
    .Z(_04340_));
 OAI21_X1 _21599_ (.A(_04339_),
    .B1(_16342_),
    .B2(_04340_),
    .ZN(_15822_));
 OR3_X1 _21600_ (.A1(_00630_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04341_));
 OAI21_X1 _21601_ (.A(_04341_),
    .B1(_16350_),
    .B2(_04340_),
    .ZN(_15826_));
 OR3_X1 _21602_ (.A1(_00661_),
    .A2(_04319_),
    .A3(_04321_),
    .ZN(_04342_));
 OAI21_X1 _21603_ (.A(_04342_),
    .B1(_16358_),
    .B2(_04340_),
    .ZN(_15830_));
 XNOR2_X1 _21604_ (.A(_04196_),
    .B(_16370_),
    .ZN(_04343_));
 MUX2_X2 _21605_ (.A(_12771_),
    .B(_12789_),
    .S(_10983_),
    .Z(_04344_));
 OAI222_X2 _21606_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .B2(_04199_),
    .C1(_04344_),
    .C2(_04200_),
    .ZN(_04345_));
 NAND2_X1 _21607_ (.A1(_04193_),
    .A2(_04345_),
    .ZN(_04346_));
 OAI21_X1 _21608_ (.A(_04346_),
    .B1(_04190_),
    .B2(net282),
    .ZN(_04347_));
 MUX2_X1 _21609_ (.A(_04343_),
    .B(_04347_),
    .S(_04177_),
    .Z(_15834_));
 CLKBUF_X2 _21610_ (.A(_04171_),
    .Z(_04348_));
 OR3_X1 _21611_ (.A1(_03940_),
    .A2(_04348_),
    .A3(_04321_),
    .ZN(_04349_));
 OAI21_X1 _21612_ (.A(_04349_),
    .B1(_16377_),
    .B2(_04340_),
    .ZN(_15838_));
 CLKBUF_X2 _21613_ (.A(_04173_),
    .Z(_04350_));
 OR3_X1 _21614_ (.A1(_03944_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04351_));
 OAI21_X1 _21615_ (.A(_04351_),
    .B1(_16385_),
    .B2(_04340_),
    .ZN(_15842_));
 OR3_X1 _21616_ (.A1(_03946_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04352_));
 OAI21_X1 _21617_ (.A(_04352_),
    .B1(_16393_),
    .B2(_04340_),
    .ZN(_15846_));
 XNOR2_X1 _21618_ (.A(_04196_),
    .B(_16397_),
    .ZN(_04353_));
 OAI222_X2 _21619_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .B2(_04199_),
    .C1(_03836_),
    .C2(_04200_),
    .ZN(_04354_));
 NAND2_X1 _21620_ (.A1(_04193_),
    .A2(_04354_),
    .ZN(_04355_));
 OAI21_X1 _21621_ (.A(_04355_),
    .B1(_04190_),
    .B2(net369),
    .ZN(_04356_));
 MUX2_X1 _21622_ (.A(_04353_),
    .B(_04356_),
    .S(_04177_),
    .Z(_15850_));
 OR3_X1 _21623_ (.A1(_03950_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04357_));
 OAI21_X1 _21624_ (.A(_04357_),
    .B1(_16406_),
    .B2(_04340_),
    .ZN(_15854_));
 OR3_X1 _21625_ (.A1(_00878_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04358_));
 OAI21_X1 _21626_ (.A(_04358_),
    .B1(_16414_),
    .B2(_04340_),
    .ZN(_15858_));
 OR3_X1 _21627_ (.A1(_03955_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04359_));
 OAI21_X1 _21628_ (.A(_04359_),
    .B1(_16425_),
    .B2(_04340_),
    .ZN(_15862_));
 OR3_X1 _21629_ (.A1(_03957_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04360_));
 OAI21_X1 _21630_ (.A(_04360_),
    .B1(_16433_),
    .B2(_04340_),
    .ZN(_15866_));
 OR3_X1 _21631_ (.A1(_03959_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04361_));
 OAI21_X1 _21632_ (.A(_04361_),
    .B1(_16441_),
    .B2(_04179_),
    .ZN(_15870_));
 OR3_X1 _21633_ (.A1(_01002_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04362_));
 OAI21_X1 _21634_ (.A(_04362_),
    .B1(_16449_),
    .B2(_04179_),
    .ZN(_15874_));
 OR3_X1 _21635_ (.A1(_01033_),
    .A2(_04348_),
    .A3(_04350_),
    .ZN(_04363_));
 OAI21_X1 _21636_ (.A(_04363_),
    .B1(_16457_),
    .B2(_04179_),
    .ZN(_15878_));
 OR3_X1 _21637_ (.A1(_03967_),
    .A2(_04171_),
    .A3(_04350_),
    .ZN(_04364_));
 OAI21_X1 _21638_ (.A(_04364_),
    .B1(_16465_),
    .B2(_04179_),
    .ZN(_15882_));
 OR3_X1 _21639_ (.A1(_01095_),
    .A2(_04171_),
    .A3(_04173_),
    .ZN(_04365_));
 OAI21_X1 _21640_ (.A(_04365_),
    .B1(_16473_),
    .B2(_04179_),
    .ZN(_15886_));
 XNOR2_X1 _21641_ (.A(_04196_),
    .B(_16477_),
    .ZN(_04366_));
 OAI222_X2 _21642_ (.A1(_04198_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .B2(_04199_),
    .C1(_03922_),
    .C2(_04200_),
    .ZN(_04367_));
 NAND2_X1 _21643_ (.A1(_04193_),
    .A2(_04367_),
    .ZN(_04368_));
 OAI21_X1 _21644_ (.A(_04368_),
    .B1(_04190_),
    .B2(_03372_),
    .ZN(_04369_));
 MUX2_X1 _21645_ (.A(_04366_),
    .B(_04369_),
    .S(_04177_),
    .Z(_15890_));
 INV_X1 _21646_ (.A(_15928_),
    .ZN(_15925_));
 INV_X1 _21647_ (.A(_14477_),
    .ZN(_15960_));
 INV_X1 _21648_ (.A(_14471_),
    .ZN(_15959_));
 INV_X1 _21649_ (.A(_14482_),
    .ZN(_15972_));
 INV_X1 _21650_ (.A(_14476_),
    .ZN(_15971_));
 INV_X1 _21651_ (.A(_14492_),
    .ZN(_14495_));
 INV_X1 _21652_ (.A(_14481_),
    .ZN(_14493_));
 INV_X1 _21653_ (.A(_14515_),
    .ZN(_15994_));
 INV_X1 _21654_ (.A(_14501_),
    .ZN(_14523_));
 INV_X1 _21655_ (.A(_14538_),
    .ZN(_16011_));
 INV_X1 _21656_ (.A(_14514_),
    .ZN(_16010_));
 INV_X1 _21657_ (.A(_14519_),
    .ZN(_16019_));
 INV_X1 _21658_ (.A(_14548_),
    .ZN(_14555_));
 INV_X1 _21659_ (.A(_14537_),
    .ZN(_16025_));
 INV_X1 _21660_ (.A(_14570_),
    .ZN(_16028_));
 INV_X1 _21661_ (.A(_14542_),
    .ZN(_16031_));
 INV_X1 _21662_ (.A(_14588_),
    .ZN(_16034_));
 INV_X1 _21663_ (.A(_14569_),
    .ZN(_14603_));
 INV_X1 _21664_ (.A(_14574_),
    .ZN(_16044_));
 INV_X1 _21665_ (.A(_14587_),
    .ZN(_16052_));
 INV_X1 _21666_ (.A(_14595_),
    .ZN(_16056_));
 INV_X1 _21667_ (.A(_14632_),
    .ZN(_14635_));
 INV_X1 _21668_ (.A(_14600_),
    .ZN(_14639_));
 INV_X1 _21669_ (.A(_14646_),
    .ZN(_16061_));
 INV_X1 _21670_ (.A(_14618_),
    .ZN(_16065_));
 INV_X1 _21671_ (.A(_14626_),
    .ZN(_16069_));
 INV_X1 _21672_ (.A(_14672_),
    .ZN(_14675_));
 INV_X1 _21673_ (.A(_14686_),
    .ZN(_16076_));
 INV_X1 _21674_ (.A(_14666_),
    .ZN(_16083_));
 INV_X1 _21675_ (.A(_14715_),
    .ZN(_14718_));
 INV_X1 _21676_ (.A(_14680_),
    .ZN(_16086_));
 INV_X1 _21677_ (.A(_14685_),
    .ZN(_16094_));
 INV_X1 _21678_ (.A(_14709_),
    .ZN(_16098_));
 INV_X1 _21679_ (.A(_14701_),
    .ZN(_14760_));
 INV_X1 _21680_ (.A(_14723_),
    .ZN(_16100_));
 INV_X1 _21681_ (.A(_14783_),
    .ZN(_16103_));
 INV_X2 _21682_ (.A(_14826_),
    .ZN(_16107_));
 INV_X1 _21683_ (.A(_14839_),
    .ZN(_16113_));
 INV_X2 _21684_ (.A(_14854_),
    .ZN(_14856_));
 INV_X2 _21685_ (.A(_14880_),
    .ZN(_16117_));
 INV_X1 _21686_ (.A(_14912_),
    .ZN(_14913_));
 INV_X1 _21687_ (.A(_14866_),
    .ZN(_16124_));
 INV_X1 _21688_ (.A(_14853_),
    .ZN(_14926_));
 INV_X1 _21689_ (.A(_14879_),
    .ZN(_16126_));
 INV_X1 _21690_ (.A(_14942_),
    .ZN(_14949_));
 INV_X1 _21691_ (.A(_14923_),
    .ZN(_14994_));
 INV_X1 _21692_ (.A(_15007_),
    .ZN(_16130_));
 INV_X1 _21693_ (.A(_15006_),
    .ZN(_16139_));
 INV_X1 _21694_ (.A(_15057_),
    .ZN(_16143_));
 INV_X1 _21695_ (.A(_15045_),
    .ZN(_15117_));
 INV_X1 _21696_ (.A(_15066_),
    .ZN(_16145_));
 INV_X1 _21697_ (.A(_15183_),
    .ZN(_16151_));
 INV_X1 _21698_ (.A(_15171_),
    .ZN(_16155_));
 INV_X1 _21699_ (.A(_15161_),
    .ZN(_15232_));
 INV_X1 _21700_ (.A(_15182_),
    .ZN(_16157_));
 INV_X1 _21701_ (.A(_15228_),
    .ZN(_16161_));
 INV_X1 _21702_ (.A(_15219_),
    .ZN(_15284_));
 INV_X1 _21703_ (.A(_15239_),
    .ZN(_16163_));
 INV_X1 _21704_ (.A(_15267_),
    .ZN(_15322_));
 INV_X1 _21705_ (.A(_15281_),
    .ZN(_16167_));
 INV_X1 _21706_ (.A(_15292_),
    .ZN(_16169_));
 INV_X1 _21707_ (.A(_15335_),
    .ZN(_16173_));
 INV_X1 _21708_ (.A(_15326_),
    .ZN(_15391_));
 INV_X1 _21709_ (.A(_15346_),
    .ZN(_16175_));
 INV_X1 _21710_ (.A(_15388_),
    .ZN(_16179_));
 INV_X1 _21711_ (.A(_15379_),
    .ZN(_15437_));
 INV_X1 _21712_ (.A(_15399_),
    .ZN(_16181_));
 INV_X1 _21713_ (.A(_15478_),
    .ZN(_16185_));
 INV_X1 _21714_ (.A(_15445_),
    .ZN(_16187_));
 INV_X1 _21715_ (.A(_15477_),
    .ZN(_16191_));
 INV_X1 _21716_ (.A(_15488_),
    .ZN(_16193_));
 INV_X1 _21717_ (.A(_15521_),
    .ZN(_16197_));
 INV_X1 _21718_ (.A(_15532_),
    .ZN(_16199_));
 INV_X1 _21719_ (.A(_15560_),
    .ZN(_16203_));
 INV_X1 _21720_ (.A(_15571_),
    .ZN(_16205_));
 INV_X1 _21721_ (.A(_15597_),
    .ZN(_16209_));
 INV_X1 _21722_ (.A(_15588_),
    .ZN(_15639_));
 INV_X1 _21723_ (.A(_15608_),
    .ZN(_16211_));
 INV_X1 _21724_ (.A(_15613_),
    .ZN(_15655_));
 INV_X1 _21725_ (.A(_15636_),
    .ZN(_16215_));
 INV_X1 _21726_ (.A(_15627_),
    .ZN(_15678_));
 INV_X1 _21727_ (.A(_15647_),
    .ZN(_16217_));
 INV_X1 _21728_ (.A(_15652_),
    .ZN(_15693_));
 INV_X1 _21729_ (.A(_15712_),
    .ZN(_16221_));
 INV_X1 _21730_ (.A(_15675_),
    .ZN(_16220_));
 INV_X1 _21731_ (.A(_15686_),
    .ZN(_16223_));
 INV_X1 _21732_ (.A(_15690_),
    .ZN(_15727_));
 INV_X1 _21733_ (.A(_15698_),
    .ZN(_15735_));
 INV_X1 _21734_ (.A(_15711_),
    .ZN(_16226_));
 INV_X1 _21735_ (.A(_15721_),
    .ZN(_16229_));
 INV_X1 _21736_ (.A(_16298_),
    .ZN(_16294_));
 INV_X1 _21737_ (.A(_15988_),
    .ZN(_14499_));
 INV_X1 _21738_ (.A(_16000_),
    .ZN(_14516_));
 INV_X1 _21739_ (.A(_16017_),
    .ZN(_14540_));
 INV_X1 _21740_ (.A(_16027_),
    .ZN(_14566_));
 INV_X1 _21741_ (.A(_16029_),
    .ZN(_14571_));
 INV_X1 _21742_ (.A(_16042_),
    .ZN(_14599_));
 INV_X1 _21743_ (.A(_16058_),
    .ZN(_14629_));
 INV_X1 _21744_ (.A(_16071_),
    .ZN(_14669_));
 INV_X1 _21745_ (.A(_16084_),
    .ZN(_14712_));
 INV_X1 _21746_ (.A(_16137_),
    .ZN(_15059_));
 INV_X1 _21747_ (.A(_16062_),
    .ZN(_14700_));
 INV_X1 _21748_ (.A(_16077_),
    .ZN(_14743_));
 INV_X1 _21749_ (.A(_16091_),
    .ZN(_14781_));
 INV_X1 _21750_ (.A(_16095_),
    .ZN(_14797_));
 NOR2_X4 _21751_ (.A1(_04000_),
    .A2(_03996_),
    .ZN(_04370_));
 CLKBUF_X3 _21752_ (.A(_04370_),
    .Z(_04371_));
 NAND2_X1 _21753_ (.A1(net2),
    .A2(_04371_),
    .ZN(_04372_));
 NOR2_X4 _21754_ (.A1(_03591_),
    .A2(_16330_),
    .ZN(_04373_));
 NAND2_X1 _21755_ (.A1(_15909_),
    .A2(_03587_),
    .ZN(_04374_));
 NOR2_X1 _21756_ (.A1(_11489_),
    .A2(_03556_),
    .ZN(_04375_));
 AOI21_X1 _21757_ (.A(_03591_),
    .B1(_11478_),
    .B2(_16282_),
    .ZN(_04376_));
 NAND3_X1 _21758_ (.A1(_03636_),
    .A2(_11478_),
    .A3(_16282_),
    .ZN(_04377_));
 OAI221_X2 _21759_ (.A(_04374_),
    .B1(_04375_),
    .B2(_04376_),
    .C1(_04377_),
    .C2(_11491_),
    .ZN(_04378_));
 NAND3_X4 _21760_ (.A1(_04373_),
    .A2(_04378_),
    .A3(_03584_),
    .ZN(_04379_));
 BUF_X4 _21761_ (.A(_04379_),
    .Z(_04380_));
 BUF_X8 _21762_ (.A(_04380_),
    .Z(_04381_));
 BUF_X2 _21763_ (.A(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .Z(_04382_));
 BUF_X4 _21764_ (.A(_03592_),
    .Z(_04383_));
 NAND2_X1 _21765_ (.A1(_04383_),
    .A2(_03557_),
    .ZN(_04384_));
 NOR2_X1 _21766_ (.A1(_03552_),
    .A2(_03633_),
    .ZN(_04385_));
 NAND2_X1 _21767_ (.A1(_11492_),
    .A2(_04385_),
    .ZN(_04386_));
 AOI21_X4 _21768_ (.A(_15910_),
    .B1(_04384_),
    .B2(_04386_),
    .ZN(_04387_));
 BUF_X8 _21769_ (.A(_04387_),
    .Z(_04388_));
 BUF_X8 _21770_ (.A(_04388_),
    .Z(_04389_));
 NAND2_X4 _21771_ (.A1(_03554_),
    .A2(_11492_),
    .ZN(_04390_));
 NOR2_X4 _21772_ (.A1(_15909_),
    .A2(_04390_),
    .ZN(_04391_));
 BUF_X8 _21773_ (.A(_04391_),
    .Z(_04392_));
 BUF_X8 _21774_ (.A(_04392_),
    .Z(_04393_));
 BUF_X2 _21775_ (.A(\cs_registers_i.mhpmcounter[2][43] ),
    .Z(_04394_));
 AOI22_X4 _21776_ (.A1(_04382_),
    .A2(_04389_),
    .B1(_04393_),
    .B2(_04394_),
    .ZN(_04395_));
 BUF_X2 _21777_ (.A(\cs_registers_i.mhpmcounter[2][11] ),
    .Z(_04396_));
 AOI22_X4 _21778_ (.A1(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .A2(_04389_),
    .B1(_04393_),
    .B2(_04396_),
    .ZN(_04397_));
 NOR2_X4 _21779_ (.A1(_16286_),
    .A2(_16294_),
    .ZN(_04398_));
 AND4_X2 _21780_ (.A1(_16282_),
    .A2(_04373_),
    .A3(_04398_),
    .A4(_03607_),
    .ZN(_04399_));
 AOI21_X4 _21781_ (.A(_03589_),
    .B1(_11478_),
    .B2(_11491_),
    .ZN(_04400_));
 OAI21_X4 _21782_ (.A(_04399_),
    .B1(_04400_),
    .B2(_03578_),
    .ZN(_04401_));
 BUF_X8 _21783_ (.A(_04401_),
    .Z(_04402_));
 OAI22_X4 _21784_ (.A1(_04381_),
    .A2(_04395_),
    .B1(_04397_),
    .B2(_04402_),
    .ZN(_04403_));
 OR4_X4 _21785_ (.A1(_11478_),
    .A2(_16326_),
    .A3(_03560_),
    .A4(_03561_),
    .ZN(_04404_));
 NOR3_X4 _21786_ (.A1(_04383_),
    .A2(_03546_),
    .A3(_04404_),
    .ZN(_04405_));
 AND2_X1 _21787_ (.A1(_03636_),
    .A2(_04405_),
    .ZN(_04406_));
 BUF_X4 _21788_ (.A(_04406_),
    .Z(_04407_));
 BUF_X4 _21789_ (.A(_04407_),
    .Z(_04408_));
 BUF_X4 _21790_ (.A(_03553_),
    .Z(_04409_));
 NAND3_X4 _21791_ (.A1(_11328_),
    .A2(_16309_),
    .A3(net11),
    .ZN(_04410_));
 OR3_X4 _21792_ (.A1(_16270_),
    .A2(_16278_),
    .A3(_04410_),
    .ZN(_04411_));
 NOR4_X4 _21793_ (.A1(_04409_),
    .A2(_04383_),
    .A3(_04411_),
    .A4(_03621_),
    .ZN(_04412_));
 BUF_X4 _21794_ (.A(_04412_),
    .Z(_04413_));
 BUF_X4 _21795_ (.A(_04413_),
    .Z(_04414_));
 AND2_X2 _21796_ (.A1(_03554_),
    .A2(_04405_),
    .ZN(_04415_));
 BUF_X4 _21797_ (.A(_04415_),
    .Z(_04416_));
 BUF_X4 _21798_ (.A(_04416_),
    .Z(_04417_));
 AOI222_X2 _21799_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(_04408_),
    .B1(_04414_),
    .B2(\cs_registers_i.mtval_q[11] ),
    .C1(_04417_),
    .C2(\cs_registers_i.dscratch0_q[11] ),
    .ZN(_04418_));
 OR2_X1 _21800_ (.A1(_04411_),
    .A2(_03621_),
    .ZN(_04419_));
 BUF_X4 _21801_ (.A(_04419_),
    .Z(_04420_));
 NAND2_X4 _21802_ (.A1(_03636_),
    .A2(_11492_),
    .ZN(_04421_));
 NOR2_X4 _21803_ (.A1(_04420_),
    .A2(_04421_),
    .ZN(_04422_));
 BUF_X4 _21804_ (.A(_04422_),
    .Z(_04423_));
 BUF_X4 _21805_ (.A(_04423_),
    .Z(_04424_));
 AND2_X2 _21806_ (.A1(_03552_),
    .A2(_04405_),
    .ZN(_04425_));
 BUF_X4 _21807_ (.A(_04425_),
    .Z(_04426_));
 BUF_X4 _21808_ (.A(_04426_),
    .Z(_04427_));
 AOI22_X2 _21809_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_04424_),
    .B1(_04427_),
    .B2(\cs_registers_i.dscratch1_q[11] ),
    .ZN(_04428_));
 OR2_X4 _21810_ (.A1(_03576_),
    .A2(_03640_),
    .ZN(_04429_));
 NOR2_X4 _21811_ (.A1(_04429_),
    .A2(_04420_),
    .ZN(_04430_));
 BUF_X4 _21812_ (.A(_04430_),
    .Z(_04431_));
 AND2_X1 _21813_ (.A1(_11490_),
    .A2(_04405_),
    .ZN(_04432_));
 BUF_X4 _21814_ (.A(_04432_),
    .Z(_04433_));
 AOI22_X2 _21815_ (.A1(net125),
    .A2(_04431_),
    .B1(_04433_),
    .B2(\cs_registers_i.dcsr_q[11] ),
    .ZN(_04434_));
 NAND3_X2 _21816_ (.A1(_04418_),
    .A2(_04428_),
    .A3(_04434_),
    .ZN(_04435_));
 AND3_X1 _21817_ (.A1(_11328_),
    .A2(_16309_),
    .A3(net14),
    .ZN(_04436_));
 CLKBUF_X3 _21818_ (.A(_04436_),
    .Z(_04437_));
 INV_X1 _21819_ (.A(_04437_),
    .ZN(_04438_));
 NOR4_X4 _21820_ (.A1(_03591_),
    .A2(_11476_),
    .A3(_16278_),
    .A4(_16330_),
    .ZN(_04439_));
 NAND2_X2 _21821_ (.A1(_04398_),
    .A2(_04439_),
    .ZN(_04440_));
 NOR3_X4 _21822_ (.A1(_04438_),
    .A2(_04429_),
    .A3(_04440_),
    .ZN(_04441_));
 BUF_X4 _21823_ (.A(_04441_),
    .Z(_04442_));
 NOR4_X4 _21824_ (.A1(_03576_),
    .A2(_03591_),
    .A3(_11379_),
    .A4(_16262_),
    .ZN(_04443_));
 NAND2_X1 _21825_ (.A1(_11329_),
    .A2(_03566_),
    .ZN(_04444_));
 NOR2_X1 _21826_ (.A1(_04373_),
    .A2(_04411_),
    .ZN(_04445_));
 AND3_X1 _21827_ (.A1(_04443_),
    .A2(_04444_),
    .A3(_04445_),
    .ZN(_04446_));
 BUF_X4 _21828_ (.A(_04446_),
    .Z(_04447_));
 BUF_X4 _21829_ (.A(_04447_),
    .Z(_04448_));
 AOI22_X4 _21830_ (.A1(net63),
    .A2(_04442_),
    .B1(_04448_),
    .B2(\cs_registers_i.mie_q[15] ),
    .ZN(_04449_));
 NOR3_X4 _21831_ (.A1(_16326_),
    .A2(_03566_),
    .A3(_04410_),
    .ZN(_04450_));
 AND2_X2 _21832_ (.A1(_04450_),
    .A2(_03588_),
    .ZN(_04451_));
 NOR2_X2 _21833_ (.A1(_04411_),
    .A2(_03621_),
    .ZN(_04452_));
 AOI22_X1 _21834_ (.A1(\cs_registers_i.mstack_d[0] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(\cs_registers_i.mscratch_q[11] ),
    .ZN(_04453_));
 OAI21_X2 _21835_ (.A(_04449_),
    .B1(_04453_),
    .B2(_11493_),
    .ZN(_04454_));
 NOR4_X4 _21836_ (.A1(_16326_),
    .A2(_03561_),
    .A3(_03566_),
    .A4(_04410_),
    .ZN(_04455_));
 NAND4_X4 _21837_ (.A1(_11490_),
    .A2(_16274_),
    .A3(_11492_),
    .A4(_04455_),
    .ZN(_04456_));
 BUF_X4 _21838_ (.A(_04456_),
    .Z(_04457_));
 NOR4_X4 _21839_ (.A1(_03589_),
    .A2(_03591_),
    .A3(_11379_),
    .A4(_16262_),
    .ZN(_04458_));
 NAND3_X4 _21840_ (.A1(_04450_),
    .A2(_03588_),
    .A3(_04458_),
    .ZN(_04459_));
 CLKBUF_X3 _21841_ (.A(_04459_),
    .Z(_04460_));
 BUF_X4 _21842_ (.A(_04460_),
    .Z(_04461_));
 OAI21_X2 _21843_ (.A(_04457_),
    .B1(_04461_),
    .B2(_00551_),
    .ZN(_04462_));
 NOR4_X4 _21844_ (.A1(_04403_),
    .A2(_04435_),
    .A3(_04454_),
    .A4(_04462_),
    .ZN(_04463_));
 NAND2_X1 _21845_ (.A1(_16329_),
    .A2(_04463_),
    .ZN(_04464_));
 BUF_X1 _21846_ (.A(_15932_),
    .Z(_04465_));
 CLKBUF_X2 _21847_ (.A(_04465_),
    .Z(_04466_));
 CLKBUF_X2 _21848_ (.A(_11772_),
    .Z(_04467_));
 MUX2_X1 _21849_ (.A(_04466_),
    .B(_04467_),
    .S(_16325_),
    .Z(_04468_));
 BUF_X4 _21850_ (.A(_15926_),
    .Z(_04469_));
 BUF_X8 _21851_ (.A(_04469_),
    .Z(_04470_));
 OAI21_X2 _21852_ (.A(_04464_),
    .B1(_04468_),
    .B2(_04470_),
    .ZN(_04471_));
 BUF_X4 _21853_ (.A(_04471_),
    .Z(_04472_));
 NAND2_X1 _21854_ (.A1(_11328_),
    .A2(_03687_),
    .ZN(_04473_));
 NOR2_X1 _21855_ (.A1(_03646_),
    .A2(_04473_),
    .ZN(_04474_));
 NAND2_X1 _21856_ (.A1(_03645_),
    .A2(_04474_),
    .ZN(_04475_));
 NAND4_X4 _21857_ (.A1(_04398_),
    .A2(_04437_),
    .A3(_04443_),
    .A4(_04439_),
    .ZN(_04476_));
 OAI21_X1 _21858_ (.A(_11478_),
    .B1(_16262_),
    .B2(_16253_),
    .ZN(_04477_));
 NAND3_X1 _21859_ (.A1(_03562_),
    .A2(_03607_),
    .A3(_04477_),
    .ZN(_04478_));
 AND3_X1 _21860_ (.A1(_03563_),
    .A2(_04476_),
    .A3(_04478_),
    .ZN(_04479_));
 OR4_X1 _21861_ (.A1(_16270_),
    .A2(_16326_),
    .A3(_03566_),
    .A4(_04410_),
    .ZN(_04480_));
 OAI21_X1 _21862_ (.A(_03627_),
    .B1(_16266_),
    .B2(_03591_),
    .ZN(_04481_));
 NOR3_X2 _21863_ (.A1(_03625_),
    .A2(_04480_),
    .A3(_04481_),
    .ZN(_04482_));
 NOR4_X1 _21864_ (.A1(_04411_),
    .A2(_03619_),
    .A3(_03620_),
    .A4(_03621_),
    .ZN(_04483_));
 NOR4_X2 _21865_ (.A1(_10957_),
    .A2(_03591_),
    .A3(net10),
    .A4(_16298_),
    .ZN(_04484_));
 NAND4_X1 _21866_ (.A1(_16274_),
    .A2(_16282_),
    .A3(_04437_),
    .A4(_04484_),
    .ZN(_04485_));
 NOR4_X1 _21867_ (.A1(_04383_),
    .A2(_16326_),
    .A3(_03596_),
    .A4(_04485_),
    .ZN(_04486_));
 NOR3_X1 _21868_ (.A1(_04482_),
    .A2(_04483_),
    .A3(_04486_),
    .ZN(_04487_));
 AND4_X1 _21869_ (.A1(_04379_),
    .A2(_04401_),
    .A3(_04479_),
    .A4(_04487_),
    .ZN(_04488_));
 NAND2_X2 _21870_ (.A1(_03642_),
    .A2(_04455_),
    .ZN(_04489_));
 AOI211_X2 _21871_ (.A(_03565_),
    .B(_04475_),
    .C1(_04488_),
    .C2(_04489_),
    .ZN(_04490_));
 NAND3_X4 _21872_ (.A1(_04451_),
    .A2(_04458_),
    .A3(net12),
    .ZN(_04491_));
 CLKBUF_X3 _21873_ (.A(_04491_),
    .Z(_04492_));
 OAI21_X4 _21874_ (.A(_04491_),
    .B1(_03996_),
    .B2(_04000_),
    .ZN(_04493_));
 CLKBUF_X3 _21875_ (.A(_04493_),
    .Z(_04494_));
 INV_X1 _21876_ (.A(\cs_registers_i.csr_mtvec_o[11] ),
    .ZN(_04495_));
 OAI221_X1 _21877_ (.A(_04372_),
    .B1(_04472_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04495_),
    .ZN(_01186_));
 NAND2_X1 _21878_ (.A1(net3),
    .A2(_04371_),
    .ZN(_04496_));
 MUX2_X1 _21879_ (.A(_04466_),
    .B(_04467_),
    .S(_16333_),
    .Z(_04497_));
 BUF_X8 _21880_ (.A(_04381_),
    .Z(_04498_));
 BUF_X8 _21881_ (.A(_04388_),
    .Z(_04499_));
 BUF_X8 _21882_ (.A(_04499_),
    .Z(_04500_));
 BUF_X8 _21883_ (.A(_04392_),
    .Z(_04501_));
 AOI22_X4 _21884_ (.A1(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .A2(_04500_),
    .B1(_04501_),
    .B2(\cs_registers_i.mhpmcounter[2][44] ),
    .ZN(_04502_));
 BUF_X2 _21885_ (.A(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .Z(_04503_));
 BUF_X2 _21886_ (.A(\cs_registers_i.mhpmcounter[2][12] ),
    .Z(_04504_));
 AOI22_X4 _21887_ (.A1(_04503_),
    .A2(_04500_),
    .B1(_04501_),
    .B2(_04504_),
    .ZN(_04505_));
 OAI22_X4 _21888_ (.A1(_04498_),
    .A2(_04502_),
    .B1(_04505_),
    .B2(_04402_),
    .ZN(_04506_));
 NOR2_X2 _21889_ (.A1(_11493_),
    .A2(_04420_),
    .ZN(_04507_));
 BUF_X4 _21890_ (.A(_04507_),
    .Z(_04508_));
 BUF_X4 _21891_ (.A(_04508_),
    .Z(_04509_));
 AOI22_X2 _21892_ (.A1(\cs_registers_i.csr_mepc_o[12] ),
    .A2(_04424_),
    .B1(_04509_),
    .B2(\cs_registers_i.mscratch_q[12] ),
    .ZN(_04510_));
 AND2_X1 _21893_ (.A1(_16274_),
    .A2(_04450_),
    .ZN(_04511_));
 NAND2_X2 _21894_ (.A1(_11379_),
    .A2(_11434_),
    .ZN(_04512_));
 OAI33_X1 _21895_ (.A1(_03589_),
    .A2(_04383_),
    .A3(_16278_),
    .B1(_03561_),
    .B2(_04512_),
    .B3(_03576_),
    .ZN(_04513_));
 NAND2_X2 _21896_ (.A1(_04511_),
    .A2(_04513_),
    .ZN(_04514_));
 INV_X1 _21897_ (.A(\cs_registers_i.mstack_d[1] ),
    .ZN(_04515_));
 OAI33_X1 _21898_ (.A1(_03576_),
    .A2(_04515_),
    .A3(_04383_),
    .B1(_03640_),
    .B2(_03589_),
    .B3(_00550_),
    .ZN(_04516_));
 NAND2_X1 _21899_ (.A1(_04451_),
    .A2(_04516_),
    .ZN(_04517_));
 BUF_X4 _21900_ (.A(_04408_),
    .Z(_04518_));
 AOI22_X2 _21901_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(_04518_),
    .B1(_04417_),
    .B2(\cs_registers_i.dscratch0_q[12] ),
    .ZN(_04519_));
 NAND4_X1 _21902_ (.A1(_04510_),
    .A2(_04514_),
    .A3(_04517_),
    .A4(_04519_),
    .ZN(_04520_));
 INV_X1 _21903_ (.A(_00549_),
    .ZN(_04521_));
 AOI222_X2 _21904_ (.A1(net64),
    .A2(_04442_),
    .B1(_04414_),
    .B2(\cs_registers_i.mtval_q[12] ),
    .C1(_04521_),
    .C2(_04433_),
    .ZN(_04522_));
 BUF_X4 _21905_ (.A(_04426_),
    .Z(_04523_));
 NAND2_X1 _21906_ (.A1(\cs_registers_i.dscratch1_q[12] ),
    .A2(_04523_),
    .ZN(_04524_));
 NAND2_X1 _21907_ (.A1(_04522_),
    .A2(_04524_),
    .ZN(_04525_));
 OR3_X4 _21908_ (.A1(_04506_),
    .A2(_04520_),
    .A3(_04525_),
    .ZN(_04526_));
 OAI22_X4 _21909_ (.A1(_04470_),
    .A2(_04497_),
    .B1(_04526_),
    .B2(_16333_),
    .ZN(_04527_));
 BUF_X4 _21910_ (.A(_04527_),
    .Z(_04528_));
 INV_X1 _21911_ (.A(\cs_registers_i.csr_mtvec_o[12] ),
    .ZN(_04529_));
 OAI221_X1 _21912_ (.A(_04496_),
    .B1(_04528_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04529_),
    .ZN(_01187_));
 INV_X1 _21913_ (.A(_03565_),
    .ZN(_04530_));
 AND2_X2 _21914_ (.A1(_03645_),
    .A2(_04474_),
    .ZN(_04531_));
 AND3_X1 _21915_ (.A1(_11492_),
    .A2(_03547_),
    .A3(_03562_),
    .ZN(_04532_));
 AND4_X1 _21916_ (.A1(_04398_),
    .A2(_04437_),
    .A3(_04443_),
    .A4(_04439_),
    .ZN(_04533_));
 AND3_X1 _21917_ (.A1(_03562_),
    .A2(_03607_),
    .A3(_04477_),
    .ZN(_04534_));
 NOR3_X2 _21918_ (.A1(_04532_),
    .A2(_04533_),
    .A3(_04534_),
    .ZN(_04535_));
 NOR2_X1 _21919_ (.A1(_03619_),
    .A2(_03620_),
    .ZN(_04536_));
 NAND4_X1 _21920_ (.A1(_11478_),
    .A2(_16282_),
    .A3(_04437_),
    .A4(_04484_),
    .ZN(_04537_));
 NOR3_X1 _21921_ (.A1(_16326_),
    .A2(_03596_),
    .A3(_04537_),
    .ZN(_04538_));
 AOI221_X2 _21922_ (.A(_04482_),
    .B1(_04452_),
    .B2(_04536_),
    .C1(_04538_),
    .C2(_11492_),
    .ZN(_04539_));
 NAND4_X4 _21923_ (.A1(_04379_),
    .A2(_04401_),
    .A3(_04535_),
    .A4(_04539_),
    .ZN(_04540_));
 AND2_X1 _21924_ (.A1(_03642_),
    .A2(_04455_),
    .ZN(_04541_));
 OAI211_X4 _21925_ (.A(_04530_),
    .B(_04531_),
    .C1(_04540_),
    .C2(_04541_),
    .ZN(_04542_));
 MUX2_X1 _21926_ (.A(_04466_),
    .B(_04467_),
    .S(_16346_),
    .Z(_04543_));
 AND3_X2 _21927_ (.A1(_16274_),
    .A2(_15908_),
    .A3(_04455_),
    .ZN(_04544_));
 BUF_X4 _21928_ (.A(_04544_),
    .Z(_04545_));
 BUF_X2 _21929_ (.A(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .Z(_04546_));
 BUF_X2 _21930_ (.A(\cs_registers_i.mhpmcounter[2][45] ),
    .Z(_04547_));
 AOI22_X2 _21931_ (.A1(_04546_),
    .A2(_04388_),
    .B1(_04391_),
    .B2(_04547_),
    .ZN(_04548_));
 CLKBUF_X2 _21932_ (.A(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .Z(_04549_));
 BUF_X2 _21933_ (.A(\cs_registers_i.mhpmcounter[2][13] ),
    .Z(_04550_));
 AOI22_X2 _21934_ (.A1(_04549_),
    .A2(_04388_),
    .B1(_04391_),
    .B2(_04550_),
    .ZN(_04551_));
 OAI22_X2 _21935_ (.A1(_04380_),
    .A2(_04548_),
    .B1(_04551_),
    .B2(_04401_),
    .ZN(_04552_));
 NAND2_X1 _21936_ (.A1(\cs_registers_i.mtval_q[13] ),
    .A2(_04414_),
    .ZN(_04553_));
 NOR2_X1 _21937_ (.A1(_01172_),
    .A2(_04459_),
    .ZN(_04554_));
 AOI221_X2 _21938_ (.A(_04554_),
    .B1(_04441_),
    .B2(net65),
    .C1(\cs_registers_i.dscratch1_q[13] ),
    .C2(_04425_),
    .ZN(_04555_));
 AOI22_X2 _21939_ (.A1(\cs_registers_i.dscratch0_q[13] ),
    .A2(_04416_),
    .B1(_04433_),
    .B2(\cs_registers_i.dcsr_q[13] ),
    .ZN(_04556_));
 AOI22_X2 _21940_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_04407_),
    .B1(_04423_),
    .B2(\cs_registers_i.csr_mepc_o[13] ),
    .ZN(_04557_));
 NAND4_X2 _21941_ (.A1(_04553_),
    .A2(_04555_),
    .A3(_04556_),
    .A4(_04557_),
    .ZN(_04558_));
 BUF_X4 _21942_ (.A(_04508_),
    .Z(_04559_));
 AND2_X1 _21943_ (.A1(\cs_registers_i.mscratch_q[13] ),
    .A2(_04559_),
    .ZN(_04560_));
 OR4_X4 _21944_ (.A1(_04545_),
    .A2(_04552_),
    .A3(_04558_),
    .A4(_04560_),
    .ZN(_04561_));
 OAI22_X4 _21945_ (.A1(_04470_),
    .A2(_04543_),
    .B1(_04561_),
    .B2(_16346_),
    .ZN(_04562_));
 INV_X1 _21946_ (.A(_04562_),
    .ZN(_04563_));
 OAI33_X1 _21947_ (.A1(_04000_),
    .A2(net4),
    .A3(_03996_),
    .B1(_04461_),
    .B2(_04542_),
    .B3(_04563_),
    .ZN(_04564_));
 NOR2_X1 _21948_ (.A1(\cs_registers_i.csr_mtvec_o[13] ),
    .A2(_04493_),
    .ZN(_04565_));
 NOR2_X1 _21949_ (.A1(_04564_),
    .A2(_04565_),
    .ZN(_01188_));
 NAND2_X1 _21950_ (.A1(net5),
    .A2(_04371_),
    .ZN(_04566_));
 MUX2_X1 _21951_ (.A(_04466_),
    .B(_04467_),
    .S(_16354_),
    .Z(_04567_));
 OR3_X4 _21952_ (.A1(_16274_),
    .A2(_03546_),
    .A3(_03610_),
    .ZN(_04568_));
 NOR2_X2 _21953_ (.A1(_04421_),
    .A2(_04568_),
    .ZN(_04569_));
 NOR4_X4 _21954_ (.A1(_04409_),
    .A2(_03595_),
    .A3(_03621_),
    .A4(_03622_),
    .ZN(_04570_));
 NOR3_X4 _21955_ (.A1(_03621_),
    .A2(_03622_),
    .A3(_04421_),
    .ZN(_04571_));
 AOI222_X2 _21956_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(_04569_),
    .B1(_04570_),
    .B2(\cs_registers_i.mtval_q[14] ),
    .C1(_04571_),
    .C2(\cs_registers_i.csr_mepc_o[14] ),
    .ZN(_04572_));
 NOR4_X4 _21957_ (.A1(_16270_),
    .A2(_11493_),
    .A3(_03609_),
    .A4(_03626_),
    .ZN(_04573_));
 NOR3_X4 _21958_ (.A1(_03601_),
    .A2(_03604_),
    .A3(_03605_),
    .ZN(_04574_));
 NOR3_X4 _21959_ (.A1(_11493_),
    .A2(_03621_),
    .A3(_03622_),
    .ZN(_04575_));
 AOI221_X2 _21960_ (.A(_04573_),
    .B1(_04574_),
    .B2(net66),
    .C1(\cs_registers_i.mscratch_q[14] ),
    .C2(_04575_),
    .ZN(_04576_));
 NOR2_X2 _21961_ (.A1(_03580_),
    .A2(_03603_),
    .ZN(_04577_));
 AOI21_X1 _21962_ (.A(_03580_),
    .B1(_16282_),
    .B2(_16274_),
    .ZN(_04578_));
 NOR2_X1 _21963_ (.A1(_03626_),
    .A2(_04578_),
    .ZN(_04579_));
 NAND4_X2 _21964_ (.A1(_03636_),
    .A2(_16266_),
    .A3(_04577_),
    .A4(_04579_),
    .ZN(_04580_));
 OR2_X1 _21965_ (.A1(_01173_),
    .A2(_04580_),
    .ZN(_04581_));
 NAND3_X1 _21966_ (.A1(_04572_),
    .A2(_04576_),
    .A3(_04581_),
    .ZN(_04582_));
 NOR2_X4 _21967_ (.A1(_04390_),
    .A2(_04568_),
    .ZN(_04583_));
 NOR3_X4 _21968_ (.A1(_04409_),
    .A2(_03595_),
    .A3(_04568_),
    .ZN(_04584_));
 AOI221_X2 _21969_ (.A(_04582_),
    .B1(_04583_),
    .B2(\cs_registers_i.dscratch0_q[14] ),
    .C1(\cs_registers_i.dscratch1_q[14] ),
    .C2(_04584_),
    .ZN(_04585_));
 BUF_X2 _21970_ (.A(\cs_registers_i.mhpmcounter[2][14] ),
    .Z(_04586_));
 AOI22_X2 _21971_ (.A1(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .A2(_04500_),
    .B1(_04501_),
    .B2(_04586_),
    .ZN(_04587_));
 OR2_X4 _21972_ (.A1(_03593_),
    .A2(_03586_),
    .ZN(_04588_));
 BUF_X4 _21973_ (.A(_04388_),
    .Z(_04589_));
 BUF_X8 _21974_ (.A(_04589_),
    .Z(_04590_));
 BUF_X4 _21975_ (.A(_04391_),
    .Z(_04591_));
 BUF_X8 _21976_ (.A(_04591_),
    .Z(_04592_));
 BUF_X2 _21977_ (.A(\cs_registers_i.mhpmcounter[2][46] ),
    .Z(_04593_));
 AOI22_X2 _21978_ (.A1(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .A2(_04590_),
    .B1(_04592_),
    .B2(_04593_),
    .ZN(_04594_));
 OAI221_X2 _21979_ (.A(_04585_),
    .B1(_04587_),
    .B2(_03583_),
    .C1(_04588_),
    .C2(_04594_),
    .ZN(_04595_));
 OAI22_X4 _21980_ (.A1(_04470_),
    .A2(_04567_),
    .B1(_04595_),
    .B2(_16354_),
    .ZN(_04596_));
 BUF_X4 _21981_ (.A(_04596_),
    .Z(_04597_));
 INV_X1 _21982_ (.A(\cs_registers_i.csr_mtvec_o[14] ),
    .ZN(_04598_));
 OAI221_X1 _21983_ (.A(_04566_),
    .B1(_04597_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04598_),
    .ZN(_01189_));
 NAND2_X1 _21984_ (.A1(net6),
    .A2(_04371_),
    .ZN(_04599_));
 BUF_X8 _21985_ (.A(_04470_),
    .Z(_04600_));
 CLKBUF_X2 _21986_ (.A(_04466_),
    .Z(_04601_));
 MUX2_X1 _21987_ (.A(_04601_),
    .B(_15928_),
    .S(_16362_),
    .Z(_04602_));
 CLKBUF_X3 _21988_ (.A(\cs_registers_i.mhpmcounter[2][47] ),
    .Z(_04603_));
 AOI22_X2 _21989_ (.A1(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .A2(_04589_),
    .B1(_04591_),
    .B2(_04603_),
    .ZN(_04604_));
 BUF_X2 _21990_ (.A(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .Z(_04605_));
 BUF_X2 _21991_ (.A(\cs_registers_i.mhpmcounter[2][15] ),
    .Z(_04606_));
 AOI22_X2 _21992_ (.A1(_04605_),
    .A2(_04589_),
    .B1(_04591_),
    .B2(_04606_),
    .ZN(_04607_));
 BUF_X4 _21993_ (.A(_04401_),
    .Z(_04608_));
 OAI22_X2 _21994_ (.A1(_04381_),
    .A2(_04604_),
    .B1(_04607_),
    .B2(_04608_),
    .ZN(_04609_));
 INV_X1 _21995_ (.A(net67),
    .ZN(_04610_));
 OAI22_X2 _21996_ (.A1(_04610_),
    .A2(_04476_),
    .B1(_04459_),
    .B2(_01174_),
    .ZN(_04611_));
 AOI221_X1 _21997_ (.A(_04611_),
    .B1(_04413_),
    .B2(\cs_registers_i.mtval_q[15] ),
    .C1(\cs_registers_i.dscratch1_q[15] ),
    .C2(_04426_),
    .ZN(_04612_));
 INV_X1 _21998_ (.A(_00556_),
    .ZN(_04613_));
 AOI22_X1 _21999_ (.A1(\cs_registers_i.dscratch0_q[15] ),
    .A2(_04417_),
    .B1(_04433_),
    .B2(_04613_),
    .ZN(_04614_));
 BUF_X4 _22000_ (.A(_04423_),
    .Z(_04615_));
 AOI22_X2 _22001_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(_04408_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[15] ),
    .ZN(_04616_));
 NAND3_X1 _22002_ (.A1(_04612_),
    .A2(_04614_),
    .A3(_04616_),
    .ZN(_04617_));
 AND2_X1 _22003_ (.A1(\cs_registers_i.mscratch_q[15] ),
    .A2(_04509_),
    .ZN(_04618_));
 OR4_X4 _22004_ (.A1(_04545_),
    .A2(_04609_),
    .A3(_04617_),
    .A4(_04618_),
    .ZN(_04619_));
 OAI22_X4 _22005_ (.A1(_04600_),
    .A2(_04602_),
    .B1(_04619_),
    .B2(_16362_),
    .ZN(_04620_));
 INV_X1 _22006_ (.A(\cs_registers_i.csr_mtvec_o[15] ),
    .ZN(_04621_));
 OAI221_X1 _22007_ (.A(_04599_),
    .B1(_04620_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04621_),
    .ZN(_01190_));
 NAND2_X1 _22008_ (.A1(net15),
    .A2(_04371_),
    .ZN(_04622_));
 CLKBUF_X3 _22009_ (.A(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .Z(_04623_));
 CLKBUF_X3 _22010_ (.A(\cs_registers_i.mhpmcounter[2][48] ),
    .Z(_04624_));
 AOI22_X4 _22011_ (.A1(_04623_),
    .A2(_04590_),
    .B1(_04592_),
    .B2(_04624_),
    .ZN(_04625_));
 BUF_X2 _22012_ (.A(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .Z(_04626_));
 BUF_X2 _22013_ (.A(\cs_registers_i.mhpmcounter[2][16] ),
    .Z(_04627_));
 AOI22_X4 _22014_ (.A1(_04626_),
    .A2(_04590_),
    .B1(_04592_),
    .B2(_04627_),
    .ZN(_04628_));
 BUF_X4 _22015_ (.A(_04608_),
    .Z(_04629_));
 OAI22_X4 _22016_ (.A1(_04498_),
    .A2(_04625_),
    .B1(_04628_),
    .B2(_04629_),
    .ZN(_04630_));
 AOI22_X2 _22017_ (.A1(\cs_registers_i.csr_mepc_o[16] ),
    .A2(_04424_),
    .B1(_04431_),
    .B2(net126),
    .ZN(_04631_));
 BUF_X4 _22018_ (.A(_04417_),
    .Z(_04632_));
 AOI22_X4 _22019_ (.A1(\cs_registers_i.dscratch0_q[16] ),
    .A2(_04632_),
    .B1(_04523_),
    .B2(\cs_registers_i.dscratch1_q[16] ),
    .ZN(_04633_));
 BUF_X4 _22020_ (.A(_04413_),
    .Z(_04634_));
 AOI222_X2 _22021_ (.A1(\cs_registers_i.csr_depc_o[16] ),
    .A2(_04518_),
    .B1(_04634_),
    .B2(\cs_registers_i.mtval_q[16] ),
    .C1(_04559_),
    .C2(\cs_registers_i.mscratch_q[16] ),
    .ZN(_04635_));
 OAI21_X2 _22022_ (.A(_04457_),
    .B1(_04460_),
    .B2(_01175_),
    .ZN(_04636_));
 BUF_X4 _22023_ (.A(_04441_),
    .Z(_04637_));
 AOI221_X2 _22024_ (.A(_04636_),
    .B1(_04637_),
    .B2(net68),
    .C1(\cs_registers_i.mie_q[0] ),
    .C2(_04448_),
    .ZN(_04638_));
 NAND4_X4 _22025_ (.A1(_04631_),
    .A2(_04633_),
    .A3(_04635_),
    .A4(_04638_),
    .ZN(_04639_));
 NOR2_X4 _22026_ (.A1(_04630_),
    .A2(_04639_),
    .ZN(_04640_));
 NAND2_X1 _22027_ (.A1(_16369_),
    .A2(_04640_),
    .ZN(_04641_));
 CLKBUF_X2 _22028_ (.A(_04466_),
    .Z(_04642_));
 CLKBUF_X2 _22029_ (.A(_11772_),
    .Z(_04643_));
 MUX2_X1 _22030_ (.A(_04642_),
    .B(_04643_),
    .S(_16365_),
    .Z(_04644_));
 OAI21_X4 _22031_ (.A(_04641_),
    .B1(_04644_),
    .B2(_04600_),
    .ZN(_04645_));
 INV_X1 _22032_ (.A(\cs_registers_i.csr_mtvec_o[16] ),
    .ZN(_04646_));
 OAI221_X1 _22033_ (.A(_04622_),
    .B1(_04645_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04646_),
    .ZN(_01191_));
 NAND2_X1 _22034_ (.A1(net16),
    .A2(_04371_),
    .ZN(_04647_));
 MUX2_X1 _22035_ (.A(_04601_),
    .B(_15928_),
    .S(_16373_),
    .Z(_04648_));
 AOI22_X1 _22036_ (.A1(\cs_registers_i.csr_mepc_o[17] ),
    .A2(_04615_),
    .B1(_04559_),
    .B2(\cs_registers_i.mscratch_q[17] ),
    .ZN(_04649_));
 NOR2_X1 _22037_ (.A1(_01176_),
    .A2(_04460_),
    .ZN(_04650_));
 AOI21_X1 _22038_ (.A(_04650_),
    .B1(_04448_),
    .B2(\cs_registers_i.mie_q[1] ),
    .ZN(_04651_));
 AOI22_X1 _22039_ (.A1(net69),
    .A2(_04637_),
    .B1(_04430_),
    .B2(net132),
    .ZN(_04652_));
 AOI21_X1 _22040_ (.A(_04544_),
    .B1(_04414_),
    .B2(\cs_registers_i.mtval_q[17] ),
    .ZN(_04653_));
 NAND4_X1 _22041_ (.A1(_04649_),
    .A2(_04651_),
    .A3(_04652_),
    .A4(_04653_),
    .ZN(_04654_));
 AOI22_X1 _22042_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(_04408_),
    .B1(_04417_),
    .B2(\cs_registers_i.dscratch0_q[17] ),
    .ZN(_04655_));
 NAND2_X4 _22043_ (.A1(_04450_),
    .A2(_03588_),
    .ZN(_04656_));
 NOR2_X4 _22044_ (.A1(_11493_),
    .A2(_04656_),
    .ZN(_04657_));
 AOI22_X1 _22045_ (.A1(\cs_registers_i.dscratch1_q[17] ),
    .A2(_04427_),
    .B1(_04657_),
    .B2(\cs_registers_i.mstatus_q[1] ),
    .ZN(_04658_));
 NAND2_X1 _22046_ (.A1(_04655_),
    .A2(_04658_),
    .ZN(_04659_));
 NOR2_X2 _22047_ (.A1(_04654_),
    .A2(_04659_),
    .ZN(_04660_));
 AOI22_X2 _22048_ (.A1(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .A2(_04389_),
    .B1(_04393_),
    .B2(\cs_registers_i.mhpmcounter[2][17] ),
    .ZN(_04661_));
 CLKBUF_X3 _22049_ (.A(\cs_registers_i.mhpmcounter[2][49] ),
    .Z(_04662_));
 AOI22_X2 _22050_ (.A1(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .A2(_04500_),
    .B1(_04501_),
    .B2(_04662_),
    .ZN(_04663_));
 OAI221_X2 _22051_ (.A(_04660_),
    .B1(_04661_),
    .B2(_04402_),
    .C1(_04381_),
    .C2(_04663_),
    .ZN(_04664_));
 OAI22_X4 _22052_ (.A1(_04600_),
    .A2(_04648_),
    .B1(_04664_),
    .B2(_16373_),
    .ZN(_04665_));
 INV_X1 _22053_ (.A(\cs_registers_i.csr_mtvec_o[17] ),
    .ZN(_04666_));
 OAI221_X1 _22054_ (.A(_04647_),
    .B1(_04665_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04666_),
    .ZN(_01192_));
 NAND2_X1 _22055_ (.A1(net17),
    .A2(_04371_),
    .ZN(_04667_));
 BUF_X8 _22056_ (.A(_04469_),
    .Z(_04668_));
 MUX2_X1 _22057_ (.A(_04642_),
    .B(_04643_),
    .S(_16381_),
    .Z(_04669_));
 BUF_X2 _22058_ (.A(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .Z(_04670_));
 BUF_X2 _22059_ (.A(\cs_registers_i.mhpmcounter[2][50] ),
    .Z(_04671_));
 AOI22_X2 _22060_ (.A1(_04670_),
    .A2(_04589_),
    .B1(_04591_),
    .B2(_04671_),
    .ZN(_04672_));
 BUF_X2 _22061_ (.A(\cs_registers_i.mhpmcounter[2][18] ),
    .Z(_04673_));
 AOI22_X2 _22062_ (.A1(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .A2(_04589_),
    .B1(_04591_),
    .B2(_04673_),
    .ZN(_04674_));
 OAI22_X2 _22063_ (.A1(_04381_),
    .A2(_04672_),
    .B1(_04674_),
    .B2(_04608_),
    .ZN(_04675_));
 NOR2_X1 _22064_ (.A1(_01177_),
    .A2(_04461_),
    .ZN(_04676_));
 AOI21_X2 _22065_ (.A(_04676_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[18] ),
    .ZN(_04677_));
 AOI22_X2 _22066_ (.A1(\cs_registers_i.csr_depc_o[18] ),
    .A2(_04408_),
    .B1(_04427_),
    .B2(\cs_registers_i.dscratch1_q[18] ),
    .ZN(_04678_));
 NAND2_X2 _22067_ (.A1(_04677_),
    .A2(_04678_),
    .ZN(_04679_));
 AOI222_X2 _22068_ (.A1(\cs_registers_i.dscratch0_q[18] ),
    .A2(_04416_),
    .B1(_04413_),
    .B2(\cs_registers_i.mtval_q[18] ),
    .C1(_04447_),
    .C2(\cs_registers_i.mie_q[2] ),
    .ZN(_04680_));
 AOI22_X1 _22069_ (.A1(net70),
    .A2(_04637_),
    .B1(_04430_),
    .B2(net133),
    .ZN(_04681_));
 AOI21_X1 _22070_ (.A(_04545_),
    .B1(_04559_),
    .B2(\cs_registers_i.mscratch_q[18] ),
    .ZN(_04682_));
 NAND3_X1 _22071_ (.A1(_04680_),
    .A2(_04681_),
    .A3(_04682_),
    .ZN(_04683_));
 OR3_X4 _22072_ (.A1(_04675_),
    .A2(_04679_),
    .A3(_04683_),
    .ZN(_04684_));
 OAI22_X4 _22073_ (.A1(_04668_),
    .A2(_04669_),
    .B1(_04684_),
    .B2(_16381_),
    .ZN(_04685_));
 INV_X1 _22074_ (.A(\cs_registers_i.csr_mtvec_o[18] ),
    .ZN(_04686_));
 OAI221_X1 _22075_ (.A(_04667_),
    .B1(_04685_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04686_),
    .ZN(_01193_));
 NAND2_X1 _22076_ (.A1(net18),
    .A2(_04371_),
    .ZN(_04687_));
 MUX2_X1 _22077_ (.A(_04642_),
    .B(_04467_),
    .S(_16389_),
    .Z(_04688_));
 AOI22_X1 _22078_ (.A1(\cs_registers_i.dscratch0_q[19] ),
    .A2(_04415_),
    .B1(_04425_),
    .B2(\cs_registers_i.dscratch1_q[19] ),
    .ZN(_04689_));
 AOI22_X1 _22079_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_04407_),
    .B1(_04430_),
    .B2(net134),
    .ZN(_04690_));
 AOI222_X2 _22080_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_04412_),
    .B1(_04422_),
    .B2(\cs_registers_i.csr_mepc_o[19] ),
    .C1(_04507_),
    .C2(\cs_registers_i.mscratch_q[19] ),
    .ZN(_04691_));
 OAI21_X1 _22081_ (.A(_04456_),
    .B1(_04459_),
    .B2(_01178_),
    .ZN(_04692_));
 AOI221_X1 _22082_ (.A(_04692_),
    .B1(_04441_),
    .B2(net71),
    .C1(\cs_registers_i.mie_q[3] ),
    .C2(_04447_),
    .ZN(_04693_));
 AND4_X1 _22083_ (.A1(_04689_),
    .A2(_04690_),
    .A3(_04691_),
    .A4(_04693_),
    .ZN(_04694_));
 AOI22_X2 _22084_ (.A1(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .A2(_04387_),
    .B1(_04391_),
    .B2(\cs_registers_i.mhpmcounter[2][19] ),
    .ZN(_04695_));
 BUF_X2 _22085_ (.A(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .Z(_04696_));
 BUF_X2 _22086_ (.A(\cs_registers_i.mhpmcounter[2][51] ),
    .Z(_04697_));
 AOI22_X2 _22087_ (.A1(_04696_),
    .A2(_04388_),
    .B1(_04391_),
    .B2(_04697_),
    .ZN(_04698_));
 OAI221_X2 _22088_ (.A(_04694_),
    .B1(_04695_),
    .B2(_04401_),
    .C1(_04379_),
    .C2(_04698_),
    .ZN(_04699_));
 OAI22_X4 _22089_ (.A1(_04668_),
    .A2(_04688_),
    .B1(_04699_),
    .B2(_16389_),
    .ZN(_04700_));
 INV_X1 _22090_ (.A(\cs_registers_i.csr_mtvec_o[19] ),
    .ZN(_04701_));
 OAI221_X1 _22091_ (.A(_04687_),
    .B1(_04700_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04701_),
    .ZN(_01194_));
 NAND2_X1 _22092_ (.A1(net19),
    .A2(_04371_),
    .ZN(_04702_));
 CLKBUF_X3 _22093_ (.A(\cs_registers_i.mhpmcounter[2][52] ),
    .Z(_04703_));
 AOI22_X4 _22094_ (.A1(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .A2(_04500_),
    .B1(_04501_),
    .B2(_04703_),
    .ZN(_04704_));
 BUF_X2 _22095_ (.A(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .Z(_04705_));
 BUF_X2 _22096_ (.A(\cs_registers_i.mhpmcounter[2][20] ),
    .Z(_04706_));
 AOI22_X4 _22097_ (.A1(_04705_),
    .A2(_04500_),
    .B1(_04501_),
    .B2(_04706_),
    .ZN(_04707_));
 OAI22_X4 _22098_ (.A1(_04498_),
    .A2(_04704_),
    .B1(_04707_),
    .B2(_04402_),
    .ZN(_04708_));
 AOI22_X2 _22099_ (.A1(\cs_registers_i.dscratch0_q[20] ),
    .A2(_04632_),
    .B1(_04448_),
    .B2(\cs_registers_i.mie_q[4] ),
    .ZN(_04709_));
 AOI22_X2 _22100_ (.A1(\cs_registers_i.mtval_q[20] ),
    .A2(_04634_),
    .B1(_04431_),
    .B2(net135),
    .ZN(_04710_));
 NOR2_X2 _22101_ (.A1(_01179_),
    .A2(_04461_),
    .ZN(_04711_));
 AOI21_X1 _22102_ (.A(_04711_),
    .B1(_04442_),
    .B2(net73),
    .ZN(_04712_));
 NAND4_X2 _22103_ (.A1(_04514_),
    .A2(_04709_),
    .A3(_04710_),
    .A4(_04712_),
    .ZN(_04713_));
 AOI22_X1 _22104_ (.A1(\cs_registers_i.csr_depc_o[20] ),
    .A2(_04518_),
    .B1(_04509_),
    .B2(\cs_registers_i.mscratch_q[20] ),
    .ZN(_04714_));
 AOI22_X2 _22105_ (.A1(\cs_registers_i.csr_mepc_o[20] ),
    .A2(_04424_),
    .B1(_04523_),
    .B2(\cs_registers_i.dscratch1_q[20] ),
    .ZN(_04715_));
 NAND2_X2 _22106_ (.A1(_04714_),
    .A2(_04715_),
    .ZN(_04716_));
 NOR3_X4 _22107_ (.A1(_04708_),
    .A2(_04713_),
    .A3(_04716_),
    .ZN(_04717_));
 NAND2_X1 _22108_ (.A1(_16398_),
    .A2(_04717_),
    .ZN(_04718_));
 MUX2_X1 _22109_ (.A(_04642_),
    .B(_04643_),
    .S(_16402_),
    .Z(_04719_));
 OAI21_X2 _22110_ (.A(_04718_),
    .B1(_04719_),
    .B2(_04668_),
    .ZN(_04720_));
 BUF_X4 _22111_ (.A(_04720_),
    .Z(_04721_));
 INV_X1 _22112_ (.A(\cs_registers_i.csr_mtvec_o[20] ),
    .ZN(_04722_));
 OAI221_X1 _22113_ (.A(_04702_),
    .B1(_04721_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04722_),
    .ZN(_01195_));
 BUF_X2 _22114_ (.A(_04370_),
    .Z(_04723_));
 NAND2_X1 _22115_ (.A1(net20),
    .A2(_04723_),
    .ZN(_04724_));
 MUX2_X1 _22116_ (.A(_04601_),
    .B(_15928_),
    .S(_16410_),
    .Z(_04725_));
 NOR2_X1 _22117_ (.A1(_01180_),
    .A2(_04460_),
    .ZN(_04726_));
 AOI21_X1 _22118_ (.A(_04726_),
    .B1(_04416_),
    .B2(\cs_registers_i.dscratch0_q[21] ),
    .ZN(_04727_));
 AOI22_X1 _22119_ (.A1(\cs_registers_i.dscratch1_q[21] ),
    .A2(_04426_),
    .B1(_04430_),
    .B2(net136),
    .ZN(_04728_));
 AOI22_X1 _22120_ (.A1(net74),
    .A2(_04441_),
    .B1(_04447_),
    .B2(\cs_registers_i.mie_q[5] ),
    .ZN(_04729_));
 AOI21_X1 _22121_ (.A(_04544_),
    .B1(_04413_),
    .B2(\cs_registers_i.mtval_q[21] ),
    .ZN(_04730_));
 NAND4_X1 _22122_ (.A1(_04727_),
    .A2(_04728_),
    .A3(_04729_),
    .A4(_04730_),
    .ZN(_04731_));
 NAND2_X1 _22123_ (.A1(\cs_registers_i.mscratch_q[21] ),
    .A2(_04508_),
    .ZN(_04732_));
 AOI222_X2 _22124_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(_04407_),
    .B1(_04423_),
    .B2(\cs_registers_i.csr_mepc_o[21] ),
    .C1(_04657_),
    .C2(\cs_registers_i.csr_mstatus_tw_o ),
    .ZN(_04733_));
 NAND2_X1 _22125_ (.A1(_04732_),
    .A2(_04733_),
    .ZN(_04734_));
 NOR2_X2 _22126_ (.A1(_04731_),
    .A2(_04734_),
    .ZN(_04735_));
 CLKBUF_X2 _22127_ (.A(\cs_registers_i.mhpmcounter[2][21] ),
    .Z(_04736_));
 AOI22_X2 _22128_ (.A1(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .A2(_04589_),
    .B1(_04591_),
    .B2(_04736_),
    .ZN(_04737_));
 CLKBUF_X3 _22129_ (.A(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .Z(_04738_));
 BUF_X2 _22130_ (.A(\cs_registers_i.mhpmcounter[2][53] ),
    .Z(_04739_));
 AOI22_X2 _22131_ (.A1(_04738_),
    .A2(_04589_),
    .B1(_04591_),
    .B2(_04739_),
    .ZN(_04740_));
 OAI221_X2 _22132_ (.A(_04735_),
    .B1(_04737_),
    .B2(_04608_),
    .C1(_04381_),
    .C2(_04740_),
    .ZN(_04741_));
 OAI22_X4 _22133_ (.A1(_04600_),
    .A2(_04725_),
    .B1(_04741_),
    .B2(_16410_),
    .ZN(_04742_));
 INV_X1 _22134_ (.A(\cs_registers_i.csr_mtvec_o[21] ),
    .ZN(_04743_));
 OAI221_X1 _22135_ (.A(_04724_),
    .B1(_04742_),
    .B2(_04492_),
    .C1(_04494_),
    .C2(_04743_),
    .ZN(_01196_));
 INV_X1 _22136_ (.A(\cs_registers_i.csr_mtvec_o[22] ),
    .ZN(_04744_));
 MUX2_X1 _22137_ (.A(_04642_),
    .B(_04643_),
    .S(_16418_),
    .Z(_04745_));
 NAND2_X1 _22138_ (.A1(\cs_registers_i.mtval_q[22] ),
    .A2(_04413_),
    .ZN(_04746_));
 OAI21_X1 _22139_ (.A(_04746_),
    .B1(_04460_),
    .B2(_01181_),
    .ZN(_04747_));
 AOI221_X1 _22140_ (.A(_04747_),
    .B1(_04416_),
    .B2(\cs_registers_i.dscratch0_q[22] ),
    .C1(\cs_registers_i.dscratch1_q[22] ),
    .C2(_04426_),
    .ZN(_04748_));
 AOI222_X2 _22141_ (.A1(\cs_registers_i.csr_mepc_o[22] ),
    .A2(_04615_),
    .B1(_04559_),
    .B2(\cs_registers_i.mscratch_q[22] ),
    .C1(_04448_),
    .C2(\cs_registers_i.mie_q[6] ),
    .ZN(_04749_));
 AOI222_X2 _22142_ (.A1(net75),
    .A2(_04442_),
    .B1(_04408_),
    .B2(\cs_registers_i.csr_depc_o[22] ),
    .C1(net137),
    .C2(_04430_),
    .ZN(_04750_));
 AND4_X1 _22143_ (.A1(_04457_),
    .A2(_04748_),
    .A3(_04749_),
    .A4(_04750_),
    .ZN(_04751_));
 BUF_X4 _22144_ (.A(_04389_),
    .Z(_04752_));
 BUF_X4 _22145_ (.A(_04393_),
    .Z(_04753_));
 CLKBUF_X2 _22146_ (.A(\cs_registers_i.mhpmcounter[2][22] ),
    .Z(_04754_));
 AOI22_X2 _22147_ (.A1(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04754_),
    .ZN(_04755_));
 BUF_X4 _22148_ (.A(_04498_),
    .Z(_04756_));
 BUF_X2 _22149_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .Z(_04757_));
 CLKBUF_X2 _22150_ (.A(\cs_registers_i.mhpmcounter[2][54] ),
    .Z(_04758_));
 AOI22_X2 _22151_ (.A1(_04757_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04758_),
    .ZN(_04759_));
 OAI221_X2 _22152_ (.A(_04751_),
    .B1(_04755_),
    .B2(_04629_),
    .C1(_04756_),
    .C2(_04759_),
    .ZN(_04760_));
 OAI22_X4 _22153_ (.A1(_04668_),
    .A2(_04745_),
    .B1(_04760_),
    .B2(_16418_),
    .ZN(_04761_));
 BUF_X4 _22154_ (.A(_04761_),
    .Z(_04762_));
 OAI22_X1 _22155_ (.A1(_04744_),
    .A2(_04493_),
    .B1(_04762_),
    .B2(_04491_),
    .ZN(_04763_));
 AOI21_X1 _22156_ (.A(_04763_),
    .B1(_04371_),
    .B2(net21),
    .ZN(_04764_));
 INV_X1 _22157_ (.A(_04764_),
    .ZN(_01197_));
 NAND2_X1 _22158_ (.A1(net22),
    .A2(_04723_),
    .ZN(_04765_));
 MUX2_X1 _22159_ (.A(_04601_),
    .B(_04643_),
    .S(_16421_),
    .Z(_04766_));
 NOR2_X1 _22160_ (.A1(_03580_),
    .A2(_04398_),
    .ZN(_04767_));
 NOR4_X2 _22161_ (.A1(_03585_),
    .A2(_03604_),
    .A3(_03622_),
    .A4(_04767_),
    .ZN(_04768_));
 NOR3_X1 _22162_ (.A1(_03621_),
    .A2(_03604_),
    .A3(_03622_),
    .ZN(_04769_));
 AOI222_X2 _22163_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(_04768_),
    .B1(_04769_),
    .B2(net138),
    .C1(_04571_),
    .C2(\cs_registers_i.csr_mepc_o[23] ),
    .ZN(_04770_));
 NAND2_X1 _22164_ (.A1(\cs_registers_i.mtval_q[23] ),
    .A2(_04570_),
    .ZN(_04771_));
 OAI21_X1 _22165_ (.A(_04771_),
    .B1(_04580_),
    .B2(_01182_),
    .ZN(_04772_));
 AOI221_X2 _22166_ (.A(_04772_),
    .B1(_04575_),
    .B2(\cs_registers_i.mscratch_q[23] ),
    .C1(\cs_registers_i.csr_depc_o[23] ),
    .C2(_04569_),
    .ZN(_04773_));
 AOI221_X2 _22167_ (.A(_04573_),
    .B1(_04583_),
    .B2(\cs_registers_i.dscratch0_q[23] ),
    .C1(net76),
    .C2(_04574_),
    .ZN(_04774_));
 NAND2_X2 _22168_ (.A1(\cs_registers_i.dscratch1_q[23] ),
    .A2(_04584_),
    .ZN(_04775_));
 NAND4_X4 _22169_ (.A1(_04770_),
    .A2(_04773_),
    .A3(_04774_),
    .A4(_04775_),
    .ZN(_04776_));
 CLKBUF_X3 _22170_ (.A(\cs_registers_i.mhpmcounter[2][55] ),
    .Z(_04777_));
 AOI22_X4 _22171_ (.A1(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .A2(_04590_),
    .B1(_04592_),
    .B2(_04777_),
    .ZN(_04778_));
 CLKBUF_X3 _22172_ (.A(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .Z(_04779_));
 AOI22_X4 _22173_ (.A1(_04779_),
    .A2(_04590_),
    .B1(_04592_),
    .B2(\cs_registers_i.mhpmcounter[2][23] ),
    .ZN(_04780_));
 OAI22_X4 _22174_ (.A1(_04588_),
    .A2(_04778_),
    .B1(_04780_),
    .B2(_03583_),
    .ZN(_04781_));
 OR2_X1 _22175_ (.A1(_04776_),
    .A2(_04781_),
    .ZN(_04782_));
 OAI22_X4 _22176_ (.A1(_04600_),
    .A2(_04766_),
    .B1(_04782_),
    .B2(_16421_),
    .ZN(_04783_));
 CLKBUF_X3 _22177_ (.A(_04491_),
    .Z(_04784_));
 CLKBUF_X3 _22178_ (.A(_04493_),
    .Z(_04785_));
 INV_X1 _22179_ (.A(\cs_registers_i.csr_mtvec_o[23] ),
    .ZN(_04786_));
 OAI221_X1 _22180_ (.A(_04765_),
    .B1(_04783_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04786_),
    .ZN(_01198_));
 NAND2_X1 _22181_ (.A1(net23),
    .A2(_04723_),
    .ZN(_04787_));
 BUF_X2 _22182_ (.A(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .Z(_04788_));
 CLKBUF_X3 _22183_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .Z(_04789_));
 AOI22_X4 _22184_ (.A1(_04788_),
    .A2(_04590_),
    .B1(_04592_),
    .B2(_04789_),
    .ZN(_04790_));
 AOI22_X4 _22185_ (.A1(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .A2(_04590_),
    .B1(_04592_),
    .B2(\cs_registers_i.mhpmcounter[2][24] ),
    .ZN(_04791_));
 OAI22_X4 _22186_ (.A1(_04498_),
    .A2(_04790_),
    .B1(_04791_),
    .B2(_04629_),
    .ZN(_04792_));
 AOI22_X1 _22187_ (.A1(\cs_registers_i.dscratch0_q[24] ),
    .A2(_04632_),
    .B1(_04523_),
    .B2(\cs_registers_i.dscratch1_q[24] ),
    .ZN(_04793_));
 NOR2_X1 _22188_ (.A1(_01183_),
    .A2(_04461_),
    .ZN(_04794_));
 AOI21_X2 _22189_ (.A(_04794_),
    .B1(_04634_),
    .B2(\cs_registers_i.mtval_q[24] ),
    .ZN(_04795_));
 NAND2_X1 _22190_ (.A1(_04793_),
    .A2(_04795_),
    .ZN(_04796_));
 AOI222_X2 _22191_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(_04518_),
    .B1(_04509_),
    .B2(\cs_registers_i.mscratch_q[24] ),
    .C1(_04448_),
    .C2(\cs_registers_i.mie_q[8] ),
    .ZN(_04797_));
 AOI22_X2 _22192_ (.A1(net77),
    .A2(_04442_),
    .B1(_04431_),
    .B2(net139),
    .ZN(_04798_));
 AOI21_X1 _22193_ (.A(_04545_),
    .B1(_04424_),
    .B2(\cs_registers_i.csr_mepc_o[24] ),
    .ZN(_04799_));
 NAND3_X2 _22194_ (.A1(_04797_),
    .A2(_04798_),
    .A3(_04799_),
    .ZN(_04800_));
 NOR3_X4 _22195_ (.A1(_04792_),
    .A2(_04796_),
    .A3(_04800_),
    .ZN(_04801_));
 NAND2_X1 _22196_ (.A1(_16433_),
    .A2(_04801_),
    .ZN(_04802_));
 MUX2_X1 _22197_ (.A(_04466_),
    .B(_04467_),
    .S(_16429_),
    .Z(_04803_));
 OAI21_X4 _22198_ (.A(_04802_),
    .B1(_04803_),
    .B2(_04470_),
    .ZN(_04804_));
 BUF_X4 _22199_ (.A(_04804_),
    .Z(_04805_));
 INV_X1 _22200_ (.A(\cs_registers_i.csr_mtvec_o[24] ),
    .ZN(_04806_));
 OAI221_X1 _22201_ (.A(_04787_),
    .B1(_04805_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04806_),
    .ZN(_01199_));
 NAND2_X1 _22202_ (.A1(net24),
    .A2(_04723_),
    .ZN(_04807_));
 MUX2_X1 _22203_ (.A(_04601_),
    .B(_15928_),
    .S(_16437_),
    .Z(_04808_));
 AOI22_X1 _22204_ (.A1(\cs_registers_i.dscratch0_q[25] ),
    .A2(_04417_),
    .B1(_04427_),
    .B2(\cs_registers_i.dscratch1_q[25] ),
    .ZN(_04809_));
 AOI22_X1 _22205_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(_04408_),
    .B1(_04431_),
    .B2(net140),
    .ZN(_04810_));
 AOI222_X2 _22206_ (.A1(\cs_registers_i.mtval_q[25] ),
    .A2(_04414_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[25] ),
    .C1(_04508_),
    .C2(\cs_registers_i.mscratch_q[25] ),
    .ZN(_04811_));
 OAI21_X1 _22207_ (.A(_04457_),
    .B1(_04460_),
    .B2(_01184_),
    .ZN(_04812_));
 AOI221_X1 _22208_ (.A(_04812_),
    .B1(_04441_),
    .B2(net78),
    .C1(\cs_registers_i.mie_q[9] ),
    .C2(_04447_),
    .ZN(_04813_));
 AND4_X1 _22209_ (.A1(_04809_),
    .A2(_04810_),
    .A3(_04811_),
    .A4(_04813_),
    .ZN(_04814_));
 CLKBUF_X2 _22210_ (.A(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .Z(_04815_));
 CLKBUF_X2 _22211_ (.A(\cs_registers_i.mhpmcounter[2][25] ),
    .Z(_04816_));
 AOI22_X2 _22212_ (.A1(_04815_),
    .A2(_04590_),
    .B1(_04592_),
    .B2(_04816_),
    .ZN(_04817_));
 BUF_X2 _22213_ (.A(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .Z(_04818_));
 BUF_X2 _22214_ (.A(\cs_registers_i.mhpmcounter[2][57] ),
    .Z(_04819_));
 AOI22_X2 _22215_ (.A1(_04818_),
    .A2(_04590_),
    .B1(_04592_),
    .B2(_04819_),
    .ZN(_04820_));
 OAI221_X2 _22216_ (.A(_04814_),
    .B1(_04817_),
    .B2(_04629_),
    .C1(_04498_),
    .C2(_04820_),
    .ZN(_04821_));
 OAI22_X4 _22217_ (.A1(_04600_),
    .A2(_04808_),
    .B1(_04821_),
    .B2(_16437_),
    .ZN(_04822_));
 INV_X1 _22218_ (.A(\cs_registers_i.csr_mtvec_o[25] ),
    .ZN(_04823_));
 OAI221_X1 _22219_ (.A(_04807_),
    .B1(_04822_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04823_),
    .ZN(_01200_));
 NAND2_X1 _22220_ (.A1(net25),
    .A2(_04723_),
    .ZN(_04824_));
 MUX2_X1 _22221_ (.A(_04467_),
    .B(_04466_),
    .S(_16449_),
    .Z(_04825_));
 AOI22_X1 _22222_ (.A1(\cs_registers_i.dscratch0_q[26] ),
    .A2(_04632_),
    .B1(_04523_),
    .B2(\cs_registers_i.dscratch1_q[26] ),
    .ZN(_04826_));
 AOI22_X1 _22223_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(_04518_),
    .B1(_04431_),
    .B2(net127),
    .ZN(_04827_));
 AOI222_X2 _22224_ (.A1(\cs_registers_i.mtval_q[26] ),
    .A2(_04634_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[26] ),
    .C1(_04559_),
    .C2(\cs_registers_i.mscratch_q[26] ),
    .ZN(_04828_));
 OAI21_X1 _22225_ (.A(_04457_),
    .B1(_04460_),
    .B2(_01185_),
    .ZN(_04829_));
 AOI221_X1 _22226_ (.A(_04829_),
    .B1(_04637_),
    .B2(net79),
    .C1(\cs_registers_i.mie_q[10] ),
    .C2(_04448_),
    .ZN(_04830_));
 AND4_X2 _22227_ (.A1(_04826_),
    .A2(_04827_),
    .A3(_04828_),
    .A4(_04830_),
    .ZN(_04831_));
 BUF_X2 _22228_ (.A(\cs_registers_i.mhpmcounter[2][26] ),
    .Z(_04832_));
 AOI22_X2 _22229_ (.A1(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04832_),
    .ZN(_04833_));
 BUF_X2 _22230_ (.A(\cs_registers_i.mhpmcounter[2][58] ),
    .Z(_04834_));
 AOI22_X2 _22231_ (.A1(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04834_),
    .ZN(_04835_));
 OAI221_X2 _22232_ (.A(_04831_),
    .B1(_04833_),
    .B2(_04629_),
    .C1(_04756_),
    .C2(_04835_),
    .ZN(_04836_));
 OAI22_X4 _22233_ (.A1(_04470_),
    .A2(_04825_),
    .B1(_04836_),
    .B2(_16445_),
    .ZN(_04837_));
 BUF_X4 _22234_ (.A(_04837_),
    .Z(_04838_));
 INV_X1 _22235_ (.A(\cs_registers_i.csr_mtvec_o[26] ),
    .ZN(_04839_));
 OAI221_X1 _22236_ (.A(_04824_),
    .B1(_04838_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04839_),
    .ZN(_01201_));
 NAND2_X1 _22237_ (.A1(net26),
    .A2(_04723_),
    .ZN(_04840_));
 MUX2_X1 _22238_ (.A(_04642_),
    .B(_04643_),
    .S(_16453_),
    .Z(_04841_));
 AOI22_X1 _22239_ (.A1(\cs_registers_i.dscratch0_q[27] ),
    .A2(_04632_),
    .B1(_04523_),
    .B2(\cs_registers_i.dscratch1_q[27] ),
    .ZN(_04842_));
 AOI22_X1 _22240_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(_04518_),
    .B1(_04431_),
    .B2(net128),
    .ZN(_04843_));
 AOI222_X2 _22241_ (.A1(\cs_registers_i.mtval_q[27] ),
    .A2(_04634_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[27] ),
    .C1(_04559_),
    .C2(\cs_registers_i.mscratch_q[27] ),
    .ZN(_04844_));
 OAI21_X1 _22242_ (.A(_04457_),
    .B1(_04460_),
    .B2(_00007_),
    .ZN(_04845_));
 AOI221_X1 _22243_ (.A(_04845_),
    .B1(_04637_),
    .B2(net80),
    .C1(\cs_registers_i.mie_q[11] ),
    .C2(_04447_),
    .ZN(_04846_));
 AND4_X1 _22244_ (.A1(_04842_),
    .A2(_04843_),
    .A3(_04844_),
    .A4(_04846_),
    .ZN(_04847_));
 AOI22_X2 _22245_ (.A1(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\cs_registers_i.mhpmcounter[2][27] ),
    .ZN(_04848_));
 BUF_X2 _22246_ (.A(\cs_registers_i.mhpmcounter[2][59] ),
    .Z(_04849_));
 AOI22_X2 _22247_ (.A1(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04849_),
    .ZN(_04850_));
 OAI221_X2 _22248_ (.A(_04847_),
    .B1(_04848_),
    .B2(_04629_),
    .C1(_04498_),
    .C2(_04850_),
    .ZN(_04851_));
 OAI22_X4 _22249_ (.A1(_04668_),
    .A2(_04841_),
    .B1(_04851_),
    .B2(_16453_),
    .ZN(_04852_));
 BUF_X4 _22250_ (.A(_04852_),
    .Z(_04853_));
 INV_X1 _22251_ (.A(\cs_registers_i.csr_mtvec_o[27] ),
    .ZN(_04854_));
 OAI221_X1 _22252_ (.A(_04840_),
    .B1(_04853_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04854_),
    .ZN(_01202_));
 NAND2_X1 _22253_ (.A1(net27),
    .A2(_04723_),
    .ZN(_04855_));
 MUX2_X1 _22254_ (.A(_04642_),
    .B(_04643_),
    .S(_16461_),
    .Z(_04856_));
 AOI22_X1 _22255_ (.A1(\cs_registers_i.dscratch0_q[28] ),
    .A2(_04632_),
    .B1(_04523_),
    .B2(\cs_registers_i.dscratch1_q[28] ),
    .ZN(_04857_));
 AOI22_X1 _22256_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(_04518_),
    .B1(_04431_),
    .B2(net129),
    .ZN(_04858_));
 AOI222_X2 _22257_ (.A1(\cs_registers_i.mtval_q[28] ),
    .A2(_04634_),
    .B1(_04424_),
    .B2(\cs_registers_i.csr_mepc_o[28] ),
    .C1(_04509_),
    .C2(\cs_registers_i.mscratch_q[28] ),
    .ZN(_04859_));
 OAI21_X1 _22258_ (.A(_04457_),
    .B1(_04460_),
    .B2(_00008_),
    .ZN(_04860_));
 AOI221_X1 _22259_ (.A(_04860_),
    .B1(_04637_),
    .B2(net81),
    .C1(\cs_registers_i.mie_q[12] ),
    .C2(_04448_),
    .ZN(_04861_));
 AND4_X2 _22260_ (.A1(_04857_),
    .A2(_04858_),
    .A3(_04859_),
    .A4(_04861_),
    .ZN(_04862_));
 AOI22_X2 _22261_ (.A1(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(\cs_registers_i.mhpmcounter[2][28] ),
    .ZN(_04863_));
 BUF_X2 _22262_ (.A(\cs_registers_i.mhpmcounter[2][60] ),
    .Z(_04864_));
 AOI22_X2 _22263_ (.A1(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_04864_),
    .ZN(_04865_));
 OAI221_X2 _22264_ (.A(_04862_),
    .B1(_04863_),
    .B2(_04629_),
    .C1(_04756_),
    .C2(_04865_),
    .ZN(_04866_));
 OAI22_X4 _22265_ (.A1(_04668_),
    .A2(_04856_),
    .B1(_04866_),
    .B2(_16461_),
    .ZN(_04867_));
 BUF_X4 _22266_ (.A(_04867_),
    .Z(_04868_));
 INV_X1 _22267_ (.A(\cs_registers_i.csr_mtvec_o[28] ),
    .ZN(_04869_));
 OAI221_X1 _22268_ (.A(_04855_),
    .B1(_04868_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04869_),
    .ZN(_01203_));
 NAND2_X1 _22269_ (.A1(net28),
    .A2(_04723_),
    .ZN(_04870_));
 MUX2_X1 _22270_ (.A(_04601_),
    .B(_15928_),
    .S(_16469_),
    .Z(_04871_));
 AOI22_X1 _22271_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(_04407_),
    .B1(_04426_),
    .B2(\cs_registers_i.dscratch1_q[29] ),
    .ZN(_04872_));
 NOR2_X1 _22272_ (.A1(_00009_),
    .A2(_04459_),
    .ZN(_04873_));
 AOI21_X1 _22273_ (.A(_04873_),
    .B1(_04447_),
    .B2(\cs_registers_i.mie_q[13] ),
    .ZN(_04874_));
 AOI222_X2 _22274_ (.A1(\cs_registers_i.dscratch0_q[29] ),
    .A2(_04415_),
    .B1(_04422_),
    .B2(\cs_registers_i.csr_mepc_o[29] ),
    .C1(_04508_),
    .C2(\cs_registers_i.mscratch_q[29] ),
    .ZN(_04875_));
 NAND2_X1 _22275_ (.A1(\cs_registers_i.mtval_q[29] ),
    .A2(_04412_),
    .ZN(_04876_));
 NAND2_X1 _22276_ (.A1(_04457_),
    .A2(_04876_),
    .ZN(_04877_));
 AOI221_X1 _22277_ (.A(_04877_),
    .B1(_04441_),
    .B2(net82),
    .C1(net130),
    .C2(_04430_),
    .ZN(_04878_));
 AND4_X2 _22278_ (.A1(_04872_),
    .A2(_04874_),
    .A3(_04875_),
    .A4(_04878_),
    .ZN(_04879_));
 BUF_X2 _22279_ (.A(\cs_registers_i.mhpmcounter[2][29] ),
    .Z(_04880_));
 AOI22_X2 _22280_ (.A1(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .A2(_04388_),
    .B1(_04391_),
    .B2(_04880_),
    .ZN(_04881_));
 BUF_X2 _22281_ (.A(\cs_registers_i.mhpmcounter[2][61] ),
    .Z(_04882_));
 AOI22_X2 _22282_ (.A1(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .A2(_04499_),
    .B1(_04392_),
    .B2(_04882_),
    .ZN(_04883_));
 OAI221_X2 _22283_ (.A(_04879_),
    .B1(_04881_),
    .B2(_04608_),
    .C1(_04380_),
    .C2(_04883_),
    .ZN(_04884_));
 OAI22_X4 _22284_ (.A1(_04600_),
    .A2(_04871_),
    .B1(_04884_),
    .B2(_16469_),
    .ZN(_04885_));
 INV_X1 _22285_ (.A(\cs_registers_i.csr_mtvec_o[29] ),
    .ZN(_04886_));
 OAI221_X1 _22286_ (.A(_04870_),
    .B1(_04885_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04886_),
    .ZN(_01204_));
 NAND2_X1 _22287_ (.A1(net29),
    .A2(_04723_),
    .ZN(_04887_));
 BUF_X2 _22288_ (.A(\cs_registers_i.mhpmcounter[2][62] ),
    .Z(_04888_));
 AOI22_X4 _22289_ (.A1(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .A2(_04389_),
    .B1(_04393_),
    .B2(_04888_),
    .ZN(_04889_));
 AOI22_X4 _22290_ (.A1(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .A2(_04389_),
    .B1(_04393_),
    .B2(\cs_registers_i.mhpmcounter[2][30] ),
    .ZN(_04890_));
 OAI22_X4 _22291_ (.A1(_04381_),
    .A2(_04889_),
    .B1(_04890_),
    .B2(_04402_),
    .ZN(_04891_));
 AOI22_X2 _22292_ (.A1(\cs_registers_i.dscratch0_q[30] ),
    .A2(_04632_),
    .B1(_04523_),
    .B2(\cs_registers_i.dscratch1_q[30] ),
    .ZN(_04892_));
 AOI222_X2 _22293_ (.A1(\cs_registers_i.mtval_q[30] ),
    .A2(_04414_),
    .B1(_04559_),
    .B2(\cs_registers_i.mscratch_q[30] ),
    .C1(_04448_),
    .C2(\cs_registers_i.mie_q[14] ),
    .ZN(_04893_));
 NOR2_X1 _22294_ (.A1(_00010_),
    .A2(_04461_),
    .ZN(_04894_));
 AOI21_X2 _22295_ (.A(_04894_),
    .B1(_04518_),
    .B2(\cs_registers_i.csr_depc_o[30] ),
    .ZN(_04895_));
 NAND3_X2 _22296_ (.A1(_04892_),
    .A2(_04893_),
    .A3(_04895_),
    .ZN(_04896_));
 AOI22_X2 _22297_ (.A1(net84),
    .A2(_04442_),
    .B1(_04431_),
    .B2(net131),
    .ZN(_04897_));
 NAND2_X1 _22298_ (.A1(_04514_),
    .A2(_04897_),
    .ZN(_04898_));
 AND2_X1 _22299_ (.A1(\cs_registers_i.csr_mepc_o[30] ),
    .A2(_04423_),
    .ZN(_04899_));
 OR2_X1 _22300_ (.A1(_04433_),
    .A2(_04899_),
    .ZN(_04900_));
 NOR4_X4 _22301_ (.A1(_04891_),
    .A2(_04896_),
    .A3(_04898_),
    .A4(_04900_),
    .ZN(_04901_));
 NAND2_X1 _22302_ (.A1(_16478_),
    .A2(_04901_),
    .ZN(_04902_));
 MUX2_X1 _22303_ (.A(_04642_),
    .B(_04643_),
    .S(_16482_),
    .Z(_04903_));
 OAI21_X4 _22304_ (.A(_04902_),
    .B1(_04903_),
    .B2(_04470_),
    .ZN(_04904_));
 BUF_X4 _22305_ (.A(_04904_),
    .Z(_04905_));
 INV_X1 _22306_ (.A(\cs_registers_i.csr_mtvec_o[30] ),
    .ZN(_04906_));
 OAI221_X1 _22307_ (.A(_04887_),
    .B1(_04905_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04906_),
    .ZN(_01205_));
 NAND2_X1 _22308_ (.A1(net30),
    .A2(_04723_),
    .ZN(_04907_));
 MUX2_X1 _22309_ (.A(_04467_),
    .B(_04642_),
    .S(_15894_),
    .Z(_04908_));
 BUF_X2 _22310_ (.A(\cs_registers_i.mhpmcounter[2][63] ),
    .Z(_04909_));
 AOI22_X4 _22311_ (.A1(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .A2(_04389_),
    .B1(_04393_),
    .B2(_04909_),
    .ZN(_04910_));
 BUF_X2 _22312_ (.A(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .Z(_04911_));
 AOI22_X4 _22313_ (.A1(_04911_),
    .A2(_04389_),
    .B1(_04591_),
    .B2(\cs_registers_i.mhpmcounter[2][31] ),
    .ZN(_04912_));
 OAI22_X4 _22314_ (.A1(_04381_),
    .A2(_04910_),
    .B1(_04912_),
    .B2(_04402_),
    .ZN(_04913_));
 NAND2_X1 _22315_ (.A1(\cs_registers_i.mscratch_q[31] ),
    .A2(_04509_),
    .ZN(_04914_));
 NOR2_X1 _22316_ (.A1(_00011_),
    .A2(_04460_),
    .ZN(_04915_));
 AOI221_X2 _22317_ (.A(_04915_),
    .B1(_04441_),
    .B2(net85),
    .C1(\cs_registers_i.csr_depc_o[31] ),
    .C2(_04407_),
    .ZN(_04916_));
 AOI22_X2 _22318_ (.A1(\cs_registers_i.dscratch0_q[31] ),
    .A2(_04417_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[31] ),
    .ZN(_04917_));
 NOR2_X4 _22319_ (.A1(_04420_),
    .A2(_04390_),
    .ZN(_04918_));
 AOI22_X4 _22320_ (.A1(\cs_registers_i.mtval_q[31] ),
    .A2(_04634_),
    .B1(_04918_),
    .B2(\cs_registers_i.mcause_q[5] ),
    .ZN(_04919_));
 NAND4_X2 _22321_ (.A1(_04914_),
    .A2(_04916_),
    .A3(_04917_),
    .A4(_04919_),
    .ZN(_04920_));
 AND2_X1 _22322_ (.A1(\cs_registers_i.dscratch1_q[31] ),
    .A2(_04523_),
    .ZN(_04921_));
 OR4_X4 _22323_ (.A1(_04545_),
    .A2(_04913_),
    .A3(_04920_),
    .A4(_04921_),
    .ZN(_04922_));
 OAI22_X4 _22324_ (.A1(_04470_),
    .A2(_04908_),
    .B1(_04922_),
    .B2(_15898_),
    .ZN(_04923_));
 BUF_X4 _22325_ (.A(_04923_),
    .Z(_04924_));
 INV_X1 _22326_ (.A(\cs_registers_i.csr_mtvec_o[31] ),
    .ZN(_04925_));
 OAI221_X1 _22327_ (.A(_04907_),
    .B1(_04924_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04925_),
    .ZN(_01206_));
 NAND2_X1 _22328_ (.A1(net31),
    .A2(_04370_),
    .ZN(_04926_));
 MUX2_X1 _22329_ (.A(_04601_),
    .B(_15928_),
    .S(_16302_),
    .Z(_04927_));
 AOI222_X2 _22330_ (.A1(\cs_registers_i.dscratch0_q[8] ),
    .A2(_04632_),
    .B1(_04424_),
    .B2(\cs_registers_i.csr_mepc_o[8] ),
    .C1(_04427_),
    .C2(\cs_registers_i.dscratch1_q[8] ),
    .ZN(_04928_));
 CLKBUF_X3 _22331_ (.A(\cs_registers_i.mhpmcounter[2][40] ),
    .Z(_04929_));
 AOI22_X4 _22332_ (.A1(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .A2(_04499_),
    .B1(_04392_),
    .B2(_04929_),
    .ZN(_04930_));
 BUF_X2 _22333_ (.A(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .Z(_04931_));
 BUF_X2 _22334_ (.A(\cs_registers_i.mhpmcounter[2][8] ),
    .Z(_04932_));
 AOI22_X4 _22335_ (.A1(_04931_),
    .A2(_04499_),
    .B1(_04392_),
    .B2(_04932_),
    .ZN(_04933_));
 OAI22_X4 _22336_ (.A1(_04380_),
    .A2(_04930_),
    .B1(_04933_),
    .B2(_04608_),
    .ZN(_04934_));
 AOI22_X1 _22337_ (.A1(\cs_registers_i.csr_depc_o[8] ),
    .A2(_04408_),
    .B1(_04433_),
    .B2(\cs_registers_i.dcsr_q[8] ),
    .ZN(_04935_));
 AOI22_X1 _22338_ (.A1(\cs_registers_i.mtval_q[8] ),
    .A2(_04414_),
    .B1(_04508_),
    .B2(\cs_registers_i.mscratch_q[8] ),
    .ZN(_04936_));
 NAND3_X1 _22339_ (.A1(_04514_),
    .A2(_04935_),
    .A3(_04936_),
    .ZN(_04937_));
 INV_X1 _22340_ (.A(net91),
    .ZN(_04938_));
 OAI22_X2 _22341_ (.A1(_04938_),
    .A2(_04476_),
    .B1(_04461_),
    .B2(_01169_),
    .ZN(_04939_));
 NOR3_X2 _22342_ (.A1(_04934_),
    .A2(_04937_),
    .A3(_04939_),
    .ZN(_04940_));
 NAND2_X4 _22343_ (.A1(_04928_),
    .A2(_04940_),
    .ZN(_04941_));
 OAI22_X4 _22344_ (.A1(_04600_),
    .A2(_04927_),
    .B1(_04941_),
    .B2(_16302_),
    .ZN(_04942_));
 INV_X1 _22345_ (.A(\cs_registers_i.csr_mtvec_o[8] ),
    .ZN(_04943_));
 OAI221_X1 _22346_ (.A(_04926_),
    .B1(_04942_),
    .B2(_04784_),
    .C1(_04785_),
    .C2(_04943_),
    .ZN(_01207_));
 NAND2_X1 _22347_ (.A1(net32),
    .A2(_04370_),
    .ZN(_04944_));
 BUF_X2 _22348_ (.A(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .Z(_04945_));
 CLKBUF_X3 _22349_ (.A(\cs_registers_i.mhpmcounter[2][41] ),
    .Z(_04946_));
 AOI22_X4 _22350_ (.A1(_04945_),
    .A2(_04500_),
    .B1(_04393_),
    .B2(_04946_),
    .ZN(_04947_));
 CLKBUF_X3 _22351_ (.A(\cs_registers_i.mhpmcounter[2][9] ),
    .Z(_04948_));
 AOI22_X4 _22352_ (.A1(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .A2(_04389_),
    .B1(_04393_),
    .B2(_04948_),
    .ZN(_04949_));
 OAI22_X4 _22353_ (.A1(_04381_),
    .A2(_04947_),
    .B1(_04949_),
    .B2(_04402_),
    .ZN(_04950_));
 AOI222_X2 _22354_ (.A1(\cs_registers_i.csr_depc_o[9] ),
    .A2(_04408_),
    .B1(_04414_),
    .B2(\cs_registers_i.mtval_q[9] ),
    .C1(_04427_),
    .C2(\cs_registers_i.dscratch1_q[9] ),
    .ZN(_04951_));
 AOI22_X2 _22355_ (.A1(\cs_registers_i.dscratch0_q[9] ),
    .A2(_04632_),
    .B1(_04509_),
    .B2(\cs_registers_i.mscratch_q[9] ),
    .ZN(_04952_));
 NOR2_X1 _22356_ (.A1(_01170_),
    .A2(_04461_),
    .ZN(_04953_));
 AOI21_X1 _22357_ (.A(_04953_),
    .B1(_04442_),
    .B2(net92),
    .ZN(_04954_));
 NAND3_X2 _22358_ (.A1(_04951_),
    .A2(_04952_),
    .A3(_04954_),
    .ZN(_04955_));
 AND2_X1 _22359_ (.A1(\cs_registers_i.csr_mepc_o[9] ),
    .A2(_04424_),
    .ZN(_04956_));
 NOR4_X4 _22360_ (.A1(_04545_),
    .A2(_04950_),
    .A3(_04955_),
    .A4(_04956_),
    .ZN(_04957_));
 NAND2_X1 _22361_ (.A1(_16314_),
    .A2(_04957_),
    .ZN(_04958_));
 MUX2_X1 _22362_ (.A(_04601_),
    .B(_15928_),
    .S(_16310_),
    .Z(_04959_));
 OAI21_X4 _22363_ (.A(_04958_),
    .B1(_04959_),
    .B2(_04600_),
    .ZN(_04960_));
 INV_X1 _22364_ (.A(\cs_registers_i.csr_mtvec_o[9] ),
    .ZN(_04961_));
 OAI221_X1 _22365_ (.A(_04944_),
    .B1(_04960_),
    .B2(_04491_),
    .C1(_04493_),
    .C2(_04961_),
    .ZN(_01208_));
 NOR3_X4 _22366_ (.A1(_10882_),
    .A2(_03686_),
    .A3(_03747_),
    .ZN(_04962_));
 NAND3_X1 _22367_ (.A1(_03701_),
    .A2(_03689_),
    .A3(_04962_),
    .ZN(_04963_));
 MUX2_X1 _22368_ (.A(_03745_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .S(_04963_),
    .Z(_01209_));
 BUF_X4 _22369_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Z(_04964_));
 NOR2_X1 _22370_ (.A1(_04964_),
    .A2(_03702_),
    .ZN(_04965_));
 NOR4_X1 _22371_ (.A1(_03734_),
    .A2(_03701_),
    .A3(_03683_),
    .A4(_15940_),
    .ZN(_04966_));
 AOI21_X1 _22372_ (.A(_04965_),
    .B1(_04966_),
    .B2(_03702_),
    .ZN(_01210_));
 CLKBUF_X3 _22373_ (.A(_15943_),
    .Z(_04967_));
 BUF_X4 _22374_ (.A(_04967_),
    .Z(_04968_));
 NOR3_X1 _22375_ (.A1(_03734_),
    .A2(_03701_),
    .A3(_03683_),
    .ZN(_04969_));
 NAND2_X1 _22376_ (.A1(_04968_),
    .A2(_04969_),
    .ZN(_04970_));
 MUX2_X1 _22377_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(_04970_),
    .S(_03702_),
    .Z(_01211_));
 NOR2_X1 _22378_ (.A1(_03695_),
    .A2(_03702_),
    .ZN(_04971_));
 BUF_X4 _22379_ (.A(_00066_),
    .Z(_04972_));
 XNOR2_X2 _22380_ (.A(_15944_),
    .B(_04972_),
    .ZN(_04973_));
 NOR4_X1 _22381_ (.A1(_03734_),
    .A2(_03701_),
    .A3(_03683_),
    .A4(_04973_),
    .ZN(_04974_));
 AOI21_X1 _22382_ (.A(_04971_),
    .B1(_04974_),
    .B2(_03702_),
    .ZN(_01212_));
 NOR2_X1 _22383_ (.A1(_03694_),
    .A2(_03702_),
    .ZN(_04975_));
 BUF_X4 _22384_ (.A(_00067_),
    .Z(_04976_));
 NOR3_X2 _22385_ (.A1(_03695_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A3(_04964_),
    .ZN(_04977_));
 XNOR2_X2 _22386_ (.A(_04976_),
    .B(_04977_),
    .ZN(_04978_));
 NOR4_X1 _22387_ (.A1(_03734_),
    .A2(_03701_),
    .A3(_03683_),
    .A4(_04978_),
    .ZN(_04979_));
 AOI21_X1 _22388_ (.A(_04975_),
    .B1(_04979_),
    .B2(_03702_),
    .ZN(_01213_));
 NAND2_X1 _22389_ (.A1(_15944_),
    .A2(_03696_),
    .ZN(_04980_));
 XNOR2_X1 _22390_ (.A(_01162_),
    .B(_04980_),
    .ZN(_04981_));
 AND3_X1 _22391_ (.A1(_03689_),
    .A2(_04969_),
    .A3(_04981_),
    .ZN(_04982_));
 INV_X1 _22392_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .ZN(_04983_));
 AOI21_X1 _22393_ (.A(_04982_),
    .B1(_03740_),
    .B2(_04983_),
    .ZN(_01214_));
 MUX2_X1 _22394_ (.A(_03796_),
    .B(_03786_),
    .S(_03930_),
    .Z(_04984_));
 NOR2_X2 _22395_ (.A1(_04185_),
    .A2(_03740_),
    .ZN(_04985_));
 CLKBUF_X3 _22396_ (.A(_04985_),
    .Z(_04986_));
 MUX2_X1 _22397_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .B(_04984_),
    .S(_04986_),
    .Z(_01215_));
 MUX2_X1 _22398_ (.A(_03889_),
    .B(\alu_adder_result_ex[10] ),
    .S(_03930_),
    .Z(_04987_));
 MUX2_X1 _22399_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .B(_04987_),
    .S(_04986_),
    .Z(_01216_));
 MUX2_X1 _22400_ (.A(_03896_),
    .B(net486),
    .S(_03930_),
    .Z(_04988_));
 MUX2_X1 _22401_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .B(_04988_),
    .S(_04986_),
    .Z(_01217_));
 MUX2_X1 _22402_ (.A(_03905_),
    .B(\alu_adder_result_ex[12] ),
    .S(_03930_),
    .Z(_04989_));
 MUX2_X1 _22403_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .B(_04989_),
    .S(_04986_),
    .Z(_01218_));
 MUX2_X1 _22404_ (.A(_03914_),
    .B(\alu_adder_result_ex[13] ),
    .S(_03930_),
    .Z(_04990_));
 MUX2_X1 _22405_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .B(_04990_),
    .S(_04986_),
    .Z(_01219_));
 MUX2_X1 _22406_ (.A(_03921_),
    .B(net7),
    .S(_03930_),
    .Z(_04991_));
 MUX2_X1 _22407_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .B(_04991_),
    .S(_04986_),
    .Z(_01220_));
 MUX2_X1 _22408_ (.A(_03928_),
    .B(net437),
    .S(_03930_),
    .Z(_04992_));
 MUX2_X1 _22409_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .B(_04992_),
    .S(_04986_),
    .Z(_01221_));
 CLKBUF_X3 _22410_ (.A(_03760_),
    .Z(_04993_));
 MUX2_X1 _22411_ (.A(_04344_),
    .B(\alu_adder_result_ex[16] ),
    .S(_04993_),
    .Z(_04994_));
 MUX2_X1 _22412_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .B(_04994_),
    .S(_04986_),
    .Z(_01222_));
 MUX2_X1 _22413_ (.A(_03812_),
    .B(\alu_adder_result_ex[17] ),
    .S(_04993_),
    .Z(_04995_));
 CLKBUF_X3 _22414_ (.A(_04985_),
    .Z(_04996_));
 MUX2_X1 _22415_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .B(_04995_),
    .S(_04996_),
    .Z(_01223_));
 MUX2_X1 _22416_ (.A(_03822_),
    .B(\alu_adder_result_ex[18] ),
    .S(_04993_),
    .Z(_04997_));
 MUX2_X1 _22417_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .B(_04997_),
    .S(_04996_),
    .Z(_01224_));
 MUX2_X1 _22418_ (.A(_03828_),
    .B(\alu_adder_result_ex[19] ),
    .S(_04993_),
    .Z(_04998_));
 MUX2_X1 _22419_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .B(_04998_),
    .S(_04996_),
    .Z(_01225_));
 MUX2_X1 _22420_ (.A(_03811_),
    .B(\alu_adder_result_ex[1] ),
    .S(_04993_),
    .Z(_04999_));
 MUX2_X1 _22421_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .B(_04999_),
    .S(_04996_),
    .Z(_01226_));
 MUX2_X1 _22422_ (.A(_03836_),
    .B(\alu_adder_result_ex[20] ),
    .S(_04993_),
    .Z(_05000_));
 MUX2_X1 _22423_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .B(_05000_),
    .S(_04996_),
    .Z(_01227_));
 MUX2_X1 _22424_ (.A(_03846_),
    .B(\alu_adder_result_ex[21] ),
    .S(_04993_),
    .Z(_05001_));
 MUX2_X1 _22425_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .B(_05001_),
    .S(_04996_),
    .Z(_01228_));
 MUX2_X1 _22426_ (.A(_03855_),
    .B(\alu_adder_result_ex[22] ),
    .S(_04993_),
    .Z(_05002_));
 MUX2_X1 _22427_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .B(_05002_),
    .S(_04996_),
    .Z(_01229_));
 MUX2_X1 _22428_ (.A(_03862_),
    .B(net356),
    .S(_04993_),
    .Z(_05003_));
 MUX2_X1 _22429_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .B(_05003_),
    .S(_04996_),
    .Z(_01230_));
 MUX2_X1 _22430_ (.A(_03873_),
    .B(\alu_adder_result_ex[24] ),
    .S(_04993_),
    .Z(_05004_));
 MUX2_X1 _22431_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .B(_05004_),
    .S(_04996_),
    .Z(_01231_));
 CLKBUF_X3 _22432_ (.A(_03760_),
    .Z(_05005_));
 MUX2_X1 _22433_ (.A(_03881_),
    .B(net389),
    .S(_05005_),
    .Z(_05006_));
 MUX2_X1 _22434_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .B(_05006_),
    .S(_04996_),
    .Z(_01232_));
 NOR2_X1 _22435_ (.A1(_13686_),
    .A2(_03930_),
    .ZN(_05007_));
 AOI21_X1 _22436_ (.A(_05007_),
    .B1(_03930_),
    .B2(net392),
    .ZN(_05008_));
 CLKBUF_X3 _22437_ (.A(_04985_),
    .Z(_05009_));
 MUX2_X1 _22438_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .B(_05008_),
    .S(_05009_),
    .Z(_01233_));
 MUX2_X1 _22439_ (.A(_03139_),
    .B(\alu_adder_result_ex[27] ),
    .S(_05005_),
    .Z(_05010_));
 MUX2_X1 _22440_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .B(_05010_),
    .S(_05009_),
    .Z(_01234_));
 MUX2_X1 _22441_ (.A(_03906_),
    .B(net386),
    .S(_05005_),
    .Z(_05011_));
 MUX2_X1 _22442_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .B(_05011_),
    .S(_05009_),
    .Z(_01235_));
 MUX2_X1 _22443_ (.A(_03915_),
    .B(net411),
    .S(_05005_),
    .Z(_05012_));
 MUX2_X1 _22444_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .B(_05012_),
    .S(_05009_),
    .Z(_01236_));
 MUX2_X1 _22445_ (.A(_03820_),
    .B(\alu_adder_result_ex[2] ),
    .S(_05005_),
    .Z(_05013_));
 MUX2_X1 _22446_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .B(_05013_),
    .S(_05009_),
    .Z(_01237_));
 MUX2_X1 _22447_ (.A(_03922_),
    .B(net346),
    .S(_05005_),
    .Z(_05014_));
 MUX2_X1 _22448_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .B(_05014_),
    .S(_05009_),
    .Z(_01238_));
 OR2_X1 _22449_ (.A1(net289),
    .A2(_03757_),
    .ZN(_05015_));
 NAND3_X1 _22450_ (.A1(_03488_),
    .A2(_04986_),
    .A3(_05015_),
    .ZN(_05016_));
 INV_X1 _22451_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .ZN(_05017_));
 OAI21_X1 _22452_ (.A(_05016_),
    .B1(_04986_),
    .B2(_05017_),
    .ZN(_01239_));
 MUX2_X1 _22453_ (.A(_11967_),
    .B(\alu_adder_result_ex[3] ),
    .S(_05005_),
    .Z(_05018_));
 MUX2_X1 _22454_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .B(_05018_),
    .S(_05009_),
    .Z(_01240_));
 MUX2_X1 _22455_ (.A(_12008_),
    .B(\alu_adder_result_ex[4] ),
    .S(_05005_),
    .Z(_05019_));
 MUX2_X1 _22456_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .B(_05019_),
    .S(_05009_),
    .Z(_01241_));
 MUX2_X1 _22457_ (.A(_12051_),
    .B(\alu_adder_result_ex[5] ),
    .S(_05005_),
    .Z(_05020_));
 MUX2_X1 _22458_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .B(_05020_),
    .S(_05009_),
    .Z(_01242_));
 MUX2_X1 _22459_ (.A(_03854_),
    .B(net8),
    .S(_05005_),
    .Z(_05021_));
 MUX2_X1 _22460_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .B(_05021_),
    .S(_05009_),
    .Z(_01243_));
 MUX2_X1 _22461_ (.A(_03861_),
    .B(\alu_adder_result_ex[7] ),
    .S(_03760_),
    .Z(_05022_));
 MUX2_X1 _22462_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .B(_05022_),
    .S(_04985_),
    .Z(_01244_));
 MUX2_X1 _22463_ (.A(_03872_),
    .B(\alu_adder_result_ex[8] ),
    .S(_03760_),
    .Z(_05023_));
 MUX2_X1 _22464_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .B(_05023_),
    .S(_04985_),
    .Z(_01245_));
 MUX2_X1 _22465_ (.A(_03880_),
    .B(\alu_adder_result_ex[9] ),
    .S(_03760_),
    .Z(_05024_));
 MUX2_X1 _22466_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .B(_05024_),
    .S(_04985_),
    .Z(_01246_));
 NAND2_X2 _22467_ (.A1(_03784_),
    .A2(_03689_),
    .ZN(_05025_));
 CLKBUF_X3 _22468_ (.A(_05025_),
    .Z(_05026_));
 INV_X1 _22469_ (.A(_00068_),
    .ZN(_05027_));
 BUF_X4 _22470_ (.A(_15942_),
    .Z(_05028_));
 XOR2_X1 _22471_ (.A(_03499_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .Z(_05029_));
 AND2_X1 _22472_ (.A1(_03503_),
    .A2(_05029_),
    .ZN(_05030_));
 INV_X1 _22473_ (.A(_05029_),
    .ZN(_05031_));
 AOI21_X4 _22474_ (.A(_05030_),
    .B1(_05031_),
    .B2(net288),
    .ZN(_05032_));
 BUF_X4 _22475_ (.A(_05032_),
    .Z(_05033_));
 NAND2_X4 _22476_ (.A1(_01162_),
    .A2(_05033_),
    .ZN(_05034_));
 NOR3_X4 _22477_ (.A1(_03694_),
    .A2(_03695_),
    .A3(_05034_),
    .ZN(_05035_));
 AOI21_X2 _22478_ (.A(_05027_),
    .B1(_05028_),
    .B2(_05035_),
    .ZN(_05036_));
 AOI21_X2 _22479_ (.A(_03740_),
    .B1(_03735_),
    .B2(_03700_),
    .ZN(_05037_));
 INV_X1 _22480_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .ZN(_05038_));
 OAI22_X1 _22481_ (.A1(_05026_),
    .A2(_05036_),
    .B1(_05037_),
    .B2(_05038_),
    .ZN(_01247_));
 INV_X1 _22482_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .ZN(_05039_));
 CLKBUF_X3 _22483_ (.A(_05037_),
    .Z(_05040_));
 INV_X1 _22484_ (.A(_00078_),
    .ZN(_05041_));
 BUF_X4 _22485_ (.A(_15946_),
    .Z(_05042_));
 NOR3_X4 _22486_ (.A1(_03695_),
    .A2(_04976_),
    .A3(_05034_),
    .ZN(_05043_));
 AOI21_X2 _22487_ (.A(_05041_),
    .B1(_05042_),
    .B2(_05043_),
    .ZN(_05044_));
 OAI22_X1 _22488_ (.A1(_05039_),
    .A2(_05040_),
    .B1(_05044_),
    .B2(_05026_),
    .ZN(_01248_));
 INV_X1 _22489_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .ZN(_05045_));
 INV_X1 _22490_ (.A(_00079_),
    .ZN(_05046_));
 BUF_X4 _22491_ (.A(_15950_),
    .Z(_05047_));
 AOI21_X2 _22492_ (.A(_05046_),
    .B1(_05047_),
    .B2(_05043_),
    .ZN(_05048_));
 OAI22_X1 _22493_ (.A1(_05045_),
    .A2(_05040_),
    .B1(_05048_),
    .B2(_05026_),
    .ZN(_01249_));
 INV_X1 _22494_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .ZN(_05049_));
 INV_X1 _22495_ (.A(_00080_),
    .ZN(_05050_));
 NOR3_X4 _22496_ (.A1(_04972_),
    .A2(_04976_),
    .A3(_05034_),
    .ZN(_05051_));
 AOI21_X2 _22497_ (.A(_05050_),
    .B1(_05028_),
    .B2(_05051_),
    .ZN(_05052_));
 OAI22_X1 _22498_ (.A1(_05049_),
    .A2(_05040_),
    .B1(_05052_),
    .B2(_05026_),
    .ZN(_01250_));
 INV_X1 _22499_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .ZN(_05053_));
 INV_X1 _22500_ (.A(_00081_),
    .ZN(_05054_));
 AOI21_X2 _22501_ (.A(_05054_),
    .B1(_03693_),
    .B2(_05051_),
    .ZN(_05055_));
 OAI22_X1 _22502_ (.A1(_05053_),
    .A2(_05040_),
    .B1(_05055_),
    .B2(_05026_),
    .ZN(_01251_));
 INV_X1 _22503_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .ZN(_05056_));
 INV_X1 _22504_ (.A(_00082_),
    .ZN(_05057_));
 AOI21_X2 _22505_ (.A(_05057_),
    .B1(_05042_),
    .B2(_05051_),
    .ZN(_05058_));
 OAI22_X1 _22506_ (.A1(_05056_),
    .A2(_05040_),
    .B1(_05058_),
    .B2(_05026_),
    .ZN(_01252_));
 INV_X1 _22507_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .ZN(_05059_));
 INV_X1 _22508_ (.A(_00083_),
    .ZN(_05060_));
 AOI21_X2 _22509_ (.A(_05060_),
    .B1(_05047_),
    .B2(_05051_),
    .ZN(_05061_));
 OAI22_X1 _22510_ (.A1(_05059_),
    .A2(_05040_),
    .B1(_05061_),
    .B2(_05026_),
    .ZN(_01253_));
 INV_X1 _22511_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .ZN(_05062_));
 INV_X1 _22512_ (.A(_00084_),
    .ZN(_05063_));
 NAND2_X2 _22513_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_05032_),
    .ZN(_05064_));
 NOR3_X4 _22514_ (.A1(_03694_),
    .A2(_03695_),
    .A3(_05064_),
    .ZN(_05065_));
 AOI21_X2 _22515_ (.A(_05063_),
    .B1(_05028_),
    .B2(_05065_),
    .ZN(_05066_));
 OAI22_X1 _22516_ (.A1(_05062_),
    .A2(_05040_),
    .B1(_05066_),
    .B2(_05026_),
    .ZN(_01254_));
 INV_X1 _22517_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .ZN(_05067_));
 INV_X1 _22518_ (.A(_00085_),
    .ZN(_05068_));
 AOI21_X2 _22519_ (.A(_05068_),
    .B1(_03693_),
    .B2(_05065_),
    .ZN(_05069_));
 OAI22_X1 _22520_ (.A1(_05067_),
    .A2(_05040_),
    .B1(_05069_),
    .B2(_05026_),
    .ZN(_01255_));
 INV_X1 _22521_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .ZN(_05070_));
 INV_X1 _22522_ (.A(_00086_),
    .ZN(_05071_));
 AOI21_X2 _22523_ (.A(_05071_),
    .B1(_05042_),
    .B2(_05065_),
    .ZN(_05072_));
 OAI22_X1 _22524_ (.A1(_05070_),
    .A2(_05040_),
    .B1(_05072_),
    .B2(_05026_),
    .ZN(_01256_));
 INV_X1 _22525_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .ZN(_05073_));
 INV_X1 _22526_ (.A(_00087_),
    .ZN(_05074_));
 AOI21_X2 _22527_ (.A(_05074_),
    .B1(_05047_),
    .B2(_05065_),
    .ZN(_05075_));
 CLKBUF_X3 _22528_ (.A(_05025_),
    .Z(_05076_));
 OAI22_X1 _22529_ (.A1(_05073_),
    .A2(_05040_),
    .B1(_05075_),
    .B2(_05076_),
    .ZN(_01257_));
 INV_X1 _22530_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .ZN(_05077_));
 CLKBUF_X3 _22531_ (.A(_05037_),
    .Z(_05078_));
 INV_X1 _22532_ (.A(_00069_),
    .ZN(_05079_));
 AOI21_X1 _22533_ (.A(_05079_),
    .B1(_03697_),
    .B2(_05033_),
    .ZN(_05080_));
 OAI22_X1 _22534_ (.A1(_05077_),
    .A2(_05078_),
    .B1(_05080_),
    .B2(_05076_),
    .ZN(_01258_));
 INV_X1 _22535_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .ZN(_05081_));
 INV_X1 _22536_ (.A(_00088_),
    .ZN(_05082_));
 NOR3_X2 _22537_ (.A1(_03694_),
    .A2(_04972_),
    .A3(_05064_),
    .ZN(_05083_));
 AOI21_X1 _22538_ (.A(_05082_),
    .B1(_05028_),
    .B2(_05083_),
    .ZN(_05084_));
 OAI22_X1 _22539_ (.A1(_05081_),
    .A2(_05078_),
    .B1(_05084_),
    .B2(_05076_),
    .ZN(_01259_));
 INV_X1 _22540_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .ZN(_05085_));
 INV_X1 _22541_ (.A(_00089_),
    .ZN(_05086_));
 AOI21_X1 _22542_ (.A(_05086_),
    .B1(_03693_),
    .B2(_05083_),
    .ZN(_05087_));
 OAI22_X1 _22543_ (.A1(_05085_),
    .A2(_05078_),
    .B1(_05087_),
    .B2(_05076_),
    .ZN(_01260_));
 INV_X1 _22544_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .ZN(_05088_));
 INV_X1 _22545_ (.A(_00090_),
    .ZN(_05089_));
 AOI21_X1 _22546_ (.A(_05089_),
    .B1(_05042_),
    .B2(_05083_),
    .ZN(_05090_));
 OAI22_X1 _22547_ (.A1(_05088_),
    .A2(_05078_),
    .B1(_05090_),
    .B2(_05076_),
    .ZN(_01261_));
 INV_X1 _22548_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .ZN(_05091_));
 INV_X1 _22549_ (.A(_00091_),
    .ZN(_05092_));
 AOI21_X1 _22550_ (.A(_05092_),
    .B1(_05047_),
    .B2(_05083_),
    .ZN(_05093_));
 OAI22_X1 _22551_ (.A1(_05091_),
    .A2(_05078_),
    .B1(_05093_),
    .B2(_05076_),
    .ZN(_01262_));
 INV_X1 _22552_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .ZN(_05094_));
 INV_X1 _22553_ (.A(_00092_),
    .ZN(_05095_));
 NOR3_X4 _22554_ (.A1(_03695_),
    .A2(_04976_),
    .A3(_05064_),
    .ZN(_05096_));
 AOI21_X2 _22555_ (.A(_05095_),
    .B1(_05028_),
    .B2(_05096_),
    .ZN(_05097_));
 OAI22_X1 _22556_ (.A1(_05094_),
    .A2(_05078_),
    .B1(_05097_),
    .B2(_05076_),
    .ZN(_01263_));
 INV_X1 _22557_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .ZN(_05098_));
 INV_X1 _22558_ (.A(_00093_),
    .ZN(_05099_));
 AOI21_X2 _22559_ (.A(_05099_),
    .B1(_03693_),
    .B2(_05096_),
    .ZN(_05100_));
 OAI22_X1 _22560_ (.A1(_05098_),
    .A2(_05078_),
    .B1(_05100_),
    .B2(_05076_),
    .ZN(_01264_));
 INV_X1 _22561_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .ZN(_05101_));
 INV_X1 _22562_ (.A(_00094_),
    .ZN(_05102_));
 AOI21_X2 _22563_ (.A(_05102_),
    .B1(_05042_),
    .B2(_05096_),
    .ZN(_05103_));
 OAI22_X1 _22564_ (.A1(_05101_),
    .A2(_05078_),
    .B1(_05103_),
    .B2(_05076_),
    .ZN(_01265_));
 INV_X1 _22565_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .ZN(_05104_));
 INV_X1 _22566_ (.A(_00095_),
    .ZN(_05105_));
 AOI21_X1 _22567_ (.A(_05105_),
    .B1(_05047_),
    .B2(_05096_),
    .ZN(_05106_));
 OAI22_X1 _22568_ (.A1(_05104_),
    .A2(_05078_),
    .B1(_05106_),
    .B2(_05076_),
    .ZN(_01266_));
 INV_X1 _22569_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .ZN(_05107_));
 INV_X1 _22570_ (.A(_00096_),
    .ZN(_05108_));
 MUX2_X1 _22571_ (.A(_03503_),
    .B(_03517_),
    .S(_05031_),
    .Z(_05109_));
 BUF_X4 _22572_ (.A(_05109_),
    .Z(_05110_));
 NOR4_X4 _22573_ (.A1(_04972_),
    .A2(_04976_),
    .A3(_04983_),
    .A4(_05110_),
    .ZN(_05111_));
 AOI21_X2 _22574_ (.A(_05108_),
    .B1(_05028_),
    .B2(_05111_),
    .ZN(_05112_));
 CLKBUF_X3 _22575_ (.A(_05025_),
    .Z(_05113_));
 OAI22_X1 _22576_ (.A1(_05107_),
    .A2(_05078_),
    .B1(_05112_),
    .B2(_05113_),
    .ZN(_01267_));
 INV_X1 _22577_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .ZN(_05114_));
 CLKBUF_X3 _22578_ (.A(_05037_),
    .Z(_05115_));
 INV_X1 _22579_ (.A(_00097_),
    .ZN(_05116_));
 AOI21_X2 _22580_ (.A(_05116_),
    .B1(_03693_),
    .B2(_05111_),
    .ZN(_05117_));
 OAI22_X1 _22581_ (.A1(_05114_),
    .A2(_05115_),
    .B1(_05117_),
    .B2(_05113_),
    .ZN(_01268_));
 INV_X1 _22582_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .ZN(_05118_));
 INV_X1 _22583_ (.A(_00070_),
    .ZN(_05119_));
 AOI21_X2 _22584_ (.A(_05119_),
    .B1(_05042_),
    .B2(_05035_),
    .ZN(_05120_));
 OAI22_X1 _22585_ (.A1(_05118_),
    .A2(_05115_),
    .B1(_05120_),
    .B2(_05113_),
    .ZN(_01269_));
 INV_X1 _22586_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .ZN(_05121_));
 INV_X1 _22587_ (.A(_00098_),
    .ZN(_05122_));
 AOI21_X2 _22588_ (.A(_05122_),
    .B1(_05042_),
    .B2(_05111_),
    .ZN(_05123_));
 OAI22_X1 _22589_ (.A1(_05121_),
    .A2(_05115_),
    .B1(_05123_),
    .B2(_05113_),
    .ZN(_01270_));
 INV_X1 _22590_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .ZN(_05124_));
 INV_X1 _22591_ (.A(_00099_),
    .ZN(_05125_));
 AND2_X1 _22592_ (.A1(_05047_),
    .A2(_05111_),
    .ZN(_05126_));
 NOR2_X1 _22593_ (.A1(_05125_),
    .A2(_05126_),
    .ZN(_05127_));
 OAI22_X1 _22594_ (.A1(_05124_),
    .A2(_05115_),
    .B1(_05127_),
    .B2(_05113_),
    .ZN(_01271_));
 INV_X1 _22595_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .ZN(_05128_));
 INV_X1 _22596_ (.A(_00071_),
    .ZN(_05129_));
 AOI21_X2 _22597_ (.A(_05129_),
    .B1(_05047_),
    .B2(_05035_),
    .ZN(_05130_));
 OAI22_X1 _22598_ (.A1(_05128_),
    .A2(_05115_),
    .B1(_05130_),
    .B2(_05113_),
    .ZN(_01272_));
 INV_X1 _22599_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .ZN(_05131_));
 INV_X1 _22600_ (.A(_00072_),
    .ZN(_05132_));
 NOR3_X4 _22601_ (.A1(_03694_),
    .A2(_04972_),
    .A3(_05034_),
    .ZN(_05133_));
 AOI21_X2 _22602_ (.A(_05132_),
    .B1(_05028_),
    .B2(_05133_),
    .ZN(_05134_));
 OAI22_X1 _22603_ (.A1(_05131_),
    .A2(_05115_),
    .B1(_05134_),
    .B2(_05113_),
    .ZN(_01273_));
 INV_X1 _22604_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .ZN(_05135_));
 INV_X1 _22605_ (.A(_00073_),
    .ZN(_05136_));
 AOI21_X2 _22606_ (.A(_05136_),
    .B1(_03693_),
    .B2(_05133_),
    .ZN(_05137_));
 OAI22_X1 _22607_ (.A1(_05135_),
    .A2(_05115_),
    .B1(_05137_),
    .B2(_05113_),
    .ZN(_01274_));
 INV_X1 _22608_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .ZN(_05138_));
 INV_X1 _22609_ (.A(_00074_),
    .ZN(_05139_));
 AOI21_X2 _22610_ (.A(_05139_),
    .B1(_05042_),
    .B2(_05133_),
    .ZN(_05140_));
 OAI22_X1 _22611_ (.A1(_05138_),
    .A2(_05115_),
    .B1(_05140_),
    .B2(_05113_),
    .ZN(_01275_));
 INV_X1 _22612_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .ZN(_05141_));
 INV_X1 _22613_ (.A(_00075_),
    .ZN(_05142_));
 AOI21_X2 _22614_ (.A(_05142_),
    .B1(_05047_),
    .B2(_05133_),
    .ZN(_05143_));
 OAI22_X1 _22615_ (.A1(_05141_),
    .A2(_05115_),
    .B1(_05143_),
    .B2(_05113_),
    .ZN(_01276_));
 INV_X1 _22616_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .ZN(_05144_));
 INV_X1 _22617_ (.A(_00076_),
    .ZN(_05145_));
 AOI21_X2 _22618_ (.A(_05145_),
    .B1(_05028_),
    .B2(_05043_),
    .ZN(_05146_));
 OAI22_X1 _22619_ (.A1(_05144_),
    .A2(_05115_),
    .B1(_05146_),
    .B2(_05025_),
    .ZN(_01277_));
 INV_X1 _22620_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .ZN(_05147_));
 INV_X1 _22621_ (.A(_00077_),
    .ZN(_05148_));
 AOI21_X2 _22622_ (.A(_05148_),
    .B1(_03693_),
    .B2(_05043_),
    .ZN(_05149_));
 OAI22_X1 _22623_ (.A1(_05147_),
    .A2(_05037_),
    .B1(_05149_),
    .B2(_05025_),
    .ZN(_01278_));
 OR2_X1 _22624_ (.A1(fetch_enable_q),
    .A2(net60),
    .ZN(_01279_));
 OR3_X2 _22625_ (.A1(_03776_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A3(_03750_),
    .ZN(_05150_));
 NAND2_X1 _22626_ (.A1(_15955_),
    .A2(_05150_),
    .ZN(_05151_));
 OAI21_X2 _22627_ (.A(_05151_),
    .B1(_05150_),
    .B2(_00217_),
    .ZN(_05152_));
 OAI221_X2 _22628_ (.A(_12276_),
    .B1(_03737_),
    .B2(_05152_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .C2(_10912_),
    .ZN(_05153_));
 NAND2_X1 _22629_ (.A1(_10973_),
    .A2(_05153_),
    .ZN(_05154_));
 NAND2_X4 _22630_ (.A1(_11874_),
    .A2(_11924_),
    .ZN(_05155_));
 NAND2_X2 _22631_ (.A1(_11897_),
    .A2(_11921_),
    .ZN(_05156_));
 CLKBUF_X2 _22632_ (.A(_15761_),
    .Z(_05157_));
 BUF_X4 _22633_ (.A(_05157_),
    .Z(_05158_));
 AOI21_X2 _22634_ (.A(_05158_),
    .B1(_11926_),
    .B2(_11916_),
    .ZN(_05159_));
 AOI21_X4 _22635_ (.A(_05155_),
    .B1(_05156_),
    .B2(_05159_),
    .ZN(_05160_));
 BUF_X4 _22636_ (.A(_05160_),
    .Z(_05161_));
 AND3_X2 _22637_ (.A1(_05158_),
    .A2(_11903_),
    .A3(_11924_),
    .ZN(_05162_));
 BUF_X4 _22638_ (.A(_05162_),
    .Z(_05163_));
 OR3_X1 _22639_ (.A1(_11883_),
    .A2(_11885_),
    .A3(_11922_),
    .ZN(_05164_));
 NAND2_X1 _22640_ (.A1(_11926_),
    .A2(_05164_),
    .ZN(_05165_));
 CLKBUF_X3 _22641_ (.A(_15764_),
    .Z(_05166_));
 NOR2_X2 _22642_ (.A1(_10910_),
    .A2(_11875_),
    .ZN(_05167_));
 AOI22_X1 _22643_ (.A1(_05166_),
    .A2(_05167_),
    .B1(_05164_),
    .B2(_05158_),
    .ZN(_05168_));
 NAND2_X1 _22644_ (.A1(_05167_),
    .A2(_11921_),
    .ZN(_05169_));
 INV_X1 _22645_ (.A(_11897_),
    .ZN(_05170_));
 OAI221_X1 _22646_ (.A(_05165_),
    .B1(_05168_),
    .B2(_11921_),
    .C1(_05169_),
    .C2(_05170_),
    .ZN(_05171_));
 NAND2_X1 _22647_ (.A1(_11874_),
    .A2(_05171_),
    .ZN(_05172_));
 INV_X1 _22648_ (.A(_05166_),
    .ZN(_05173_));
 NAND2_X4 _22649_ (.A1(_11903_),
    .A2(_11921_),
    .ZN(_05174_));
 OR2_X1 _22650_ (.A1(_05158_),
    .A2(_11926_),
    .ZN(_05175_));
 NOR2_X1 _22651_ (.A1(_11897_),
    .A2(_05175_),
    .ZN(_05176_));
 NAND2_X1 _22652_ (.A1(_11874_),
    .A2(_11916_),
    .ZN(_05177_));
 OAI22_X1 _22653_ (.A1(_05173_),
    .A2(_05174_),
    .B1(_05176_),
    .B2(_05177_),
    .ZN(_05178_));
 NAND2_X1 _22654_ (.A1(_11919_),
    .A2(_05178_),
    .ZN(_05179_));
 NAND2_X2 _22655_ (.A1(_05172_),
    .A2(_05179_),
    .ZN(_05180_));
 NAND2_X1 _22656_ (.A1(_05174_),
    .A2(_05177_),
    .ZN(_05181_));
 AOI221_X2 _22657_ (.A(_05166_),
    .B1(_11926_),
    .B2(_11921_),
    .C1(_05181_),
    .C2(_11897_),
    .ZN(_05182_));
 NOR4_X4 _22658_ (.A1(_10943_),
    .A2(_11883_),
    .A3(_11885_),
    .A4(_05182_),
    .ZN(_05183_));
 NOR4_X4 _22659_ (.A1(_05161_),
    .A2(_05163_),
    .A3(_05180_),
    .A4(_05183_),
    .ZN(_05184_));
 NOR2_X4 _22660_ (.A1(_12276_),
    .A2(_05184_),
    .ZN(_05185_));
 NOR2_X1 _22661_ (.A1(_05154_),
    .A2(_05185_),
    .ZN(_05186_));
 NOR2_X2 _22662_ (.A1(_11874_),
    .A2(_11916_),
    .ZN(_05187_));
 NAND3_X1 _22663_ (.A1(_11919_),
    .A2(_05187_),
    .A3(_05175_),
    .ZN(_05188_));
 NAND2_X1 _22664_ (.A1(_05172_),
    .A2(_05188_),
    .ZN(_05189_));
 MUX2_X1 _22665_ (.A(_05166_),
    .B(_05175_),
    .S(_11874_),
    .Z(_05190_));
 AOI22_X1 _22666_ (.A1(_11897_),
    .A2(_05187_),
    .B1(_05190_),
    .B2(_11916_),
    .ZN(_05191_));
 NOR2_X1 _22667_ (.A1(_11876_),
    .A2(_05191_),
    .ZN(_05192_));
 AOI22_X1 _22668_ (.A1(_11897_),
    .A2(_11921_),
    .B1(_05181_),
    .B2(_11926_),
    .ZN(_05193_));
 OAI22_X2 _22669_ (.A1(_11903_),
    .A2(_05165_),
    .B1(_05193_),
    .B2(_11876_),
    .ZN(_05194_));
 XNOR2_X1 _22670_ (.A(_15894_),
    .B(_05194_),
    .ZN(_05195_));
 NAND2_X1 _22671_ (.A1(_15896_),
    .A2(_05195_),
    .ZN(_05196_));
 OAI21_X1 _22672_ (.A(_05196_),
    .B1(net313),
    .B2(_15896_),
    .ZN(_05197_));
 MUX2_X1 _22673_ (.A(_05189_),
    .B(_05192_),
    .S(_05197_),
    .Z(_05198_));
 AND3_X1 _22674_ (.A1(_05166_),
    .A2(_11919_),
    .A3(_05187_),
    .ZN(_05199_));
 NOR3_X2 _22675_ (.A1(_05192_),
    .A2(_05189_),
    .A3(_05199_),
    .ZN(_05200_));
 MUX2_X1 _22676_ (.A(_05199_),
    .B(_05200_),
    .S(_03745_),
    .Z(_05201_));
 OAI21_X1 _22677_ (.A(_05180_),
    .B1(_05198_),
    .B2(_05201_),
    .ZN(_05202_));
 NOR2_X1 _22678_ (.A1(_11897_),
    .A2(_05166_),
    .ZN(_05203_));
 OR3_X4 _22679_ (.A1(_11921_),
    .A2(_05155_),
    .A3(_05203_),
    .ZN(_05204_));
 NAND2_X1 _22680_ (.A1(_05158_),
    .A2(_11916_),
    .ZN(_05205_));
 AOI21_X2 _22681_ (.A(_05155_),
    .B1(_05156_),
    .B2(_05205_),
    .ZN(_05206_));
 OR2_X2 _22682_ (.A1(_05204_),
    .A2(_05206_),
    .ZN(_05207_));
 NOR2_X1 _22683_ (.A1(_16244_),
    .A2(_05207_),
    .ZN(_05208_));
 BUF_X4 _22684_ (.A(_05206_),
    .Z(_05209_));
 AOI21_X1 _22685_ (.A(_05208_),
    .B1(_05209_),
    .B2(_16240_),
    .ZN(_05210_));
 OAI21_X1 _22686_ (.A(_05160_),
    .B1(_05209_),
    .B2(_16241_),
    .ZN(_05211_));
 NAND2_X1 _22687_ (.A1(_05204_),
    .A2(_05211_),
    .ZN(_05212_));
 NOR2_X1 _22688_ (.A1(_05166_),
    .A2(_11926_),
    .ZN(_05213_));
 NOR3_X4 _22689_ (.A1(_11916_),
    .A2(_05155_),
    .A3(_05213_),
    .ZN(_05214_));
 AOI221_X2 _22690_ (.A(_05154_),
    .B1(_05210_),
    .B2(_05212_),
    .C1(_05214_),
    .C2(_03786_),
    .ZN(_05215_));
 AND4_X2 _22691_ (.A1(_10806_),
    .A2(_10868_),
    .A3(_11169_),
    .A4(_11379_),
    .ZN(_05216_));
 NOR2_X2 _22692_ (.A1(_10824_),
    .A2(_05216_),
    .ZN(_05217_));
 XNOR2_X2 _22693_ (.A(_16266_),
    .B(_05217_),
    .ZN(_05218_));
 INV_X1 _22694_ (.A(_16237_),
    .ZN(_05219_));
 OAI21_X2 _22695_ (.A(_10847_),
    .B1(_04512_),
    .B2(_05219_),
    .ZN(_05220_));
 XNOR2_X2 _22696_ (.A(_16270_),
    .B(_05220_),
    .ZN(_05221_));
 NOR2_X4 _22697_ (.A1(_05218_),
    .A2(_05221_),
    .ZN(_05222_));
 MUX2_X2 _22698_ (.A(_15894_),
    .B(_16239_),
    .S(_05158_),
    .Z(_05223_));
 NAND3_X2 _22699_ (.A1(_05166_),
    .A2(_10910_),
    .A3(_05187_),
    .ZN(_05224_));
 NOR2_X4 _22700_ (.A1(_05223_),
    .A2(_05224_),
    .ZN(_05225_));
 INV_X1 _22701_ (.A(_05225_),
    .ZN(_05226_));
 NOR2_X1 _22702_ (.A1(_05222_),
    .A2(_05226_),
    .ZN(_05227_));
 NOR2_X2 _22703_ (.A1(_16237_),
    .A2(_10824_),
    .ZN(_05228_));
 XNOR2_X2 _22704_ (.A(_11379_),
    .B(_05228_),
    .ZN(_05229_));
 AOI21_X1 _22705_ (.A(_11136_),
    .B1(_10774_),
    .B2(_10855_),
    .ZN(_05230_));
 AND4_X1 _22706_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_10774_),
    .A3(_10855_),
    .A4(_10859_),
    .ZN(_05231_));
 OAI21_X1 _22707_ (.A(_10865_),
    .B1(_05230_),
    .B2(_05231_),
    .ZN(_05232_));
 NAND3_X1 _22708_ (.A1(_10862_),
    .A2(_11486_),
    .A3(_11487_),
    .ZN(_05233_));
 AOI221_X2 _22709_ (.A(_10847_),
    .B1(_05232_),
    .B2(_05233_),
    .C1(_10804_),
    .C2(_10838_),
    .ZN(_05234_));
 NAND2_X1 _22710_ (.A1(_16238_),
    .A2(_10847_),
    .ZN(_05235_));
 NAND2_X1 _22711_ (.A1(_10824_),
    .A2(_11168_),
    .ZN(_05236_));
 OAI21_X4 _22712_ (.A(_05235_),
    .B1(_05236_),
    .B2(net301),
    .ZN(_05237_));
 OR2_X2 _22713_ (.A1(_05234_),
    .A2(_05237_),
    .ZN(_05238_));
 CLKBUF_X3 _22714_ (.A(_05238_),
    .Z(_05239_));
 CLKBUF_X3 _22715_ (.A(_05239_),
    .Z(_05240_));
 NOR2_X2 _22716_ (.A1(_05229_),
    .A2(_05240_),
    .ZN(_05241_));
 NOR2_X2 _22717_ (.A1(_05241_),
    .A2(_05225_),
    .ZN(_05242_));
 NAND4_X4 _22718_ (.A1(_05157_),
    .A2(_10910_),
    .A3(_11903_),
    .A4(_11921_),
    .ZN(_05243_));
 CLKBUF_X3 _22719_ (.A(_05243_),
    .Z(_05244_));
 MUX2_X1 _22720_ (.A(_16239_),
    .B(_15894_),
    .S(_05244_),
    .Z(_05245_));
 AOI21_X1 _22721_ (.A(_05245_),
    .B1(_05224_),
    .B2(_11170_),
    .ZN(_05246_));
 INV_X1 _22722_ (.A(_05246_),
    .ZN(_05247_));
 XNOR2_X2 _22723_ (.A(_16253_),
    .B(_05228_),
    .ZN(_05248_));
 BUF_X4 _22724_ (.A(_05248_),
    .Z(_05249_));
 AOI21_X4 _22725_ (.A(_05242_),
    .B1(_05247_),
    .B2(_05249_),
    .ZN(_05250_));
 AOI21_X1 _22726_ (.A(_05227_),
    .B1(_05250_),
    .B2(_05222_),
    .ZN(_05251_));
 NAND3_X4 _22727_ (.A1(_05158_),
    .A2(_11903_),
    .A3(_11924_),
    .ZN(_05252_));
 OAI21_X1 _22728_ (.A(_05215_),
    .B1(_05251_),
    .B2(_05252_),
    .ZN(_05253_));
 NOR3_X2 _22729_ (.A1(_11897_),
    .A2(_05166_),
    .A3(_11926_),
    .ZN(_05254_));
 OR4_X2 _22730_ (.A1(_05158_),
    .A2(_10943_),
    .A3(_05174_),
    .A4(_05254_),
    .ZN(_05255_));
 BUF_X4 _22731_ (.A(_05255_),
    .Z(_05256_));
 NOR2_X4 _22732_ (.A1(_05256_),
    .A2(_05221_),
    .ZN(_05257_));
 AND4_X2 _22733_ (.A1(_05157_),
    .A2(_10910_),
    .A3(_11903_),
    .A4(_11921_),
    .ZN(_05258_));
 MUX2_X1 _22734_ (.A(_16273_),
    .B(_16457_),
    .S(_05258_),
    .Z(_05259_));
 CLKBUF_X3 _22735_ (.A(_05258_),
    .Z(_05260_));
 MUX2_X1 _22736_ (.A(_16289_),
    .B(_16441_),
    .S(_05260_),
    .Z(_05261_));
 MUX2_X1 _22737_ (.A(_05259_),
    .B(_05261_),
    .S(_05239_),
    .Z(_05262_));
 INV_X1 _22738_ (.A(_05262_),
    .ZN(_05263_));
 NAND3_X4 _22739_ (.A1(_05158_),
    .A2(_11903_),
    .A3(_11924_),
    .ZN(_05264_));
 MUX2_X1 _22740_ (.A(_16445_),
    .B(_16277_),
    .S(_05264_),
    .Z(_05265_));
 MUX2_X1 _22741_ (.A(_16293_),
    .B(_16429_),
    .S(_05260_),
    .Z(_05266_));
 MUX2_X1 _22742_ (.A(_05265_),
    .B(_05266_),
    .S(_05239_),
    .Z(_05267_));
 MUX2_X1 _22743_ (.A(_05263_),
    .B(_05267_),
    .S(_11170_),
    .Z(_05268_));
 NOR2_X4 _22744_ (.A1(_05234_),
    .A2(_05237_),
    .ZN(_05269_));
 BUF_X4 _22745_ (.A(_05269_),
    .Z(_05270_));
 BUF_X4 _22746_ (.A(_05270_),
    .Z(_05271_));
 BUF_X4 _22747_ (.A(_05258_),
    .Z(_05272_));
 NOR2_X1 _22748_ (.A1(_16254_),
    .A2(_05272_),
    .ZN(_05273_));
 BUF_X4 _22749_ (.A(_05244_),
    .Z(_05274_));
 OAI21_X1 _22750_ (.A(_11172_),
    .B1(_16469_),
    .B2(_05274_),
    .ZN(_05275_));
 NAND2_X1 _22751_ (.A1(_16465_),
    .A2(_05162_),
    .ZN(_05276_));
 OAI21_X1 _22752_ (.A(_05276_),
    .B1(_05272_),
    .B2(_16261_),
    .ZN(_05277_));
 OAI22_X1 _22753_ (.A1(_05273_),
    .A2(_05275_),
    .B1(_05277_),
    .B2(_11172_),
    .ZN(_05278_));
 NOR2_X1 _22754_ (.A1(_05271_),
    .A2(_05278_),
    .ZN(_05279_));
 MUX2_X1 _22755_ (.A(_16250_),
    .B(_16478_),
    .S(_05272_),
    .Z(_05280_));
 MUX2_X1 _22756_ (.A(_16239_),
    .B(_15894_),
    .S(_05162_),
    .Z(_05281_));
 MUX2_X1 _22757_ (.A(_05280_),
    .B(_05281_),
    .S(_11172_),
    .Z(_05282_));
 AOI21_X1 _22758_ (.A(_05279_),
    .B1(_05282_),
    .B2(_05271_),
    .ZN(_05283_));
 MUX2_X1 _22759_ (.A(_05268_),
    .B(_05283_),
    .S(_05248_),
    .Z(_05284_));
 MUX2_X1 _22760_ (.A(_16333_),
    .B(_16389_),
    .S(_05258_),
    .Z(_05285_));
 MUX2_X1 _22761_ (.A(_16354_),
    .B(_16373_),
    .S(_05258_),
    .Z(_05286_));
 MUX2_X1 _22762_ (.A(_05285_),
    .B(_05286_),
    .S(_05239_),
    .Z(_05287_));
 MUX2_X1 _22763_ (.A(_16346_),
    .B(_16381_),
    .S(_05260_),
    .Z(_05288_));
 MUX2_X1 _22764_ (.A(_16362_),
    .B(_16365_),
    .S(_05260_),
    .Z(_05289_));
 MUX2_X1 _22765_ (.A(_05288_),
    .B(_05289_),
    .S(_05239_),
    .Z(_05290_));
 MUX2_X1 _22766_ (.A(_05287_),
    .B(_05290_),
    .S(_11170_),
    .Z(_05291_));
 MUX2_X1 _22767_ (.A(_16302_),
    .B(_16421_),
    .S(_05260_),
    .Z(_05292_));
 MUX2_X1 _22768_ (.A(_16317_),
    .B(_16410_),
    .S(_05260_),
    .Z(_05293_));
 MUX2_X1 _22769_ (.A(_05292_),
    .B(_05293_),
    .S(_05239_),
    .Z(_05294_));
 NOR2_X1 _22770_ (.A1(_11170_),
    .A2(_05294_),
    .ZN(_05295_));
 MUX2_X1 _22771_ (.A(_16329_),
    .B(_16398_),
    .S(_05260_),
    .Z(_05296_));
 NOR2_X1 _22772_ (.A1(_05270_),
    .A2(_05296_),
    .ZN(_05297_));
 MUX2_X1 _22773_ (.A(_16310_),
    .B(_16418_),
    .S(_05260_),
    .Z(_05298_));
 AOI21_X2 _22774_ (.A(_05297_),
    .B1(_05298_),
    .B2(_05271_),
    .ZN(_05299_));
 AOI21_X1 _22775_ (.A(_05295_),
    .B1(_05299_),
    .B2(_11171_),
    .ZN(_05300_));
 MUX2_X1 _22776_ (.A(_05291_),
    .B(_05300_),
    .S(_05248_),
    .Z(_05301_));
 MUX2_X1 _22777_ (.A(_05284_),
    .B(_05301_),
    .S(_05218_),
    .Z(_05302_));
 XNOR2_X2 _22778_ (.A(_11478_),
    .B(_05220_),
    .ZN(_05303_));
 NOR2_X4 _22779_ (.A1(_05255_),
    .A2(_05303_),
    .ZN(_05304_));
 XNOR2_X2 _22780_ (.A(_16262_),
    .B(_05217_),
    .ZN(_05305_));
 MUX2_X1 _22781_ (.A(_16325_),
    .B(_16402_),
    .S(_05243_),
    .Z(_05306_));
 MUX2_X1 _22782_ (.A(_16310_),
    .B(_16418_),
    .S(_05243_),
    .Z(_05307_));
 MUX2_X1 _22783_ (.A(_05306_),
    .B(_05307_),
    .S(_05238_),
    .Z(_05308_));
 MUX2_X1 _22784_ (.A(_16317_),
    .B(_16410_),
    .S(_05243_),
    .Z(_05309_));
 MUX2_X1 _22785_ (.A(_16302_),
    .B(_16421_),
    .S(_05243_),
    .Z(_05310_));
 MUX2_X1 _22786_ (.A(_05309_),
    .B(_05310_),
    .S(_05239_),
    .Z(_05311_));
 MUX2_X1 _22787_ (.A(_05308_),
    .B(_05311_),
    .S(_11170_),
    .Z(_05312_));
 NAND2_X1 _22788_ (.A1(_05305_),
    .A2(_05312_),
    .ZN(_05313_));
 MUX2_X1 _22789_ (.A(_16254_),
    .B(_16469_),
    .S(_05244_),
    .Z(_05314_));
 NAND2_X1 _22790_ (.A1(_05271_),
    .A2(_05314_),
    .ZN(_05315_));
 OR2_X1 _22791_ (.A1(_05270_),
    .A2(_05245_),
    .ZN(_05316_));
 AOI21_X2 _22792_ (.A(_11173_),
    .B1(_05315_),
    .B2(_05316_),
    .ZN(_05317_));
 MUX2_X1 _22793_ (.A(_16461_),
    .B(_16482_),
    .S(_05238_),
    .Z(_05318_));
 MUX2_X1 _22794_ (.A(_16246_),
    .B(_16261_),
    .S(_05269_),
    .Z(_05319_));
 MUX2_X2 _22795_ (.A(_05318_),
    .B(_05319_),
    .S(_05272_),
    .Z(_05320_));
 AOI21_X4 _22796_ (.A(_05317_),
    .B1(_05320_),
    .B2(_11173_),
    .ZN(_05321_));
 OAI21_X1 _22797_ (.A(_05313_),
    .B1(_05321_),
    .B2(_05305_),
    .ZN(_05322_));
 MUX2_X1 _22798_ (.A(_16354_),
    .B(_16373_),
    .S(_05243_),
    .Z(_05323_));
 MUX2_X1 _22799_ (.A(_16333_),
    .B(_16389_),
    .S(_05243_),
    .Z(_05324_));
 MUX2_X1 _22800_ (.A(_05323_),
    .B(_05324_),
    .S(_05238_),
    .Z(_05325_));
 MUX2_X1 _22801_ (.A(_16362_),
    .B(_16365_),
    .S(_05243_),
    .Z(_05326_));
 MUX2_X1 _22802_ (.A(_16346_),
    .B(_16381_),
    .S(_05244_),
    .Z(_05327_));
 MUX2_X1 _22803_ (.A(_05326_),
    .B(_05327_),
    .S(_05239_),
    .Z(_05328_));
 MUX2_X1 _22804_ (.A(_05325_),
    .B(_05328_),
    .S(_11172_),
    .Z(_05329_));
 MUX2_X1 _22805_ (.A(_16281_),
    .B(_16449_),
    .S(_05244_),
    .Z(_05330_));
 MUX2_X1 _22806_ (.A(_16297_),
    .B(_16433_),
    .S(_05244_),
    .Z(_05331_));
 MUX2_X1 _22807_ (.A(_05330_),
    .B(_05331_),
    .S(_05269_),
    .Z(_05332_));
 NAND2_X1 _22808_ (.A1(_16457_),
    .A2(_05274_),
    .ZN(_05333_));
 OAI221_X2 _22809_ (.A(_05333_),
    .B1(_05237_),
    .B2(_05234_),
    .C1(_16269_),
    .C2(_05274_),
    .ZN(_05334_));
 MUX2_X1 _22810_ (.A(_16285_),
    .B(_16437_),
    .S(_05244_),
    .Z(_05335_));
 AOI21_X1 _22811_ (.A(_11172_),
    .B1(_05270_),
    .B2(_05335_),
    .ZN(_05336_));
 AOI22_X2 _22812_ (.A1(_11172_),
    .A2(_05332_),
    .B1(_05334_),
    .B2(_05336_),
    .ZN(_05337_));
 MUX2_X1 _22813_ (.A(_05329_),
    .B(_05337_),
    .S(_05218_),
    .Z(_05338_));
 BUF_X4 _22814_ (.A(_05249_),
    .Z(_05339_));
 MUX2_X2 _22815_ (.A(_05322_),
    .B(_05338_),
    .S(_05339_),
    .Z(_05340_));
 AOI221_X2 _22816_ (.A(_05253_),
    .B1(_05257_),
    .B2(_05302_),
    .C1(_05304_),
    .C2(_05340_),
    .ZN(_05341_));
 INV_X1 _22817_ (.A(_04589_),
    .ZN(_05342_));
 NOR2_X2 _22818_ (.A1(_04489_),
    .A2(_05342_),
    .ZN(_05343_));
 INV_X1 _22819_ (.A(_00552_),
    .ZN(_05344_));
 INV_X1 _22820_ (.A(_00553_),
    .ZN(_05345_));
 AOI22_X4 _22821_ (.A1(_05344_),
    .A2(_04388_),
    .B1(_04391_),
    .B2(_05345_),
    .ZN(_05346_));
 BUF_X2 _22822_ (.A(\cs_registers_i.mhpmcounter[2][32] ),
    .Z(_05347_));
 AOI22_X4 _22823_ (.A1(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .A2(_04388_),
    .B1(_04391_),
    .B2(_05347_),
    .ZN(_05348_));
 OAI22_X4 _22824_ (.A1(_04608_),
    .A2(_05346_),
    .B1(_05348_),
    .B2(_04380_),
    .ZN(_05349_));
 AOI22_X2 _22825_ (.A1(net61),
    .A2(_04637_),
    .B1(_04426_),
    .B2(\cs_registers_i.dscratch1_q[0] ),
    .ZN(_05350_));
 AOI22_X2 _22826_ (.A1(\cs_registers_i.dscratch0_q[0] ),
    .A2(_04416_),
    .B1(_04918_),
    .B2(\cs_registers_i.mcause_q[0] ),
    .ZN(_05351_));
 NAND2_X1 _22827_ (.A1(\cs_registers_i.csr_mepc_o[0] ),
    .A2(_04423_),
    .ZN(_05352_));
 AOI222_X2 _22828_ (.A1(\cs_registers_i.mtval_q[0] ),
    .A2(_04413_),
    .B1(_04508_),
    .B2(\cs_registers_i.mscratch_q[0] ),
    .C1(_04433_),
    .C2(\cs_registers_i.dcsr_q[0] ),
    .ZN(_05353_));
 NAND4_X2 _22829_ (.A1(_05350_),
    .A2(_05351_),
    .A3(_05352_),
    .A4(_05353_),
    .ZN(_05354_));
 OAI21_X2 _22830_ (.A(_04461_),
    .B1(_04457_),
    .B2(_00554_),
    .ZN(_05355_));
 NOR4_X4 _22831_ (.A1(_05343_),
    .A2(_05349_),
    .A3(_05354_),
    .A4(_05355_),
    .ZN(_05356_));
 BUF_X4 _22832_ (.A(_11282_),
    .Z(_05357_));
 AOI221_X2 _22833_ (.A(_05186_),
    .B1(_05202_),
    .B2(_05341_),
    .C1(_05356_),
    .C2(_05357_),
    .ZN(_05358_));
 BUF_X2 _22834_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_05359_));
 BUF_X4 _22835_ (.A(_05359_),
    .Z(_05360_));
 BUF_X4 _22836_ (.A(_05360_),
    .Z(_05361_));
 CLKBUF_X2 _22837_ (.A(\load_store_unit_i.data_type_q[2] ),
    .Z(_05362_));
 BUF_X4 _22838_ (.A(_05362_),
    .Z(_05363_));
 CLKBUF_X3 _22839_ (.A(\load_store_unit_i.data_type_q[1] ),
    .Z(_05364_));
 OR2_X2 _22840_ (.A1(_05363_),
    .A2(_05364_),
    .ZN(_05365_));
 BUF_X4 _22841_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(_05366_));
 INV_X2 _22842_ (.A(_05366_),
    .ZN(_05367_));
 NOR2_X1 _22843_ (.A1(_05359_),
    .A2(_05367_),
    .ZN(_05368_));
 BUF_X4 _22844_ (.A(_05368_),
    .Z(_05369_));
 INV_X2 _22845_ (.A(_05359_),
    .ZN(_05370_));
 NOR2_X4 _22846_ (.A1(_05370_),
    .A2(_05366_),
    .ZN(_05371_));
 AOI221_X1 _22847_ (.A(_05365_),
    .B1(_05369_),
    .B2(\load_store_unit_i.rdata_q[16] ),
    .C1(_05371_),
    .C2(\load_store_unit_i.rdata_q[8] ),
    .ZN(_05372_));
 BUF_X4 _22848_ (.A(_05371_),
    .Z(_05373_));
 BUF_X1 _22849_ (.A(data_rdata_i[8]),
    .Z(_05374_));
 AOI22_X1 _22850_ (.A1(net36),
    .A2(_05369_),
    .B1(_05373_),
    .B2(_05374_),
    .ZN(_05375_));
 BUF_X4 _22851_ (.A(_05365_),
    .Z(_05376_));
 AOI21_X1 _22852_ (.A(_05372_),
    .B1(_05375_),
    .B2(_05376_),
    .ZN(_05377_));
 CLKBUF_X3 _22853_ (.A(_05367_),
    .Z(_05378_));
 BUF_X4 _22854_ (.A(_05364_),
    .Z(_05379_));
 INV_X1 _22855_ (.A(_05362_),
    .ZN(_05380_));
 NAND2_X4 _22856_ (.A1(_05380_),
    .A2(_05379_),
    .ZN(_05381_));
 AOI22_X1 _22857_ (.A1(_05379_),
    .A2(net45),
    .B1(_05381_),
    .B2(\load_store_unit_i.rdata_q[24] ),
    .ZN(_05382_));
 NOR2_X1 _22858_ (.A1(_05378_),
    .A2(_05382_),
    .ZN(_05383_));
 OAI21_X1 _22859_ (.A(_05361_),
    .B1(_05377_),
    .B2(_05383_),
    .ZN(_05384_));
 CLKBUF_X3 _22860_ (.A(_05366_),
    .Z(_05385_));
 CLKBUF_X3 _22861_ (.A(_05385_),
    .Z(_05386_));
 CLKBUF_X3 _22862_ (.A(_05386_),
    .Z(_05387_));
 CLKBUF_X3 _22863_ (.A(_05366_),
    .Z(_05388_));
 NOR2_X1 _22864_ (.A1(_05359_),
    .A2(_05388_),
    .ZN(_05389_));
 AOI22_X1 _22865_ (.A1(_05387_),
    .A2(_05377_),
    .B1(_05389_),
    .B2(net34),
    .ZN(_05390_));
 NAND2_X1 _22866_ (.A1(_05384_),
    .A2(_05390_),
    .ZN(_05391_));
 AND2_X1 _22867_ (.A1(_03751_),
    .A2(_03777_),
    .ZN(_05392_));
 NOR4_X4 _22868_ (.A1(_03776_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .A3(_11864_),
    .A4(_05392_),
    .ZN(_05393_));
 INV_X1 _22869_ (.A(_05393_),
    .ZN(_05394_));
 OAI33_X1 _22870_ (.A1(_10823_),
    .A2(_10824_),
    .A3(_10854_),
    .B1(_10962_),
    .B2(_10968_),
    .B3(net306),
    .ZN(_05395_));
 OAI21_X4 _22871_ (.A(_05394_),
    .B1(_05395_),
    .B2(net366),
    .ZN(_05396_));
 AOI21_X1 _22872_ (.A(_03565_),
    .B1(_04489_),
    .B2(_04488_),
    .ZN(_05397_));
 OR2_X1 _22873_ (.A1(_03646_),
    .A2(_03645_),
    .ZN(_05398_));
 AOI21_X2 _22874_ (.A(_03631_),
    .B1(_05397_),
    .B2(_05398_),
    .ZN(_05399_));
 OR3_X2 _22875_ (.A1(_03688_),
    .A2(_05396_),
    .A3(_05399_),
    .ZN(_05400_));
 BUF_X4 _22876_ (.A(_05400_),
    .Z(_05401_));
 MUX2_X2 _22877_ (.A(_05358_),
    .B(_05391_),
    .S(_05401_),
    .Z(_05402_));
 BUF_X2 _22878_ (.A(_05402_),
    .Z(_05403_));
 OAI221_X1 _22879_ (.A(_04530_),
    .B1(_04541_),
    .B2(_04540_),
    .C1(_03645_),
    .C2(_03646_),
    .ZN(_05404_));
 AOI211_X4 _22880_ (.A(_03688_),
    .B(_05396_),
    .C1(_05404_),
    .C2(_11329_),
    .ZN(_05405_));
 AND2_X1 _22881_ (.A1(_01159_),
    .A2(_03529_),
    .ZN(_05406_));
 INV_X2 _22882_ (.A(net59),
    .ZN(_05407_));
 NOR3_X4 _22883_ (.A1(_03523_),
    .A2(_05407_),
    .A3(_03526_),
    .ZN(_05408_));
 AOI21_X4 _22884_ (.A(_05405_),
    .B1(_05406_),
    .B2(_05408_),
    .ZN(_05409_));
 NOR3_X4 _22885_ (.A1(_10862_),
    .A2(_11307_),
    .A3(_05409_),
    .ZN(_05410_));
 AND2_X2 _22886_ (.A1(_11311_),
    .A2(_05410_),
    .ZN(_05411_));
 BUF_X4 _22887_ (.A(_05411_),
    .Z(_05412_));
 MUX2_X1 _22888_ (.A(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .B(_05403_),
    .S(_05412_),
    .Z(_01280_));
 BUF_X4 _22889_ (.A(_05401_),
    .Z(_05413_));
 AOI221_X1 _22890_ (.A(_05376_),
    .B1(_05369_),
    .B2(\load_store_unit_i.rdata_q[20] ),
    .C1(_05373_),
    .C2(\load_store_unit_i.rdata_q[12] ),
    .ZN(_05414_));
 BUF_X4 _22891_ (.A(_05360_),
    .Z(_05415_));
 CLKBUF_X3 _22892_ (.A(_05388_),
    .Z(_05416_));
 NAND2_X1 _22893_ (.A1(_05416_),
    .A2(net41),
    .ZN(_05417_));
 NOR2_X1 _22894_ (.A1(_05415_),
    .A2(_05417_),
    .ZN(_05418_));
 BUF_X1 _22895_ (.A(data_rdata_i[12]),
    .Z(_05419_));
 AOI21_X1 _22896_ (.A(_05418_),
    .B1(_05373_),
    .B2(_05419_),
    .ZN(_05420_));
 AOI21_X1 _22897_ (.A(_05414_),
    .B1(_05420_),
    .B2(_05376_),
    .ZN(_05421_));
 NAND2_X1 _22898_ (.A1(_05378_),
    .A2(net55),
    .ZN(_05422_));
 NAND2_X2 _22899_ (.A1(_05415_),
    .A2(_05387_),
    .ZN(_05423_));
 AOI22_X2 _22900_ (.A1(_05379_),
    .A2(net49),
    .B1(_05381_),
    .B2(\load_store_unit_i.rdata_q[28] ),
    .ZN(_05424_));
 OAI22_X2 _22901_ (.A1(_05361_),
    .A2(_05422_),
    .B1(_05423_),
    .B2(_05424_),
    .ZN(_05425_));
 OAI21_X2 _22902_ (.A(_05413_),
    .B1(_05421_),
    .B2(_05425_),
    .ZN(_05426_));
 BUF_X4 _22903_ (.A(_05185_),
    .Z(_05427_));
 CLKBUF_X3 _22904_ (.A(_05150_),
    .Z(_05428_));
 NAND2_X1 _22905_ (.A1(_15990_),
    .A2(_05428_),
    .ZN(_05429_));
 BUF_X4 _22906_ (.A(_05428_),
    .Z(_05430_));
 OAI21_X2 _22907_ (.A(_05429_),
    .B1(_05430_),
    .B2(_00560_),
    .ZN(_05431_));
 OAI221_X2 _22908_ (.A(_03755_),
    .B1(_03737_),
    .B2(_05431_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .C2(_10912_),
    .ZN(_05432_));
 NAND2_X1 _22909_ (.A1(_10973_),
    .A2(_05432_),
    .ZN(_05433_));
 OR2_X1 _22910_ (.A1(_05427_),
    .A2(_05433_),
    .ZN(_05434_));
 NOR4_X4 _22911_ (.A1(_05158_),
    .A2(_10943_),
    .A3(_05174_),
    .A4(_05254_),
    .ZN(_05435_));
 MUX2_X1 _22912_ (.A(_05329_),
    .B(_05291_),
    .S(_05248_),
    .Z(_05436_));
 CLKBUF_X3 _22913_ (.A(_05229_),
    .Z(_05437_));
 MUX2_X1 _22914_ (.A(_05268_),
    .B(_05300_),
    .S(_05437_),
    .Z(_05438_));
 CLKBUF_X3 _22915_ (.A(_05305_),
    .Z(_05439_));
 CLKBUF_X3 _22916_ (.A(_05439_),
    .Z(_05440_));
 MUX2_X1 _22917_ (.A(_05436_),
    .B(_05438_),
    .S(_05440_),
    .Z(_05441_));
 MUX2_X1 _22918_ (.A(_05312_),
    .B(_05337_),
    .S(_05229_),
    .Z(_05442_));
 NAND2_X1 _22919_ (.A1(_05437_),
    .A2(_05225_),
    .ZN(_05443_));
 OAI21_X1 _22920_ (.A(_05443_),
    .B1(_05321_),
    .B2(_05437_),
    .ZN(_05444_));
 BUF_X4 _22921_ (.A(_05218_),
    .Z(_05445_));
 MUX2_X1 _22922_ (.A(_05442_),
    .B(_05444_),
    .S(_05445_),
    .Z(_05446_));
 MUX2_X1 _22923_ (.A(_05441_),
    .B(_05446_),
    .S(_05221_),
    .Z(_05447_));
 AND2_X1 _22924_ (.A1(_05435_),
    .A2(_05447_),
    .ZN(_05448_));
 CLKBUF_X3 _22925_ (.A(_05207_),
    .Z(_05449_));
 CLKBUF_X3 _22926_ (.A(_05449_),
    .Z(_05450_));
 CLKBUF_X3 _22927_ (.A(_05450_),
    .Z(_05451_));
 NOR2_X1 _22928_ (.A1(_16271_),
    .A2(_05451_),
    .ZN(_05452_));
 CLKBUF_X3 _22929_ (.A(_05161_),
    .Z(_05453_));
 CLKBUF_X3 _22930_ (.A(_05453_),
    .Z(_05454_));
 BUF_X4 _22931_ (.A(_05209_),
    .Z(_05455_));
 BUF_X4 _22932_ (.A(_05455_),
    .Z(_05456_));
 OAI21_X1 _22933_ (.A(_05454_),
    .B1(_05456_),
    .B2(_16272_),
    .ZN(_05457_));
 BUF_X4 _22934_ (.A(_05204_),
    .Z(_05458_));
 BUF_X4 _22935_ (.A(_05458_),
    .Z(_05459_));
 BUF_X4 _22936_ (.A(_05459_),
    .Z(_05460_));
 BUF_X4 _22937_ (.A(_05455_),
    .Z(_05461_));
 BUF_X4 _22938_ (.A(_05461_),
    .Z(_05462_));
 AOI221_X2 _22939_ (.A(_05452_),
    .B1(_05457_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16275_),
    .ZN(_05463_));
 NOR2_X1 _22940_ (.A1(_05433_),
    .A2(_05463_),
    .ZN(_05464_));
 NAND2_X1 _22941_ (.A1(_05439_),
    .A2(_05303_),
    .ZN(_05465_));
 MUX2_X1 _22942_ (.A(_16453_),
    .B(_16469_),
    .S(_05238_),
    .Z(_05466_));
 MUX2_X1 _22943_ (.A(_16254_),
    .B(_16269_),
    .S(_05269_),
    .Z(_05467_));
 MUX2_X1 _22944_ (.A(_05466_),
    .B(_05467_),
    .S(_05272_),
    .Z(_05468_));
 MUX2_X1 _22945_ (.A(_05320_),
    .B(_05468_),
    .S(_11173_),
    .Z(_05469_));
 NOR2_X1 _22946_ (.A1(_05271_),
    .A2(_05225_),
    .ZN(_05470_));
 NOR2_X1 _22947_ (.A1(_05247_),
    .A2(_05470_),
    .ZN(_05471_));
 MUX2_X1 _22948_ (.A(_05469_),
    .B(_05471_),
    .S(_05437_),
    .Z(_05472_));
 NOR2_X2 _22949_ (.A1(_05465_),
    .A2(_05472_),
    .ZN(_05473_));
 BUF_X4 _22950_ (.A(_05225_),
    .Z(_05474_));
 OAI21_X1 _22951_ (.A(_05272_),
    .B1(_05222_),
    .B2(_05474_),
    .ZN(_05475_));
 BUF_X4 _22952_ (.A(_05214_),
    .Z(_05476_));
 BUF_X4 _22953_ (.A(_05476_),
    .Z(_05477_));
 INV_X1 _22954_ (.A(_05477_),
    .ZN(_05478_));
 OAI221_X2 _22955_ (.A(_05464_),
    .B1(_05473_),
    .B2(_05475_),
    .C1(_05478_),
    .C2(_03725_),
    .ZN(_05479_));
 AOI22_X1 _22956_ (.A1(\cs_registers_i.dscratch0_q[4] ),
    .A2(_04417_),
    .B1(_04559_),
    .B2(\cs_registers_i.mscratch_q[4] ),
    .ZN(_05480_));
 INV_X1 _22957_ (.A(_01166_),
    .ZN(_05481_));
 AOI22_X1 _22958_ (.A1(net87),
    .A2(_04442_),
    .B1(_04408_),
    .B2(_05481_),
    .ZN(_05482_));
 AOI222_X2 _22959_ (.A1(\cs_registers_i.mtval_q[4] ),
    .A2(_04414_),
    .B1(_04918_),
    .B2(\cs_registers_i.mcause_q[4] ),
    .C1(_04426_),
    .C2(\cs_registers_i.dscratch1_q[4] ),
    .ZN(_05483_));
 AOI21_X1 _22960_ (.A(_04545_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .ZN(_05484_));
 AND4_X1 _22961_ (.A1(_05480_),
    .A2(_05482_),
    .A3(_05483_),
    .A4(_05484_),
    .ZN(_05485_));
 AOI22_X2 _22962_ (.A1(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .A2(_04500_),
    .B1(_04501_),
    .B2(\cs_registers_i.mhpmcounter[2][4] ),
    .ZN(_05486_));
 AOI22_X2 _22963_ (.A1(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .A2(_04500_),
    .B1(_04501_),
    .B2(\cs_registers_i.mhpmcounter[2][36] ),
    .ZN(_05487_));
 OAI221_X2 _22964_ (.A(_05485_),
    .B1(_05486_),
    .B2(_04402_),
    .C1(_04498_),
    .C2(_05487_),
    .ZN(_05488_));
 CLKBUF_X3 _22965_ (.A(_10973_),
    .Z(_05489_));
 OAI221_X2 _22966_ (.A(_05434_),
    .B1(_05448_),
    .B2(_05479_),
    .C1(_05488_),
    .C2(_05489_),
    .ZN(_05490_));
 OAI21_X4 _22967_ (.A(_05426_),
    .B1(_05490_),
    .B2(_05413_),
    .ZN(_05491_));
 BUF_X2 _22968_ (.A(_05491_),
    .Z(_05492_));
 NAND2_X2 _22969_ (.A1(_11428_),
    .A2(_11309_),
    .ZN(_05493_));
 NOR2_X4 _22970_ (.A1(_11310_),
    .A2(_05493_),
    .ZN(_05494_));
 NOR3_X4 _22971_ (.A1(_10862_),
    .A2(_11306_),
    .A3(_05409_),
    .ZN(_05495_));
 AND2_X1 _22972_ (.A1(_05494_),
    .A2(_05495_),
    .ZN(_05496_));
 BUF_X4 _22973_ (.A(_05496_),
    .Z(_05497_));
 BUF_X4 _22974_ (.A(_05497_),
    .Z(_05498_));
 MUX2_X1 _22975_ (.A(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .B(_05492_),
    .S(_05498_),
    .Z(_01281_));
 NOR2_X4 _22976_ (.A1(_05363_),
    .A2(_05364_),
    .ZN(_05499_));
 BUF_X1 _22977_ (.A(data_rdata_i[13]),
    .Z(_05500_));
 INV_X1 _22978_ (.A(net42),
    .ZN(_05501_));
 NOR2_X1 _22979_ (.A1(_05367_),
    .A2(_05501_),
    .ZN(_05502_));
 BUF_X4 _22980_ (.A(_05370_),
    .Z(_05503_));
 AOI221_X2 _22981_ (.A(_05499_),
    .B1(_05373_),
    .B2(_05500_),
    .C1(_05502_),
    .C2(_05503_),
    .ZN(_05504_));
 AOI221_X2 _22982_ (.A(_05376_),
    .B1(_05369_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .C1(_05373_),
    .C2(\load_store_unit_i.rdata_q[13] ),
    .ZN(_05505_));
 AOI22_X2 _22983_ (.A1(_05379_),
    .A2(net50),
    .B1(_05381_),
    .B2(\load_store_unit_i.rdata_q[29] ),
    .ZN(_05506_));
 NAND2_X1 _22984_ (.A1(_05367_),
    .A2(net56),
    .ZN(_05507_));
 OAI222_X2 _22985_ (.A1(_05504_),
    .A2(_05505_),
    .B1(_05506_),
    .B2(_05423_),
    .C1(_05361_),
    .C2(_05507_),
    .ZN(_05508_));
 NAND2_X1 _22986_ (.A1(_14525_),
    .A2(_05428_),
    .ZN(_05509_));
 OAI21_X2 _22987_ (.A(_05509_),
    .B1(_05428_),
    .B2(_00561_),
    .ZN(_05510_));
 OAI221_X2 _22988_ (.A(_12276_),
    .B1(_03737_),
    .B2(_05510_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .C2(_10912_),
    .ZN(_05511_));
 NAND2_X1 _22989_ (.A1(_10973_),
    .A2(_05511_),
    .ZN(_05512_));
 INV_X1 _22990_ (.A(_01167_),
    .ZN(_05513_));
 AOI22_X1 _22991_ (.A1(net88),
    .A2(_04637_),
    .B1(_04407_),
    .B2(_05513_),
    .ZN(_05514_));
 AOI22_X1 _22992_ (.A1(\cs_registers_i.csr_mepc_o[5] ),
    .A2(_04423_),
    .B1(_04426_),
    .B2(\cs_registers_i.dscratch1_q[5] ),
    .ZN(_05515_));
 AOI22_X1 _22993_ (.A1(\cs_registers_i.dscratch0_q[5] ),
    .A2(_04416_),
    .B1(_04413_),
    .B2(\cs_registers_i.mtval_q[5] ),
    .ZN(_05516_));
 AOI21_X1 _22994_ (.A(_04544_),
    .B1(_04508_),
    .B2(\cs_registers_i.mscratch_q[5] ),
    .ZN(_05517_));
 AND4_X1 _22995_ (.A1(_05514_),
    .A2(_05515_),
    .A3(_05516_),
    .A4(_05517_),
    .ZN(_05518_));
 CLKBUF_X2 _22996_ (.A(\cs_registers_i.mhpmcounter[2][5] ),
    .Z(_05519_));
 AOI22_X2 _22997_ (.A1(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .A2(_04589_),
    .B1(_04591_),
    .B2(_05519_),
    .ZN(_05520_));
 BUF_X2 _22998_ (.A(\cs_registers_i.mhpmcounter[2][37] ),
    .Z(_05521_));
 AOI22_X2 _22999_ (.A1(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .A2(_04389_),
    .B1(_04393_),
    .B2(_05521_),
    .ZN(_05522_));
 OAI221_X2 _23000_ (.A(_05518_),
    .B1(_05520_),
    .B2(_04402_),
    .C1(_04381_),
    .C2(_05522_),
    .ZN(_05523_));
 OAI22_X1 _23001_ (.A1(_05427_),
    .A2(_05512_),
    .B1(_05523_),
    .B2(_05489_),
    .ZN(_05524_));
 MUX2_X1 _23002_ (.A(_16437_),
    .B(_16453_),
    .S(_05240_),
    .Z(_05525_));
 MUX2_X1 _23003_ (.A(_16269_),
    .B(_16285_),
    .S(_05270_),
    .Z(_05526_));
 MUX2_X1 _23004_ (.A(_05525_),
    .B(_05526_),
    .S(_05163_),
    .Z(_05527_));
 MUX2_X1 _23005_ (.A(_16445_),
    .B(_16461_),
    .S(_05239_),
    .Z(_05528_));
 MUX2_X1 _23006_ (.A(_16261_),
    .B(_16277_),
    .S(_05269_),
    .Z(_05529_));
 MUX2_X1 _23007_ (.A(_05528_),
    .B(_05529_),
    .S(_05272_),
    .Z(_05530_));
 MUX2_X2 _23008_ (.A(_05527_),
    .B(_05530_),
    .S(_16242_),
    .Z(_05531_));
 MUX2_X1 _23009_ (.A(_16293_),
    .B(_16429_),
    .S(_05244_),
    .Z(_05532_));
 MUX2_X1 _23010_ (.A(_05307_),
    .B(_05532_),
    .S(_05240_),
    .Z(_05533_));
 MUX2_X1 _23011_ (.A(_05311_),
    .B(_05533_),
    .S(_16242_),
    .Z(_05534_));
 MUX2_X1 _23012_ (.A(_05531_),
    .B(_05534_),
    .S(_05339_),
    .Z(_05535_));
 CLKBUF_X3 _23013_ (.A(_05339_),
    .Z(_05536_));
 MUX2_X1 _23014_ (.A(_16246_),
    .B(_16482_),
    .S(_05244_),
    .Z(_05537_));
 MUX2_X1 _23015_ (.A(_05314_),
    .B(_05537_),
    .S(_11170_),
    .Z(_05538_));
 MUX2_X2 _23016_ (.A(_05246_),
    .B(_05538_),
    .S(_05271_),
    .Z(_05539_));
 NAND2_X1 _23017_ (.A1(_05536_),
    .A2(_05539_),
    .ZN(_05540_));
 NAND2_X1 _23018_ (.A1(_05443_),
    .A2(_05540_),
    .ZN(_05541_));
 BUF_X4 _23019_ (.A(_05445_),
    .Z(_05542_));
 MUX2_X1 _23020_ (.A(_05535_),
    .B(_05541_),
    .S(_05542_),
    .Z(_05543_));
 NAND2_X1 _23021_ (.A1(_05304_),
    .A2(_05543_),
    .ZN(_05544_));
 OAI21_X1 _23022_ (.A(_05453_),
    .B1(_05455_),
    .B2(_16280_),
    .ZN(_05545_));
 NAND2_X1 _23023_ (.A1(_05459_),
    .A2(_05545_),
    .ZN(_05546_));
 NOR2_X1 _23024_ (.A1(_16279_),
    .A2(_05449_),
    .ZN(_05547_));
 BUF_X4 _23025_ (.A(_05209_),
    .Z(_05548_));
 BUF_X4 _23026_ (.A(_05548_),
    .Z(_05549_));
 AOI21_X2 _23027_ (.A(_05547_),
    .B1(_05549_),
    .B2(_16283_),
    .ZN(_05550_));
 AOI221_X2 _23028_ (.A(_05512_),
    .B1(_05546_),
    .B2(_05550_),
    .C1(\alu_adder_result_ex[5] ),
    .C2(_05476_),
    .ZN(_05551_));
 NAND3_X4 _23029_ (.A1(_05163_),
    .A2(_05221_),
    .A3(_05474_),
    .ZN(_05552_));
 NAND2_X1 _23030_ (.A1(_05551_),
    .A2(_05552_),
    .ZN(_05553_));
 NOR2_X2 _23031_ (.A1(_05439_),
    .A2(_05225_),
    .ZN(_05554_));
 NOR2_X1 _23032_ (.A1(_11172_),
    .A2(_05245_),
    .ZN(_05555_));
 AOI21_X2 _23033_ (.A(_05555_),
    .B1(_05537_),
    .B2(_11173_),
    .ZN(_05556_));
 AOI211_X2 _23034_ (.A(_05248_),
    .B(_05470_),
    .C1(_05556_),
    .C2(_05271_),
    .ZN(_05557_));
 MUX2_X2 _23035_ (.A(_05468_),
    .B(_05530_),
    .S(_11173_),
    .Z(_05558_));
 AOI21_X4 _23036_ (.A(_05557_),
    .B1(_05558_),
    .B2(_05249_),
    .ZN(_05559_));
 CLKBUF_X3 _23037_ (.A(_05440_),
    .Z(_05560_));
 AOI21_X2 _23038_ (.A(_05554_),
    .B1(_05559_),
    .B2(_05560_),
    .ZN(_05561_));
 NOR2_X4 _23039_ (.A1(_05274_),
    .A2(_05221_),
    .ZN(_05562_));
 NOR2_X1 _23040_ (.A1(_16242_),
    .A2(_05325_),
    .ZN(_05563_));
 MUX2_X1 _23041_ (.A(_16329_),
    .B(_16398_),
    .S(_05244_),
    .Z(_05564_));
 MUX2_X1 _23042_ (.A(_16342_),
    .B(_16385_),
    .S(_05274_),
    .Z(_05565_));
 MUX2_X1 _23043_ (.A(_05564_),
    .B(_05565_),
    .S(_05270_),
    .Z(_05566_));
 AOI21_X2 _23044_ (.A(_05563_),
    .B1(_05566_),
    .B2(_16242_),
    .ZN(_05567_));
 XNOR2_X1 _23045_ (.A(_11172_),
    .B(_05162_),
    .ZN(_05568_));
 MUX2_X1 _23046_ (.A(_16362_),
    .B(_16365_),
    .S(_05568_),
    .Z(_05569_));
 NAND2_X1 _23047_ (.A1(_05240_),
    .A2(_05569_),
    .ZN(_05570_));
 MUX2_X1 _23048_ (.A(_05286_),
    .B(_05288_),
    .S(_11172_),
    .Z(_05571_));
 NAND2_X1 _23049_ (.A1(_05271_),
    .A2(_05571_),
    .ZN(_05572_));
 NAND2_X1 _23050_ (.A1(_05570_),
    .A2(_05572_),
    .ZN(_05573_));
 MUX2_X1 _23051_ (.A(_05567_),
    .B(_05573_),
    .S(_05249_),
    .Z(_05574_));
 MUX2_X1 _23052_ (.A(_16337_),
    .B(_16393_),
    .S(_05260_),
    .Z(_05575_));
 MUX2_X1 _23053_ (.A(_16321_),
    .B(_16406_),
    .S(_05272_),
    .Z(_05576_));
 MUX2_X1 _23054_ (.A(_05575_),
    .B(_05576_),
    .S(_05270_),
    .Z(_05577_));
 AND2_X1 _23055_ (.A1(_11171_),
    .A2(_05577_),
    .ZN(_05578_));
 AOI21_X2 _23056_ (.A(_05578_),
    .B1(_05299_),
    .B2(_11173_),
    .ZN(_05579_));
 NAND2_X1 _23057_ (.A1(_05240_),
    .A2(_05292_),
    .ZN(_05580_));
 OAI21_X1 _23058_ (.A(_05580_),
    .B1(_05261_),
    .B2(_05240_),
    .ZN(_05581_));
 MUX2_X1 _23059_ (.A(_05267_),
    .B(_05581_),
    .S(_16242_),
    .Z(_05582_));
 MUX2_X1 _23060_ (.A(_05579_),
    .B(_05582_),
    .S(_05249_),
    .Z(_05583_));
 MUX2_X1 _23061_ (.A(_05574_),
    .B(_05583_),
    .S(_05440_),
    .Z(_05584_));
 BUF_X4 _23062_ (.A(_05257_),
    .Z(_05585_));
 AOI221_X2 _23063_ (.A(_05553_),
    .B1(_05561_),
    .B2(_05562_),
    .C1(_05584_),
    .C2(_05585_),
    .ZN(_05586_));
 AOI21_X1 _23064_ (.A(_05524_),
    .B1(_05544_),
    .B2(_05586_),
    .ZN(_05587_));
 BUF_X4 _23065_ (.A(_05405_),
    .Z(_05588_));
 MUX2_X2 _23066_ (.A(_05508_),
    .B(_05587_),
    .S(_05588_),
    .Z(_05589_));
 BUF_X2 _23067_ (.A(_05589_),
    .Z(_05590_));
 MUX2_X1 _23068_ (.A(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .B(_05590_),
    .S(_05498_),
    .Z(_01282_));
 BUF_X4 _23069_ (.A(_05495_),
    .Z(_05591_));
 NAND2_X2 _23070_ (.A1(_05494_),
    .A2(_05591_),
    .ZN(_05592_));
 CLKBUF_X3 _23071_ (.A(_05592_),
    .Z(_05593_));
 NAND2_X1 _23072_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .A2(_05593_),
    .ZN(_05594_));
 OR2_X1 _23073_ (.A1(_12276_),
    .A2(_05184_),
    .ZN(_05595_));
 BUF_X4 _23074_ (.A(_05595_),
    .Z(_05596_));
 XNOR2_X1 _23075_ (.A(_14524_),
    .B(_16021_),
    .ZN(_05597_));
 MUX2_X1 _23076_ (.A(_00562_),
    .B(_05597_),
    .S(_05428_),
    .Z(_05598_));
 INV_X1 _23077_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .ZN(_05599_));
 AOI221_X2 _23078_ (.A(_11865_),
    .B1(_03685_),
    .B2(_05598_),
    .C1(_05599_),
    .C2(net414),
    .ZN(_05600_));
 NOR2_X1 _23079_ (.A1(_11282_),
    .A2(_05600_),
    .ZN(_05601_));
 NAND2_X1 _23080_ (.A1(_05596_),
    .A2(_05601_),
    .ZN(_05602_));
 BUF_X2 _23081_ (.A(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .Z(_05603_));
 CLKBUF_X2 _23082_ (.A(\cs_registers_i.mhpmcounter[2][38] ),
    .Z(_05604_));
 AOI22_X2 _23083_ (.A1(_05603_),
    .A2(_04499_),
    .B1(_04392_),
    .B2(_05604_),
    .ZN(_05605_));
 BUF_X2 _23084_ (.A(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .Z(_05606_));
 AOI22_X2 _23085_ (.A1(_05606_),
    .A2(_04499_),
    .B1(_04392_),
    .B2(\cs_registers_i.mhpmcounter[2][6] ),
    .ZN(_05607_));
 OAI22_X2 _23086_ (.A1(_04380_),
    .A2(_05605_),
    .B1(_05607_),
    .B2(_04608_),
    .ZN(_05608_));
 NAND2_X2 _23087_ (.A1(_03636_),
    .A2(_04405_),
    .ZN(_05609_));
 NOR2_X1 _23088_ (.A1(_01168_),
    .A2(_05609_),
    .ZN(_05610_));
 AOI221_X2 _23089_ (.A(_05610_),
    .B1(_04413_),
    .B2(\cs_registers_i.mtval_q[6] ),
    .C1(\cs_registers_i.dscratch0_q[6] ),
    .C2(_04416_),
    .ZN(_05611_));
 AOI22_X2 _23090_ (.A1(\cs_registers_i.csr_mepc_o[6] ),
    .A2(_04423_),
    .B1(_04433_),
    .B2(\cs_registers_i.dcsr_q[6] ),
    .ZN(_05612_));
 AOI22_X1 _23091_ (.A1(net89),
    .A2(_04637_),
    .B1(_04427_),
    .B2(\cs_registers_i.dscratch1_q[6] ),
    .ZN(_05613_));
 NAND3_X1 _23092_ (.A1(_05611_),
    .A2(_05612_),
    .A3(_05613_),
    .ZN(_05614_));
 AND2_X1 _23093_ (.A1(\cs_registers_i.mscratch_q[6] ),
    .A2(_04509_),
    .ZN(_05615_));
 OR4_X4 _23094_ (.A1(_04545_),
    .A2(_05608_),
    .A3(_05614_),
    .A4(_05615_),
    .ZN(_05616_));
 OAI21_X2 _23095_ (.A(_05602_),
    .B1(_05616_),
    .B2(_05489_),
    .ZN(_05617_));
 NOR2_X1 _23096_ (.A1(_16287_),
    .A2(_05450_),
    .ZN(_05618_));
 OAI21_X1 _23097_ (.A(_05453_),
    .B1(_05549_),
    .B2(_16288_),
    .ZN(_05619_));
 AOI221_X2 _23098_ (.A(_05618_),
    .B1(_05619_),
    .B2(_05459_),
    .C1(_05456_),
    .C2(_16291_),
    .ZN(_05620_));
 AOI21_X1 _23099_ (.A(_05620_),
    .B1(_05477_),
    .B2(net8),
    .ZN(_05621_));
 AND2_X1 _23100_ (.A1(_05601_),
    .A2(_05621_),
    .ZN(_05622_));
 AND2_X1 _23101_ (.A1(_05437_),
    .A2(_05539_),
    .ZN(_05623_));
 AOI211_X2 _23102_ (.A(_05465_),
    .B(_05623_),
    .C1(_05531_),
    .C2(_05339_),
    .ZN(_05624_));
 OAI21_X1 _23103_ (.A(_05622_),
    .B1(_05624_),
    .B2(_05475_),
    .ZN(_05625_));
 AND2_X1 _23104_ (.A1(_11173_),
    .A2(_05577_),
    .ZN(_05626_));
 MUX2_X1 _23105_ (.A(_16342_),
    .B(_16385_),
    .S(_05260_),
    .Z(_05627_));
 MUX2_X1 _23106_ (.A(_05627_),
    .B(_05296_),
    .S(_05269_),
    .Z(_05628_));
 AND2_X1 _23107_ (.A1(_11171_),
    .A2(_05628_),
    .ZN(_05629_));
 OR3_X1 _23108_ (.A1(_05445_),
    .A2(_05626_),
    .A3(_05629_),
    .ZN(_05630_));
 MUX2_X1 _23109_ (.A(_16321_),
    .B(_16406_),
    .S(_05274_),
    .Z(_05631_));
 MUX2_X1 _23110_ (.A(_16337_),
    .B(_16393_),
    .S(_05274_),
    .Z(_05632_));
 MUX2_X1 _23111_ (.A(_05631_),
    .B(_05632_),
    .S(_05270_),
    .Z(_05633_));
 MUX2_X1 _23112_ (.A(_05566_),
    .B(_05633_),
    .S(_11171_),
    .Z(_05634_));
 OR2_X1 _23113_ (.A1(_05440_),
    .A2(_05634_),
    .ZN(_05635_));
 NAND2_X1 _23114_ (.A1(_05630_),
    .A2(_05635_),
    .ZN(_05636_));
 MUX2_X1 _23115_ (.A(_05266_),
    .B(_05298_),
    .S(_05240_),
    .Z(_05637_));
 MUX2_X1 _23116_ (.A(_05581_),
    .B(_05637_),
    .S(_11171_),
    .Z(_05638_));
 MUX2_X1 _23117_ (.A(_05323_),
    .B(_05289_),
    .S(_05269_),
    .Z(_05639_));
 MUX2_X1 _23118_ (.A(_05326_),
    .B(_05286_),
    .S(_05270_),
    .Z(_05640_));
 MUX2_X1 _23119_ (.A(_05639_),
    .B(_05640_),
    .S(_11173_),
    .Z(_05641_));
 MUX2_X1 _23120_ (.A(_05638_),
    .B(_05641_),
    .S(_05445_),
    .Z(_05642_));
 MUX2_X1 _23121_ (.A(_05636_),
    .B(_05642_),
    .S(_05536_),
    .Z(_05643_));
 AOI21_X2 _23122_ (.A(_05242_),
    .B1(_05556_),
    .B2(_05241_),
    .ZN(_05644_));
 NAND2_X1 _23123_ (.A1(_05542_),
    .A2(_05644_),
    .ZN(_05645_));
 MUX2_X1 _23124_ (.A(_05310_),
    .B(_05335_),
    .S(_05239_),
    .Z(_05646_));
 MUX2_X1 _23125_ (.A(_05533_),
    .B(_05646_),
    .S(_11171_),
    .Z(_05647_));
 AND2_X1 _23126_ (.A1(_05249_),
    .A2(_05647_),
    .ZN(_05648_));
 AOI21_X2 _23127_ (.A(_05648_),
    .B1(_05558_),
    .B2(_05437_),
    .ZN(_05649_));
 OAI21_X2 _23128_ (.A(_05645_),
    .B1(_05649_),
    .B2(_05542_),
    .ZN(_05650_));
 CLKBUF_X3 _23129_ (.A(_05221_),
    .Z(_05651_));
 MUX2_X1 _23130_ (.A(_05643_),
    .B(_05650_),
    .S(_05651_),
    .Z(_05652_));
 AOI21_X2 _23131_ (.A(_05625_),
    .B1(_05652_),
    .B2(_05435_),
    .ZN(_05653_));
 NOR3_X4 _23132_ (.A1(_05413_),
    .A2(_05617_),
    .A3(_05653_),
    .ZN(_05654_));
 INV_X1 _23133_ (.A(net43),
    .ZN(_05655_));
 NOR2_X1 _23134_ (.A1(_05378_),
    .A2(_05655_),
    .ZN(_05656_));
 AOI221_X2 _23135_ (.A(_05499_),
    .B1(_05373_),
    .B2(net35),
    .C1(_05656_),
    .C2(_05503_),
    .ZN(_05657_));
 AOI221_X2 _23136_ (.A(_05376_),
    .B1(_05369_),
    .B2(\load_store_unit_i.rdata_q[22] ),
    .C1(_05373_),
    .C2(\load_store_unit_i.rdata_q[14] ),
    .ZN(_05658_));
 AOI22_X2 _23137_ (.A1(_05379_),
    .A2(net52),
    .B1(_05381_),
    .B2(\load_store_unit_i.rdata_q[30] ),
    .ZN(_05659_));
 NAND2_X1 _23138_ (.A1(_05378_),
    .A2(net57),
    .ZN(_05660_));
 OAI222_X2 _23139_ (.A1(_05657_),
    .A2(_05658_),
    .B1(_05659_),
    .B2(_05423_),
    .C1(_05361_),
    .C2(_05660_),
    .ZN(_05661_));
 AOI21_X4 _23140_ (.A(_05654_),
    .B1(_05661_),
    .B2(_05413_),
    .ZN(_05662_));
 BUF_X4 _23141_ (.A(_05662_),
    .Z(_05663_));
 OAI21_X1 _23142_ (.A(_05594_),
    .B1(_05663_),
    .B2(_05593_),
    .ZN(_01283_));
 NOR3_X2 _23143_ (.A1(_03571_),
    .A2(_03688_),
    .A3(_05396_),
    .ZN(_05664_));
 NOR2_X1 _23144_ (.A1(_03646_),
    .A2(_03645_),
    .ZN(_05665_));
 NOR3_X2 _23145_ (.A1(_03688_),
    .A2(_05396_),
    .A3(_05665_),
    .ZN(_05666_));
 NOR2_X2 _23146_ (.A1(_03565_),
    .A2(_03644_),
    .ZN(_05667_));
 AOI21_X4 _23147_ (.A(_05664_),
    .B1(_05666_),
    .B2(_05667_),
    .ZN(_05668_));
 AND2_X1 _23148_ (.A1(\load_store_unit_i.rdata_q[23] ),
    .A2(_05499_),
    .ZN(_05669_));
 AOI21_X1 _23149_ (.A(_05669_),
    .B1(_05376_),
    .B2(net44),
    .ZN(_05670_));
 AOI21_X1 _23150_ (.A(_05503_),
    .B1(\load_store_unit_i.rdata_q[15] ),
    .B2(_05499_),
    .ZN(_05671_));
 OAI22_X2 _23151_ (.A1(_05360_),
    .A2(_05670_),
    .B1(_05671_),
    .B2(_05387_),
    .ZN(_05672_));
 OAI21_X1 _23152_ (.A(_05672_),
    .B1(net58),
    .B2(_05387_),
    .ZN(_05673_));
 BUF_X1 _23153_ (.A(data_rdata_i[15]),
    .Z(_05674_));
 NAND3_X1 _23154_ (.A1(_05367_),
    .A2(_05674_),
    .A3(_05376_),
    .ZN(_05675_));
 AND2_X1 _23155_ (.A1(_05364_),
    .A2(net53),
    .ZN(_05676_));
 OAI22_X1 _23156_ (.A1(net53),
    .A2(_05381_),
    .B1(_05676_),
    .B2(\load_store_unit_i.rdata_q[31] ),
    .ZN(_05677_));
 OAI21_X1 _23157_ (.A(_05675_),
    .B1(_05677_),
    .B2(_05378_),
    .ZN(_05678_));
 OAI21_X1 _23158_ (.A(_05361_),
    .B1(_05672_),
    .B2(_05678_),
    .ZN(_05679_));
 AND3_X1 _23159_ (.A1(_05668_),
    .A2(_05673_),
    .A3(_05679_),
    .ZN(_05680_));
 INV_X1 _23160_ (.A(_16033_),
    .ZN(_05681_));
 INV_X1 _23161_ (.A(_16020_),
    .ZN(_05682_));
 AOI21_X1 _23162_ (.A(_16001_),
    .B1(_16002_),
    .B2(_14521_),
    .ZN(_05683_));
 INV_X1 _23163_ (.A(_16021_),
    .ZN(_05684_));
 OAI21_X2 _23164_ (.A(_05682_),
    .B1(_05683_),
    .B2(_05684_),
    .ZN(_05685_));
 XNOR2_X2 _23165_ (.A(_05681_),
    .B(_05685_),
    .ZN(_05686_));
 NAND2_X1 _23166_ (.A1(_05430_),
    .A2(_05686_),
    .ZN(_05687_));
 OAI21_X2 _23167_ (.A(_05687_),
    .B1(_05430_),
    .B2(_00563_),
    .ZN(_05688_));
 OAI221_X2 _23168_ (.A(_03755_),
    .B1(_03737_),
    .B2(_05688_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .C2(_10912_),
    .ZN(_05689_));
 BUF_X2 _23169_ (.A(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .Z(_05690_));
 CLKBUF_X3 _23170_ (.A(\cs_registers_i.mhpmcounter[2][39] ),
    .Z(_05691_));
 AOI22_X4 _23171_ (.A1(_05690_),
    .A2(_04499_),
    .B1(_04392_),
    .B2(_05691_),
    .ZN(_05692_));
 BUF_X2 _23172_ (.A(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .Z(_05693_));
 BUF_X2 _23173_ (.A(\cs_registers_i.mhpmcounter[2][7] ),
    .Z(_05694_));
 AOI22_X4 _23174_ (.A1(_05693_),
    .A2(_04499_),
    .B1(_04392_),
    .B2(_05694_),
    .ZN(_05695_));
 OAI22_X4 _23175_ (.A1(_04380_),
    .A2(_05692_),
    .B1(_05695_),
    .B2(_04608_),
    .ZN(_05696_));
 AOI222_X2 _23176_ (.A1(\cs_registers_i.dscratch0_q[7] ),
    .A2(_04416_),
    .B1(_04423_),
    .B2(\cs_registers_i.csr_mepc_o[7] ),
    .C1(_04447_),
    .C2(\cs_registers_i.mie_q[16] ),
    .ZN(_05697_));
 NAND2_X1 _23177_ (.A1(\cs_registers_i.dscratch1_q[7] ),
    .A2(_04427_),
    .ZN(_05698_));
 AOI222_X2 _23178_ (.A1(net90),
    .A2(_04441_),
    .B1(_04407_),
    .B2(\cs_registers_i.csr_depc_o[7] ),
    .C1(net143),
    .C2(_04430_),
    .ZN(_05699_));
 NAND4_X2 _23179_ (.A1(_04457_),
    .A2(_05697_),
    .A3(_05698_),
    .A4(_05699_),
    .ZN(_05700_));
 AOI222_X2 _23180_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_04433_),
    .B1(_04508_),
    .B2(\cs_registers_i.mscratch_q[7] ),
    .C1(_04657_),
    .C2(\cs_registers_i.mstack_d[2] ),
    .ZN(_05701_));
 NAND2_X1 _23181_ (.A1(\cs_registers_i.mtval_q[7] ),
    .A2(_04414_),
    .ZN(_05702_));
 NAND2_X1 _23182_ (.A1(_05701_),
    .A2(_05702_),
    .ZN(_05703_));
 NOR3_X4 _23183_ (.A1(_05696_),
    .A2(_05700_),
    .A3(_05703_),
    .ZN(_05704_));
 NAND2_X1 _23184_ (.A1(_05689_),
    .A2(_05704_),
    .ZN(_05705_));
 NOR2_X1 _23185_ (.A1(_11173_),
    .A2(_05287_),
    .ZN(_05706_));
 AOI21_X1 _23186_ (.A(_05706_),
    .B1(_05628_),
    .B2(_11173_),
    .ZN(_05707_));
 MUX2_X1 _23187_ (.A(_05309_),
    .B(_05324_),
    .S(_05270_),
    .Z(_05708_));
 MUX2_X1 _23188_ (.A(_05308_),
    .B(_05708_),
    .S(_11173_),
    .Z(_05709_));
 MUX2_X1 _23189_ (.A(_05707_),
    .B(_05709_),
    .S(_05218_),
    .Z(_05710_));
 MUX2_X1 _23190_ (.A(_05294_),
    .B(_05637_),
    .S(_11173_),
    .Z(_05711_));
 MUX2_X1 _23191_ (.A(_05323_),
    .B(_05327_),
    .S(_11171_),
    .Z(_05712_));
 MUX2_X1 _23192_ (.A(_05569_),
    .B(_05712_),
    .S(_05240_),
    .Z(_05713_));
 MUX2_X1 _23193_ (.A(_05711_),
    .B(_05713_),
    .S(_05218_),
    .Z(_05714_));
 MUX2_X1 _23194_ (.A(_05710_),
    .B(_05714_),
    .S(_05339_),
    .Z(_05715_));
 NOR2_X1 _23195_ (.A1(_11171_),
    .A2(_05646_),
    .ZN(_05716_));
 AND2_X1 _23196_ (.A1(_11171_),
    .A2(_05332_),
    .ZN(_05717_));
 NOR2_X1 _23197_ (.A1(_05716_),
    .A2(_05717_),
    .ZN(_05718_));
 MUX2_X1 _23198_ (.A(_05469_),
    .B(_05718_),
    .S(_05248_),
    .Z(_05719_));
 MUX2_X2 _23199_ (.A(_05250_),
    .B(_05719_),
    .S(_05439_),
    .Z(_05720_));
 MUX2_X2 _23200_ (.A(_05715_),
    .B(_05720_),
    .S(_05651_),
    .Z(_05721_));
 NOR2_X1 _23201_ (.A1(_16295_),
    .A2(_05451_),
    .ZN(_05722_));
 OAI21_X1 _23202_ (.A(_05454_),
    .B1(_05461_),
    .B2(_16296_),
    .ZN(_05723_));
 AOI221_X2 _23203_ (.A(_05722_),
    .B1(_05723_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16299_),
    .ZN(_05724_));
 BUF_X4 _23204_ (.A(_05477_),
    .Z(_05725_));
 AOI21_X1 _23205_ (.A(_05724_),
    .B1(_05725_),
    .B2(\alu_adder_result_ex[7] ),
    .ZN(_05726_));
 NOR2_X2 _23206_ (.A1(_05264_),
    .A2(_05221_),
    .ZN(_05727_));
 NOR2_X1 _23207_ (.A1(_05437_),
    .A2(_05337_),
    .ZN(_05728_));
 AOI21_X1 _23208_ (.A(_05728_),
    .B1(_05321_),
    .B2(_05437_),
    .ZN(_05729_));
 MUX2_X1 _23209_ (.A(_05474_),
    .B(_05729_),
    .S(_05440_),
    .Z(_05730_));
 NAND2_X1 _23210_ (.A1(_05727_),
    .A2(_05730_),
    .ZN(_05731_));
 NAND3_X1 _23211_ (.A1(_05552_),
    .A2(_05726_),
    .A3(_05731_),
    .ZN(_05732_));
 AOI221_X2 _23212_ (.A(_05705_),
    .B1(_05721_),
    .B2(_05435_),
    .C1(_05732_),
    .C2(_05185_),
    .ZN(_05733_));
 BUF_X8 _23213_ (.A(_05588_),
    .Z(_05734_));
 AOI21_X4 _23214_ (.A(_05680_),
    .B1(_05733_),
    .B2(_05734_),
    .ZN(_05735_));
 BUF_X2 _23215_ (.A(_05735_),
    .Z(_05736_));
 NOR3_X4 _23216_ (.A1(_10862_),
    .A2(_11306_),
    .A3(_05409_),
    .ZN(_05737_));
 NAND2_X4 _23217_ (.A1(_05494_),
    .A2(_05737_),
    .ZN(_05738_));
 MUX2_X1 _23218_ (.A(_05736_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .S(_05738_),
    .Z(_01284_));
 CLKBUF_X3 _23219_ (.A(_05303_),
    .Z(_05739_));
 NAND2_X1 _23220_ (.A1(_05435_),
    .A2(_05739_),
    .ZN(_05740_));
 NAND2_X1 _23221_ (.A1(_05437_),
    .A2(_05312_),
    .ZN(_05741_));
 NAND2_X1 _23222_ (.A1(_05339_),
    .A2(_05329_),
    .ZN(_05742_));
 AOI21_X1 _23223_ (.A(_05440_),
    .B1(_05741_),
    .B2(_05742_),
    .ZN(_05743_));
 AOI21_X1 _23224_ (.A(_05743_),
    .B1(_05301_),
    .B2(_05560_),
    .ZN(_05744_));
 NOR2_X1 _23225_ (.A1(_05740_),
    .A2(_05744_),
    .ZN(_05745_));
 AND2_X1 _23226_ (.A1(_05727_),
    .A2(_05720_),
    .ZN(_05746_));
 NOR3_X1 _23227_ (.A1(_05256_),
    .A2(_05303_),
    .A3(_05554_),
    .ZN(_05747_));
 OAI21_X1 _23228_ (.A(_05747_),
    .B1(_05729_),
    .B2(_05542_),
    .ZN(_05748_));
 NAND2_X1 _23229_ (.A1(\alu_adder_result_ex[8] ),
    .A2(_05725_),
    .ZN(_05749_));
 BUF_X1 _23230_ (.A(_16046_),
    .Z(_05750_));
 INV_X1 _23231_ (.A(_16032_),
    .ZN(_05751_));
 AOI21_X1 _23232_ (.A(_16020_),
    .B1(_16021_),
    .B2(_14524_),
    .ZN(_05752_));
 OAI21_X2 _23233_ (.A(_05751_),
    .B1(_05752_),
    .B2(_05681_),
    .ZN(_05753_));
 XNOR2_X1 _23234_ (.A(_05750_),
    .B(_05753_),
    .ZN(_05754_));
 MUX2_X1 _23235_ (.A(_00564_),
    .B(_05754_),
    .S(_05428_),
    .Z(_05755_));
 INV_X1 _23236_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .ZN(_05756_));
 AOI221_X2 _23237_ (.A(_11865_),
    .B1(_03685_),
    .B2(_05755_),
    .C1(_05756_),
    .C2(net414),
    .ZN(_05757_));
 OR2_X1 _23238_ (.A1(_11282_),
    .A2(_05757_),
    .ZN(_05758_));
 NOR2_X1 _23239_ (.A1(_16303_),
    .A2(_05451_),
    .ZN(_05759_));
 OAI21_X1 _23240_ (.A(_05454_),
    .B1(_05461_),
    .B2(_16304_),
    .ZN(_05760_));
 AOI221_X2 _23241_ (.A(_05759_),
    .B1(_05760_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16307_),
    .ZN(_05761_));
 NOR2_X1 _23242_ (.A1(_05758_),
    .A2(_05761_),
    .ZN(_05762_));
 NAND4_X1 _23243_ (.A1(_05552_),
    .A2(_05748_),
    .A3(_05749_),
    .A4(_05762_),
    .ZN(_05763_));
 NOR3_X1 _23244_ (.A1(_05745_),
    .A2(_05746_),
    .A3(_05763_),
    .ZN(_05764_));
 OAI22_X1 _23245_ (.A1(_05489_),
    .A2(_04941_),
    .B1(_05185_),
    .B2(_05758_),
    .ZN(_05765_));
 OR3_X2 _23246_ (.A1(_05401_),
    .A2(_05764_),
    .A3(_05765_),
    .ZN(_05766_));
 MUX2_X1 _23247_ (.A(_05674_),
    .B(net53),
    .S(_05366_),
    .Z(_05767_));
 MUX2_X1 _23248_ (.A(net58),
    .B(net44),
    .S(_05366_),
    .Z(_05768_));
 MUX2_X2 _23249_ (.A(_05767_),
    .B(_05768_),
    .S(_05370_),
    .Z(_05769_));
 AND3_X2 _23250_ (.A1(_05379_),
    .A2(\load_store_unit_i.data_sign_ext_q ),
    .A3(_05769_),
    .ZN(_05770_));
 MUX2_X1 _23251_ (.A(net36),
    .B(net34),
    .S(_05366_),
    .Z(_05771_));
 MUX2_X1 _23252_ (.A(_05374_),
    .B(net45),
    .S(_05385_),
    .Z(_05772_));
 MUX2_X1 _23253_ (.A(_05771_),
    .B(_05772_),
    .S(_05503_),
    .Z(_05773_));
 MUX2_X1 _23254_ (.A(_05374_),
    .B(\load_store_unit_i.rdata_q[24] ),
    .S(_05385_),
    .Z(_05774_));
 MUX2_X1 _23255_ (.A(\load_store_unit_i.rdata_q[16] ),
    .B(net34),
    .S(_05388_),
    .Z(_05775_));
 MUX2_X1 _23256_ (.A(_05774_),
    .B(_05775_),
    .S(_05360_),
    .Z(_05776_));
 AOI221_X2 _23257_ (.A(_05770_),
    .B1(_05773_),
    .B2(_05363_),
    .C1(_05776_),
    .C2(_05499_),
    .ZN(_05777_));
 OAI21_X4 _23258_ (.A(_05766_),
    .B1(_05777_),
    .B2(_05734_),
    .ZN(_05778_));
 BUF_X2 _23259_ (.A(_05778_),
    .Z(_05779_));
 MUX2_X1 _23260_ (.A(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .B(_05779_),
    .S(_05498_),
    .Z(_01285_));
 INV_X1 _23261_ (.A(_16045_),
    .ZN(_05780_));
 AOI21_X1 _23262_ (.A(_16032_),
    .B1(_05685_),
    .B2(_16033_),
    .ZN(_05781_));
 INV_X1 _23263_ (.A(_05750_),
    .ZN(_05782_));
 OAI21_X1 _23264_ (.A(_05780_),
    .B1(_05781_),
    .B2(_05782_),
    .ZN(_05783_));
 XNOR2_X2 _23265_ (.A(_16060_),
    .B(_05783_),
    .ZN(_05784_));
 MUX2_X1 _23266_ (.A(_00565_),
    .B(_05784_),
    .S(_05428_),
    .Z(_05785_));
 AND2_X1 _23267_ (.A1(_03685_),
    .A2(_05785_),
    .ZN(_05786_));
 OAI21_X1 _23268_ (.A(_12276_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B2(_10912_),
    .ZN(_05787_));
 OAI21_X2 _23269_ (.A(_10973_),
    .B1(_05786_),
    .B2(_05787_),
    .ZN(_05788_));
 OAI21_X1 _23270_ (.A(_05454_),
    .B1(_05456_),
    .B2(_16312_),
    .ZN(_05789_));
 NAND2_X1 _23271_ (.A1(_05460_),
    .A2(_05789_),
    .ZN(_05790_));
 NOR2_X1 _23272_ (.A1(_16311_),
    .A2(_05451_),
    .ZN(_05791_));
 AOI21_X2 _23273_ (.A(_05791_),
    .B1(_05456_),
    .B2(_16315_),
    .ZN(_05792_));
 AOI221_X2 _23274_ (.A(_05788_),
    .B1(_05790_),
    .B2(_05792_),
    .C1(\alu_adder_result_ex[9] ),
    .C2(_05477_),
    .ZN(_05793_));
 NAND2_X1 _23275_ (.A1(_05552_),
    .A2(_05793_),
    .ZN(_05794_));
 AOI21_X1 _23276_ (.A(_05794_),
    .B1(_05650_),
    .B2(_05562_),
    .ZN(_05795_));
 MUX2_X1 _23277_ (.A(_05573_),
    .B(_05534_),
    .S(_05542_),
    .Z(_05796_));
 MUX2_X1 _23278_ (.A(_05567_),
    .B(_05579_),
    .S(_05440_),
    .Z(_05797_));
 MUX2_X1 _23279_ (.A(_05796_),
    .B(_05797_),
    .S(_05536_),
    .Z(_05798_));
 AOI21_X1 _23280_ (.A(_05623_),
    .B1(_05531_),
    .B2(_05536_),
    .ZN(_05799_));
 NAND2_X1 _23281_ (.A1(_05560_),
    .A2(_05799_),
    .ZN(_05800_));
 NOR2_X1 _23282_ (.A1(_05739_),
    .A2(_05554_),
    .ZN(_05801_));
 AOI22_X1 _23283_ (.A1(_05739_),
    .A2(_05798_),
    .B1(_05800_),
    .B2(_05801_),
    .ZN(_05802_));
 OAI21_X1 _23284_ (.A(_05795_),
    .B1(_05802_),
    .B2(_05256_),
    .ZN(_05803_));
 NOR2_X1 _23285_ (.A1(_05427_),
    .A2(_05788_),
    .ZN(_05804_));
 AOI21_X1 _23286_ (.A(_05804_),
    .B1(_04957_),
    .B2(_05357_),
    .ZN(_05805_));
 NAND3_X2 _23287_ (.A1(_05734_),
    .A2(_05803_),
    .A3(_05805_),
    .ZN(_05806_));
 MUX2_X1 _23288_ (.A(net37),
    .B(net40),
    .S(_05366_),
    .Z(_05807_));
 BUF_X1 _23289_ (.A(data_rdata_i[9]),
    .Z(_05808_));
 MUX2_X1 _23290_ (.A(_05808_),
    .B(net46),
    .S(_05385_),
    .Z(_05809_));
 MUX2_X1 _23291_ (.A(_05807_),
    .B(_05809_),
    .S(_05503_),
    .Z(_05810_));
 MUX2_X1 _23292_ (.A(_05808_),
    .B(\load_store_unit_i.rdata_q[25] ),
    .S(_05385_),
    .Z(_05811_));
 MUX2_X1 _23293_ (.A(\load_store_unit_i.rdata_q[17] ),
    .B(net40),
    .S(_05385_),
    .Z(_05812_));
 MUX2_X1 _23294_ (.A(_05811_),
    .B(_05812_),
    .S(_05360_),
    .Z(_05813_));
 AOI221_X2 _23295_ (.A(_05770_),
    .B1(_05810_),
    .B2(_05363_),
    .C1(_05813_),
    .C2(_05499_),
    .ZN(_05814_));
 OAI21_X4 _23296_ (.A(_05806_),
    .B1(_05814_),
    .B2(_05734_),
    .ZN(_05815_));
 BUF_X2 _23297_ (.A(_05815_),
    .Z(_05816_));
 MUX2_X1 _23298_ (.A(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .B(_05816_),
    .S(_05498_),
    .Z(_01286_));
 BUF_X4 _23299_ (.A(_05738_),
    .Z(_05817_));
 NAND2_X1 _23300_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .A2(_05817_),
    .ZN(_05818_));
 NAND3_X4 _23301_ (.A1(_05364_),
    .A2(\load_store_unit_i.data_sign_ext_q ),
    .A3(_05769_),
    .ZN(_05819_));
 MUX2_X1 _23302_ (.A(net38),
    .B(net51),
    .S(_05388_),
    .Z(_05820_));
 CLKBUF_X2 _23303_ (.A(data_rdata_i[10]),
    .Z(_05821_));
 MUX2_X1 _23304_ (.A(_05821_),
    .B(net47),
    .S(_05386_),
    .Z(_05822_));
 MUX2_X1 _23305_ (.A(_05820_),
    .B(_05822_),
    .S(_05503_),
    .Z(_05823_));
 MUX2_X1 _23306_ (.A(_05821_),
    .B(\load_store_unit_i.rdata_q[26] ),
    .S(_05388_),
    .Z(_05824_));
 MUX2_X1 _23307_ (.A(\load_store_unit_i.rdata_q[18] ),
    .B(net51),
    .S(_05388_),
    .Z(_05825_));
 MUX2_X1 _23308_ (.A(_05824_),
    .B(_05825_),
    .S(_05360_),
    .Z(_05826_));
 BUF_X4 _23309_ (.A(_05499_),
    .Z(_05827_));
 AOI22_X2 _23310_ (.A1(_05363_),
    .A2(_05823_),
    .B1(_05826_),
    .B2(_05827_),
    .ZN(_05828_));
 AOI21_X2 _23311_ (.A(_05588_),
    .B1(_05819_),
    .B2(_05828_),
    .ZN(_05829_));
 CLKBUF_X3 _23312_ (.A(\cs_registers_i.mhpmcounter[2][42] ),
    .Z(_05830_));
 AOI22_X4 _23313_ (.A1(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .A2(_04590_),
    .B1(_04501_),
    .B2(_05830_),
    .ZN(_05831_));
 AOI22_X4 _23314_ (.A1(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .A2(_04500_),
    .B1(_04501_),
    .B2(\cs_registers_i.mhpmcounter[2][10] ),
    .ZN(_05832_));
 OAI22_X4 _23315_ (.A1(_04498_),
    .A2(_05831_),
    .B1(_05832_),
    .B2(_04629_),
    .ZN(_05833_));
 AOI222_X2 _23316_ (.A1(\cs_registers_i.csr_depc_o[10] ),
    .A2(_04518_),
    .B1(_04424_),
    .B2(\cs_registers_i.csr_mepc_o[10] ),
    .C1(_04427_),
    .C2(\cs_registers_i.dscratch1_q[10] ),
    .ZN(_05834_));
 AOI22_X2 _23317_ (.A1(\cs_registers_i.dscratch0_q[10] ),
    .A2(_04632_),
    .B1(_04509_),
    .B2(\cs_registers_i.mscratch_q[10] ),
    .ZN(_05835_));
 NOR2_X1 _23318_ (.A1(_01171_),
    .A2(_04461_),
    .ZN(_05836_));
 AOI21_X1 _23319_ (.A(_05836_),
    .B1(_04442_),
    .B2(net62),
    .ZN(_05837_));
 NAND3_X2 _23320_ (.A1(_05834_),
    .A2(_05835_),
    .A3(_05837_),
    .ZN(_05838_));
 AND2_X1 _23321_ (.A1(\cs_registers_i.mtval_q[10] ),
    .A2(_04634_),
    .ZN(_05839_));
 NOR4_X4 _23322_ (.A1(_04545_),
    .A2(_05833_),
    .A3(_05838_),
    .A4(_05839_),
    .ZN(_05840_));
 NAND2_X1 _23323_ (.A1(_05560_),
    .A2(_05559_),
    .ZN(_05841_));
 AND2_X1 _23324_ (.A1(_05841_),
    .A2(_05747_),
    .ZN(_05842_));
 NOR2_X1 _23325_ (.A1(_16319_),
    .A2(_05451_),
    .ZN(_05843_));
 OAI21_X1 _23326_ (.A(_05454_),
    .B1(_05456_),
    .B2(_16320_),
    .ZN(_05844_));
 AOI221_X2 _23327_ (.A(_05843_),
    .B1(_05844_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16323_),
    .ZN(_05845_));
 AOI21_X1 _23328_ (.A(_05845_),
    .B1(_05725_),
    .B2(\alu_adder_result_ex[10] ),
    .ZN(_05846_));
 NAND3_X1 _23329_ (.A1(_05536_),
    .A2(_05630_),
    .A3(_05635_),
    .ZN(_05847_));
 MUX2_X1 _23330_ (.A(_05641_),
    .B(_05647_),
    .S(_05542_),
    .Z(_05848_));
 OAI21_X1 _23331_ (.A(_05847_),
    .B1(_05848_),
    .B2(_05536_),
    .ZN(_05849_));
 OAI21_X1 _23332_ (.A(_05846_),
    .B1(_05849_),
    .B2(_05740_),
    .ZN(_05850_));
 OAI21_X1 _23333_ (.A(_05427_),
    .B1(_05842_),
    .B2(_05850_),
    .ZN(_05851_));
 CLKBUF_X3 _23334_ (.A(_05430_),
    .Z(_05852_));
 CLKBUF_X3 _23335_ (.A(_05852_),
    .Z(_05853_));
 INV_X1 _23336_ (.A(_16059_),
    .ZN(_05854_));
 AOI21_X1 _23337_ (.A(_16045_),
    .B1(_05753_),
    .B2(_05750_),
    .ZN(_05855_));
 INV_X1 _23338_ (.A(_16060_),
    .ZN(_05856_));
 OAI21_X1 _23339_ (.A(_05854_),
    .B1(_05855_),
    .B2(_05856_),
    .ZN(_05857_));
 XOR2_X2 _23340_ (.A(net376),
    .B(_05857_),
    .Z(_05858_));
 NAND2_X1 _23341_ (.A1(_05853_),
    .A2(_05858_),
    .ZN(_05859_));
 OAI21_X2 _23342_ (.A(_05859_),
    .B1(_05853_),
    .B2(_00566_),
    .ZN(_05860_));
 OAI221_X2 _23343_ (.A(_04176_),
    .B1(_03738_),
    .B2(_05860_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .C2(_10913_),
    .ZN(_05861_));
 NAND2_X1 _23344_ (.A1(_05651_),
    .A2(_05474_),
    .ZN(_05862_));
 OAI21_X1 _23345_ (.A(_05443_),
    .B1(_05540_),
    .B2(_05221_),
    .ZN(_05863_));
 AOI22_X1 _23346_ (.A1(_05222_),
    .A2(_05535_),
    .B1(_05863_),
    .B2(_05542_),
    .ZN(_05864_));
 NAND2_X1 _23347_ (.A1(_05862_),
    .A2(_05864_),
    .ZN(_05865_));
 NAND2_X1 _23348_ (.A1(_05163_),
    .A2(_05865_),
    .ZN(_05866_));
 NAND4_X2 _23349_ (.A1(_05840_),
    .A2(_05851_),
    .A3(_05861_),
    .A4(_05866_),
    .ZN(_05867_));
 AOI21_X4 _23350_ (.A(_05829_),
    .B1(_05867_),
    .B2(_05734_),
    .ZN(_05868_));
 CLKBUF_X3 _23351_ (.A(_05868_),
    .Z(_05869_));
 OAI21_X1 _23352_ (.A(_05818_),
    .B1(_05869_),
    .B2(_05817_),
    .ZN(_01287_));
 NOR2_X1 _23353_ (.A1(_16327_),
    .A2(_05450_),
    .ZN(_05870_));
 OAI21_X1 _23354_ (.A(_05453_),
    .B1(_05549_),
    .B2(_16328_),
    .ZN(_05871_));
 AOI221_X2 _23355_ (.A(_05870_),
    .B1(_05871_),
    .B2(_05459_),
    .C1(_05456_),
    .C2(_16331_),
    .ZN(_05872_));
 AOI21_X1 _23356_ (.A(_05872_),
    .B1(_05477_),
    .B2(\alu_adder_result_ex[11] ),
    .ZN(_05873_));
 AOI21_X1 _23357_ (.A(_05596_),
    .B1(_05552_),
    .B2(_05873_),
    .ZN(_05874_));
 AOI21_X1 _23358_ (.A(_05874_),
    .B1(_05562_),
    .B2(_05446_),
    .ZN(_05875_));
 NOR3_X1 _23359_ (.A1(_05339_),
    .A2(_05716_),
    .A3(_05717_),
    .ZN(_05876_));
 AND2_X1 _23360_ (.A1(_05249_),
    .A2(_05709_),
    .ZN(_05877_));
 OAI21_X1 _23361_ (.A(_05739_),
    .B1(_05876_),
    .B2(_05877_),
    .ZN(_05878_));
 AOI21_X1 _23362_ (.A(_05560_),
    .B1(_05862_),
    .B2(_05878_),
    .ZN(_05879_));
 MUX2_X1 _23363_ (.A(_05707_),
    .B(_05713_),
    .S(_05437_),
    .Z(_05880_));
 MUX2_X1 _23364_ (.A(_05472_),
    .B(_05880_),
    .S(_05739_),
    .Z(_05881_));
 AOI21_X2 _23365_ (.A(_05879_),
    .B1(_05881_),
    .B2(_05560_),
    .ZN(_05882_));
 OAI21_X1 _23366_ (.A(_05875_),
    .B1(_05882_),
    .B2(_05256_),
    .ZN(_05883_));
 NOR3_X4 _23367_ (.A1(_03776_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A3(_03750_),
    .ZN(_05884_));
 INV_X1 _23368_ (.A(_16073_),
    .ZN(_05885_));
 OAI21_X2 _23369_ (.A(_16074_),
    .B1(_16059_),
    .B2(_16060_),
    .ZN(_05886_));
 NAND2_X1 _23370_ (.A1(_05885_),
    .A2(_05886_),
    .ZN(_05887_));
 NOR3_X4 _23371_ (.A1(_16045_),
    .A2(_16059_),
    .A3(_16073_),
    .ZN(_05888_));
 OAI21_X1 _23372_ (.A(_05888_),
    .B1(_05781_),
    .B2(_05782_),
    .ZN(_05889_));
 NAND2_X1 _23373_ (.A1(_05887_),
    .A2(_05889_),
    .ZN(_05890_));
 XNOR2_X2 _23374_ (.A(_16088_),
    .B(_05890_),
    .ZN(_05891_));
 NOR2_X1 _23375_ (.A1(_05884_),
    .A2(_05891_),
    .ZN(_05892_));
 AOI21_X2 _23376_ (.A(_05892_),
    .B1(_05884_),
    .B2(_00567_),
    .ZN(_05893_));
 OAI221_X2 _23377_ (.A(_03755_),
    .B1(_03737_),
    .B2(_05893_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .C2(_10913_),
    .ZN(_05894_));
 NAND2_X1 _23378_ (.A1(_04463_),
    .A2(_05894_),
    .ZN(_05895_));
 NOR3_X2 _23379_ (.A1(_05401_),
    .A2(_05883_),
    .A3(_05895_),
    .ZN(_05896_));
 NOR2_X4 _23380_ (.A1(_05588_),
    .A2(_05770_),
    .ZN(_05897_));
 CLKBUF_X3 _23381_ (.A(_05385_),
    .Z(_05898_));
 MUX2_X1 _23382_ (.A(net39),
    .B(net54),
    .S(_05898_),
    .Z(_05899_));
 BUF_X1 _23383_ (.A(data_rdata_i[11]),
    .Z(_05900_));
 MUX2_X1 _23384_ (.A(_05900_),
    .B(net48),
    .S(_05898_),
    .Z(_05901_));
 CLKBUF_X3 _23385_ (.A(_05503_),
    .Z(_05902_));
 MUX2_X1 _23386_ (.A(_05899_),
    .B(_05901_),
    .S(_05902_),
    .Z(_05903_));
 MUX2_X1 _23387_ (.A(_05900_),
    .B(\load_store_unit_i.rdata_q[27] ),
    .S(_05386_),
    .Z(_05904_));
 MUX2_X1 _23388_ (.A(\load_store_unit_i.rdata_q[19] ),
    .B(net54),
    .S(_05898_),
    .Z(_05905_));
 MUX2_X1 _23389_ (.A(_05904_),
    .B(_05905_),
    .S(_05415_),
    .Z(_05906_));
 AOI22_X4 _23390_ (.A1(_05363_),
    .A2(_05903_),
    .B1(_05906_),
    .B2(_05827_),
    .ZN(_05907_));
 AOI21_X4 _23391_ (.A(_05896_),
    .B1(_05897_),
    .B2(_05907_),
    .ZN(_05908_));
 BUF_X2 _23392_ (.A(_05908_),
    .Z(_05909_));
 MUX2_X1 _23393_ (.A(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .B(_05909_),
    .S(_05498_),
    .Z(_01288_));
 OAI21_X1 _23394_ (.A(_03755_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B2(_10913_),
    .ZN(_05910_));
 NAND2_X1 _23395_ (.A1(_05750_),
    .A2(_05753_),
    .ZN(_05911_));
 AOI22_X4 _23396_ (.A1(_05885_),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_05911_),
    .ZN(_05912_));
 AOI21_X1 _23397_ (.A(_16087_),
    .B1(_05912_),
    .B2(_16088_),
    .ZN(_05913_));
 XOR2_X2 _23398_ (.A(net279),
    .B(_05913_),
    .Z(_05914_));
 MUX2_X1 _23399_ (.A(_00568_),
    .B(_05914_),
    .S(_05852_),
    .Z(_05915_));
 AOI21_X2 _23400_ (.A(_05910_),
    .B1(_05915_),
    .B2(_03686_),
    .ZN(_05916_));
 INV_X1 _23401_ (.A(_05862_),
    .ZN(_05917_));
 OR2_X1 _23402_ (.A1(_05876_),
    .A2(_05877_),
    .ZN(_05918_));
 MUX2_X2 _23403_ (.A(_05472_),
    .B(_05918_),
    .S(_05440_),
    .Z(_05919_));
 AOI21_X1 _23404_ (.A(_05917_),
    .B1(_05919_),
    .B2(_05739_),
    .ZN(_05920_));
 NOR2_X2 _23405_ (.A1(_05264_),
    .A2(_05920_),
    .ZN(_05921_));
 NOR2_X1 _23406_ (.A1(_16335_),
    .A2(_05450_),
    .ZN(_05922_));
 OAI21_X1 _23407_ (.A(_05453_),
    .B1(_05455_),
    .B2(_16336_),
    .ZN(_05923_));
 AOI221_X2 _23408_ (.A(_05922_),
    .B1(_05923_),
    .B2(_05459_),
    .C1(_05456_),
    .C2(_16339_),
    .ZN(_05924_));
 OAI21_X2 _23409_ (.A(_05225_),
    .B1(_05218_),
    .B2(_05229_),
    .ZN(_05925_));
 NAND2_X1 _23410_ (.A1(_05249_),
    .A2(_05439_),
    .ZN(_05926_));
 OAI21_X1 _23411_ (.A(_05925_),
    .B1(_05926_),
    .B2(_05321_),
    .ZN(_05927_));
 MUX2_X1 _23412_ (.A(_05436_),
    .B(_05442_),
    .S(_05218_),
    .Z(_05928_));
 MUX2_X1 _23413_ (.A(_05927_),
    .B(_05928_),
    .S(_05303_),
    .Z(_05929_));
 AOI221_X2 _23414_ (.A(_05924_),
    .B1(_05929_),
    .B2(_05435_),
    .C1(\alu_adder_result_ex[12] ),
    .C2(_05477_),
    .ZN(_05930_));
 OAI21_X2 _23415_ (.A(_05405_),
    .B1(_05596_),
    .B2(_05930_),
    .ZN(_05931_));
 NOR4_X4 _23416_ (.A1(_04526_),
    .A2(_05916_),
    .A3(_05921_),
    .A4(_05931_),
    .ZN(_05932_));
 MUX2_X1 _23417_ (.A(net41),
    .B(net55),
    .S(_05898_),
    .Z(_05933_));
 MUX2_X1 _23418_ (.A(_05419_),
    .B(net49),
    .S(_05898_),
    .Z(_05934_));
 MUX2_X1 _23419_ (.A(_05933_),
    .B(_05934_),
    .S(_05902_),
    .Z(_05935_));
 MUX2_X1 _23420_ (.A(_05419_),
    .B(\load_store_unit_i.rdata_q[28] ),
    .S(_05898_),
    .Z(_05936_));
 MUX2_X1 _23421_ (.A(\load_store_unit_i.rdata_q[20] ),
    .B(net55),
    .S(_05898_),
    .Z(_05937_));
 MUX2_X1 _23422_ (.A(_05936_),
    .B(_05937_),
    .S(_05415_),
    .Z(_05938_));
 AOI22_X4 _23423_ (.A1(_05363_),
    .A2(_05935_),
    .B1(_05938_),
    .B2(_05827_),
    .ZN(_05939_));
 AOI21_X4 _23424_ (.A(_05932_),
    .B1(_05939_),
    .B2(_05897_),
    .ZN(_05940_));
 BUF_X2 _23425_ (.A(_05940_),
    .Z(_05941_));
 MUX2_X1 _23426_ (.A(_05941_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .S(_05738_),
    .Z(_01289_));
 NOR2_X1 _23427_ (.A1(_16347_),
    .A2(_05449_),
    .ZN(_05942_));
 OAI21_X1 _23428_ (.A(_05161_),
    .B1(_05548_),
    .B2(_16344_),
    .ZN(_05943_));
 AOI221_X1 _23429_ (.A(_05942_),
    .B1(_05943_),
    .B2(_05458_),
    .C1(_05549_),
    .C2(_16343_),
    .ZN(_05944_));
 AOI21_X1 _23430_ (.A(_05944_),
    .B1(_05476_),
    .B2(\alu_adder_result_ex[13] ),
    .ZN(_05945_));
 AOI21_X1 _23431_ (.A(_05595_),
    .B1(_05552_),
    .B2(_05945_),
    .ZN(_05946_));
 NOR2_X1 _23432_ (.A1(_05229_),
    .A2(_05634_),
    .ZN(_05947_));
 AND2_X1 _23433_ (.A1(_05229_),
    .A2(_05647_),
    .ZN(_05948_));
 NOR3_X2 _23434_ (.A1(_05445_),
    .A2(_05947_),
    .A3(_05948_),
    .ZN(_05949_));
 AOI21_X4 _23435_ (.A(_05949_),
    .B1(_05559_),
    .B2(_05445_),
    .ZN(_05950_));
 AOI21_X1 _23436_ (.A(_05946_),
    .B1(_05950_),
    .B2(_05562_),
    .ZN(_05951_));
 NAND3_X1 _23437_ (.A1(_05249_),
    .A2(_05439_),
    .A3(_05539_),
    .ZN(_05952_));
 NAND3_X1 _23438_ (.A1(_05651_),
    .A2(_05925_),
    .A3(_05952_),
    .ZN(_05953_));
 MUX2_X1 _23439_ (.A(_05574_),
    .B(_05535_),
    .S(_05542_),
    .Z(_05954_));
 OAI21_X1 _23440_ (.A(_05953_),
    .B1(_05954_),
    .B2(_05651_),
    .ZN(_05955_));
 OAI21_X1 _23441_ (.A(_05951_),
    .B1(_05955_),
    .B2(_05256_),
    .ZN(_05956_));
 INV_X1 _23442_ (.A(_16087_),
    .ZN(_05957_));
 INV_X1 _23443_ (.A(_16088_),
    .ZN(_05958_));
 OAI21_X1 _23444_ (.A(_05957_),
    .B1(_05890_),
    .B2(_05958_),
    .ZN(_05959_));
 AOI21_X1 _23445_ (.A(_16101_),
    .B1(_05959_),
    .B2(_16102_),
    .ZN(_05960_));
 XOR2_X2 _23446_ (.A(net280),
    .B(_05960_),
    .Z(_05961_));
 NAND3_X1 _23447_ (.A1(_03685_),
    .A2(_05852_),
    .A3(_05961_),
    .ZN(_05962_));
 OAI21_X1 _23448_ (.A(_04163_),
    .B1(_05884_),
    .B2(_10922_),
    .ZN(_05963_));
 AND3_X1 _23449_ (.A1(_03755_),
    .A2(_05962_),
    .A3(_05963_),
    .ZN(_05964_));
 OR3_X1 _23450_ (.A1(_04561_),
    .A2(_05956_),
    .A3(_05964_),
    .ZN(_05965_));
 MUX2_X1 _23451_ (.A(net42),
    .B(net56),
    .S(_05385_),
    .Z(_05966_));
 MUX2_X1 _23452_ (.A(_05500_),
    .B(net50),
    .S(_05388_),
    .Z(_05967_));
 MUX2_X1 _23453_ (.A(_05966_),
    .B(_05967_),
    .S(_05503_),
    .Z(_05968_));
 MUX2_X1 _23454_ (.A(_05500_),
    .B(\load_store_unit_i.rdata_q[29] ),
    .S(_05385_),
    .Z(_05969_));
 MUX2_X1 _23455_ (.A(\load_store_unit_i.rdata_q[21] ),
    .B(net56),
    .S(_05385_),
    .Z(_05970_));
 MUX2_X1 _23456_ (.A(_05969_),
    .B(_05970_),
    .S(_05360_),
    .Z(_05971_));
 AOI22_X1 _23457_ (.A1(_05363_),
    .A2(_05968_),
    .B1(_05971_),
    .B2(_05499_),
    .ZN(_05972_));
 NAND2_X1 _23458_ (.A1(_05819_),
    .A2(_05972_),
    .ZN(_05973_));
 MUX2_X2 _23459_ (.A(_05965_),
    .B(_05973_),
    .S(_05401_),
    .Z(_05974_));
 BUF_X2 _23460_ (.A(_05974_),
    .Z(_05975_));
 MUX2_X1 _23461_ (.A(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .B(_05975_),
    .S(_05498_),
    .Z(_01290_));
 BUF_X4 _23462_ (.A(_05410_),
    .Z(_05976_));
 NAND2_X1 _23463_ (.A1(_11311_),
    .A2(_05976_),
    .ZN(_05977_));
 CLKBUF_X3 _23464_ (.A(_05977_),
    .Z(_05978_));
 NAND2_X1 _23465_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .A2(_05978_),
    .ZN(_05979_));
 CLKBUF_X3 _23466_ (.A(_05977_),
    .Z(_05980_));
 OAI21_X1 _23467_ (.A(_05979_),
    .B1(_05869_),
    .B2(_05980_),
    .ZN(_01291_));
 NOR3_X1 _23468_ (.A1(_05489_),
    .A2(_04595_),
    .A3(_05668_),
    .ZN(_05981_));
 INV_X1 _23469_ (.A(_16108_),
    .ZN(_05982_));
 NAND2_X1 _23470_ (.A1(_16109_),
    .A2(_16101_),
    .ZN(_05983_));
 NAND3_X1 _23471_ (.A1(_16102_),
    .A2(_16109_),
    .A3(_16087_),
    .ZN(_05984_));
 NAND2_X2 _23472_ (.A1(_05983_),
    .A2(_05984_),
    .ZN(_05985_));
 AND3_X4 _23473_ (.A1(_16088_),
    .A2(_16109_),
    .A3(_16102_),
    .ZN(_05986_));
 AOI21_X4 _23474_ (.A(_05985_),
    .B1(_05986_),
    .B2(_05912_),
    .ZN(_05987_));
 NAND2_X1 _23475_ (.A1(_05982_),
    .A2(_05987_),
    .ZN(_05988_));
 XNOR2_X2 _23476_ (.A(_16119_),
    .B(_05988_),
    .ZN(_05989_));
 NAND3_X1 _23477_ (.A1(_03685_),
    .A2(_05852_),
    .A3(_05989_),
    .ZN(_05990_));
 OAI21_X1 _23478_ (.A(_00630_),
    .B1(_05884_),
    .B2(_10922_),
    .ZN(_05991_));
 AND3_X1 _23479_ (.A1(_03755_),
    .A2(_05990_),
    .A3(_05991_),
    .ZN(_05992_));
 NOR3_X1 _23480_ (.A1(_05357_),
    .A2(_05668_),
    .A3(_05992_),
    .ZN(_05993_));
 NOR4_X4 _23481_ (.A1(_05173_),
    .A2(_10943_),
    .A3(_05174_),
    .A4(_05223_),
    .ZN(_05994_));
 AOI21_X1 _23482_ (.A(_05560_),
    .B1(_05221_),
    .B2(_05994_),
    .ZN(_05995_));
 OAI21_X1 _23483_ (.A(_05995_),
    .B1(_05649_),
    .B2(_05651_),
    .ZN(_05996_));
 NOR2_X1 _23484_ (.A1(_05303_),
    .A2(_05644_),
    .ZN(_05997_));
 NOR2_X1 _23485_ (.A1(_05249_),
    .A2(_05634_),
    .ZN(_05998_));
 AOI211_X2 _23486_ (.A(_05221_),
    .B(_05998_),
    .C1(_05641_),
    .C2(_05339_),
    .ZN(_05999_));
 OAI21_X1 _23487_ (.A(_05560_),
    .B1(_05997_),
    .B2(_05999_),
    .ZN(_06000_));
 NAND2_X1 _23488_ (.A1(_05996_),
    .A2(_06000_),
    .ZN(_06001_));
 NOR2_X1 _23489_ (.A1(_05256_),
    .A2(_06001_),
    .ZN(_06002_));
 NOR2_X1 _23490_ (.A1(_16355_),
    .A2(_05450_),
    .ZN(_06003_));
 OAI21_X1 _23491_ (.A(_05161_),
    .B1(_05455_),
    .B2(_16352_),
    .ZN(_06004_));
 AOI221_X2 _23492_ (.A(_06003_),
    .B1(_06004_),
    .B2(_05458_),
    .C1(_05461_),
    .C2(_16351_),
    .ZN(_06005_));
 NOR2_X2 _23493_ (.A1(_05274_),
    .A2(_05303_),
    .ZN(_06006_));
 AOI221_X2 _23494_ (.A(_06005_),
    .B1(_06006_),
    .B2(_05994_),
    .C1(net7),
    .C2(_05477_),
    .ZN(_06007_));
 NAND2_X1 _23495_ (.A1(_05440_),
    .A2(_05534_),
    .ZN(_06008_));
 NAND2_X1 _23496_ (.A1(_05445_),
    .A2(_05539_),
    .ZN(_06009_));
 AOI21_X1 _23497_ (.A(_05339_),
    .B1(_06008_),
    .B2(_06009_),
    .ZN(_06010_));
 MUX2_X1 _23498_ (.A(_05567_),
    .B(_05531_),
    .S(_05445_),
    .Z(_06011_));
 AOI21_X2 _23499_ (.A(_06010_),
    .B1(_06011_),
    .B2(_05536_),
    .ZN(_06012_));
 NAND2_X1 _23500_ (.A1(_05163_),
    .A2(_05739_),
    .ZN(_06013_));
 OAI21_X1 _23501_ (.A(_06007_),
    .B1(_06012_),
    .B2(_06013_),
    .ZN(_06014_));
 AOI21_X1 _23502_ (.A(_06002_),
    .B1(_06014_),
    .B2(_05185_),
    .ZN(_06015_));
 NAND2_X1 _23503_ (.A1(net35),
    .A2(_05389_),
    .ZN(_06016_));
 AOI221_X1 _23504_ (.A(_05362_),
    .B1(\load_store_unit_i.rdata_q[30] ),
    .B2(_05369_),
    .C1(\load_store_unit_i.rdata_q[22] ),
    .C2(_05367_),
    .ZN(_06017_));
 NOR2_X1 _23505_ (.A1(_05366_),
    .A2(_05655_),
    .ZN(_06018_));
 AOI221_X1 _23506_ (.A(_05380_),
    .B1(net52),
    .B2(_05368_),
    .C1(_06018_),
    .C2(_05359_),
    .ZN(_06019_));
 OR2_X1 _23507_ (.A1(_06017_),
    .A2(_06019_),
    .ZN(_06020_));
 OAI21_X1 _23508_ (.A(_06016_),
    .B1(_06020_),
    .B2(_05367_),
    .ZN(_06021_));
 NAND2_X1 _23509_ (.A1(_05898_),
    .A2(net57),
    .ZN(_06022_));
 AOI21_X1 _23510_ (.A(_05503_),
    .B1(_06020_),
    .B2(_06022_),
    .ZN(_06023_));
 OAI21_X1 _23511_ (.A(_05381_),
    .B1(_06021_),
    .B2(_06023_),
    .ZN(_06024_));
 AND2_X1 _23512_ (.A1(_05819_),
    .A2(_06024_),
    .ZN(_06025_));
 AOI221_X2 _23513_ (.A(_05981_),
    .B1(_05993_),
    .B2(_06015_),
    .C1(_05668_),
    .C2(_06025_),
    .ZN(_06026_));
 BUF_X2 _23514_ (.A(_06026_),
    .Z(_06027_));
 MUX2_X1 _23515_ (.A(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .B(_06027_),
    .S(_05498_),
    .Z(_01292_));
 MUX2_X1 _23516_ (.A(net44),
    .B(net58),
    .S(_05366_),
    .Z(_06028_));
 MUX2_X2 _23517_ (.A(_05767_),
    .B(_06028_),
    .S(_05359_),
    .Z(_06029_));
 MUX2_X1 _23518_ (.A(_05674_),
    .B(\load_store_unit_i.rdata_q[31] ),
    .S(_05386_),
    .Z(_06030_));
 MUX2_X1 _23519_ (.A(\load_store_unit_i.rdata_q[23] ),
    .B(net58),
    .S(_05386_),
    .Z(_06031_));
 MUX2_X1 _23520_ (.A(_06030_),
    .B(_06031_),
    .S(_05415_),
    .Z(_06032_));
 AOI22_X4 _23521_ (.A1(_05363_),
    .A2(_06029_),
    .B1(_06032_),
    .B2(_05827_),
    .ZN(_06033_));
 NOR2_X1 _23522_ (.A1(_16363_),
    .A2(_05449_),
    .ZN(_06034_));
 OAI21_X1 _23523_ (.A(_05161_),
    .B1(_05548_),
    .B2(_16360_),
    .ZN(_06035_));
 AOI221_X2 _23524_ (.A(_06034_),
    .B1(_06035_),
    .B2(_05458_),
    .C1(_05549_),
    .C2(_16359_),
    .ZN(_06036_));
 AOI21_X1 _23525_ (.A(_06036_),
    .B1(_05476_),
    .B2(net439),
    .ZN(_06037_));
 OAI21_X1 _23526_ (.A(_05747_),
    .B1(_05250_),
    .B2(_05542_),
    .ZN(_06038_));
 NAND3_X1 _23527_ (.A1(_05552_),
    .A2(_06037_),
    .A3(_06038_),
    .ZN(_06039_));
 MUX2_X1 _23528_ (.A(_05469_),
    .B(_05709_),
    .S(_05439_),
    .Z(_06040_));
 MUX2_X1 _23529_ (.A(_05713_),
    .B(_05718_),
    .S(_05445_),
    .Z(_06041_));
 MUX2_X1 _23530_ (.A(_06040_),
    .B(_06041_),
    .S(_05536_),
    .Z(_06042_));
 AOI221_X1 _23531_ (.A(_06039_),
    .B1(_06042_),
    .B2(_05585_),
    .C1(_05340_),
    .C2(_05562_),
    .ZN(_06043_));
 OR2_X1 _23532_ (.A1(_05596_),
    .A2(_06043_),
    .ZN(_06044_));
 NAND3_X4 _23533_ (.A1(_05887_),
    .A2(_05889_),
    .A3(_05986_),
    .ZN(_06045_));
 INV_X2 _23534_ (.A(_05985_),
    .ZN(_06046_));
 NAND3_X1 _23535_ (.A1(_05982_),
    .A2(_06045_),
    .A3(_06046_),
    .ZN(_06047_));
 AOI21_X2 _23536_ (.A(_16118_),
    .B1(_06047_),
    .B2(_16119_),
    .ZN(_06048_));
 XOR2_X2 _23537_ (.A(_16128_),
    .B(_06048_),
    .Z(_06049_));
 NAND3_X1 _23538_ (.A1(_10912_),
    .A2(_05853_),
    .A3(_06049_),
    .ZN(_06050_));
 OAI21_X1 _23539_ (.A(_00661_),
    .B1(_05884_),
    .B2(_10922_),
    .ZN(_06051_));
 AND3_X1 _23540_ (.A1(_03755_),
    .A2(_06050_),
    .A3(_06051_),
    .ZN(_06052_));
 NOR3_X2 _23541_ (.A1(_04619_),
    .A2(_05401_),
    .A3(_06052_),
    .ZN(_06053_));
 AOI22_X4 _23542_ (.A1(_05897_),
    .A2(_06033_),
    .B1(_06044_),
    .B2(_06053_),
    .ZN(_06054_));
 BUF_X2 _23543_ (.A(_06054_),
    .Z(_06055_));
 MUX2_X1 _23544_ (.A(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .B(_06055_),
    .S(_05498_),
    .Z(_01293_));
 NAND2_X1 _23545_ (.A1(_05362_),
    .A2(_06029_),
    .ZN(_06056_));
 INV_X1 _23546_ (.A(\load_store_unit_i.data_sign_ext_q ),
    .ZN(_06057_));
 OAI21_X4 _23547_ (.A(_05819_),
    .B1(_06056_),
    .B2(_06057_),
    .ZN(_06058_));
 OR2_X1 _23548_ (.A1(_05405_),
    .A2(_06058_),
    .ZN(_06059_));
 BUF_X4 _23549_ (.A(_06059_),
    .Z(_06060_));
 MUX2_X1 _23550_ (.A(\load_store_unit_i.rdata_q[24] ),
    .B(_05374_),
    .S(_05416_),
    .Z(_06061_));
 MUX2_X1 _23551_ (.A(_05771_),
    .B(_06061_),
    .S(_05415_),
    .Z(_06062_));
 BUF_X4 _23552_ (.A(_05827_),
    .Z(_06063_));
 AOI21_X2 _23553_ (.A(_06060_),
    .B1(_06062_),
    .B2(_06063_),
    .ZN(_06064_));
 NOR2_X1 _23554_ (.A1(_16367_),
    .A2(_05449_),
    .ZN(_06065_));
 OAI21_X1 _23555_ (.A(_05161_),
    .B1(_05548_),
    .B2(_16368_),
    .ZN(_06066_));
 AOI221_X2 _23556_ (.A(_06065_),
    .B1(_06066_),
    .B2(_05458_),
    .C1(_05549_),
    .C2(_16371_),
    .ZN(_06067_));
 AOI21_X1 _23557_ (.A(_06067_),
    .B1(_05476_),
    .B2(\alu_adder_result_ex[16] ),
    .ZN(_06068_));
 INV_X1 _23558_ (.A(_06068_),
    .ZN(_06069_));
 AOI221_X2 _23559_ (.A(_06069_),
    .B1(_05474_),
    .B2(_05304_),
    .C1(_05340_),
    .C2(_05585_),
    .ZN(_06070_));
 NAND2_X1 _23560_ (.A1(_05560_),
    .A2(_05250_),
    .ZN(_06071_));
 NAND2_X1 _23561_ (.A1(_05542_),
    .A2(_05474_),
    .ZN(_06072_));
 NAND3_X1 _23562_ (.A1(_05651_),
    .A2(_06071_),
    .A3(_06072_),
    .ZN(_06073_));
 OAI21_X1 _23563_ (.A(_06073_),
    .B1(_06042_),
    .B2(_05651_),
    .ZN(_06074_));
 OAI22_X2 _23564_ (.A1(_05596_),
    .A2(_06070_),
    .B1(_06074_),
    .B2(_05264_),
    .ZN(_06075_));
 AOI21_X1 _23565_ (.A(_04170_),
    .B1(_03800_),
    .B2(_10923_),
    .ZN(_06076_));
 INV_X1 _23566_ (.A(_16132_),
    .ZN(_06077_));
 OR2_X2 _23567_ (.A1(_16119_),
    .A2(_16118_),
    .ZN(_06078_));
 AOI21_X4 _23568_ (.A(_16127_),
    .B1(_06078_),
    .B2(_16128_),
    .ZN(_06079_));
 NOR3_X4 _23569_ (.A1(_16108_),
    .A2(_16118_),
    .A3(_16127_),
    .ZN(_06080_));
 AOI21_X4 _23570_ (.A(_06079_),
    .B1(_06080_),
    .B2(_05987_),
    .ZN(_06081_));
 XNOR2_X2 _23571_ (.A(_06077_),
    .B(_06081_),
    .ZN(_06082_));
 MUX2_X1 _23572_ (.A(_15955_),
    .B(_06082_),
    .S(_05852_),
    .Z(_06083_));
 OAI21_X1 _23573_ (.A(_06076_),
    .B1(_06083_),
    .B2(_03737_),
    .ZN(_06084_));
 NAND2_X1 _23574_ (.A1(_04640_),
    .A2(_06084_),
    .ZN(_06085_));
 NOR3_X2 _23575_ (.A1(_05413_),
    .A2(_06075_),
    .A3(_06085_),
    .ZN(_06086_));
 NOR2_X4 _23576_ (.A1(_06064_),
    .A2(_06086_),
    .ZN(_06087_));
 BUF_X2 _23577_ (.A(_06087_),
    .Z(_06088_));
 MUX2_X1 _23578_ (.A(_06088_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .S(_05738_),
    .Z(_01294_));
 NAND2_X1 _23579_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .A2(_05593_),
    .ZN(_06089_));
 MUX2_X1 _23580_ (.A(\load_store_unit_i.rdata_q[25] ),
    .B(_05808_),
    .S(_05416_),
    .Z(_06090_));
 MUX2_X1 _23581_ (.A(_05807_),
    .B(_06090_),
    .S(_05361_),
    .Z(_06091_));
 AOI21_X1 _23582_ (.A(_06058_),
    .B1(_06091_),
    .B2(_06063_),
    .ZN(_06092_));
 NOR2_X1 _23583_ (.A1(_16375_),
    .A2(_05449_),
    .ZN(_06093_));
 OAI21_X1 _23584_ (.A(_05161_),
    .B1(_05548_),
    .B2(_16376_),
    .ZN(_06094_));
 AOI221_X2 _23585_ (.A(_06093_),
    .B1(_06094_),
    .B2(_05458_),
    .C1(_05455_),
    .C2(_16379_),
    .ZN(_06095_));
 AOI221_X2 _23586_ (.A(_06095_),
    .B1(_05474_),
    .B2(_05304_),
    .C1(\alu_adder_result_ex[17] ),
    .C2(_05476_),
    .ZN(_06096_));
 OAI221_X2 _23587_ (.A(_06096_),
    .B1(_06012_),
    .B2(_05740_),
    .C1(_05252_),
    .C2(_06001_),
    .ZN(_06097_));
 CLKBUF_X2 _23588_ (.A(_16141_),
    .Z(_06098_));
 AND3_X4 _23589_ (.A1(_06045_),
    .A2(_06046_),
    .A3(_06080_),
    .ZN(_06099_));
 NOR3_X1 _23590_ (.A1(_06077_),
    .A2(_06079_),
    .A3(_06099_),
    .ZN(_06100_));
 NOR2_X1 _23591_ (.A1(_16131_),
    .A2(_06100_),
    .ZN(_06101_));
 XOR2_X2 _23592_ (.A(_06098_),
    .B(_06101_),
    .Z(_06102_));
 NAND2_X1 _23593_ (.A1(_05853_),
    .A2(_06102_),
    .ZN(_06103_));
 OAI21_X1 _23594_ (.A(_06103_),
    .B1(_05853_),
    .B2(_15958_),
    .ZN(_06104_));
 NAND2_X1 _23595_ (.A1(_03686_),
    .A2(_06104_),
    .ZN(_06105_));
 AOI21_X1 _23596_ (.A(_04170_),
    .B1(_03940_),
    .B2(_10923_),
    .ZN(_06106_));
 AOI221_X2 _23597_ (.A(_04664_),
    .B1(_05185_),
    .B2(_06097_),
    .C1(_06105_),
    .C2(_06106_),
    .ZN(_06107_));
 MUX2_X2 _23598_ (.A(_06092_),
    .B(_06107_),
    .S(_05734_),
    .Z(_06108_));
 CLKBUF_X3 _23599_ (.A(_06108_),
    .Z(_06109_));
 OAI21_X1 _23600_ (.A(_06089_),
    .B1(_06109_),
    .B2(_05817_),
    .ZN(_01295_));
 MUX2_X1 _23601_ (.A(\load_store_unit_i.rdata_q[26] ),
    .B(_05821_),
    .S(_05416_),
    .Z(_06110_));
 MUX2_X1 _23602_ (.A(_05820_),
    .B(_06110_),
    .S(_05415_),
    .Z(_06111_));
 AOI21_X2 _23603_ (.A(_06060_),
    .B1(_06111_),
    .B2(_06063_),
    .ZN(_06112_));
 BUF_X2 _23604_ (.A(_16147_),
    .Z(_06113_));
 INV_X1 _23605_ (.A(_16140_),
    .ZN(_06114_));
 AND2_X1 _23606_ (.A1(_16132_),
    .A2(_06081_),
    .ZN(_06115_));
 OAI21_X1 _23607_ (.A(_06098_),
    .B1(_16131_),
    .B2(_06115_),
    .ZN(_06116_));
 NAND2_X1 _23608_ (.A1(_06114_),
    .A2(_06116_),
    .ZN(_06117_));
 XNOR2_X2 _23609_ (.A(_06113_),
    .B(_06117_),
    .ZN(_06118_));
 NAND2_X1 _23610_ (.A1(_05428_),
    .A2(_06118_),
    .ZN(_06119_));
 OAI21_X2 _23611_ (.A(_06119_),
    .B1(_05430_),
    .B2(_15967_),
    .ZN(_06120_));
 AOI221_X2 _23612_ (.A(_11865_),
    .B1(_06120_),
    .B2(_03685_),
    .C1(_03944_),
    .C2(net307),
    .ZN(_06121_));
 OR2_X2 _23613_ (.A1(_06121_),
    .A2(_04684_),
    .ZN(_06122_));
 NOR3_X2 _23614_ (.A1(_05256_),
    .A2(_05303_),
    .A3(_05226_),
    .ZN(_06123_));
 NOR2_X1 _23615_ (.A1(_16383_),
    .A2(_05450_),
    .ZN(_06124_));
 OAI21_X1 _23616_ (.A(_05453_),
    .B1(_05455_),
    .B2(_16384_),
    .ZN(_06125_));
 AOI221_X1 _23617_ (.A(_06124_),
    .B1(_06125_),
    .B2(_05459_),
    .C1(_05461_),
    .C2(_16387_),
    .ZN(_06126_));
 OR2_X1 _23618_ (.A1(_06123_),
    .A2(_06126_),
    .ZN(_06127_));
 AOI221_X2 _23619_ (.A(_06127_),
    .B1(_05950_),
    .B2(_05585_),
    .C1(\alu_adder_result_ex[18] ),
    .C2(_05725_),
    .ZN(_06128_));
 OAI21_X1 _23620_ (.A(_06128_),
    .B1(_05955_),
    .B2(_05252_),
    .ZN(_06129_));
 AOI21_X4 _23621_ (.A(_06122_),
    .B1(_06129_),
    .B2(_05427_),
    .ZN(_06130_));
 AOI21_X4 _23622_ (.A(_06112_),
    .B1(_05734_),
    .B2(_06130_),
    .ZN(_06131_));
 BUF_X4 _23623_ (.A(_06131_),
    .Z(_06132_));
 MUX2_X1 _23624_ (.A(_06132_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .S(_05738_),
    .Z(_01296_));
 MUX2_X1 _23625_ (.A(\load_store_unit_i.rdata_q[27] ),
    .B(_05900_),
    .S(_05416_),
    .Z(_06133_));
 MUX2_X1 _23626_ (.A(_05899_),
    .B(_06133_),
    .S(_05415_),
    .Z(_06134_));
 AOI21_X2 _23627_ (.A(_06060_),
    .B1(_06134_),
    .B2(_06063_),
    .ZN(_06135_));
 AOI21_X1 _23628_ (.A(_04171_),
    .B1(_03946_),
    .B2(_10924_),
    .ZN(_06136_));
 NAND3_X1 _23629_ (.A1(_06098_),
    .A2(_06113_),
    .A3(_16131_),
    .ZN(_06137_));
 INV_X1 _23630_ (.A(_06113_),
    .ZN(_06138_));
 OAI21_X2 _23631_ (.A(_06137_),
    .B1(_06114_),
    .B2(_06138_),
    .ZN(_06139_));
 NAND3_X1 _23632_ (.A1(_16132_),
    .A2(_06098_),
    .A3(_06113_),
    .ZN(_06140_));
 NOR3_X4 _23633_ (.A1(_06099_),
    .A2(_06079_),
    .A3(_06140_),
    .ZN(_06141_));
 NOR3_X2 _23634_ (.A1(_16146_),
    .A2(_06139_),
    .A3(_06141_),
    .ZN(_06142_));
 XNOR2_X2 _23635_ (.A(_16153_),
    .B(_06142_),
    .ZN(_06143_));
 CLKBUF_X3 _23636_ (.A(_05852_),
    .Z(_06144_));
 MUX2_X1 _23637_ (.A(_15982_),
    .B(_06143_),
    .S(_06144_),
    .Z(_06145_));
 OAI21_X2 _23638_ (.A(_06136_),
    .B1(_06145_),
    .B2(_03738_),
    .ZN(_06146_));
 NOR2_X1 _23639_ (.A1(_16391_),
    .A2(_05207_),
    .ZN(_06147_));
 OAI21_X1 _23640_ (.A(_05160_),
    .B1(_05209_),
    .B2(_16392_),
    .ZN(_06148_));
 AOI221_X1 _23641_ (.A(_06147_),
    .B1(_06148_),
    .B2(_05204_),
    .C1(_05548_),
    .C2(_16395_),
    .ZN(_06149_));
 AOI21_X1 _23642_ (.A(_06149_),
    .B1(_05476_),
    .B2(\alu_adder_result_ex[19] ),
    .ZN(_06150_));
 NOR2_X1 _23643_ (.A1(_05595_),
    .A2(_06150_),
    .ZN(_06151_));
 OR3_X1 _23644_ (.A1(_04699_),
    .A2(_06123_),
    .A3(_06151_),
    .ZN(_06152_));
 AOI221_X2 _23645_ (.A(_06152_),
    .B1(_05919_),
    .B2(_05585_),
    .C1(_05163_),
    .C2(_05929_),
    .ZN(_06153_));
 AND2_X1 _23646_ (.A1(_05588_),
    .A2(_06153_),
    .ZN(_06154_));
 AOI21_X4 _23647_ (.A(_06135_),
    .B1(_06146_),
    .B2(_06154_),
    .ZN(_06155_));
 BUF_X2 _23648_ (.A(_06155_),
    .Z(_06156_));
 MUX2_X1 _23649_ (.A(_06156_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .S(_05738_),
    .Z(_01297_));
 MUX2_X1 _23650_ (.A(\load_store_unit_i.rdata_q[28] ),
    .B(_05419_),
    .S(_05416_),
    .Z(_06157_));
 MUX2_X1 _23651_ (.A(_05933_),
    .B(_06157_),
    .S(_05415_),
    .Z(_06158_));
 AOI21_X2 _23652_ (.A(_06060_),
    .B1(_06158_),
    .B2(_06063_),
    .ZN(_06159_));
 NOR2_X1 _23653_ (.A1(_10913_),
    .A2(_03948_),
    .ZN(_06160_));
 INV_X1 _23654_ (.A(_16152_),
    .ZN(_06161_));
 AND4_X4 _23655_ (.A1(_16132_),
    .A2(_06098_),
    .A3(_06113_),
    .A4(_06081_),
    .ZN(_06162_));
 NOR3_X1 _23656_ (.A1(_16146_),
    .A2(_06162_),
    .A3(_06139_),
    .ZN(_06163_));
 INV_X1 _23657_ (.A(_16153_),
    .ZN(_06164_));
 OAI21_X1 _23658_ (.A(_06161_),
    .B1(_06163_),
    .B2(_06164_),
    .ZN(_06165_));
 XOR2_X2 _23659_ (.A(_16159_),
    .B(_06165_),
    .Z(_06166_));
 MUX2_X1 _23660_ (.A(_15990_),
    .B(_06166_),
    .S(_05853_),
    .Z(_06167_));
 AOI21_X2 _23661_ (.A(_06160_),
    .B1(_06167_),
    .B2(_10913_),
    .ZN(_06168_));
 OR2_X2 _23662_ (.A1(_04171_),
    .A2(_06168_),
    .ZN(_06169_));
 NAND2_X1 _23663_ (.A1(_04717_),
    .A2(_05405_),
    .ZN(_06170_));
 NOR2_X1 _23664_ (.A1(_16403_),
    .A2(_05451_),
    .ZN(_06171_));
 OAI21_X1 _23665_ (.A(_05454_),
    .B1(_05461_),
    .B2(_16400_),
    .ZN(_06172_));
 AOI221_X2 _23666_ (.A(_06171_),
    .B1(_06172_),
    .B2(_05460_),
    .C1(_05456_),
    .C2(_16399_),
    .ZN(_06173_));
 AOI221_X2 _23667_ (.A(_06173_),
    .B1(_05446_),
    .B2(_05585_),
    .C1(_05304_),
    .C2(_05474_),
    .ZN(_06174_));
 OAI221_X2 _23668_ (.A(_06174_),
    .B1(_05882_),
    .B2(_05252_),
    .C1(net435),
    .C2(_05478_),
    .ZN(_06175_));
 AOI21_X4 _23669_ (.A(_06170_),
    .B1(_06175_),
    .B2(_05427_),
    .ZN(_06176_));
 AOI21_X4 _23670_ (.A(_06159_),
    .B1(_06169_),
    .B2(_06176_),
    .ZN(_06177_));
 BUF_X2 _23671_ (.A(_06177_),
    .Z(_06178_));
 MUX2_X1 _23672_ (.A(_06178_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .S(_05738_),
    .Z(_01298_));
 NAND2_X1 _23673_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .A2(_05593_),
    .ZN(_06179_));
 MUX2_X1 _23674_ (.A(\load_store_unit_i.rdata_q[29] ),
    .B(_05500_),
    .S(_05416_),
    .Z(_06180_));
 MUX2_X1 _23675_ (.A(_05966_),
    .B(_06180_),
    .S(_05415_),
    .Z(_06181_));
 AOI21_X1 _23676_ (.A(_06058_),
    .B1(_06181_),
    .B2(_06063_),
    .ZN(_06182_));
 NAND2_X1 _23677_ (.A1(_05668_),
    .A2(_06182_),
    .ZN(_06183_));
 AOI21_X1 _23678_ (.A(_04171_),
    .B1(_03950_),
    .B2(_10923_),
    .ZN(_06184_));
 NAND2_X1 _23679_ (.A1(_06164_),
    .A2(_06161_),
    .ZN(_06185_));
 AOI21_X4 _23680_ (.A(_16158_),
    .B1(_06185_),
    .B2(_16159_),
    .ZN(_06186_));
 NOR3_X4 _23681_ (.A1(_16146_),
    .A2(_16152_),
    .A3(_16158_),
    .ZN(_06187_));
 NOR2_X4 _23682_ (.A1(_06139_),
    .A2(_06141_),
    .ZN(_06188_));
 AOI21_X4 _23683_ (.A(_06186_),
    .B1(_06188_),
    .B2(_06187_),
    .ZN(_06189_));
 XOR2_X1 _23684_ (.A(_16165_),
    .B(_06189_),
    .Z(_06190_));
 MUX2_X1 _23685_ (.A(_14525_),
    .B(_06190_),
    .S(_05853_),
    .Z(_06191_));
 OAI21_X1 _23686_ (.A(_06184_),
    .B1(_06191_),
    .B2(_10924_),
    .ZN(_06192_));
 NOR2_X1 _23687_ (.A1(_16411_),
    .A2(_05451_),
    .ZN(_06193_));
 OAI21_X1 _23688_ (.A(_05454_),
    .B1(_05462_),
    .B2(_16408_),
    .ZN(_06194_));
 AOI221_X2 _23689_ (.A(_06193_),
    .B1(_06194_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16407_),
    .ZN(_06195_));
 AOI21_X1 _23690_ (.A(_06195_),
    .B1(_05725_),
    .B2(\alu_adder_result_ex[21] ),
    .ZN(_06196_));
 OAI21_X1 _23691_ (.A(_06196_),
    .B1(_05849_),
    .B2(_06013_),
    .ZN(_06197_));
 NAND2_X1 _23692_ (.A1(_05427_),
    .A2(_06197_),
    .ZN(_06198_));
 NOR2_X2 _23693_ (.A1(_05264_),
    .A2(_05739_),
    .ZN(_06199_));
 AOI221_X2 _23694_ (.A(_04741_),
    .B1(_06199_),
    .B2(_05561_),
    .C1(_05865_),
    .C2(_05435_),
    .ZN(_06200_));
 NAND3_X1 _23695_ (.A1(_06192_),
    .A2(_06198_),
    .A3(_06200_),
    .ZN(_06201_));
 OAI21_X2 _23696_ (.A(_06183_),
    .B1(_06201_),
    .B2(_05413_),
    .ZN(_06202_));
 CLKBUF_X3 _23697_ (.A(_06202_),
    .Z(_06203_));
 OAI21_X1 _23698_ (.A(_06179_),
    .B1(_06203_),
    .B2(_05817_),
    .ZN(_01299_));
 NAND2_X1 _23699_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .A2(_05593_),
    .ZN(_06204_));
 OAI21_X1 _23700_ (.A(_06022_),
    .B1(_05655_),
    .B2(_05416_),
    .ZN(_06205_));
 MUX2_X1 _23701_ (.A(\load_store_unit_i.rdata_q[30] ),
    .B(net35),
    .S(_05386_),
    .Z(_06206_));
 MUX2_X1 _23702_ (.A(_06205_),
    .B(_06206_),
    .S(_05360_),
    .Z(_06207_));
 AOI21_X1 _23703_ (.A(_06058_),
    .B1(_06207_),
    .B2(_05827_),
    .ZN(_06208_));
 NOR2_X2 _23704_ (.A1(_05588_),
    .A2(_06208_),
    .ZN(_06209_));
 NOR2_X1 _23705_ (.A1(_05489_),
    .A2(_04760_),
    .ZN(_06210_));
 NOR2_X1 _23706_ (.A1(_05413_),
    .A2(_06210_),
    .ZN(_06211_));
 NOR2_X2 _23707_ (.A1(_05357_),
    .A2(_05427_),
    .ZN(_06212_));
 NOR2_X1 _23708_ (.A1(_16419_),
    .A2(_05449_),
    .ZN(_06213_));
 OAI21_X1 _23709_ (.A(_05161_),
    .B1(_05209_),
    .B2(_16416_),
    .ZN(_06214_));
 AOI221_X2 _23710_ (.A(_06213_),
    .B1(_06214_),
    .B2(_05458_),
    .C1(_05455_),
    .C2(_16415_),
    .ZN(_06215_));
 OR3_X1 _23711_ (.A1(_11282_),
    .A2(_06123_),
    .A3(_06215_),
    .ZN(_06216_));
 AOI221_X1 _23712_ (.A(_06216_),
    .B1(_05650_),
    .B2(_05585_),
    .C1(\alu_adder_result_ex[22] ),
    .C2(_05477_),
    .ZN(_06217_));
 NAND2_X1 _23713_ (.A1(_05562_),
    .A2(_05798_),
    .ZN(_06218_));
 NAND3_X1 _23714_ (.A1(_05272_),
    .A2(_05800_),
    .A3(_05801_),
    .ZN(_06219_));
 AND3_X1 _23715_ (.A1(_06217_),
    .A2(_06218_),
    .A3(_06219_),
    .ZN(_06220_));
 NOR2_X1 _23716_ (.A1(_06144_),
    .A2(_05597_),
    .ZN(_06221_));
 NOR2_X4 _23717_ (.A1(_06162_),
    .A2(_06139_),
    .ZN(_06222_));
 AOI21_X4 _23718_ (.A(_06186_),
    .B1(_06222_),
    .B2(_06187_),
    .ZN(_06223_));
 AOI21_X1 _23719_ (.A(_16164_),
    .B1(_06223_),
    .B2(_16165_),
    .ZN(_06224_));
 XOR2_X1 _23720_ (.A(_16171_),
    .B(_06224_),
    .Z(_06225_));
 NOR2_X1 _23721_ (.A1(_05884_),
    .A2(_06225_),
    .ZN(_06226_));
 NOR3_X4 _23722_ (.A1(_10923_),
    .A2(_06221_),
    .A3(_06226_),
    .ZN(_06227_));
 OAI21_X2 _23723_ (.A(_04176_),
    .B1(_03953_),
    .B2(_10913_),
    .ZN(_06228_));
 OAI22_X4 _23724_ (.A1(_06212_),
    .A2(_06220_),
    .B1(_06227_),
    .B2(_06228_),
    .ZN(_06229_));
 AOI21_X4 _23725_ (.A(_06209_),
    .B1(_06211_),
    .B2(_06229_),
    .ZN(_06230_));
 BUF_X4 _23726_ (.A(_06230_),
    .Z(_06231_));
 OAI21_X1 _23727_ (.A(_06204_),
    .B1(_06231_),
    .B2(_05817_),
    .ZN(_01300_));
 MUX2_X1 _23728_ (.A(\load_store_unit_i.rdata_q[31] ),
    .B(_05674_),
    .S(_05388_),
    .Z(_06232_));
 MUX2_X1 _23729_ (.A(_06028_),
    .B(_06232_),
    .S(_05360_),
    .Z(_06233_));
 AOI21_X1 _23730_ (.A(_06060_),
    .B1(_06233_),
    .B2(_05827_),
    .ZN(_06234_));
 NOR2_X1 _23731_ (.A1(_05357_),
    .A2(_06123_),
    .ZN(_06235_));
 NOR2_X1 _23732_ (.A1(_16423_),
    .A2(_05450_),
    .ZN(_06236_));
 OAI21_X1 _23733_ (.A(_05453_),
    .B1(_05455_),
    .B2(_16424_),
    .ZN(_06237_));
 AOI221_X2 _23734_ (.A(_06236_),
    .B1(_06237_),
    .B2(_05459_),
    .C1(_05461_),
    .C2(_16427_),
    .ZN(_06238_));
 AOI221_X2 _23735_ (.A(_06238_),
    .B1(_05720_),
    .B2(_05257_),
    .C1(net359),
    .C2(_05477_),
    .ZN(_06239_));
 NAND2_X1 _23736_ (.A1(_06235_),
    .A2(_06239_),
    .ZN(_06240_));
 NAND2_X1 _23737_ (.A1(_05651_),
    .A2(_05730_),
    .ZN(_06241_));
 OR2_X1 _23738_ (.A1(_05651_),
    .A2(_05744_),
    .ZN(_06242_));
 AOI21_X1 _23739_ (.A(_05252_),
    .B1(_06241_),
    .B2(_06242_),
    .ZN(_06243_));
 OAI22_X2 _23740_ (.A1(_05357_),
    .A2(_05185_),
    .B1(_06240_),
    .B2(_06243_),
    .ZN(_06244_));
 NAND2_X1 _23741_ (.A1(_05884_),
    .A2(_05686_),
    .ZN(_06245_));
 AOI21_X1 _23742_ (.A(_16164_),
    .B1(_06189_),
    .B2(_16165_),
    .ZN(_06246_));
 INV_X1 _23743_ (.A(_06246_),
    .ZN(_06247_));
 AOI21_X1 _23744_ (.A(_16170_),
    .B1(_06247_),
    .B2(_16171_),
    .ZN(_06248_));
 XNOR2_X1 _23745_ (.A(_06248_),
    .B(_16177_),
    .ZN(_06249_));
 NAND2_X2 _23746_ (.A1(_06249_),
    .A2(_05853_),
    .ZN(_06250_));
 NAND3_X4 _23747_ (.A1(_10913_),
    .A2(_06245_),
    .A3(_06250_),
    .ZN(_06251_));
 AOI21_X1 _23748_ (.A(_04170_),
    .B1(_03955_),
    .B2(_10923_),
    .ZN(_06252_));
 AOI21_X4 _23749_ (.A(_05668_),
    .B1(_06251_),
    .B2(_06252_),
    .ZN(_06253_));
 NOR3_X4 _23750_ (.A1(_04776_),
    .A2(_04781_),
    .A3(_05668_),
    .ZN(_06254_));
 AOI221_X2 _23751_ (.A(_06234_),
    .B1(_06253_),
    .B2(_06244_),
    .C1(_06254_),
    .C2(_05357_),
    .ZN(_06255_));
 BUF_X8 _23752_ (.A(net461),
    .Z(_06256_));
 MUX2_X1 _23753_ (.A(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .B(_06256_),
    .S(_05498_),
    .Z(_01301_));
 MUX2_X1 _23754_ (.A(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .B(_05909_),
    .S(_05412_),
    .Z(_01302_));
 NAND2_X1 _23755_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .A2(_05593_),
    .ZN(_06257_));
 MUX2_X1 _23756_ (.A(net45),
    .B(_05374_),
    .S(_05386_),
    .Z(_06258_));
 MUX2_X1 _23757_ (.A(net34),
    .B(net36),
    .S(_05386_),
    .Z(_06259_));
 MUX2_X1 _23758_ (.A(_06258_),
    .B(_06259_),
    .S(_05360_),
    .Z(_06260_));
 AOI21_X1 _23759_ (.A(_06058_),
    .B1(_06260_),
    .B2(_05827_),
    .ZN(_06261_));
 NOR2_X2 _23760_ (.A1(_05588_),
    .A2(_06261_),
    .ZN(_06262_));
 AOI21_X2 _23761_ (.A(_05401_),
    .B1(_04801_),
    .B2(_05357_),
    .ZN(_06263_));
 INV_X1 _23762_ (.A(_16183_),
    .ZN(_06264_));
 INV_X1 _23763_ (.A(_16176_),
    .ZN(_06265_));
 AOI21_X2 _23764_ (.A(_16170_),
    .B1(_16171_),
    .B2(_16164_),
    .ZN(_06266_));
 INV_X1 _23765_ (.A(_16177_),
    .ZN(_06267_));
 OAI21_X2 _23766_ (.A(_06265_),
    .B1(_06266_),
    .B2(_06267_),
    .ZN(_06268_));
 AND3_X1 _23767_ (.A1(_16165_),
    .A2(_16171_),
    .A3(_16177_),
    .ZN(_06269_));
 AOI21_X4 _23768_ (.A(_06268_),
    .B1(_06269_),
    .B2(_06223_),
    .ZN(_06270_));
 XNOR2_X1 _23769_ (.A(_06264_),
    .B(_06270_),
    .ZN(_06271_));
 MUX2_X1 _23770_ (.A(_05754_),
    .B(_06271_),
    .S(_05853_),
    .Z(_06272_));
 NAND2_X1 _23771_ (.A1(_03686_),
    .A2(_06272_),
    .ZN(_06273_));
 AOI21_X1 _23772_ (.A(_04171_),
    .B1(_03957_),
    .B2(_10923_),
    .ZN(_06274_));
 NAND2_X1 _23773_ (.A1(_06273_),
    .A2(_06274_),
    .ZN(_06275_));
 AND2_X1 _23774_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_05476_),
    .ZN(_06276_));
 NOR2_X1 _23775_ (.A1(_16431_),
    .A2(_05450_),
    .ZN(_06277_));
 OAI21_X1 _23776_ (.A(_05453_),
    .B1(_05455_),
    .B2(_16432_),
    .ZN(_06278_));
 AOI221_X2 _23777_ (.A(_06277_),
    .B1(_06278_),
    .B2(_05459_),
    .C1(_05461_),
    .C2(_16435_),
    .ZN(_06279_));
 OR4_X1 _23778_ (.A1(_11282_),
    .A2(_06123_),
    .A3(_06276_),
    .A4(_06279_),
    .ZN(_06280_));
 AOI221_X2 _23779_ (.A(_06280_),
    .B1(_05730_),
    .B2(_05585_),
    .C1(_05163_),
    .C2(_05721_),
    .ZN(_06281_));
 OAI21_X2 _23780_ (.A(_06275_),
    .B1(_06281_),
    .B2(_06212_),
    .ZN(_06282_));
 AOI21_X4 _23781_ (.A(_06262_),
    .B1(_06263_),
    .B2(_06282_),
    .ZN(_06283_));
 CLKBUF_X3 _23782_ (.A(_06283_),
    .Z(_06284_));
 OAI21_X1 _23783_ (.A(_06257_),
    .B1(_06284_),
    .B2(_05817_),
    .ZN(_01303_));
 NAND2_X1 _23784_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .A2(_05593_),
    .ZN(_06285_));
 MUX2_X1 _23785_ (.A(net46),
    .B(_05808_),
    .S(_05387_),
    .Z(_06286_));
 MUX2_X1 _23786_ (.A(net40),
    .B(net37),
    .S(_05387_),
    .Z(_06287_));
 MUX2_X1 _23787_ (.A(_06286_),
    .B(_06287_),
    .S(_05361_),
    .Z(_06288_));
 AOI21_X1 _23788_ (.A(_06060_),
    .B1(_06288_),
    .B2(_06063_),
    .ZN(_06289_));
 OR2_X1 _23789_ (.A1(_05489_),
    .A2(_04821_),
    .ZN(_06290_));
 NOR2_X1 _23790_ (.A1(_16439_),
    .A2(_05449_),
    .ZN(_06291_));
 OAI21_X1 _23791_ (.A(_05160_),
    .B1(_05209_),
    .B2(_16440_),
    .ZN(_06292_));
 AOI221_X2 _23792_ (.A(_06291_),
    .B1(_06292_),
    .B2(_05458_),
    .C1(_05548_),
    .C2(_16443_),
    .ZN(_06293_));
 AOI221_X2 _23793_ (.A(_06293_),
    .B1(_05476_),
    .B2(\alu_adder_result_ex[25] ),
    .C1(_10971_),
    .C2(_10972_),
    .ZN(_06294_));
 OAI21_X1 _23794_ (.A(_05435_),
    .B1(_05222_),
    .B2(_05474_),
    .ZN(_06295_));
 OAI21_X1 _23795_ (.A(_06294_),
    .B1(_06295_),
    .B2(_05624_),
    .ZN(_06296_));
 AOI221_X2 _23796_ (.A(_06296_),
    .B1(_05643_),
    .B2(_05727_),
    .C1(_06199_),
    .C2(_05650_),
    .ZN(_06297_));
 AND2_X1 _23797_ (.A1(_03959_),
    .A2(_03684_),
    .ZN(_06298_));
 NOR2_X1 _23798_ (.A1(_05430_),
    .A2(_05784_),
    .ZN(_06299_));
 INV_X1 _23799_ (.A(_16189_),
    .ZN(_06300_));
 INV_X1 _23800_ (.A(_16182_),
    .ZN(_06301_));
 AOI21_X2 _23801_ (.A(_06268_),
    .B1(_06189_),
    .B2(_06269_),
    .ZN(_06302_));
 OAI21_X2 _23802_ (.A(_06301_),
    .B1(_06264_),
    .B2(_06302_),
    .ZN(_06303_));
 XNOR2_X2 _23803_ (.A(_06303_),
    .B(_06300_),
    .ZN(_06304_));
 AOI211_X2 _23804_ (.A(_10922_),
    .B(_06299_),
    .C1(_05852_),
    .C2(_06304_),
    .ZN(_06305_));
 OR2_X2 _23805_ (.A1(_06305_),
    .A2(_04170_),
    .ZN(_06306_));
 OAI22_X4 _23806_ (.A1(_06212_),
    .A2(_06297_),
    .B1(_06306_),
    .B2(_06298_),
    .ZN(_06307_));
 AOI21_X4 _23807_ (.A(_05413_),
    .B1(_06307_),
    .B2(_06290_),
    .ZN(_06308_));
 OR2_X4 _23808_ (.A1(_06308_),
    .A2(_06289_),
    .ZN(_06309_));
 BUF_X16 _23809_ (.A(_06309_),
    .Z(_06310_));
 OAI21_X2 _23810_ (.A(_06285_),
    .B1(net488),
    .B2(_05817_),
    .ZN(_01304_));
 MUX2_X1 _23811_ (.A(net51),
    .B(net38),
    .S(_05898_),
    .Z(_06311_));
 MUX2_X1 _23812_ (.A(net47),
    .B(_05821_),
    .S(_05416_),
    .Z(_06312_));
 MUX2_X1 _23813_ (.A(_06311_),
    .B(_06312_),
    .S(_05902_),
    .Z(_06313_));
 AOI21_X2 _23814_ (.A(_06060_),
    .B1(_06313_),
    .B2(_06063_),
    .ZN(_06314_));
 OAI21_X4 _23815_ (.A(_06301_),
    .B1(_06270_),
    .B2(_06264_),
    .ZN(_06315_));
 AOI21_X2 _23816_ (.A(_16188_),
    .B1(_06315_),
    .B2(_16189_),
    .ZN(_06316_));
 XNOR2_X1 _23817_ (.A(_16195_),
    .B(_06316_),
    .ZN(_06317_));
 MUX2_X1 _23818_ (.A(_05858_),
    .B(_06317_),
    .S(_06144_),
    .Z(_06318_));
 OAI221_X2 _23819_ (.A(_04176_),
    .B1(_03736_),
    .B2(_03961_),
    .C1(_06318_),
    .C2(_10924_),
    .ZN(_06319_));
 NOR2_X1 _23820_ (.A1(_16447_),
    .A2(_05449_),
    .ZN(_06320_));
 OAI21_X1 _23821_ (.A(_05161_),
    .B1(_05548_),
    .B2(_16448_),
    .ZN(_06321_));
 AOI221_X2 _23822_ (.A(_06320_),
    .B1(_06321_),
    .B2(_05458_),
    .C1(_05549_),
    .C2(_16451_),
    .ZN(_06322_));
 OR2_X1 _23823_ (.A1(_06123_),
    .A2(_06322_),
    .ZN(_06323_));
 AOI221_X2 _23824_ (.A(_06323_),
    .B1(_05562_),
    .B2(_05584_),
    .C1(\alu_adder_result_ex[26] ),
    .C2(_05725_),
    .ZN(_06324_));
 AOI22_X1 _23825_ (.A1(_05543_),
    .A2(_06199_),
    .B1(_05561_),
    .B2(_05585_),
    .ZN(_06325_));
 AOI21_X1 _23826_ (.A(_05596_),
    .B1(_06324_),
    .B2(_06325_),
    .ZN(_06326_));
 NOR3_X2 _23827_ (.A1(_04836_),
    .A2(_05401_),
    .A3(_06326_),
    .ZN(_06327_));
 AOI21_X4 _23828_ (.A(_06314_),
    .B1(_06319_),
    .B2(_06327_),
    .ZN(_06328_));
 BUF_X4 _23829_ (.A(_06328_),
    .Z(_06329_));
 MUX2_X1 _23830_ (.A(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .B(_06329_),
    .S(_05497_),
    .Z(_01305_));
 NAND2_X1 _23831_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .A2(_05593_),
    .ZN(_06330_));
 MUX2_X1 _23832_ (.A(net54),
    .B(net39),
    .S(_05386_),
    .Z(_06331_));
 MUX2_X1 _23833_ (.A(net48),
    .B(_05900_),
    .S(_05386_),
    .Z(_06332_));
 MUX2_X1 _23834_ (.A(_06331_),
    .B(_06332_),
    .S(_05902_),
    .Z(_06333_));
 AOI21_X1 _23835_ (.A(_06058_),
    .B1(_06333_),
    .B2(_05827_),
    .ZN(_06334_));
 NOR2_X1 _23836_ (.A1(_05588_),
    .A2(_06334_),
    .ZN(_06335_));
 NOR2_X1 _23837_ (.A1(_05489_),
    .A2(_04851_),
    .ZN(_06336_));
 NOR2_X2 _23838_ (.A1(_05413_),
    .A2(_06336_),
    .ZN(_06337_));
 BUF_X1 _23839_ (.A(_16201_),
    .Z(_06338_));
 INV_X1 _23840_ (.A(_16188_),
    .ZN(_06339_));
 AOI21_X1 _23841_ (.A(_16182_),
    .B1(_06268_),
    .B2(_16183_),
    .ZN(_06340_));
 OAI21_X1 _23842_ (.A(_06339_),
    .B1(_06340_),
    .B2(_06300_),
    .ZN(_06341_));
 AOI21_X1 _23843_ (.A(_16194_),
    .B1(_06341_),
    .B2(_16195_),
    .ZN(_06342_));
 INV_X1 _23844_ (.A(_06342_),
    .ZN(_06343_));
 NAND2_X1 _23845_ (.A1(_16195_),
    .A2(_06269_),
    .ZN(_06344_));
 OAI21_X1 _23846_ (.A(_16189_),
    .B1(_16182_),
    .B2(_16183_),
    .ZN(_06345_));
 AOI21_X2 _23847_ (.A(_06344_),
    .B1(_06345_),
    .B2(_06339_),
    .ZN(_06346_));
 AOI21_X1 _23848_ (.A(_06343_),
    .B1(_06346_),
    .B2(_06189_),
    .ZN(_06347_));
 XNOR2_X1 _23849_ (.A(_06338_),
    .B(_06347_),
    .ZN(_06348_));
 NAND2_X1 _23850_ (.A1(_06144_),
    .A2(_06348_),
    .ZN(_06349_));
 AOI21_X1 _23851_ (.A(_10923_),
    .B1(_05884_),
    .B2(_05891_),
    .ZN(_06350_));
 AOI21_X2 _23852_ (.A(_04170_),
    .B1(_06349_),
    .B2(_06350_),
    .ZN(_06351_));
 OAI21_X1 _23853_ (.A(_06351_),
    .B1(_03736_),
    .B2(_03964_),
    .ZN(_06352_));
 NOR2_X1 _23854_ (.A1(_16455_),
    .A2(_05450_),
    .ZN(_06353_));
 OAI21_X1 _23855_ (.A(_05453_),
    .B1(_05549_),
    .B2(_16456_),
    .ZN(_06354_));
 AOI221_X2 _23856_ (.A(_06353_),
    .B1(_06354_),
    .B2(_05459_),
    .C1(_05456_),
    .C2(_16459_),
    .ZN(_06355_));
 AOI21_X1 _23857_ (.A(_06355_),
    .B1(_05725_),
    .B2(\alu_adder_result_ex[27] ),
    .ZN(_06356_));
 OAI21_X1 _23858_ (.A(_06356_),
    .B1(_06295_),
    .B2(_05473_),
    .ZN(_06357_));
 AOI221_X2 _23859_ (.A(_05357_),
    .B1(_05163_),
    .B2(_05447_),
    .C1(_06357_),
    .C2(_05185_),
    .ZN(_06358_));
 NAND2_X1 _23860_ (.A1(_06352_),
    .A2(_06358_),
    .ZN(_06359_));
 AOI21_X4 _23861_ (.A(_06335_),
    .B1(_06337_),
    .B2(_06359_),
    .ZN(_06360_));
 BUF_X4 _23862_ (.A(_06360_),
    .Z(_06361_));
 OAI21_X1 _23863_ (.A(_06330_),
    .B1(_06361_),
    .B2(_05817_),
    .ZN(_01306_));
 NAND2_X1 _23864_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .A2(_05593_),
    .ZN(_06362_));
 NAND2_X1 _23865_ (.A1(_05417_),
    .A2(_05422_),
    .ZN(_06363_));
 MUX2_X1 _23866_ (.A(net49),
    .B(_05419_),
    .S(_05416_),
    .Z(_06364_));
 MUX2_X1 _23867_ (.A(_06363_),
    .B(_06364_),
    .S(_05902_),
    .Z(_06365_));
 AOI21_X1 _23868_ (.A(_06058_),
    .B1(_06365_),
    .B2(_06063_),
    .ZN(_06366_));
 NOR2_X1 _23869_ (.A1(_05339_),
    .A2(_05711_),
    .ZN(_06367_));
 MUX2_X1 _23870_ (.A(_16449_),
    .B(_16281_),
    .S(_05264_),
    .Z(_06368_));
 MUX2_X1 _23871_ (.A(_06368_),
    .B(_05277_),
    .S(_05271_),
    .Z(_06369_));
 MUX2_X1 _23872_ (.A(_05262_),
    .B(_06369_),
    .S(_11173_),
    .Z(_06370_));
 AOI21_X1 _23873_ (.A(_06367_),
    .B1(_06370_),
    .B2(_05536_),
    .ZN(_06371_));
 MUX2_X1 _23874_ (.A(_05880_),
    .B(_06371_),
    .S(_05560_),
    .Z(_06372_));
 AOI22_X2 _23875_ (.A1(_06006_),
    .A2(_05919_),
    .B1(_06372_),
    .B2(_05562_),
    .ZN(_06373_));
 INV_X1 _23876_ (.A(_16207_),
    .ZN(_06374_));
 AND2_X1 _23877_ (.A1(_06338_),
    .A2(_06346_),
    .ZN(_06375_));
 AOI221_X2 _23878_ (.A(_16200_),
    .B1(_06223_),
    .B2(_06375_),
    .C1(_06343_),
    .C2(_06338_),
    .ZN(_06376_));
 XNOR2_X1 _23879_ (.A(_06374_),
    .B(_06376_),
    .ZN(_06377_));
 MUX2_X1 _23880_ (.A(_05914_),
    .B(_06377_),
    .S(_05852_),
    .Z(_06378_));
 AOI21_X4 _23881_ (.A(_04170_),
    .B1(_06378_),
    .B2(_10913_),
    .ZN(_06379_));
 NAND2_X1 _23882_ (.A1(_03967_),
    .A2(_03684_),
    .ZN(_06380_));
 NOR2_X1 _23883_ (.A1(_16463_),
    .A2(_05451_),
    .ZN(_06381_));
 OAI21_X1 _23884_ (.A(_05454_),
    .B1(_05461_),
    .B2(_16464_),
    .ZN(_06382_));
 AOI221_X2 _23885_ (.A(_06381_),
    .B1(_06382_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16467_),
    .ZN(_06383_));
 AOI21_X1 _23886_ (.A(_06383_),
    .B1(_05725_),
    .B2(\alu_adder_result_ex[28] ),
    .ZN(_06384_));
 NAND3_X1 _23887_ (.A1(_05248_),
    .A2(_05305_),
    .A3(_05303_),
    .ZN(_06385_));
 MUX2_X1 _23888_ (.A(_05321_),
    .B(_05226_),
    .S(_06385_),
    .Z(_06386_));
 OAI21_X1 _23889_ (.A(_06384_),
    .B1(_06386_),
    .B2(_05256_),
    .ZN(_06387_));
 AOI22_X2 _23890_ (.A1(_06379_),
    .A2(_06380_),
    .B1(_06387_),
    .B2(_05427_),
    .ZN(_06388_));
 NAND3_X1 _23891_ (.A1(_05489_),
    .A2(_06373_),
    .A3(_06388_),
    .ZN(_06389_));
 OAI21_X1 _23892_ (.A(_06389_),
    .B1(_04866_),
    .B2(_05489_),
    .ZN(_06390_));
 MUX2_X2 _23893_ (.A(_06366_),
    .B(_06390_),
    .S(_05734_),
    .Z(_06391_));
 BUF_X4 _23894_ (.A(_06391_),
    .Z(_06392_));
 OAI21_X1 _23895_ (.A(_06362_),
    .B1(_06392_),
    .B2(_05817_),
    .ZN(_01307_));
 OAI21_X1 _23896_ (.A(_05507_),
    .B1(_05501_),
    .B2(_05378_),
    .ZN(_06393_));
 MUX2_X1 _23897_ (.A(net50),
    .B(_05500_),
    .S(_05898_),
    .Z(_06394_));
 MUX2_X1 _23898_ (.A(_06393_),
    .B(_06394_),
    .S(_05902_),
    .Z(_06395_));
 AOI21_X1 _23899_ (.A(_06060_),
    .B1(_06395_),
    .B2(_05827_),
    .ZN(_06396_));
 NOR2_X1 _23900_ (.A1(_16471_),
    .A2(_05207_),
    .ZN(_06397_));
 OAI21_X1 _23901_ (.A(_05160_),
    .B1(_05209_),
    .B2(_16472_),
    .ZN(_06398_));
 AOI221_X2 _23902_ (.A(_06397_),
    .B1(_06398_),
    .B2(_05204_),
    .C1(_05548_),
    .C2(_16475_),
    .ZN(_06399_));
 MUX2_X1 _23903_ (.A(_05539_),
    .B(_05225_),
    .S(_06385_),
    .Z(_06400_));
 AOI221_X1 _23904_ (.A(_06399_),
    .B1(_06400_),
    .B2(_05435_),
    .C1(\alu_adder_result_ex[29] ),
    .C2(_05476_),
    .ZN(_06401_));
 NOR2_X1 _23905_ (.A1(_05595_),
    .A2(_06401_),
    .ZN(_06402_));
 OR2_X1 _23906_ (.A1(_04884_),
    .A2(_06402_),
    .ZN(_06403_));
 AOI21_X2 _23907_ (.A(_04170_),
    .B1(_01095_),
    .B2(net307),
    .ZN(_06404_));
 AND4_X4 _23908_ (.A1(_06338_),
    .A2(_16207_),
    .A3(_06189_),
    .A4(_06346_),
    .ZN(_06405_));
 NAND3_X1 _23909_ (.A1(_06338_),
    .A2(_16207_),
    .A3(_06343_),
    .ZN(_06406_));
 INV_X1 _23910_ (.A(_16200_),
    .ZN(_06407_));
 OAI21_X1 _23911_ (.A(_06406_),
    .B1(_06407_),
    .B2(_06374_),
    .ZN(_06408_));
 NOR3_X2 _23912_ (.A1(_16206_),
    .A2(_06405_),
    .A3(_06408_),
    .ZN(_06409_));
 XOR2_X1 _23913_ (.A(_06409_),
    .B(_16213_),
    .Z(_06410_));
 MUX2_X1 _23914_ (.A(_05961_),
    .B(_06410_),
    .S(_05430_),
    .Z(_06411_));
 NAND2_X2 _23915_ (.A1(_03686_),
    .A2(_06411_),
    .ZN(_06412_));
 NOR2_X1 _23916_ (.A1(_05626_),
    .A2(_05629_),
    .ZN(_06413_));
 MUX2_X1 _23917_ (.A(_06413_),
    .B(_05641_),
    .S(_05229_),
    .Z(_06414_));
 NAND2_X1 _23918_ (.A1(_11170_),
    .A2(_05265_),
    .ZN(_06415_));
 OAI21_X1 _23919_ (.A(_06415_),
    .B1(_05259_),
    .B2(_11170_),
    .ZN(_06416_));
 MUX2_X1 _23920_ (.A(_05278_),
    .B(_06416_),
    .S(_05240_),
    .Z(_06417_));
 MUX2_X1 _23921_ (.A(_05638_),
    .B(_06417_),
    .S(_05248_),
    .Z(_06418_));
 MUX2_X1 _23922_ (.A(_06414_),
    .B(_06418_),
    .S(_05439_),
    .Z(_06419_));
 MUX2_X1 _23923_ (.A(_05950_),
    .B(_06419_),
    .S(_05739_),
    .Z(_06420_));
 AOI221_X2 _23924_ (.A(_06403_),
    .B1(_06412_),
    .B2(_06404_),
    .C1(_06420_),
    .C2(_05163_),
    .ZN(_06421_));
 AOI21_X4 _23925_ (.A(_06396_),
    .B1(_05734_),
    .B2(_06421_),
    .ZN(_06422_));
 BUF_X4 _23926_ (.A(_06422_),
    .Z(_06423_));
 MUX2_X1 _23927_ (.A(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .B(net458),
    .S(_05497_),
    .Z(_01308_));
 NAND2_X1 _23928_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .A2(_05593_),
    .ZN(_06424_));
 OAI21_X1 _23929_ (.A(_03686_),
    .B1(_05853_),
    .B2(_05989_),
    .ZN(_06425_));
 INV_X1 _23930_ (.A(_16206_),
    .ZN(_06426_));
 OAI21_X2 _23931_ (.A(_06426_),
    .B1(_06376_),
    .B2(_06374_),
    .ZN(_06427_));
 AOI21_X4 _23932_ (.A(_16212_),
    .B1(_16213_),
    .B2(_06427_),
    .ZN(_06428_));
 XNOR2_X2 _23933_ (.A(_16219_),
    .B(_06428_),
    .ZN(_06429_));
 AOI21_X4 _23934_ (.A(_06425_),
    .B1(_06429_),
    .B2(_06144_),
    .ZN(_06430_));
 AND2_X1 _23935_ (.A1(_10923_),
    .A2(_03971_),
    .ZN(_06431_));
 NOR3_X4 _23936_ (.A1(_06430_),
    .A2(_04171_),
    .A3(_06431_),
    .ZN(_06432_));
 NOR2_X1 _23937_ (.A1(_16483_),
    .A2(_05451_),
    .ZN(_06433_));
 OAI21_X1 _23938_ (.A(_05454_),
    .B1(_05461_),
    .B2(_16480_),
    .ZN(_06434_));
 AOI221_X2 _23939_ (.A(_06433_),
    .B1(_06434_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16479_),
    .ZN(_06435_));
 MUX2_X1 _23940_ (.A(_05474_),
    .B(_05644_),
    .S(_05222_),
    .Z(_06436_));
 AOI221_X2 _23941_ (.A(_06435_),
    .B1(_06436_),
    .B2(_05435_),
    .C1(_05725_),
    .C2(net345),
    .ZN(_06437_));
 NOR2_X1 _23942_ (.A1(_05596_),
    .A2(_06437_),
    .ZN(_06438_));
 AOI21_X1 _23943_ (.A(_05439_),
    .B1(_05570_),
    .B2(_05572_),
    .ZN(_06439_));
 AOI21_X1 _23944_ (.A(_06439_),
    .B1(_05582_),
    .B2(_05440_),
    .ZN(_06440_));
 OAI21_X1 _23945_ (.A(_16242_),
    .B1(_16469_),
    .B2(_05274_),
    .ZN(_06441_));
 OAI221_X1 _23946_ (.A(_05271_),
    .B1(_05273_),
    .B2(_06441_),
    .C1(_05280_),
    .C2(_16242_),
    .ZN(_06442_));
 NOR2_X1 _23947_ (.A1(_16261_),
    .A2(_05272_),
    .ZN(_06443_));
 OAI21_X1 _23948_ (.A(_11173_),
    .B1(_16461_),
    .B2(_05274_),
    .ZN(_06444_));
 OAI221_X1 _23949_ (.A(_05240_),
    .B1(_06443_),
    .B2(_06444_),
    .C1(_05259_),
    .C2(_11173_),
    .ZN(_06445_));
 AND3_X1 _23950_ (.A1(_05439_),
    .A2(_06442_),
    .A3(_06445_),
    .ZN(_06446_));
 AOI21_X1 _23951_ (.A(_06446_),
    .B1(_05579_),
    .B2(_05445_),
    .ZN(_06447_));
 MUX2_X1 _23952_ (.A(_06440_),
    .B(_06447_),
    .S(_05536_),
    .Z(_06448_));
 MUX2_X1 _23953_ (.A(_06012_),
    .B(_06448_),
    .S(_05739_),
    .Z(_06449_));
 OAI21_X1 _23954_ (.A(_04901_),
    .B1(_05252_),
    .B2(_06449_),
    .ZN(_06450_));
 NOR4_X4 _23955_ (.A1(_06432_),
    .A2(_05413_),
    .A3(_06438_),
    .A4(_06450_),
    .ZN(_06451_));
 OAI21_X1 _23956_ (.A(_05660_),
    .B1(_05655_),
    .B2(_05378_),
    .ZN(_06452_));
 MUX2_X1 _23957_ (.A(net52),
    .B(net35),
    .S(_05387_),
    .Z(_06453_));
 MUX2_X1 _23958_ (.A(_06452_),
    .B(_06453_),
    .S(_05902_),
    .Z(_06454_));
 AOI21_X1 _23959_ (.A(_06060_),
    .B1(_06454_),
    .B2(_06063_),
    .ZN(_06455_));
 OR2_X4 _23960_ (.A1(_06455_),
    .A2(_06451_),
    .ZN(_06456_));
 BUF_X16 _23961_ (.A(_06456_),
    .Z(_06457_));
 OAI21_X4 _23962_ (.A(_06424_),
    .B1(net457),
    .B2(_05817_),
    .ZN(_01309_));
 NAND2_X1 _23963_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A2(_05592_),
    .ZN(_06458_));
 NOR3_X1 _23964_ (.A1(_16213_),
    .A2(_16212_),
    .A3(_16218_),
    .ZN(_06459_));
 NOR3_X1 _23965_ (.A1(_16206_),
    .A2(_16212_),
    .A3(_16218_),
    .ZN(_06460_));
 NOR2_X4 _23966_ (.A1(_06405_),
    .A2(_06408_),
    .ZN(_06461_));
 INV_X1 _23967_ (.A(_16219_),
    .ZN(_06462_));
 INV_X1 _23968_ (.A(_16218_),
    .ZN(_06463_));
 AOI221_X2 _23969_ (.A(_06459_),
    .B1(_06461_),
    .B2(_06460_),
    .C1(_06462_),
    .C2(_06463_),
    .ZN(_06464_));
 XNOR2_X1 _23970_ (.A(_06464_),
    .B(_16225_),
    .ZN(_06465_));
 MUX2_X1 _23971_ (.A(_06049_),
    .B(_06465_),
    .S(_05430_),
    .Z(_06466_));
 AOI221_X2 _23972_ (.A(_04170_),
    .B1(_06466_),
    .B2(_03685_),
    .C1(_03503_),
    .C2(net307),
    .ZN(_06467_));
 NOR2_X1 _23973_ (.A1(_15899_),
    .A2(_05450_),
    .ZN(_06468_));
 OAI21_X1 _23974_ (.A(_05453_),
    .B1(_05549_),
    .B2(_15896_),
    .ZN(_06469_));
 AOI221_X2 _23975_ (.A(_06468_),
    .B1(_06469_),
    .B2(_05459_),
    .C1(_05456_),
    .C2(_15895_),
    .ZN(_06470_));
 INV_X1 _23976_ (.A(_06470_),
    .ZN(_06471_));
 OAI21_X1 _23977_ (.A(_06471_),
    .B1(_05251_),
    .B2(_05256_),
    .ZN(_06472_));
 AOI21_X1 _23978_ (.A(_06472_),
    .B1(_05562_),
    .B2(_05302_),
    .ZN(_06473_));
 AOI22_X2 _23979_ (.A1(net289),
    .A2(_05725_),
    .B1(_06006_),
    .B2(_05340_),
    .ZN(_06474_));
 AOI21_X2 _23980_ (.A(_05596_),
    .B1(_06473_),
    .B2(_06474_),
    .ZN(_06475_));
 NOR4_X4 _23981_ (.A1(_04922_),
    .A2(_05401_),
    .A3(_06467_),
    .A4(_06475_),
    .ZN(_06476_));
 BUF_X16 _23982_ (.A(net372),
    .Z(_06477_));
 MUX2_X1 _23983_ (.A(net53),
    .B(_05674_),
    .S(_05387_),
    .Z(_06478_));
 NOR2_X1 _23984_ (.A1(_05361_),
    .A2(_06478_),
    .ZN(_06479_));
 NOR2_X1 _23985_ (.A1(_05902_),
    .A2(_05768_),
    .ZN(_06480_));
 NOR3_X1 _23986_ (.A1(_05376_),
    .A2(_06479_),
    .A3(_06480_),
    .ZN(_06481_));
 OR2_X2 _23987_ (.A1(_06060_),
    .A2(_06481_),
    .ZN(_06482_));
 CLKBUF_X3 _23988_ (.A(_06482_),
    .Z(_06483_));
 NAND2_X1 _23989_ (.A1(_05498_),
    .A2(_06483_),
    .ZN(_06484_));
 OAI21_X2 _23990_ (.A(_06458_),
    .B1(net314),
    .B2(_06484_),
    .ZN(_01310_));
 AND2_X1 _23991_ (.A1(_05410_),
    .A2(_05494_),
    .ZN(_06485_));
 CLKBUF_X3 _23992_ (.A(_06485_),
    .Z(_06486_));
 BUF_X4 _23993_ (.A(_06486_),
    .Z(_06487_));
 MUX2_X1 _23994_ (.A(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .B(_05403_),
    .S(_06487_),
    .Z(_01311_));
 NAND2_X1 _23995_ (.A1(_15958_),
    .A2(_05430_),
    .ZN(_06488_));
 OAI21_X1 _23996_ (.A(_06488_),
    .B1(_05852_),
    .B2(_00185_),
    .ZN(_06489_));
 NOR2_X1 _23997_ (.A1(_03737_),
    .A2(_06489_),
    .ZN(_06490_));
 OAI21_X1 _23998_ (.A(_03755_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .B2(_10912_),
    .ZN(_06491_));
 OAI21_X2 _23999_ (.A(_10973_),
    .B1(_06490_),
    .B2(_06491_),
    .ZN(_06492_));
 CLKBUF_X2 _24000_ (.A(\cs_registers_i.mhpmcounter[2][33] ),
    .Z(_06493_));
 AOI22_X1 _24001_ (.A1(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .A2(_04499_),
    .B1(_04392_),
    .B2(_06493_),
    .ZN(_06494_));
 NOR2_X1 _24002_ (.A1(_04380_),
    .A2(_06494_),
    .ZN(_06495_));
 AOI22_X1 _24003_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(_04589_),
    .B1(_04591_),
    .B2(\cs_registers_i.mhpmcounter[2][1] ),
    .ZN(_06496_));
 INV_X1 _24004_ (.A(_06496_),
    .ZN(_06497_));
 NOR2_X2 _24005_ (.A1(_03578_),
    .A2(_04400_),
    .ZN(_06498_));
 NAND4_X2 _24006_ (.A1(_16282_),
    .A2(_04373_),
    .A3(_04398_),
    .A4(_03607_),
    .ZN(_06499_));
 NOR2_X4 _24007_ (.A1(_06498_),
    .A2(_06499_),
    .ZN(_06500_));
 AOI21_X2 _24008_ (.A(_06495_),
    .B1(_06497_),
    .B2(_06500_),
    .ZN(_06501_));
 AOI222_X2 _24009_ (.A1(\cs_registers_i.dscratch0_q[1] ),
    .A2(_04417_),
    .B1(_04433_),
    .B2(\cs_registers_i.dcsr_q[1] ),
    .C1(_04559_),
    .C2(\cs_registers_i.mscratch_q[1] ),
    .ZN(_06502_));
 NAND2_X1 _24010_ (.A1(\cs_registers_i.mcause_q[1] ),
    .A2(_04918_),
    .ZN(_06503_));
 OAI21_X1 _24011_ (.A(_06503_),
    .B1(_05609_),
    .B2(_00555_),
    .ZN(_06504_));
 AOI221_X2 _24012_ (.A(_06504_),
    .B1(_04637_),
    .B2(net72),
    .C1(\cs_registers_i.dscratch1_q[1] ),
    .C2(_04427_),
    .ZN(_06505_));
 AOI22_X4 _24013_ (.A1(\cs_registers_i.mtval_q[1] ),
    .A2(_04634_),
    .B1(_04424_),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .ZN(_06506_));
 NAND4_X4 _24014_ (.A1(_06501_),
    .A2(_06502_),
    .A3(_06505_),
    .A4(_06506_),
    .ZN(_06507_));
 OAI22_X1 _24015_ (.A1(_05427_),
    .A2(_06492_),
    .B1(_06507_),
    .B2(_10973_),
    .ZN(_06508_));
 OR2_X1 _24016_ (.A1(_05256_),
    .A2(_06449_),
    .ZN(_06509_));
 NOR2_X1 _24017_ (.A1(_16248_),
    .A2(_05451_),
    .ZN(_06510_));
 OAI21_X1 _24018_ (.A(_05454_),
    .B1(_05462_),
    .B2(_16249_),
    .ZN(_06511_));
 AOI221_X2 _24019_ (.A(_06510_),
    .B1(_06511_),
    .B2(_05460_),
    .C1(_05462_),
    .C2(_16251_),
    .ZN(_06512_));
 NOR2_X1 _24020_ (.A1(_16491_),
    .A2(_05478_),
    .ZN(_06513_));
 AND2_X1 _24021_ (.A1(_05163_),
    .A2(_06436_),
    .ZN(_06514_));
 NOR4_X2 _24022_ (.A1(_06492_),
    .A2(_06512_),
    .A3(_06513_),
    .A4(_06514_),
    .ZN(_06515_));
 AOI21_X2 _24023_ (.A(_06508_),
    .B1(_06509_),
    .B2(_06515_),
    .ZN(_06516_));
 AOI221_X1 _24024_ (.A(_05365_),
    .B1(_05369_),
    .B2(\load_store_unit_i.rdata_q[17] ),
    .C1(_05371_),
    .C2(\load_store_unit_i.rdata_q[9] ),
    .ZN(_06517_));
 AOI22_X1 _24025_ (.A1(net37),
    .A2(_05369_),
    .B1(_05373_),
    .B2(_05808_),
    .ZN(_06518_));
 AOI21_X1 _24026_ (.A(_06517_),
    .B1(_06518_),
    .B2(_05376_),
    .ZN(_06519_));
 AOI22_X1 _24027_ (.A1(_05379_),
    .A2(net46),
    .B1(_05381_),
    .B2(\load_store_unit_i.rdata_q[25] ),
    .ZN(_06520_));
 NOR2_X1 _24028_ (.A1(_05378_),
    .A2(_06520_),
    .ZN(_06521_));
 OAI21_X1 _24029_ (.A(_05361_),
    .B1(_06519_),
    .B2(_06521_),
    .ZN(_06522_));
 AOI22_X1 _24030_ (.A1(net40),
    .A2(_05389_),
    .B1(_06519_),
    .B2(_05387_),
    .ZN(_06523_));
 NAND2_X1 _24031_ (.A1(_06522_),
    .A2(_06523_),
    .ZN(_06524_));
 MUX2_X2 _24032_ (.A(_06516_),
    .B(_06524_),
    .S(_05401_),
    .Z(_06525_));
 BUF_X2 _24033_ (.A(_06525_),
    .Z(_06526_));
 MUX2_X1 _24034_ (.A(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .B(_06526_),
    .S(_06487_),
    .Z(_01312_));
 BUF_X2 _24035_ (.A(_05940_),
    .Z(_06527_));
 MUX2_X1 _24036_ (.A(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .B(_06527_),
    .S(_05412_),
    .Z(_01313_));
 NAND3_X1 _24037_ (.A1(_05902_),
    .A2(_05378_),
    .A3(net51),
    .ZN(_06528_));
 AOI221_X2 _24038_ (.A(_05376_),
    .B1(_05369_),
    .B2(\load_store_unit_i.rdata_q[18] ),
    .C1(_05373_),
    .C2(\load_store_unit_i.rdata_q[10] ),
    .ZN(_06529_));
 AND2_X1 _24039_ (.A1(_05388_),
    .A2(net38),
    .ZN(_06530_));
 AOI221_X2 _24040_ (.A(_05499_),
    .B1(_05371_),
    .B2(_05821_),
    .C1(_06530_),
    .C2(_05503_),
    .ZN(_06531_));
 AOI22_X2 _24041_ (.A1(_05379_),
    .A2(net47),
    .B1(_05381_),
    .B2(\load_store_unit_i.rdata_q[26] ),
    .ZN(_06532_));
 OAI221_X2 _24042_ (.A(_06528_),
    .B1(_06529_),
    .B2(_06531_),
    .C1(_05423_),
    .C2(_06532_),
    .ZN(_06533_));
 NAND2_X1 _24043_ (.A1(_15967_),
    .A2(_05428_),
    .ZN(_06534_));
 OAI21_X2 _24044_ (.A(_06534_),
    .B1(_05428_),
    .B2(_00558_),
    .ZN(_06535_));
 OAI221_X1 _24045_ (.A(_12276_),
    .B1(_03737_),
    .B2(_06535_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .C2(_10912_),
    .ZN(_06536_));
 AND2_X1 _24046_ (.A1(_10973_),
    .A2(_06536_),
    .ZN(_06537_));
 NOR2_X1 _24047_ (.A1(_16255_),
    .A2(_05207_),
    .ZN(_06538_));
 OAI21_X1 _24048_ (.A(_05160_),
    .B1(_05209_),
    .B2(_16256_),
    .ZN(_06539_));
 AOI221_X2 _24049_ (.A(_06538_),
    .B1(_06539_),
    .B2(_05204_),
    .C1(_05209_),
    .C2(_16259_),
    .ZN(_06540_));
 INV_X1 _24050_ (.A(_06540_),
    .ZN(_06541_));
 NAND2_X1 _24051_ (.A1(_06537_),
    .A2(_06541_),
    .ZN(_06542_));
 AOI21_X1 _24052_ (.A(_06542_),
    .B1(_05214_),
    .B2(\alu_adder_result_ex[2] ),
    .ZN(_06543_));
 NAND2_X1 _24053_ (.A1(_05925_),
    .A2(_05952_),
    .ZN(_06544_));
 NAND2_X1 _24054_ (.A1(_05727_),
    .A2(_06544_),
    .ZN(_06545_));
 NAND3_X1 _24055_ (.A1(_05552_),
    .A2(_06543_),
    .A3(_06545_),
    .ZN(_06546_));
 AOI221_X2 _24056_ (.A(_06546_),
    .B1(_06419_),
    .B2(_05257_),
    .C1(_05304_),
    .C2(_05950_),
    .ZN(_06547_));
 CLKBUF_X2 _24057_ (.A(\cs_registers_i.mhpmcounter[2][34] ),
    .Z(_06548_));
 AOI22_X1 _24058_ (.A1(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .A2(_04388_),
    .B1(_04391_),
    .B2(_06548_),
    .ZN(_06549_));
 OR2_X1 _24059_ (.A1(_04380_),
    .A2(_06549_),
    .ZN(_06550_));
 OAI22_X2 _24060_ (.A1(_04656_),
    .A2(_04421_),
    .B1(_04456_),
    .B2(_01158_),
    .ZN(_06551_));
 INV_X1 _24061_ (.A(_01164_),
    .ZN(_06552_));
 AOI221_X2 _24062_ (.A(_06551_),
    .B1(_04413_),
    .B2(\cs_registers_i.mtval_q[2] ),
    .C1(_06552_),
    .C2(_04432_),
    .ZN(_06553_));
 AOI22_X1 _24063_ (.A1(\cs_registers_i.csr_mepc_o[2] ),
    .A2(_04423_),
    .B1(_04508_),
    .B2(\cs_registers_i.mscratch_q[2] ),
    .ZN(_06554_));
 AOI22_X1 _24064_ (.A1(net83),
    .A2(_04441_),
    .B1(_04416_),
    .B2(\cs_registers_i.dscratch0_q[2] ),
    .ZN(_06555_));
 AND3_X1 _24065_ (.A1(_06553_),
    .A2(_06554_),
    .A3(_06555_),
    .ZN(_06556_));
 NAND3_X2 _24066_ (.A1(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .A2(_06500_),
    .A3(_04499_),
    .ZN(_06557_));
 AOI222_X2 _24067_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_04407_),
    .B1(_04918_),
    .B2(\cs_registers_i.mcause_q[2] ),
    .C1(_04426_),
    .C2(\cs_registers_i.dscratch1_q[2] ),
    .ZN(_06558_));
 NAND4_X2 _24068_ (.A1(_06550_),
    .A2(_06556_),
    .A3(_06557_),
    .A4(_06558_),
    .ZN(_06559_));
 BUF_X2 _24069_ (.A(\cs_registers_i.mhpmcounter[2][2] ),
    .Z(_06560_));
 INV_X1 _24070_ (.A(_06560_),
    .ZN(_06561_));
 OAI21_X2 _24071_ (.A(_04489_),
    .B1(_04402_),
    .B2(_06561_),
    .ZN(_06562_));
 AOI21_X4 _24072_ (.A(_06559_),
    .B1(_06562_),
    .B2(_04592_),
    .ZN(_06563_));
 AOI221_X2 _24073_ (.A(_06547_),
    .B1(_06537_),
    .B2(_05596_),
    .C1(_05357_),
    .C2(_06563_),
    .ZN(_06564_));
 MUX2_X2 _24074_ (.A(_06533_),
    .B(_06564_),
    .S(_05588_),
    .Z(_06565_));
 BUF_X2 _24075_ (.A(_06565_),
    .Z(_06566_));
 MUX2_X1 _24076_ (.A(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .B(_06566_),
    .S(_06487_),
    .Z(_01314_));
 NAND3_X1 _24077_ (.A1(_05902_),
    .A2(_05378_),
    .A3(net54),
    .ZN(_06567_));
 AOI221_X1 _24078_ (.A(_05365_),
    .B1(_05369_),
    .B2(\load_store_unit_i.rdata_q[19] ),
    .C1(_05373_),
    .C2(\load_store_unit_i.rdata_q[11] ),
    .ZN(_06568_));
 AND2_X1 _24079_ (.A1(_05388_),
    .A2(net39),
    .ZN(_06569_));
 AOI221_X1 _24080_ (.A(_05499_),
    .B1(_05371_),
    .B2(_05900_),
    .C1(_06569_),
    .C2(_05370_),
    .ZN(_06570_));
 AOI22_X1 _24081_ (.A1(_05379_),
    .A2(net48),
    .B1(_05381_),
    .B2(\load_store_unit_i.rdata_q[27] ),
    .ZN(_06571_));
 OAI221_X1 _24082_ (.A(_06567_),
    .B1(_06568_),
    .B2(_06570_),
    .C1(_05423_),
    .C2(_06571_),
    .ZN(_06572_));
 NOR2_X1 _24083_ (.A1(_05588_),
    .A2(_06572_),
    .ZN(_06573_));
 NAND2_X1 _24084_ (.A1(_05304_),
    .A2(_05919_),
    .ZN(_06574_));
 NOR2_X1 _24085_ (.A1(_16263_),
    .A2(_05449_),
    .ZN(_06575_));
 OAI21_X1 _24086_ (.A(_05161_),
    .B1(_05548_),
    .B2(_16264_),
    .ZN(_06576_));
 AOI221_X2 _24087_ (.A(_06575_),
    .B1(_06576_),
    .B2(_05458_),
    .C1(_05549_),
    .C2(_16267_),
    .ZN(_06577_));
 AOI21_X1 _24088_ (.A(_06577_),
    .B1(_05477_),
    .B2(\alu_adder_result_ex[3] ),
    .ZN(_06578_));
 NAND2_X1 _24089_ (.A1(_05552_),
    .A2(_06578_),
    .ZN(_06579_));
 AOI221_X2 _24090_ (.A(_06579_),
    .B1(_05927_),
    .B2(_05727_),
    .C1(_05585_),
    .C2(_06372_),
    .ZN(_06580_));
 AOI21_X1 _24091_ (.A(_05596_),
    .B1(_06574_),
    .B2(_06580_),
    .ZN(_06581_));
 NOR2_X1 _24092_ (.A1(_00559_),
    .A2(_05430_),
    .ZN(_06582_));
 AOI21_X2 _24093_ (.A(_06582_),
    .B1(_05852_),
    .B2(_15982_),
    .ZN(_06583_));
 INV_X1 _24094_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .ZN(_06584_));
 AOI221_X2 _24095_ (.A(_04170_),
    .B1(_03685_),
    .B2(_06583_),
    .C1(_06584_),
    .C2(net307),
    .ZN(_06585_));
 AOI222_X2 _24096_ (.A1(\cs_registers_i.mie_q[17] ),
    .A2(_04448_),
    .B1(_04657_),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .C1(\cs_registers_i.dscratch0_q[3] ),
    .C2(_04417_),
    .ZN(_06586_));
 NAND2_X1 _24097_ (.A1(\cs_registers_i.dscratch1_q[3] ),
    .A2(_04523_),
    .ZN(_06587_));
 AOI22_X2 _24098_ (.A1(net86),
    .A2(_04442_),
    .B1(_04431_),
    .B2(net142),
    .ZN(_06588_));
 AOI21_X2 _24099_ (.A(_04545_),
    .B1(_04918_),
    .B2(\cs_registers_i.mcause_q[3] ),
    .ZN(_06589_));
 NAND4_X2 _24100_ (.A1(_06586_),
    .A2(_06587_),
    .A3(_06588_),
    .A4(_06589_),
    .ZN(_06590_));
 AND2_X1 _24101_ (.A1(\cs_registers_i.mscratch_q[3] ),
    .A2(_04509_),
    .ZN(_06591_));
 AOI22_X1 _24102_ (.A1(\cs_registers_i.mtval_q[3] ),
    .A2(_04634_),
    .B1(_04615_),
    .B2(\cs_registers_i.csr_mepc_o[3] ),
    .ZN(_06592_));
 OAI21_X1 _24103_ (.A(_06592_),
    .B1(_05609_),
    .B2(_01165_),
    .ZN(_06593_));
 NOR3_X2 _24104_ (.A1(_06590_),
    .A2(_06591_),
    .A3(_06593_),
    .ZN(_06594_));
 BUF_X2 _24105_ (.A(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .Z(_06595_));
 BUF_X2 _24106_ (.A(\cs_registers_i.mhpmcounter[2][3] ),
    .Z(_06596_));
 AOI22_X2 _24107_ (.A1(_06595_),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_06596_),
    .ZN(_06597_));
 BUF_X2 _24108_ (.A(\cs_registers_i.mhpmcounter[2][35] ),
    .Z(_06598_));
 AOI22_X2 _24109_ (.A1(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .A2(_04752_),
    .B1(_04753_),
    .B2(_06598_),
    .ZN(_06599_));
 OAI221_X2 _24110_ (.A(_06594_),
    .B1(_06597_),
    .B2(_04629_),
    .C1(_04498_),
    .C2(_06599_),
    .ZN(_06600_));
 NOR3_X2 _24111_ (.A1(_06581_),
    .A2(_06585_),
    .A3(_06600_),
    .ZN(_06601_));
 AOI21_X4 _24112_ (.A(_06573_),
    .B1(_06601_),
    .B2(_05734_),
    .ZN(_06602_));
 BUF_X2 _24113_ (.A(_06602_),
    .Z(_06603_));
 MUX2_X1 _24114_ (.A(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .B(_06603_),
    .S(_06487_),
    .Z(_01315_));
 MUX2_X1 _24115_ (.A(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .B(_05492_),
    .S(_06487_),
    .Z(_01316_));
 MUX2_X1 _24116_ (.A(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .B(_05590_),
    .S(_06487_),
    .Z(_01317_));
 NAND2_X4 _24117_ (.A1(_05976_),
    .A2(_05494_),
    .ZN(_06604_));
 CLKBUF_X3 _24118_ (.A(_06604_),
    .Z(_06605_));
 NAND2_X1 _24119_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .A2(_06605_),
    .ZN(_06606_));
 OAI21_X1 _24120_ (.A(_06606_),
    .B1(_06605_),
    .B2(_05663_),
    .ZN(_01318_));
 BUF_X2 _24121_ (.A(_05735_),
    .Z(_06607_));
 MUX2_X1 _24122_ (.A(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .B(_06607_),
    .S(_06487_),
    .Z(_01319_));
 BUF_X4 _24123_ (.A(_06486_),
    .Z(_06608_));
 MUX2_X1 _24124_ (.A(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .B(_05779_),
    .S(_06608_),
    .Z(_01320_));
 MUX2_X1 _24125_ (.A(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .B(_05816_),
    .S(_06608_),
    .Z(_01321_));
 NOR2_X1 _24126_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .A2(_06487_),
    .ZN(_06609_));
 AOI21_X1 _24127_ (.A(_06609_),
    .B1(_06487_),
    .B2(_05869_),
    .ZN(_01322_));
 MUX2_X1 _24128_ (.A(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .B(_05909_),
    .S(_06608_),
    .Z(_01323_));
 MUX2_X1 _24129_ (.A(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .B(_05975_),
    .S(_05412_),
    .Z(_01324_));
 MUX2_X1 _24130_ (.A(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .B(_06527_),
    .S(_06608_),
    .Z(_01325_));
 MUX2_X1 _24131_ (.A(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .B(_05975_),
    .S(_06608_),
    .Z(_01326_));
 MUX2_X1 _24132_ (.A(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .B(_06027_),
    .S(_06608_),
    .Z(_01327_));
 MUX2_X1 _24133_ (.A(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .B(_06055_),
    .S(_06608_),
    .Z(_01328_));
 BUF_X2 _24134_ (.A(_06087_),
    .Z(_06610_));
 MUX2_X1 _24135_ (.A(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .B(_06610_),
    .S(_06608_),
    .Z(_01329_));
 NAND2_X1 _24136_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .A2(_06604_),
    .ZN(_06611_));
 OAI21_X1 _24137_ (.A(_06611_),
    .B1(_06605_),
    .B2(_06109_),
    .ZN(_01330_));
 BUF_X4 _24138_ (.A(_06131_),
    .Z(_06612_));
 MUX2_X1 _24139_ (.A(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .B(_06612_),
    .S(_06608_),
    .Z(_01331_));
 BUF_X2 _24140_ (.A(_06155_),
    .Z(_06613_));
 MUX2_X1 _24141_ (.A(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .B(_06613_),
    .S(_06608_),
    .Z(_01332_));
 BUF_X2 _24142_ (.A(_06177_),
    .Z(_06614_));
 MUX2_X1 _24143_ (.A(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .B(_06614_),
    .S(_06486_),
    .Z(_01333_));
 NAND2_X1 _24144_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .A2(_06604_),
    .ZN(_06615_));
 OAI21_X1 _24145_ (.A(_06615_),
    .B1(_06605_),
    .B2(_06203_),
    .ZN(_01334_));
 MUX2_X1 _24146_ (.A(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .B(_06027_),
    .S(_05412_),
    .Z(_01335_));
 NAND2_X1 _24147_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .A2(_06604_),
    .ZN(_06616_));
 OAI21_X1 _24148_ (.A(_06616_),
    .B1(_06605_),
    .B2(_06231_),
    .ZN(_01336_));
 MUX2_X1 _24149_ (.A(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .B(_06256_),
    .S(_06486_),
    .Z(_01337_));
 NAND2_X1 _24150_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .A2(_06604_),
    .ZN(_06617_));
 OAI21_X1 _24151_ (.A(_06617_),
    .B1(_06605_),
    .B2(_06284_),
    .ZN(_01338_));
 NAND2_X1 _24152_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .A2(_06604_),
    .ZN(_06618_));
 OAI21_X2 _24153_ (.A(_06618_),
    .B1(_06605_),
    .B2(_06310_),
    .ZN(_01339_));
 MUX2_X1 _24154_ (.A(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .B(_06329_),
    .S(_06486_),
    .Z(_01340_));
 NAND2_X1 _24155_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .A2(_06604_),
    .ZN(_06619_));
 OAI21_X1 _24156_ (.A(_06619_),
    .B1(_06605_),
    .B2(_06361_),
    .ZN(_01341_));
 NAND2_X1 _24157_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .A2(_06604_),
    .ZN(_06620_));
 OAI21_X1 _24158_ (.A(_06620_),
    .B1(_06605_),
    .B2(_06392_),
    .ZN(_01342_));
 MUX2_X1 _24159_ (.A(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .B(net458),
    .S(_06486_),
    .Z(_01343_));
 NAND2_X1 _24160_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .A2(_06604_),
    .ZN(_06621_));
 OAI21_X4 _24161_ (.A(_06621_),
    .B1(net457),
    .B2(_06605_),
    .ZN(_01344_));
 NAND2_X1 _24162_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(_06604_),
    .ZN(_06622_));
 CLKBUF_X3 _24163_ (.A(_06482_),
    .Z(_06623_));
 NAND2_X1 _24164_ (.A1(_06623_),
    .A2(_06487_),
    .ZN(_06624_));
 OAI21_X4 _24165_ (.A(_06622_),
    .B1(net314),
    .B2(_06624_),
    .ZN(_01345_));
 MUX2_X1 _24166_ (.A(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .B(_06055_),
    .S(_05412_),
    .Z(_01346_));
 NOR3_X4 _24167_ (.A1(_10863_),
    .A2(_11306_),
    .A3(_05409_),
    .ZN(_06625_));
 AND2_X1 _24168_ (.A1(_05494_),
    .A2(_06625_),
    .ZN(_06626_));
 BUF_X4 _24169_ (.A(_06626_),
    .Z(_06627_));
 BUF_X4 _24170_ (.A(_06627_),
    .Z(_06628_));
 MUX2_X1 _24171_ (.A(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .B(_05403_),
    .S(_06628_),
    .Z(_01347_));
 MUX2_X1 _24172_ (.A(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .B(_06526_),
    .S(_06628_),
    .Z(_01348_));
 MUX2_X1 _24173_ (.A(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .B(_06566_),
    .S(_06628_),
    .Z(_01349_));
 MUX2_X1 _24174_ (.A(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .B(_06603_),
    .S(_06628_),
    .Z(_01350_));
 MUX2_X1 _24175_ (.A(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .B(_05492_),
    .S(_06628_),
    .Z(_01351_));
 MUX2_X1 _24176_ (.A(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .B(_05590_),
    .S(_06628_),
    .Z(_01352_));
 BUF_X8 _24177_ (.A(_06625_),
    .Z(_06629_));
 NAND2_X4 _24178_ (.A1(_05494_),
    .A2(_06629_),
    .ZN(_06630_));
 CLKBUF_X3 _24179_ (.A(_06630_),
    .Z(_06631_));
 NAND2_X1 _24180_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .A2(_06631_),
    .ZN(_06632_));
 OAI21_X1 _24181_ (.A(_06632_),
    .B1(_06631_),
    .B2(_05663_),
    .ZN(_01353_));
 MUX2_X1 _24182_ (.A(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .B(_06607_),
    .S(_06628_),
    .Z(_01354_));
 BUF_X4 _24183_ (.A(_06627_),
    .Z(_06633_));
 MUX2_X1 _24184_ (.A(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .B(_05779_),
    .S(_06633_),
    .Z(_01355_));
 MUX2_X1 _24185_ (.A(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .B(_05816_),
    .S(_06633_),
    .Z(_01356_));
 MUX2_X1 _24186_ (.A(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .B(_06610_),
    .S(_05412_),
    .Z(_01357_));
 NOR2_X1 _24187_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .A2(_06628_),
    .ZN(_06634_));
 AOI21_X1 _24188_ (.A(_06634_),
    .B1(_06628_),
    .B2(_05869_),
    .ZN(_01358_));
 MUX2_X1 _24189_ (.A(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .B(_05909_),
    .S(_06633_),
    .Z(_01359_));
 MUX2_X1 _24190_ (.A(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .B(_06527_),
    .S(_06633_),
    .Z(_01360_));
 MUX2_X1 _24191_ (.A(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .B(_05975_),
    .S(_06633_),
    .Z(_01361_));
 MUX2_X1 _24192_ (.A(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .B(_06027_),
    .S(_06633_),
    .Z(_01362_));
 MUX2_X1 _24193_ (.A(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .B(_06055_),
    .S(_06633_),
    .Z(_01363_));
 MUX2_X1 _24194_ (.A(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .B(_06610_),
    .S(_06633_),
    .Z(_01364_));
 NAND2_X1 _24195_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .A2(_06630_),
    .ZN(_06635_));
 OAI21_X1 _24196_ (.A(_06635_),
    .B1(_06631_),
    .B2(_06109_),
    .ZN(_01365_));
 MUX2_X1 _24197_ (.A(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .B(_06612_),
    .S(_06633_),
    .Z(_01366_));
 MUX2_X1 _24198_ (.A(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .B(_06613_),
    .S(_06633_),
    .Z(_01367_));
 NAND2_X1 _24199_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .A2(_05978_),
    .ZN(_06636_));
 OAI21_X1 _24200_ (.A(_06636_),
    .B1(_06109_),
    .B2(_05980_),
    .ZN(_01368_));
 MUX2_X1 _24201_ (.A(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .B(_06614_),
    .S(_06627_),
    .Z(_01369_));
 NAND2_X1 _24202_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .A2(_06630_),
    .ZN(_06637_));
 OAI21_X1 _24203_ (.A(_06637_),
    .B1(_06631_),
    .B2(_06203_),
    .ZN(_01370_));
 NAND2_X1 _24204_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .A2(_06630_),
    .ZN(_06638_));
 OAI21_X1 _24205_ (.A(_06638_),
    .B1(_06631_),
    .B2(_06231_),
    .ZN(_01371_));
 MUX2_X1 _24206_ (.A(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .B(_06256_),
    .S(_06627_),
    .Z(_01372_));
 NAND2_X1 _24207_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .A2(_06630_),
    .ZN(_06639_));
 OAI21_X1 _24208_ (.A(_06639_),
    .B1(_06631_),
    .B2(_06284_),
    .ZN(_01373_));
 NAND2_X1 _24209_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .A2(_06630_),
    .ZN(_06640_));
 OAI21_X2 _24210_ (.A(_06640_),
    .B1(_06631_),
    .B2(_06310_),
    .ZN(_01374_));
 MUX2_X1 _24211_ (.A(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .B(_06329_),
    .S(_06627_),
    .Z(_01375_));
 NAND2_X1 _24212_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .A2(_06630_),
    .ZN(_06641_));
 OAI21_X1 _24213_ (.A(_06641_),
    .B1(_06631_),
    .B2(_06361_),
    .ZN(_01376_));
 NAND2_X1 _24214_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .A2(_06630_),
    .ZN(_06642_));
 OAI21_X1 _24215_ (.A(_06642_),
    .B1(_06631_),
    .B2(_06392_),
    .ZN(_01377_));
 MUX2_X1 _24216_ (.A(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .B(_06423_),
    .S(_06627_),
    .Z(_01378_));
 MUX2_X1 _24217_ (.A(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .B(_06612_),
    .S(_05412_),
    .Z(_01379_));
 NAND2_X1 _24218_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .A2(_06630_),
    .ZN(_06643_));
 OAI21_X4 _24219_ (.A(_06643_),
    .B1(net457),
    .B2(_06631_),
    .ZN(_01380_));
 NAND2_X1 _24220_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A2(_06630_),
    .ZN(_06644_));
 NAND2_X1 _24221_ (.A1(_06623_),
    .A2(_06628_),
    .ZN(_06645_));
 OAI21_X4 _24222_ (.A(_06644_),
    .B1(net314),
    .B2(_06645_),
    .ZN(_01381_));
 BUF_X2 _24223_ (.A(_05402_),
    .Z(_06646_));
 NOR3_X4 _24224_ (.A1(_10863_),
    .A2(_11307_),
    .A3(_05409_),
    .ZN(_06647_));
 NAND2_X4 _24225_ (.A1(_05494_),
    .A2(_06647_),
    .ZN(_06648_));
 BUF_X4 _24226_ (.A(_06648_),
    .Z(_06649_));
 MUX2_X1 _24227_ (.A(_06646_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S(_06649_),
    .Z(_01382_));
 BUF_X2 _24228_ (.A(_06525_),
    .Z(_06650_));
 MUX2_X1 _24229_ (.A(_06650_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S(_06649_),
    .Z(_01383_));
 BUF_X2 _24230_ (.A(_06565_),
    .Z(_06651_));
 MUX2_X1 _24231_ (.A(_06651_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S(_06649_),
    .Z(_01384_));
 BUF_X2 _24232_ (.A(_06602_),
    .Z(_06652_));
 MUX2_X1 _24233_ (.A(_06652_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(_06649_),
    .Z(_01385_));
 BUF_X2 _24234_ (.A(_05491_),
    .Z(_06653_));
 MUX2_X1 _24235_ (.A(_06653_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S(_06649_),
    .Z(_01386_));
 BUF_X2 _24236_ (.A(_05589_),
    .Z(_06654_));
 MUX2_X1 _24237_ (.A(_06654_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S(_06649_),
    .Z(_01387_));
 CLKBUF_X3 _24238_ (.A(_06648_),
    .Z(_06655_));
 NAND2_X1 _24239_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .A2(_06655_),
    .ZN(_06656_));
 OAI21_X1 _24240_ (.A(_06656_),
    .B1(_06655_),
    .B2(_05663_),
    .ZN(_01388_));
 NOR3_X4 _24241_ (.A1(_10863_),
    .A2(_11307_),
    .A3(_05409_),
    .ZN(_06657_));
 NAND2_X4 _24242_ (.A1(_05494_),
    .A2(_06657_),
    .ZN(_06658_));
 MUX2_X1 _24243_ (.A(_05736_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S(_06658_),
    .Z(_01389_));
 MUX2_X1 _24244_ (.A(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .B(_06613_),
    .S(_05412_),
    .Z(_01390_));
 BUF_X4 _24245_ (.A(_05411_),
    .Z(_06659_));
 MUX2_X1 _24246_ (.A(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .B(_06526_),
    .S(_06659_),
    .Z(_01391_));
 BUF_X2 _24247_ (.A(_05778_),
    .Z(_06660_));
 MUX2_X1 _24248_ (.A(_06660_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S(_06649_),
    .Z(_01392_));
 BUF_X2 _24249_ (.A(_05815_),
    .Z(_06661_));
 MUX2_X1 _24250_ (.A(_06661_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S(_06649_),
    .Z(_01393_));
 BUF_X4 _24251_ (.A(_06658_),
    .Z(_06662_));
 NAND2_X1 _24252_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .A2(_06662_),
    .ZN(_06663_));
 CLKBUF_X3 _24253_ (.A(_05868_),
    .Z(_06664_));
 OAI21_X1 _24254_ (.A(_06663_),
    .B1(_06662_),
    .B2(_06664_),
    .ZN(_01394_));
 BUF_X2 _24255_ (.A(_05908_),
    .Z(_06665_));
 MUX2_X1 _24256_ (.A(_06665_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S(_06649_),
    .Z(_01395_));
 MUX2_X1 _24257_ (.A(_05941_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S(_06658_),
    .Z(_01396_));
 BUF_X2 _24258_ (.A(_05974_),
    .Z(_06666_));
 MUX2_X1 _24259_ (.A(_06666_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S(_06648_),
    .Z(_01397_));
 BUF_X2 _24260_ (.A(_06026_),
    .Z(_06667_));
 MUX2_X1 _24261_ (.A(_06667_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S(_06648_),
    .Z(_01398_));
 BUF_X2 _24262_ (.A(_06054_),
    .Z(_06668_));
 MUX2_X1 _24263_ (.A(_06668_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S(_06648_),
    .Z(_01399_));
 MUX2_X1 _24264_ (.A(_06088_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S(_06658_),
    .Z(_01400_));
 NAND2_X1 _24265_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .A2(_06655_),
    .ZN(_06669_));
 OAI21_X1 _24266_ (.A(_06669_),
    .B1(_06662_),
    .B2(_06109_),
    .ZN(_01401_));
 MUX2_X1 _24267_ (.A(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .B(_06614_),
    .S(_06659_),
    .Z(_01402_));
 MUX2_X1 _24268_ (.A(_06132_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S(_06658_),
    .Z(_01403_));
 MUX2_X1 _24269_ (.A(_06156_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S(_06658_),
    .Z(_01404_));
 MUX2_X1 _24270_ (.A(_06178_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S(_06658_),
    .Z(_01405_));
 NAND2_X1 _24271_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .A2(_06655_),
    .ZN(_06670_));
 OAI21_X1 _24272_ (.A(_06670_),
    .B1(_06662_),
    .B2(_06203_),
    .ZN(_01406_));
 NAND2_X1 _24273_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .A2(_06655_),
    .ZN(_06671_));
 OAI21_X1 _24274_ (.A(_06671_),
    .B1(_06662_),
    .B2(_06231_),
    .ZN(_01407_));
 BUF_X4 _24275_ (.A(net461),
    .Z(_06672_));
 MUX2_X1 _24276_ (.A(_06672_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S(_06648_),
    .Z(_01408_));
 NAND2_X1 _24277_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .A2(_06655_),
    .ZN(_06673_));
 OAI21_X1 _24278_ (.A(_06673_),
    .B1(_06662_),
    .B2(_06284_),
    .ZN(_01409_));
 NAND2_X1 _24279_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .A2(_06655_),
    .ZN(_06674_));
 OAI21_X2 _24280_ (.A(_06674_),
    .B1(_06662_),
    .B2(_06310_),
    .ZN(_01410_));
 BUF_X4 _24281_ (.A(_06328_),
    .Z(_06675_));
 MUX2_X1 _24282_ (.A(_06675_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S(_06648_),
    .Z(_01411_));
 NAND2_X1 _24283_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .A2(_06655_),
    .ZN(_06676_));
 OAI21_X1 _24284_ (.A(_06676_),
    .B1(_06662_),
    .B2(_06361_),
    .ZN(_01412_));
 NAND2_X1 _24285_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .A2(_05978_),
    .ZN(_06677_));
 OAI21_X1 _24286_ (.A(_06677_),
    .B1(_06203_),
    .B2(_05980_),
    .ZN(_01413_));
 NAND2_X1 _24287_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .A2(_06655_),
    .ZN(_06678_));
 OAI21_X1 _24288_ (.A(_06678_),
    .B1(_06662_),
    .B2(_06392_),
    .ZN(_01414_));
 BUF_X4 _24289_ (.A(_06422_),
    .Z(_06679_));
 MUX2_X1 _24290_ (.A(_06679_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S(_06648_),
    .Z(_01415_));
 NAND2_X1 _24291_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .A2(_06655_),
    .ZN(_06680_));
 OAI21_X4 _24292_ (.A(_06680_),
    .B1(net457),
    .B2(_06662_),
    .ZN(_01416_));
 NAND2_X1 _24293_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .A2(_06649_),
    .ZN(_06681_));
 BUF_X4 _24294_ (.A(_06647_),
    .Z(_06682_));
 NAND3_X1 _24295_ (.A1(_05494_),
    .A2(_06483_),
    .A3(_06682_),
    .ZN(_06683_));
 OAI21_X4 _24296_ (.A(_06681_),
    .B1(net314),
    .B2(_06683_),
    .ZN(_01417_));
 NAND2_X1 _24297_ (.A1(_11308_),
    .A2(_11330_),
    .ZN(_06684_));
 NOR2_X1 _24298_ (.A1(_11310_),
    .A2(_06684_),
    .ZN(_06685_));
 BUF_X8 _24299_ (.A(_06685_),
    .Z(_06686_));
 NAND2_X4 _24300_ (.A1(_05591_),
    .A2(_06686_),
    .ZN(_06687_));
 BUF_X4 _24301_ (.A(_06687_),
    .Z(_06688_));
 MUX2_X1 _24302_ (.A(_06646_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .S(_06688_),
    .Z(_01418_));
 MUX2_X1 _24303_ (.A(_06650_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .S(_06688_),
    .Z(_01419_));
 MUX2_X1 _24304_ (.A(_06651_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .S(_06688_),
    .Z(_01420_));
 MUX2_X1 _24305_ (.A(_06652_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .S(_06688_),
    .Z(_01421_));
 MUX2_X1 _24306_ (.A(_06653_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .S(_06688_),
    .Z(_01422_));
 MUX2_X1 _24307_ (.A(_06654_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .S(_06688_),
    .Z(_01423_));
 NAND2_X1 _24308_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A2(_05978_),
    .ZN(_06689_));
 OAI21_X1 _24309_ (.A(_06689_),
    .B1(_06231_),
    .B2(_05980_),
    .ZN(_01424_));
 CLKBUF_X3 _24310_ (.A(_06687_),
    .Z(_06690_));
 NAND2_X1 _24311_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .A2(_06690_),
    .ZN(_06691_));
 OAI21_X1 _24312_ (.A(_06691_),
    .B1(_06690_),
    .B2(_05663_),
    .ZN(_01425_));
 NAND2_X4 _24313_ (.A1(_05737_),
    .A2(_06686_),
    .ZN(_06692_));
 MUX2_X1 _24314_ (.A(_05736_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .S(_06692_),
    .Z(_01426_));
 MUX2_X1 _24315_ (.A(_06660_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .S(_06688_),
    .Z(_01427_));
 MUX2_X1 _24316_ (.A(_06661_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .S(_06688_),
    .Z(_01428_));
 CLKBUF_X3 _24317_ (.A(_06692_),
    .Z(_06693_));
 NAND2_X1 _24318_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .A2(_06693_),
    .ZN(_06694_));
 OAI21_X1 _24319_ (.A(_06694_),
    .B1(_06693_),
    .B2(_06664_),
    .ZN(_01429_));
 MUX2_X1 _24320_ (.A(_06665_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .S(_06688_),
    .Z(_01430_));
 MUX2_X1 _24321_ (.A(_05941_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .S(_06692_),
    .Z(_01431_));
 MUX2_X1 _24322_ (.A(_06666_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .S(_06687_),
    .Z(_01432_));
 MUX2_X1 _24323_ (.A(_06667_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .S(_06687_),
    .Z(_01433_));
 MUX2_X1 _24324_ (.A(_06668_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .S(_06687_),
    .Z(_01434_));
 MUX2_X1 _24325_ (.A(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .B(_06256_),
    .S(_06659_),
    .Z(_01435_));
 MUX2_X1 _24326_ (.A(_06088_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .S(_06692_),
    .Z(_01436_));
 NAND2_X1 _24327_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .A2(_06690_),
    .ZN(_06695_));
 OAI21_X1 _24328_ (.A(_06695_),
    .B1(_06693_),
    .B2(_06109_),
    .ZN(_01437_));
 MUX2_X1 _24329_ (.A(_06132_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .S(_06692_),
    .Z(_01438_));
 MUX2_X1 _24330_ (.A(_06156_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .S(_06692_),
    .Z(_01439_));
 MUX2_X1 _24331_ (.A(_06178_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .S(_06692_),
    .Z(_01440_));
 NAND2_X1 _24332_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .A2(_06690_),
    .ZN(_06696_));
 OAI21_X1 _24333_ (.A(_06696_),
    .B1(_06693_),
    .B2(_06203_),
    .ZN(_01441_));
 NAND2_X1 _24334_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .A2(_06690_),
    .ZN(_06697_));
 OAI21_X1 _24335_ (.A(_06697_),
    .B1(_06693_),
    .B2(_06231_),
    .ZN(_01442_));
 MUX2_X1 _24336_ (.A(_06672_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .S(_06687_),
    .Z(_01443_));
 NAND2_X1 _24337_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .A2(_06690_),
    .ZN(_06698_));
 OAI21_X1 _24338_ (.A(_06698_),
    .B1(_06693_),
    .B2(_06284_),
    .ZN(_01444_));
 NAND2_X1 _24339_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .A2(_06690_),
    .ZN(_06699_));
 OAI21_X2 _24340_ (.A(_06699_),
    .B1(_06693_),
    .B2(_06310_),
    .ZN(_01445_));
 NAND2_X1 _24341_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .A2(_05978_),
    .ZN(_06700_));
 OAI21_X1 _24342_ (.A(_06700_),
    .B1(_06284_),
    .B2(_05980_),
    .ZN(_01446_));
 MUX2_X1 _24343_ (.A(net485),
    .B(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .S(_06687_),
    .Z(_01447_));
 NAND2_X1 _24344_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .A2(_06690_),
    .ZN(_06701_));
 OAI21_X1 _24345_ (.A(_06701_),
    .B1(_06693_),
    .B2(_06361_),
    .ZN(_01448_));
 NAND2_X1 _24346_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .A2(_06690_),
    .ZN(_06702_));
 OAI21_X1 _24347_ (.A(_06702_),
    .B1(_06693_),
    .B2(_06392_),
    .ZN(_01449_));
 MUX2_X1 _24348_ (.A(net450),
    .B(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .S(_06687_),
    .Z(_01450_));
 NAND2_X1 _24349_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .A2(_06690_),
    .ZN(_06703_));
 OAI21_X4 _24350_ (.A(_06703_),
    .B1(_06457_),
    .B2(_06693_),
    .ZN(_01451_));
 NAND2_X1 _24351_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A2(_06688_),
    .ZN(_06704_));
 NAND3_X1 _24352_ (.A1(_05591_),
    .A2(_06483_),
    .A3(_06686_),
    .ZN(_06705_));
 OAI21_X4 _24353_ (.A(_06704_),
    .B1(net314),
    .B2(_06705_),
    .ZN(_01452_));
 AND2_X1 _24354_ (.A1(_05410_),
    .A2(_06686_),
    .ZN(_06706_));
 CLKBUF_X3 _24355_ (.A(_06706_),
    .Z(_06707_));
 BUF_X4 _24356_ (.A(_06707_),
    .Z(_06708_));
 MUX2_X1 _24357_ (.A(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .B(_05403_),
    .S(_06708_),
    .Z(_01453_));
 MUX2_X1 _24358_ (.A(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .B(_06526_),
    .S(_06708_),
    .Z(_01454_));
 MUX2_X1 _24359_ (.A(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .B(_06566_),
    .S(_06708_),
    .Z(_01455_));
 MUX2_X1 _24360_ (.A(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .B(_06603_),
    .S(_06708_),
    .Z(_01456_));
 NAND2_X1 _24361_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .A2(_05978_),
    .ZN(_06709_));
 OAI21_X4 _24362_ (.A(_06709_),
    .B1(net488),
    .B2(_05980_),
    .ZN(_01457_));
 MUX2_X1 _24363_ (.A(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .B(_05492_),
    .S(_06708_),
    .Z(_01458_));
 MUX2_X1 _24364_ (.A(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .B(_05590_),
    .S(_06708_),
    .Z(_01459_));
 NAND2_X4 _24365_ (.A1(_05976_),
    .A2(_06686_),
    .ZN(_06710_));
 CLKBUF_X3 _24366_ (.A(_06710_),
    .Z(_06711_));
 NAND2_X1 _24367_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .A2(_06711_),
    .ZN(_06712_));
 OAI21_X1 _24368_ (.A(_06712_),
    .B1(_06711_),
    .B2(_05663_),
    .ZN(_01460_));
 MUX2_X1 _24369_ (.A(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .B(_06607_),
    .S(_06708_),
    .Z(_01461_));
 BUF_X4 _24370_ (.A(_06707_),
    .Z(_06713_));
 MUX2_X1 _24371_ (.A(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .B(_05779_),
    .S(_06713_),
    .Z(_01462_));
 MUX2_X1 _24372_ (.A(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .B(_05816_),
    .S(_06713_),
    .Z(_01463_));
 NOR2_X1 _24373_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .A2(_06708_),
    .ZN(_06714_));
 AOI21_X1 _24374_ (.A(_06714_),
    .B1(_06708_),
    .B2(_05869_),
    .ZN(_01464_));
 MUX2_X1 _24375_ (.A(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .B(_05909_),
    .S(_06713_),
    .Z(_01465_));
 MUX2_X1 _24376_ (.A(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .B(_06527_),
    .S(_06713_),
    .Z(_01466_));
 MUX2_X1 _24377_ (.A(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .B(_05975_),
    .S(_06713_),
    .Z(_01467_));
 MUX2_X1 _24378_ (.A(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .B(net484),
    .S(_06659_),
    .Z(_01468_));
 MUX2_X1 _24379_ (.A(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .B(_06027_),
    .S(_06713_),
    .Z(_01469_));
 MUX2_X1 _24380_ (.A(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .B(_06055_),
    .S(_06713_),
    .Z(_01470_));
 MUX2_X1 _24381_ (.A(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .B(_06610_),
    .S(_06713_),
    .Z(_01471_));
 NAND2_X1 _24382_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .A2(_06710_),
    .ZN(_06715_));
 OAI21_X1 _24383_ (.A(_06715_),
    .B1(_06711_),
    .B2(_06109_),
    .ZN(_01472_));
 MUX2_X1 _24384_ (.A(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .B(_06612_),
    .S(_06713_),
    .Z(_01473_));
 MUX2_X1 _24385_ (.A(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .B(_06613_),
    .S(_06713_),
    .Z(_01474_));
 MUX2_X1 _24386_ (.A(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .B(_06614_),
    .S(_06707_),
    .Z(_01475_));
 NAND2_X1 _24387_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .A2(_06710_),
    .ZN(_06716_));
 OAI21_X1 _24388_ (.A(_06716_),
    .B1(_06711_),
    .B2(_06203_),
    .ZN(_01476_));
 NAND2_X1 _24389_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .A2(_06710_),
    .ZN(_06717_));
 OAI21_X1 _24390_ (.A(_06717_),
    .B1(_06711_),
    .B2(_06231_),
    .ZN(_01477_));
 MUX2_X1 _24391_ (.A(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .B(_06256_),
    .S(_06707_),
    .Z(_01478_));
 NAND2_X1 _24392_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .A2(_05978_),
    .ZN(_06718_));
 OAI21_X1 _24393_ (.A(_06718_),
    .B1(_06361_),
    .B2(_05980_),
    .ZN(_01479_));
 NAND2_X1 _24394_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .A2(_06710_),
    .ZN(_06719_));
 OAI21_X1 _24395_ (.A(_06719_),
    .B1(_06711_),
    .B2(_06284_),
    .ZN(_01480_));
 NAND2_X1 _24396_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .A2(_06710_),
    .ZN(_06720_));
 OAI21_X2 _24397_ (.A(_06720_),
    .B1(_06711_),
    .B2(net488),
    .ZN(_01481_));
 MUX2_X1 _24398_ (.A(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .B(net484),
    .S(_06707_),
    .Z(_01482_));
 NAND2_X1 _24399_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .A2(_06710_),
    .ZN(_06721_));
 OAI21_X1 _24400_ (.A(_06721_),
    .B1(_06711_),
    .B2(_06361_),
    .ZN(_01483_));
 NAND2_X1 _24401_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .A2(_06710_),
    .ZN(_06722_));
 OAI21_X1 _24402_ (.A(_06722_),
    .B1(_06711_),
    .B2(_06392_),
    .ZN(_01484_));
 MUX2_X1 _24403_ (.A(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .B(net458),
    .S(_06707_),
    .Z(_01485_));
 NAND2_X1 _24404_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .A2(_06710_),
    .ZN(_06723_));
 OAI21_X4 _24405_ (.A(_06723_),
    .B1(_06457_),
    .B2(_06711_),
    .ZN(_01486_));
 NAND2_X1 _24406_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .A2(_06710_),
    .ZN(_06724_));
 NAND2_X1 _24407_ (.A1(_06623_),
    .A2(_06708_),
    .ZN(_06725_));
 OAI21_X4 _24408_ (.A(_06724_),
    .B1(_06477_),
    .B2(_06725_),
    .ZN(_01487_));
 AND2_X1 _24409_ (.A1(_06629_),
    .A2(_06686_),
    .ZN(_06726_));
 BUF_X4 _24410_ (.A(_06726_),
    .Z(_06727_));
 BUF_X4 _24411_ (.A(_06727_),
    .Z(_06728_));
 MUX2_X1 _24412_ (.A(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .B(_05403_),
    .S(_06728_),
    .Z(_01488_));
 MUX2_X1 _24413_ (.A(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .B(_06526_),
    .S(_06728_),
    .Z(_01489_));
 NAND2_X1 _24414_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .A2(_05978_),
    .ZN(_06729_));
 OAI21_X1 _24415_ (.A(_06729_),
    .B1(_06392_),
    .B2(_05980_),
    .ZN(_01490_));
 MUX2_X1 _24416_ (.A(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .B(_06566_),
    .S(_06728_),
    .Z(_01491_));
 MUX2_X1 _24417_ (.A(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .B(_06603_),
    .S(_06728_),
    .Z(_01492_));
 MUX2_X1 _24418_ (.A(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .B(_05492_),
    .S(_06728_),
    .Z(_01493_));
 MUX2_X1 _24419_ (.A(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .B(_05590_),
    .S(_06728_),
    .Z(_01494_));
 NAND2_X4 _24420_ (.A1(_06629_),
    .A2(_06686_),
    .ZN(_06730_));
 CLKBUF_X3 _24421_ (.A(_06730_),
    .Z(_06731_));
 NAND2_X1 _24422_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .A2(_06731_),
    .ZN(_06732_));
 OAI21_X1 _24423_ (.A(_06732_),
    .B1(_06731_),
    .B2(_05663_),
    .ZN(_01495_));
 MUX2_X1 _24424_ (.A(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .B(_06607_),
    .S(_06728_),
    .Z(_01496_));
 BUF_X4 _24425_ (.A(_06727_),
    .Z(_06733_));
 MUX2_X1 _24426_ (.A(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .B(_05779_),
    .S(_06733_),
    .Z(_01497_));
 MUX2_X1 _24427_ (.A(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .B(_05816_),
    .S(_06733_),
    .Z(_01498_));
 NOR2_X1 _24428_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .A2(_06728_),
    .ZN(_06734_));
 AOI21_X1 _24429_ (.A(_06734_),
    .B1(_06728_),
    .B2(_05869_),
    .ZN(_01499_));
 MUX2_X1 _24430_ (.A(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .B(_05909_),
    .S(_06733_),
    .Z(_01500_));
 MUX2_X1 _24431_ (.A(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .B(net458),
    .S(_06659_),
    .Z(_01501_));
 MUX2_X1 _24432_ (.A(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .B(_06566_),
    .S(_06659_),
    .Z(_01502_));
 MUX2_X1 _24433_ (.A(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .B(_06527_),
    .S(_06733_),
    .Z(_01503_));
 MUX2_X1 _24434_ (.A(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .B(_05975_),
    .S(_06733_),
    .Z(_01504_));
 MUX2_X1 _24435_ (.A(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .B(_06027_),
    .S(_06733_),
    .Z(_01505_));
 MUX2_X1 _24436_ (.A(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .B(_06055_),
    .S(_06733_),
    .Z(_01506_));
 MUX2_X1 _24437_ (.A(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .B(_06610_),
    .S(_06733_),
    .Z(_01507_));
 NAND2_X1 _24438_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .A2(_06730_),
    .ZN(_06735_));
 OAI21_X1 _24439_ (.A(_06735_),
    .B1(_06731_),
    .B2(_06109_),
    .ZN(_01508_));
 MUX2_X1 _24440_ (.A(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .B(_06612_),
    .S(_06733_),
    .Z(_01509_));
 MUX2_X1 _24441_ (.A(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .B(_06613_),
    .S(_06733_),
    .Z(_01510_));
 MUX2_X1 _24442_ (.A(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .B(_06614_),
    .S(_06727_),
    .Z(_01511_));
 NAND2_X1 _24443_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .A2(_06730_),
    .ZN(_06736_));
 OAI21_X1 _24444_ (.A(_06736_),
    .B1(_06731_),
    .B2(_06203_),
    .ZN(_01512_));
 NAND2_X1 _24445_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .A2(_05978_),
    .ZN(_06737_));
 OAI21_X4 _24446_ (.A(_06737_),
    .B1(net457),
    .B2(_05980_),
    .ZN(_01513_));
 NAND2_X1 _24447_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .A2(_06730_),
    .ZN(_06738_));
 OAI21_X1 _24448_ (.A(_06738_),
    .B1(_06731_),
    .B2(_06231_),
    .ZN(_01514_));
 MUX2_X1 _24449_ (.A(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .B(_06256_),
    .S(_06727_),
    .Z(_01515_));
 NAND2_X1 _24450_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .A2(_06730_),
    .ZN(_06739_));
 OAI21_X1 _24451_ (.A(_06739_),
    .B1(_06731_),
    .B2(_06284_),
    .ZN(_01516_));
 NAND2_X1 _24452_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .A2(_06730_),
    .ZN(_06740_));
 OAI21_X2 _24453_ (.A(_06740_),
    .B1(_06731_),
    .B2(net488),
    .ZN(_01517_));
 MUX2_X1 _24454_ (.A(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .B(net484),
    .S(_06727_),
    .Z(_01518_));
 NAND2_X1 _24455_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .A2(_06730_),
    .ZN(_06741_));
 OAI21_X1 _24456_ (.A(_06741_),
    .B1(_06731_),
    .B2(_06361_),
    .ZN(_01519_));
 NAND2_X1 _24457_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .A2(_06730_),
    .ZN(_06742_));
 OAI21_X1 _24458_ (.A(_06742_),
    .B1(_06731_),
    .B2(_06392_),
    .ZN(_01520_));
 MUX2_X1 _24459_ (.A(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .B(_06423_),
    .S(_06727_),
    .Z(_01521_));
 NAND2_X1 _24460_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .A2(_06730_),
    .ZN(_06743_));
 OAI21_X2 _24461_ (.A(_06743_),
    .B1(_06731_),
    .B2(_06457_),
    .ZN(_01522_));
 NAND2_X1 _24462_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .A2(_06730_),
    .ZN(_06744_));
 NAND2_X1 _24463_ (.A1(_06623_),
    .A2(_06728_),
    .ZN(_06745_));
 OAI21_X4 _24464_ (.A(_06744_),
    .B1(_06745_),
    .B2(_06477_),
    .ZN(_01523_));
 NAND2_X1 _24465_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .A2(_05978_),
    .ZN(_06746_));
 CLKBUF_X3 _24466_ (.A(_06482_),
    .Z(_06747_));
 NAND2_X1 _24467_ (.A1(_05412_),
    .A2(_06747_),
    .ZN(_06748_));
 OAI21_X4 _24468_ (.A(_06746_),
    .B1(_06477_),
    .B2(_06748_),
    .ZN(_01524_));
 NAND2_X4 _24469_ (.A1(_06682_),
    .A2(_06686_),
    .ZN(_06749_));
 BUF_X4 _24470_ (.A(_06749_),
    .Z(_06750_));
 MUX2_X1 _24471_ (.A(_06646_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .S(_06750_),
    .Z(_01525_));
 MUX2_X1 _24472_ (.A(_06650_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S(_06750_),
    .Z(_01526_));
 MUX2_X1 _24473_ (.A(_06651_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S(_06750_),
    .Z(_01527_));
 MUX2_X1 _24474_ (.A(_06652_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .S(_06750_),
    .Z(_01528_));
 MUX2_X1 _24475_ (.A(_06653_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S(_06750_),
    .Z(_01529_));
 MUX2_X1 _24476_ (.A(_06654_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .S(_06750_),
    .Z(_01530_));
 CLKBUF_X3 _24477_ (.A(_06749_),
    .Z(_06751_));
 NAND2_X1 _24478_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .A2(_06751_),
    .ZN(_06752_));
 OAI21_X1 _24479_ (.A(_06752_),
    .B1(_06751_),
    .B2(_05663_),
    .ZN(_01531_));
 NAND2_X4 _24480_ (.A1(_06657_),
    .A2(_06686_),
    .ZN(_06753_));
 MUX2_X1 _24481_ (.A(_05736_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S(_06753_),
    .Z(_01532_));
 MUX2_X1 _24482_ (.A(_06660_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S(_06750_),
    .Z(_01533_));
 MUX2_X1 _24483_ (.A(_06661_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .S(_06750_),
    .Z(_01534_));
 AND2_X1 _24484_ (.A1(_11311_),
    .A2(_06625_),
    .ZN(_06754_));
 CLKBUF_X3 _24485_ (.A(_06754_),
    .Z(_06755_));
 BUF_X4 _24486_ (.A(_06755_),
    .Z(_06756_));
 MUX2_X1 _24487_ (.A(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .B(_05403_),
    .S(_06756_),
    .Z(_01535_));
 CLKBUF_X3 _24488_ (.A(_06753_),
    .Z(_06757_));
 NAND2_X1 _24489_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .A2(_06757_),
    .ZN(_06758_));
 OAI21_X1 _24490_ (.A(_06758_),
    .B1(_06757_),
    .B2(_06664_),
    .ZN(_01536_));
 MUX2_X1 _24491_ (.A(_06665_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S(_06750_),
    .Z(_01537_));
 MUX2_X1 _24492_ (.A(_05941_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S(_06753_),
    .Z(_01538_));
 MUX2_X1 _24493_ (.A(_06666_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S(_06749_),
    .Z(_01539_));
 MUX2_X1 _24494_ (.A(_06667_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S(_06749_),
    .Z(_01540_));
 MUX2_X1 _24495_ (.A(_06668_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S(_06749_),
    .Z(_01541_));
 MUX2_X1 _24496_ (.A(_06088_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S(_06753_),
    .Z(_01542_));
 NAND2_X1 _24497_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .A2(_06751_),
    .ZN(_06759_));
 OAI21_X1 _24498_ (.A(_06759_),
    .B1(_06757_),
    .B2(_06109_),
    .ZN(_01543_));
 MUX2_X1 _24499_ (.A(_06132_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S(_06753_),
    .Z(_01544_));
 MUX2_X1 _24500_ (.A(_06156_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S(_06753_),
    .Z(_01545_));
 MUX2_X1 _24501_ (.A(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .B(_06526_),
    .S(_06756_),
    .Z(_01546_));
 MUX2_X1 _24502_ (.A(_06178_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S(_06753_),
    .Z(_01547_));
 NAND2_X1 _24503_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .A2(_06751_),
    .ZN(_06760_));
 OAI21_X1 _24504_ (.A(_06760_),
    .B1(_06757_),
    .B2(_06203_),
    .ZN(_01548_));
 NAND2_X1 _24505_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .A2(_06751_),
    .ZN(_06761_));
 OAI21_X1 _24506_ (.A(_06761_),
    .B1(_06757_),
    .B2(_06231_),
    .ZN(_01549_));
 MUX2_X1 _24507_ (.A(_06672_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S(_06749_),
    .Z(_01550_));
 NAND2_X1 _24508_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .A2(_06751_),
    .ZN(_06762_));
 OAI21_X1 _24509_ (.A(_06762_),
    .B1(_06757_),
    .B2(_06284_),
    .ZN(_01551_));
 NAND2_X1 _24510_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .A2(_06751_),
    .ZN(_06763_));
 OAI21_X1 _24511_ (.A(_06763_),
    .B1(_06757_),
    .B2(_06310_),
    .ZN(_01552_));
 MUX2_X1 _24512_ (.A(_06675_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S(_06749_),
    .Z(_01553_));
 NAND2_X1 _24513_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .A2(_06751_),
    .ZN(_06764_));
 OAI21_X1 _24514_ (.A(_06764_),
    .B1(_06757_),
    .B2(_06361_),
    .ZN(_01554_));
 NAND2_X1 _24515_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .A2(_06751_),
    .ZN(_06765_));
 OAI21_X1 _24516_ (.A(_06765_),
    .B1(_06757_),
    .B2(_06392_),
    .ZN(_01555_));
 MUX2_X1 _24517_ (.A(net450),
    .B(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S(_06749_),
    .Z(_01556_));
 MUX2_X1 _24518_ (.A(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .B(_06566_),
    .S(_06756_),
    .Z(_01557_));
 NAND2_X1 _24519_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .A2(_06751_),
    .ZN(_06766_));
 OAI21_X4 _24520_ (.A(_06766_),
    .B1(_06457_),
    .B2(_06757_),
    .ZN(_01558_));
 NAND2_X1 _24521_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .A2(_06750_),
    .ZN(_06767_));
 NAND3_X1 _24522_ (.A1(_06747_),
    .A2(_06682_),
    .A3(_06686_),
    .ZN(_06768_));
 OAI21_X4 _24523_ (.A(_06767_),
    .B1(_06477_),
    .B2(_06768_),
    .ZN(_01559_));
 BUF_X2 _24524_ (.A(_05402_),
    .Z(_06769_));
 NAND2_X2 _24525_ (.A1(_11308_),
    .A2(_11309_),
    .ZN(_06770_));
 NOR2_X1 _24526_ (.A1(_11310_),
    .A2(_06770_),
    .ZN(_06771_));
 BUF_X8 _24527_ (.A(_06771_),
    .Z(_06772_));
 NAND2_X4 _24528_ (.A1(_05591_),
    .A2(_06772_),
    .ZN(_06773_));
 BUF_X4 _24529_ (.A(_06773_),
    .Z(_06774_));
 MUX2_X1 _24530_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .S(_06774_),
    .Z(_01560_));
 BUF_X2 _24531_ (.A(_06525_),
    .Z(_06775_));
 MUX2_X1 _24532_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .S(_06774_),
    .Z(_01561_));
 BUF_X2 _24533_ (.A(_06565_),
    .Z(_06776_));
 MUX2_X1 _24534_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .S(_06774_),
    .Z(_01562_));
 BUF_X2 _24535_ (.A(_06602_),
    .Z(_06777_));
 MUX2_X1 _24536_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .S(_06774_),
    .Z(_01563_));
 BUF_X2 _24537_ (.A(_05491_),
    .Z(_06778_));
 MUX2_X1 _24538_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .S(_06774_),
    .Z(_01564_));
 BUF_X2 _24539_ (.A(_05589_),
    .Z(_06779_));
 MUX2_X1 _24540_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .S(_06774_),
    .Z(_01565_));
 CLKBUF_X3 _24541_ (.A(_06773_),
    .Z(_06780_));
 NAND2_X1 _24542_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .A2(_06780_),
    .ZN(_06781_));
 OAI21_X1 _24543_ (.A(_06781_),
    .B1(_06780_),
    .B2(_05663_),
    .ZN(_01566_));
 BUF_X2 _24544_ (.A(_05735_),
    .Z(_06782_));
 NAND2_X4 _24545_ (.A1(_05737_),
    .A2(_06772_),
    .ZN(_06783_));
 MUX2_X1 _24546_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .S(_06783_),
    .Z(_01567_));
 MUX2_X1 _24547_ (.A(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .B(_06603_),
    .S(_06756_),
    .Z(_01568_));
 BUF_X2 _24548_ (.A(_05778_),
    .Z(_06784_));
 MUX2_X1 _24549_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .S(_06774_),
    .Z(_01569_));
 BUF_X2 _24550_ (.A(_05815_),
    .Z(_06785_));
 MUX2_X1 _24551_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .S(_06774_),
    .Z(_01570_));
 BUF_X4 _24552_ (.A(_06783_),
    .Z(_06786_));
 NAND2_X1 _24553_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .A2(_06786_),
    .ZN(_06787_));
 OAI21_X1 _24554_ (.A(_06787_),
    .B1(_06786_),
    .B2(_06664_),
    .ZN(_01571_));
 BUF_X2 _24555_ (.A(_05908_),
    .Z(_06788_));
 MUX2_X1 _24556_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .S(_06774_),
    .Z(_01572_));
 BUF_X2 _24557_ (.A(_05940_),
    .Z(_06789_));
 MUX2_X1 _24558_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .S(_06783_),
    .Z(_01573_));
 BUF_X2 _24559_ (.A(_05974_),
    .Z(_06790_));
 MUX2_X1 _24560_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .S(_06773_),
    .Z(_01574_));
 BUF_X2 _24561_ (.A(_06026_),
    .Z(_06791_));
 MUX2_X1 _24562_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .S(_06773_),
    .Z(_01575_));
 BUF_X2 _24563_ (.A(_06054_),
    .Z(_06792_));
 MUX2_X1 _24564_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .S(_06773_),
    .Z(_01576_));
 BUF_X2 _24565_ (.A(_06087_),
    .Z(_06793_));
 MUX2_X1 _24566_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .S(_06783_),
    .Z(_01577_));
 NAND2_X1 _24567_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .A2(_06780_),
    .ZN(_06794_));
 OAI21_X1 _24568_ (.A(_06794_),
    .B1(_06786_),
    .B2(_06109_),
    .ZN(_01578_));
 MUX2_X1 _24569_ (.A(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .B(_05492_),
    .S(_06756_),
    .Z(_01579_));
 BUF_X4 _24570_ (.A(_06131_),
    .Z(_06795_));
 MUX2_X1 _24571_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .S(_06783_),
    .Z(_01580_));
 BUF_X2 _24572_ (.A(_06155_),
    .Z(_06796_));
 MUX2_X1 _24573_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .S(_06783_),
    .Z(_01581_));
 BUF_X2 _24574_ (.A(_06177_),
    .Z(_06797_));
 MUX2_X1 _24575_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .S(_06783_),
    .Z(_01582_));
 NAND2_X1 _24576_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .A2(_06780_),
    .ZN(_06798_));
 OAI21_X1 _24577_ (.A(_06798_),
    .B1(_06786_),
    .B2(_06203_),
    .ZN(_01583_));
 NAND2_X1 _24578_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .A2(_06780_),
    .ZN(_06799_));
 OAI21_X1 _24579_ (.A(_06799_),
    .B1(_06786_),
    .B2(_06231_),
    .ZN(_01584_));
 BUF_X8 _24580_ (.A(net461),
    .Z(_06800_));
 MUX2_X1 _24581_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .S(_06773_),
    .Z(_01585_));
 NAND2_X1 _24582_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .A2(_06780_),
    .ZN(_06801_));
 OAI21_X1 _24583_ (.A(_06801_),
    .B1(_06786_),
    .B2(_06284_),
    .ZN(_01586_));
 NAND2_X1 _24584_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .A2(_06780_),
    .ZN(_06802_));
 OAI21_X2 _24585_ (.A(_06802_),
    .B1(_06786_),
    .B2(net488),
    .ZN(_01587_));
 BUF_X4 _24586_ (.A(_06328_),
    .Z(_06803_));
 MUX2_X1 _24587_ (.A(_06803_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .S(_06773_),
    .Z(_01588_));
 NAND2_X1 _24588_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .A2(_06780_),
    .ZN(_06804_));
 OAI21_X1 _24589_ (.A(_06804_),
    .B1(_06786_),
    .B2(_06361_),
    .ZN(_01589_));
 MUX2_X1 _24590_ (.A(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .B(_05590_),
    .S(_06756_),
    .Z(_01590_));
 NAND2_X1 _24591_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .A2(_06780_),
    .ZN(_06805_));
 OAI21_X1 _24592_ (.A(_06805_),
    .B1(_06786_),
    .B2(_06392_),
    .ZN(_01591_));
 BUF_X4 _24593_ (.A(_06422_),
    .Z(_06806_));
 MUX2_X1 _24594_ (.A(net599),
    .B(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .S(_06773_),
    .Z(_01592_));
 NAND2_X1 _24595_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .A2(_06780_),
    .ZN(_06807_));
 OAI21_X4 _24596_ (.A(_06807_),
    .B1(_06457_),
    .B2(_06786_),
    .ZN(_01593_));
 NAND2_X1 _24597_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A2(_06774_),
    .ZN(_06808_));
 NAND3_X1 _24598_ (.A1(_05591_),
    .A2(_06483_),
    .A3(_06772_),
    .ZN(_06809_));
 OAI21_X4 _24599_ (.A(_06808_),
    .B1(_06477_),
    .B2(_06809_),
    .ZN(_01594_));
 AND2_X1 _24600_ (.A1(_05410_),
    .A2(_06772_),
    .ZN(_06810_));
 BUF_X4 _24601_ (.A(_06810_),
    .Z(_06811_));
 BUF_X4 _24602_ (.A(_06811_),
    .Z(_06812_));
 MUX2_X1 _24603_ (.A(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .B(_05403_),
    .S(_06812_),
    .Z(_01595_));
 MUX2_X1 _24604_ (.A(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .B(_06526_),
    .S(_06812_),
    .Z(_01596_));
 MUX2_X1 _24605_ (.A(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .B(_06566_),
    .S(_06812_),
    .Z(_01597_));
 MUX2_X1 _24606_ (.A(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .B(_06603_),
    .S(_06812_),
    .Z(_01598_));
 MUX2_X1 _24607_ (.A(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .B(_05492_),
    .S(_06812_),
    .Z(_01599_));
 MUX2_X1 _24608_ (.A(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .B(_05590_),
    .S(_06812_),
    .Z(_01600_));
 NAND2_X4 _24609_ (.A1(_11311_),
    .A2(_06629_),
    .ZN(_06813_));
 CLKBUF_X3 _24610_ (.A(_06813_),
    .Z(_06814_));
 NAND2_X1 _24611_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .A2(_06814_),
    .ZN(_06815_));
 CLKBUF_X3 _24612_ (.A(_05662_),
    .Z(_06816_));
 OAI21_X1 _24613_ (.A(_06815_),
    .B1(_06814_),
    .B2(_06816_),
    .ZN(_01601_));
 NAND2_X4 _24614_ (.A1(_05976_),
    .A2(_06772_),
    .ZN(_06817_));
 CLKBUF_X3 _24615_ (.A(_06817_),
    .Z(_06818_));
 NAND2_X1 _24616_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .A2(_06818_),
    .ZN(_06819_));
 OAI21_X1 _24617_ (.A(_06819_),
    .B1(_06818_),
    .B2(_06816_),
    .ZN(_01602_));
 MUX2_X1 _24618_ (.A(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .B(_06607_),
    .S(_06812_),
    .Z(_01603_));
 BUF_X4 _24619_ (.A(_06811_),
    .Z(_06820_));
 MUX2_X1 _24620_ (.A(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .B(_05779_),
    .S(_06820_),
    .Z(_01604_));
 MUX2_X1 _24621_ (.A(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .B(_05816_),
    .S(_06820_),
    .Z(_01605_));
 NOR2_X1 _24622_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .A2(_06812_),
    .ZN(_06821_));
 AOI21_X1 _24623_ (.A(_06821_),
    .B1(_06812_),
    .B2(_05869_),
    .ZN(_01606_));
 MUX2_X1 _24624_ (.A(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .B(_05909_),
    .S(_06820_),
    .Z(_01607_));
 MUX2_X1 _24625_ (.A(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .B(_06527_),
    .S(_06820_),
    .Z(_01608_));
 MUX2_X1 _24626_ (.A(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .B(_05975_),
    .S(_06820_),
    .Z(_01609_));
 MUX2_X1 _24627_ (.A(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .B(_06027_),
    .S(_06820_),
    .Z(_01610_));
 MUX2_X1 _24628_ (.A(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .B(_06055_),
    .S(_06820_),
    .Z(_01611_));
 MUX2_X1 _24629_ (.A(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .B(_06607_),
    .S(_06756_),
    .Z(_01612_));
 MUX2_X1 _24630_ (.A(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .B(_06603_),
    .S(_06659_),
    .Z(_01613_));
 MUX2_X1 _24631_ (.A(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .B(_06610_),
    .S(_06820_),
    .Z(_01614_));
 NAND2_X1 _24632_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .A2(_06817_),
    .ZN(_06822_));
 CLKBUF_X3 _24633_ (.A(_06108_),
    .Z(_06823_));
 OAI21_X1 _24634_ (.A(_06822_),
    .B1(_06818_),
    .B2(_06823_),
    .ZN(_01615_));
 MUX2_X1 _24635_ (.A(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .B(_06612_),
    .S(_06820_),
    .Z(_01616_));
 MUX2_X1 _24636_ (.A(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .B(_06613_),
    .S(_06820_),
    .Z(_01617_));
 MUX2_X1 _24637_ (.A(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .B(_06614_),
    .S(_06811_),
    .Z(_01618_));
 NAND2_X1 _24638_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .A2(_06817_),
    .ZN(_06824_));
 CLKBUF_X3 _24639_ (.A(_06202_),
    .Z(_06825_));
 OAI21_X1 _24640_ (.A(_06824_),
    .B1(_06818_),
    .B2(_06825_),
    .ZN(_01619_));
 NAND2_X1 _24641_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .A2(_06817_),
    .ZN(_06826_));
 BUF_X4 _24642_ (.A(_06230_),
    .Z(_06827_));
 OAI21_X1 _24643_ (.A(_06826_),
    .B1(_06818_),
    .B2(_06827_),
    .ZN(_01620_));
 MUX2_X1 _24644_ (.A(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .B(_06256_),
    .S(_06811_),
    .Z(_01621_));
 NAND2_X1 _24645_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .A2(_06817_),
    .ZN(_06828_));
 CLKBUF_X3 _24646_ (.A(_06283_),
    .Z(_06829_));
 OAI21_X1 _24647_ (.A(_06828_),
    .B1(_06818_),
    .B2(_06829_),
    .ZN(_01622_));
 NAND2_X1 _24648_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .A2(_06817_),
    .ZN(_06830_));
 BUF_X8 _24649_ (.A(_06309_),
    .Z(_06831_));
 OAI21_X2 _24650_ (.A(_06830_),
    .B1(_06818_),
    .B2(_06831_),
    .ZN(_01623_));
 BUF_X4 _24651_ (.A(_06755_),
    .Z(_06832_));
 MUX2_X1 _24652_ (.A(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .B(_05779_),
    .S(_06832_),
    .Z(_01624_));
 MUX2_X1 _24653_ (.A(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .B(_06329_),
    .S(_06811_),
    .Z(_01625_));
 NAND2_X1 _24654_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .A2(_06817_),
    .ZN(_06833_));
 BUF_X4 _24655_ (.A(_06360_),
    .Z(_06834_));
 OAI21_X1 _24656_ (.A(_06833_),
    .B1(_06818_),
    .B2(_06834_),
    .ZN(_01626_));
 NAND2_X1 _24657_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .A2(_06817_),
    .ZN(_06835_));
 BUF_X4 _24658_ (.A(_06391_),
    .Z(_06836_));
 OAI21_X1 _24659_ (.A(_06835_),
    .B1(_06818_),
    .B2(_06836_),
    .ZN(_01627_));
 MUX2_X1 _24660_ (.A(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .B(net458),
    .S(_06811_),
    .Z(_01628_));
 NAND2_X1 _24661_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .A2(_06817_),
    .ZN(_06837_));
 BUF_X8 _24662_ (.A(_06456_),
    .Z(_06838_));
 OAI21_X4 _24663_ (.A(_06837_),
    .B1(net459),
    .B2(_06818_),
    .ZN(_01629_));
 NAND2_X1 _24664_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .A2(_06817_),
    .ZN(_06839_));
 NAND2_X1 _24665_ (.A1(_06623_),
    .A2(_06812_),
    .ZN(_06840_));
 BUF_X16 _24666_ (.A(net372),
    .Z(_06841_));
 OAI21_X4 _24667_ (.A(_06839_),
    .B1(_06841_),
    .B2(_06840_),
    .ZN(_01630_));
 AND2_X1 _24668_ (.A1(_06625_),
    .A2(_06772_),
    .ZN(_06842_));
 BUF_X4 _24669_ (.A(_06842_),
    .Z(_06843_));
 BUF_X4 _24670_ (.A(_06843_),
    .Z(_06844_));
 MUX2_X1 _24671_ (.A(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .B(_05403_),
    .S(_06844_),
    .Z(_01631_));
 MUX2_X1 _24672_ (.A(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .B(_06526_),
    .S(_06844_),
    .Z(_01632_));
 MUX2_X1 _24673_ (.A(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .B(_06566_),
    .S(_06844_),
    .Z(_01633_));
 MUX2_X1 _24674_ (.A(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .B(_06603_),
    .S(_06844_),
    .Z(_01634_));
 MUX2_X1 _24675_ (.A(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .B(_05816_),
    .S(_06832_),
    .Z(_01635_));
 MUX2_X1 _24676_ (.A(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .B(_05492_),
    .S(_06844_),
    .Z(_01636_));
 MUX2_X1 _24677_ (.A(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .B(_05590_),
    .S(_06844_),
    .Z(_01637_));
 NAND2_X4 _24678_ (.A1(_06629_),
    .A2(_06772_),
    .ZN(_06845_));
 CLKBUF_X3 _24679_ (.A(_06845_),
    .Z(_06846_));
 NAND2_X1 _24680_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .A2(_06846_),
    .ZN(_06847_));
 OAI21_X1 _24681_ (.A(_06847_),
    .B1(_06846_),
    .B2(_06816_),
    .ZN(_01638_));
 MUX2_X1 _24682_ (.A(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .B(_06607_),
    .S(_06844_),
    .Z(_01639_));
 BUF_X4 _24683_ (.A(_06843_),
    .Z(_06848_));
 MUX2_X1 _24684_ (.A(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .B(_05779_),
    .S(_06848_),
    .Z(_01640_));
 MUX2_X1 _24685_ (.A(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .B(_05816_),
    .S(_06848_),
    .Z(_01641_));
 NOR2_X1 _24686_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .A2(_06844_),
    .ZN(_06849_));
 AOI21_X1 _24687_ (.A(_06849_),
    .B1(_06844_),
    .B2(_05869_),
    .ZN(_01642_));
 MUX2_X1 _24688_ (.A(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .B(_05909_),
    .S(_06848_),
    .Z(_01643_));
 MUX2_X1 _24689_ (.A(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .B(_06527_),
    .S(_06848_),
    .Z(_01644_));
 MUX2_X1 _24690_ (.A(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .B(_05975_),
    .S(_06848_),
    .Z(_01645_));
 NOR2_X1 _24691_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .A2(_06756_),
    .ZN(_06850_));
 AOI21_X1 _24692_ (.A(_06850_),
    .B1(_06756_),
    .B2(_05869_),
    .ZN(_01646_));
 MUX2_X1 _24693_ (.A(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .B(_06027_),
    .S(_06848_),
    .Z(_01647_));
 MUX2_X1 _24694_ (.A(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .B(_06055_),
    .S(_06848_),
    .Z(_01648_));
 MUX2_X1 _24695_ (.A(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .B(_06610_),
    .S(_06848_),
    .Z(_01649_));
 NAND2_X1 _24696_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .A2(_06845_),
    .ZN(_06851_));
 OAI21_X1 _24697_ (.A(_06851_),
    .B1(_06846_),
    .B2(_06823_),
    .ZN(_01650_));
 MUX2_X1 _24698_ (.A(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .B(_06612_),
    .S(_06848_),
    .Z(_01651_));
 MUX2_X1 _24699_ (.A(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .B(_06613_),
    .S(_06848_),
    .Z(_01652_));
 MUX2_X1 _24700_ (.A(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .B(_06614_),
    .S(_06843_),
    .Z(_01653_));
 NAND2_X1 _24701_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .A2(_06845_),
    .ZN(_06852_));
 OAI21_X1 _24702_ (.A(_06852_),
    .B1(_06846_),
    .B2(_06825_),
    .ZN(_01654_));
 NAND2_X1 _24703_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .A2(_06845_),
    .ZN(_06853_));
 OAI21_X1 _24704_ (.A(_06853_),
    .B1(_06846_),
    .B2(_06827_),
    .ZN(_01655_));
 MUX2_X1 _24705_ (.A(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .B(_06256_),
    .S(_06843_),
    .Z(_01656_));
 MUX2_X1 _24706_ (.A(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .B(_05909_),
    .S(_06832_),
    .Z(_01657_));
 NAND2_X1 _24707_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .A2(_06845_),
    .ZN(_06854_));
 OAI21_X1 _24708_ (.A(_06854_),
    .B1(_06846_),
    .B2(_06829_),
    .ZN(_01658_));
 NAND2_X1 _24709_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .A2(_06845_),
    .ZN(_06855_));
 OAI21_X2 _24710_ (.A(_06855_),
    .B1(_06846_),
    .B2(_06831_),
    .ZN(_01659_));
 MUX2_X1 _24711_ (.A(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .B(_06329_),
    .S(_06843_),
    .Z(_01660_));
 NAND2_X1 _24712_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .A2(_06845_),
    .ZN(_06856_));
 OAI21_X1 _24713_ (.A(_06856_),
    .B1(_06846_),
    .B2(_06834_),
    .ZN(_01661_));
 NAND2_X1 _24714_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .A2(_06845_),
    .ZN(_06857_));
 OAI21_X1 _24715_ (.A(_06857_),
    .B1(_06846_),
    .B2(_06836_),
    .ZN(_01662_));
 MUX2_X1 _24716_ (.A(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .B(_06423_),
    .S(_06843_),
    .Z(_01663_));
 NAND2_X1 _24717_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .A2(_06845_),
    .ZN(_06858_));
 OAI21_X4 _24718_ (.A(_06858_),
    .B1(net459),
    .B2(_06846_),
    .ZN(_01664_));
 NAND2_X1 _24719_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .A2(_06845_),
    .ZN(_06859_));
 NAND2_X1 _24720_ (.A1(_06623_),
    .A2(_06844_),
    .ZN(_06860_));
 OAI21_X4 _24721_ (.A(_06859_),
    .B1(_06841_),
    .B2(_06860_),
    .ZN(_01665_));
 NAND2_X4 _24722_ (.A1(_06682_),
    .A2(_06772_),
    .ZN(_06861_));
 BUF_X4 _24723_ (.A(_06861_),
    .Z(_06862_));
 MUX2_X1 _24724_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S(_06862_),
    .Z(_01666_));
 MUX2_X1 _24725_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S(_06862_),
    .Z(_01667_));
 MUX2_X1 _24726_ (.A(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .B(_06527_),
    .S(_06832_),
    .Z(_01668_));
 MUX2_X1 _24727_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S(_06862_),
    .Z(_01669_));
 MUX2_X1 _24728_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S(_06862_),
    .Z(_01670_));
 MUX2_X1 _24729_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S(_06862_),
    .Z(_01671_));
 MUX2_X1 _24730_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S(_06862_),
    .Z(_01672_));
 CLKBUF_X3 _24731_ (.A(_06861_),
    .Z(_06863_));
 NAND2_X1 _24732_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .A2(_06863_),
    .ZN(_06864_));
 OAI21_X1 _24733_ (.A(_06864_),
    .B1(_06863_),
    .B2(_06816_),
    .ZN(_01673_));
 NAND2_X4 _24734_ (.A1(_06657_),
    .A2(_06772_),
    .ZN(_06865_));
 MUX2_X1 _24735_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S(_06865_),
    .Z(_01674_));
 MUX2_X1 _24736_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S(_06862_),
    .Z(_01675_));
 MUX2_X1 _24737_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S(_06862_),
    .Z(_01676_));
 BUF_X4 _24738_ (.A(_06865_),
    .Z(_06866_));
 NAND2_X1 _24739_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .A2(_06866_),
    .ZN(_06867_));
 OAI21_X1 _24740_ (.A(_06867_),
    .B1(_06866_),
    .B2(_06664_),
    .ZN(_01677_));
 MUX2_X1 _24741_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S(_06862_),
    .Z(_01678_));
 MUX2_X1 _24742_ (.A(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .B(_05975_),
    .S(_06832_),
    .Z(_01679_));
 MUX2_X1 _24743_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S(_06865_),
    .Z(_01680_));
 MUX2_X1 _24744_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S(_06861_),
    .Z(_01681_));
 MUX2_X1 _24745_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S(_06861_),
    .Z(_01682_));
 MUX2_X1 _24746_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S(_06861_),
    .Z(_01683_));
 MUX2_X1 _24747_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S(_06865_),
    .Z(_01684_));
 NAND2_X1 _24748_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .A2(_06863_),
    .ZN(_06868_));
 OAI21_X1 _24749_ (.A(_06868_),
    .B1(_06866_),
    .B2(_06823_),
    .ZN(_01685_));
 MUX2_X1 _24750_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S(_06865_),
    .Z(_01686_));
 MUX2_X1 _24751_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S(_06865_),
    .Z(_01687_));
 MUX2_X1 _24752_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S(_06865_),
    .Z(_01688_));
 NAND2_X1 _24753_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .A2(_06863_),
    .ZN(_06869_));
 OAI21_X1 _24754_ (.A(_06869_),
    .B1(_06866_),
    .B2(_06825_),
    .ZN(_01689_));
 MUX2_X1 _24755_ (.A(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .B(_06027_),
    .S(_06832_),
    .Z(_01690_));
 NAND2_X1 _24756_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .A2(_06863_),
    .ZN(_06870_));
 OAI21_X1 _24757_ (.A(_06870_),
    .B1(_06866_),
    .B2(_06827_),
    .ZN(_01691_));
 MUX2_X1 _24758_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S(_06861_),
    .Z(_01692_));
 NAND2_X1 _24759_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .A2(_06863_),
    .ZN(_06871_));
 OAI21_X1 _24760_ (.A(_06871_),
    .B1(_06866_),
    .B2(_06829_),
    .ZN(_01693_));
 NAND2_X1 _24761_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .A2(_06863_),
    .ZN(_06872_));
 OAI21_X2 _24762_ (.A(_06872_),
    .B1(_06866_),
    .B2(_06831_),
    .ZN(_01694_));
 MUX2_X1 _24763_ (.A(_06803_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S(_06861_),
    .Z(_01695_));
 NAND2_X1 _24764_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .A2(_06863_),
    .ZN(_06873_));
 OAI21_X1 _24765_ (.A(_06873_),
    .B1(_06866_),
    .B2(_06834_),
    .ZN(_01696_));
 NAND2_X1 _24766_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .A2(_06863_),
    .ZN(_06874_));
 OAI21_X1 _24767_ (.A(_06874_),
    .B1(_06866_),
    .B2(_06836_),
    .ZN(_01697_));
 MUX2_X1 _24768_ (.A(net599),
    .B(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S(_06861_),
    .Z(_01698_));
 NAND2_X1 _24769_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .A2(_06863_),
    .ZN(_06875_));
 OAI21_X4 _24770_ (.A(_06875_),
    .B1(net459),
    .B2(_06866_),
    .ZN(_01699_));
 NAND2_X1 _24771_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .A2(_06862_),
    .ZN(_06876_));
 NAND3_X1 _24772_ (.A1(_06747_),
    .A2(_06682_),
    .A3(_06772_),
    .ZN(_06877_));
 OAI21_X4 _24773_ (.A(_06876_),
    .B1(_06841_),
    .B2(_06877_),
    .ZN(_01700_));
 MUX2_X1 _24774_ (.A(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .B(_06055_),
    .S(_06832_),
    .Z(_01701_));
 BUF_X4 _24775_ (.A(_00039_),
    .Z(_06878_));
 NOR3_X4 _24776_ (.A1(_11308_),
    .A2(_11309_),
    .A3(_06878_),
    .ZN(_06879_));
 NAND2_X4 _24777_ (.A1(_05591_),
    .A2(_06879_),
    .ZN(_06880_));
 BUF_X4 _24778_ (.A(_06880_),
    .Z(_06881_));
 MUX2_X1 _24779_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .S(_06881_),
    .Z(_01702_));
 MUX2_X1 _24780_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .S(_06881_),
    .Z(_01703_));
 MUX2_X1 _24781_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .S(_06881_),
    .Z(_01704_));
 MUX2_X1 _24782_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .S(_06881_),
    .Z(_01705_));
 MUX2_X1 _24783_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .S(_06881_),
    .Z(_01706_));
 MUX2_X1 _24784_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .S(_06881_),
    .Z(_01707_));
 BUF_X4 _24785_ (.A(_06880_),
    .Z(_06882_));
 NAND2_X1 _24786_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .A2(_06882_),
    .ZN(_06883_));
 OAI21_X1 _24787_ (.A(_06883_),
    .B1(_06882_),
    .B2(_06816_),
    .ZN(_01708_));
 NAND2_X4 _24788_ (.A1(_05737_),
    .A2(_06879_),
    .ZN(_06884_));
 MUX2_X1 _24789_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .S(_06884_),
    .Z(_01709_));
 MUX2_X1 _24790_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .S(_06881_),
    .Z(_01710_));
 MUX2_X1 _24791_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .S(_06881_),
    .Z(_01711_));
 MUX2_X1 _24792_ (.A(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .B(_06610_),
    .S(_06832_),
    .Z(_01712_));
 BUF_X4 _24793_ (.A(_06884_),
    .Z(_06885_));
 NAND2_X1 _24794_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .A2(_06885_),
    .ZN(_06886_));
 OAI21_X1 _24795_ (.A(_06886_),
    .B1(_06885_),
    .B2(_06664_),
    .ZN(_01713_));
 MUX2_X1 _24796_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .S(_06881_),
    .Z(_01714_));
 MUX2_X1 _24797_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .S(_06884_),
    .Z(_01715_));
 MUX2_X1 _24798_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .S(_06880_),
    .Z(_01716_));
 MUX2_X1 _24799_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .S(_06880_),
    .Z(_01717_));
 MUX2_X1 _24800_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .S(_06880_),
    .Z(_01718_));
 MUX2_X1 _24801_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .S(_06884_),
    .Z(_01719_));
 NAND2_X1 _24802_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .A2(_06882_),
    .ZN(_06887_));
 OAI21_X1 _24803_ (.A(_06887_),
    .B1(_06885_),
    .B2(_06823_),
    .ZN(_01720_));
 MUX2_X1 _24804_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .S(_06884_),
    .Z(_01721_));
 MUX2_X1 _24805_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .S(_06884_),
    .Z(_01722_));
 NAND2_X1 _24806_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .A2(_06813_),
    .ZN(_06888_));
 OAI21_X1 _24807_ (.A(_06888_),
    .B1(_06814_),
    .B2(_06823_),
    .ZN(_01723_));
 MUX2_X1 _24808_ (.A(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B(_05492_),
    .S(_06659_),
    .Z(_01724_));
 MUX2_X1 _24809_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .S(_06884_),
    .Z(_01725_));
 NAND2_X1 _24810_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .A2(_06882_),
    .ZN(_06889_));
 OAI21_X1 _24811_ (.A(_06889_),
    .B1(_06885_),
    .B2(_06825_),
    .ZN(_01726_));
 NAND2_X1 _24812_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .A2(_06882_),
    .ZN(_06890_));
 OAI21_X1 _24813_ (.A(_06890_),
    .B1(_06885_),
    .B2(_06827_),
    .ZN(_01727_));
 MUX2_X1 _24814_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .S(_06880_),
    .Z(_01728_));
 NAND2_X1 _24815_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .A2(_06882_),
    .ZN(_06891_));
 OAI21_X1 _24816_ (.A(_06891_),
    .B1(_06885_),
    .B2(_06829_),
    .ZN(_01729_));
 NAND2_X1 _24817_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .A2(_06882_),
    .ZN(_06892_));
 OAI21_X4 _24818_ (.A(_06892_),
    .B1(_06831_),
    .B2(_06885_),
    .ZN(_01730_));
 MUX2_X1 _24819_ (.A(net483),
    .B(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .S(_06880_),
    .Z(_01731_));
 NAND2_X1 _24820_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .A2(_06882_),
    .ZN(_06893_));
 OAI21_X1 _24821_ (.A(_06893_),
    .B1(_06885_),
    .B2(_06834_),
    .ZN(_01732_));
 NAND2_X1 _24822_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .A2(_06882_),
    .ZN(_06894_));
 OAI21_X1 _24823_ (.A(_06894_),
    .B1(_06885_),
    .B2(_06836_),
    .ZN(_01733_));
 MUX2_X1 _24824_ (.A(_06806_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .S(_06880_),
    .Z(_01734_));
 MUX2_X1 _24825_ (.A(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .B(_06612_),
    .S(_06832_),
    .Z(_01735_));
 NAND2_X1 _24826_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .A2(_06882_),
    .ZN(_06895_));
 OAI21_X2 _24827_ (.A(_06895_),
    .B1(_06885_),
    .B2(_06838_),
    .ZN(_01736_));
 NAND2_X1 _24828_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A2(_06881_),
    .ZN(_06896_));
 NAND3_X1 _24829_ (.A1(_05591_),
    .A2(_06483_),
    .A3(_06879_),
    .ZN(_06897_));
 OAI21_X4 _24830_ (.A(_06896_),
    .B1(_06841_),
    .B2(_06897_),
    .ZN(_01737_));
 AND2_X2 _24831_ (.A1(_05976_),
    .A2(_06879_),
    .ZN(_06898_));
 BUF_X4 _24832_ (.A(_06898_),
    .Z(_06899_));
 MUX2_X1 _24833_ (.A(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .B(_05403_),
    .S(_06899_),
    .Z(_01738_));
 MUX2_X1 _24834_ (.A(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .B(_06526_),
    .S(_06899_),
    .Z(_01739_));
 MUX2_X1 _24835_ (.A(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .B(_06566_),
    .S(_06899_),
    .Z(_01740_));
 MUX2_X1 _24836_ (.A(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .B(_06603_),
    .S(_06899_),
    .Z(_01741_));
 MUX2_X1 _24837_ (.A(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .B(_05492_),
    .S(_06899_),
    .Z(_01742_));
 MUX2_X1 _24838_ (.A(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .B(_05590_),
    .S(_06899_),
    .Z(_01743_));
 NAND2_X2 _24839_ (.A1(_05976_),
    .A2(_06879_),
    .ZN(_06900_));
 BUF_X4 _24840_ (.A(_06900_),
    .Z(_06901_));
 NAND2_X1 _24841_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .A2(_06901_),
    .ZN(_06902_));
 BUF_X4 _24842_ (.A(_06900_),
    .Z(_06903_));
 OAI21_X1 _24843_ (.A(_06902_),
    .B1(_06903_),
    .B2(_06816_),
    .ZN(_01744_));
 MUX2_X1 _24844_ (.A(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .B(_06607_),
    .S(_06899_),
    .Z(_01745_));
 MUX2_X1 _24845_ (.A(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .B(_06613_),
    .S(_06832_),
    .Z(_01746_));
 MUX2_X1 _24846_ (.A(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .B(_05779_),
    .S(_06899_),
    .Z(_01747_));
 MUX2_X1 _24847_ (.A(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .B(_05816_),
    .S(_06899_),
    .Z(_01748_));
 NAND2_X1 _24848_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .A2(_06901_),
    .ZN(_06904_));
 CLKBUF_X3 _24849_ (.A(_05868_),
    .Z(_06905_));
 OAI21_X1 _24850_ (.A(_06904_),
    .B1(_06903_),
    .B2(_06905_),
    .ZN(_01749_));
 BUF_X4 _24851_ (.A(_06898_),
    .Z(_06906_));
 MUX2_X1 _24852_ (.A(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .B(_05909_),
    .S(_06906_),
    .Z(_01750_));
 MUX2_X1 _24853_ (.A(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .B(_06527_),
    .S(_06906_),
    .Z(_01751_));
 MUX2_X1 _24854_ (.A(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .B(_05975_),
    .S(_06906_),
    .Z(_01752_));
 MUX2_X1 _24855_ (.A(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .B(_06027_),
    .S(_06906_),
    .Z(_01753_));
 MUX2_X1 _24856_ (.A(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .B(_06055_),
    .S(_06906_),
    .Z(_01754_));
 MUX2_X1 _24857_ (.A(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .B(_06610_),
    .S(_06906_),
    .Z(_01755_));
 NAND2_X1 _24858_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .A2(_06901_),
    .ZN(_06907_));
 OAI21_X1 _24859_ (.A(_06907_),
    .B1(_06903_),
    .B2(_06823_),
    .ZN(_01756_));
 MUX2_X1 _24860_ (.A(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .B(_06614_),
    .S(_06755_),
    .Z(_01757_));
 MUX2_X1 _24861_ (.A(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .B(_06612_),
    .S(_06906_),
    .Z(_01758_));
 MUX2_X1 _24862_ (.A(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .B(_06613_),
    .S(_06906_),
    .Z(_01759_));
 MUX2_X1 _24863_ (.A(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .B(_06614_),
    .S(_06906_),
    .Z(_01760_));
 NAND2_X1 _24864_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .A2(_06901_),
    .ZN(_06908_));
 OAI21_X1 _24865_ (.A(_06908_),
    .B1(_06903_),
    .B2(_06825_),
    .ZN(_01761_));
 NAND2_X1 _24866_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .A2(_06901_),
    .ZN(_06909_));
 OAI21_X1 _24867_ (.A(_06909_),
    .B1(_06903_),
    .B2(_06827_),
    .ZN(_01762_));
 MUX2_X1 _24868_ (.A(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .B(_06256_),
    .S(_06906_),
    .Z(_01763_));
 NAND2_X1 _24869_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .A2(_06901_),
    .ZN(_06910_));
 OAI21_X1 _24870_ (.A(_06910_),
    .B1(_06903_),
    .B2(_06829_),
    .ZN(_01764_));
 NAND2_X1 _24871_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .A2(_06901_),
    .ZN(_06911_));
 OAI21_X2 _24872_ (.A(_06911_),
    .B1(_06903_),
    .B2(net487),
    .ZN(_01765_));
 MUX2_X1 _24873_ (.A(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .B(net484),
    .S(_06898_),
    .Z(_01766_));
 NAND2_X1 _24874_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .A2(_06901_),
    .ZN(_06912_));
 OAI21_X1 _24875_ (.A(_06912_),
    .B1(_06903_),
    .B2(_06834_),
    .ZN(_01767_));
 NAND2_X1 _24876_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .A2(_06813_),
    .ZN(_06913_));
 OAI21_X1 _24877_ (.A(_06913_),
    .B1(_06814_),
    .B2(_06825_),
    .ZN(_01768_));
 NAND2_X1 _24878_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .A2(_06901_),
    .ZN(_06914_));
 OAI21_X1 _24879_ (.A(_06914_),
    .B1(_06903_),
    .B2(_06836_),
    .ZN(_01769_));
 MUX2_X1 _24880_ (.A(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .B(_06423_),
    .S(_06898_),
    .Z(_01770_));
 NAND2_X1 _24881_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .A2(_06901_),
    .ZN(_06915_));
 OAI21_X2 _24882_ (.A(_06915_),
    .B1(_06903_),
    .B2(_06838_),
    .ZN(_01771_));
 NAND2_X1 _24883_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .A2(_06900_),
    .ZN(_06916_));
 NAND2_X1 _24884_ (.A1(_06623_),
    .A2(_06899_),
    .ZN(_06917_));
 OAI21_X4 _24885_ (.A(_06916_),
    .B1(net358),
    .B2(_06917_),
    .ZN(_01772_));
 AND2_X1 _24886_ (.A1(_06625_),
    .A2(_06879_),
    .ZN(_06918_));
 BUF_X4 _24887_ (.A(_06918_),
    .Z(_06919_));
 BUF_X4 _24888_ (.A(_06919_),
    .Z(_06920_));
 MUX2_X1 _24889_ (.A(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .B(_05403_),
    .S(_06920_),
    .Z(_01773_));
 MUX2_X1 _24890_ (.A(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .B(_06526_),
    .S(_06920_),
    .Z(_01774_));
 MUX2_X1 _24891_ (.A(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .B(_06566_),
    .S(_06920_),
    .Z(_01775_));
 MUX2_X1 _24892_ (.A(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .B(_06603_),
    .S(_06920_),
    .Z(_01776_));
 MUX2_X1 _24893_ (.A(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .B(_06653_),
    .S(_06920_),
    .Z(_01777_));
 MUX2_X1 _24894_ (.A(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .B(_05590_),
    .S(_06920_),
    .Z(_01778_));
 NAND2_X1 _24895_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .A2(_06813_),
    .ZN(_06921_));
 OAI21_X1 _24896_ (.A(_06921_),
    .B1(_06814_),
    .B2(_06827_),
    .ZN(_01779_));
 NAND2_X4 _24897_ (.A1(_06629_),
    .A2(_06879_),
    .ZN(_06922_));
 BUF_X4 _24898_ (.A(_06922_),
    .Z(_06923_));
 NAND2_X1 _24899_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .A2(_06923_),
    .ZN(_06924_));
 OAI21_X1 _24900_ (.A(_06924_),
    .B1(_06923_),
    .B2(_06816_),
    .ZN(_01780_));
 MUX2_X1 _24901_ (.A(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .B(_06607_),
    .S(_06920_),
    .Z(_01781_));
 BUF_X4 _24902_ (.A(_06919_),
    .Z(_06925_));
 MUX2_X1 _24903_ (.A(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .B(_05779_),
    .S(_06925_),
    .Z(_01782_));
 MUX2_X1 _24904_ (.A(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .B(_05816_),
    .S(_06925_),
    .Z(_01783_));
 NOR2_X1 _24905_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .A2(_06920_),
    .ZN(_06926_));
 AOI21_X1 _24906_ (.A(_06926_),
    .B1(_06920_),
    .B2(_05869_),
    .ZN(_01784_));
 MUX2_X1 _24907_ (.A(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .B(_06665_),
    .S(_06925_),
    .Z(_01785_));
 MUX2_X1 _24908_ (.A(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .B(_06527_),
    .S(_06925_),
    .Z(_01786_));
 MUX2_X1 _24909_ (.A(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .B(_06666_),
    .S(_06925_),
    .Z(_01787_));
 MUX2_X1 _24910_ (.A(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .B(_06667_),
    .S(_06925_),
    .Z(_01788_));
 MUX2_X1 _24911_ (.A(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .B(_06668_),
    .S(_06925_),
    .Z(_01789_));
 MUX2_X1 _24912_ (.A(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .B(_06256_),
    .S(_06755_),
    .Z(_01790_));
 MUX2_X1 _24913_ (.A(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .B(_06610_),
    .S(_06925_),
    .Z(_01791_));
 NAND2_X1 _24914_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .A2(_06922_),
    .ZN(_06927_));
 OAI21_X1 _24915_ (.A(_06927_),
    .B1(_06923_),
    .B2(_06823_),
    .ZN(_01792_));
 MUX2_X1 _24916_ (.A(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .B(_06612_),
    .S(_06925_),
    .Z(_01793_));
 MUX2_X1 _24917_ (.A(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .B(_06613_),
    .S(_06925_),
    .Z(_01794_));
 MUX2_X1 _24918_ (.A(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .B(_06614_),
    .S(_06919_),
    .Z(_01795_));
 NAND2_X1 _24919_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .A2(_06922_),
    .ZN(_06928_));
 OAI21_X1 _24920_ (.A(_06928_),
    .B1(_06923_),
    .B2(_06825_),
    .ZN(_01796_));
 NAND2_X1 _24921_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .A2(_06922_),
    .ZN(_06929_));
 OAI21_X1 _24922_ (.A(_06929_),
    .B1(_06923_),
    .B2(_06827_),
    .ZN(_01797_));
 MUX2_X1 _24923_ (.A(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .B(net460),
    .S(_06919_),
    .Z(_01798_));
 NAND2_X1 _24924_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .A2(_06922_),
    .ZN(_06930_));
 OAI21_X1 _24925_ (.A(_06930_),
    .B1(_06923_),
    .B2(_06829_),
    .ZN(_01799_));
 NAND2_X1 _24926_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .A2(_06922_),
    .ZN(_06931_));
 OAI21_X2 _24927_ (.A(_06931_),
    .B1(_06923_),
    .B2(net487),
    .ZN(_01800_));
 NAND2_X1 _24928_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .A2(_06813_),
    .ZN(_06932_));
 OAI21_X1 _24929_ (.A(_06932_),
    .B1(_06814_),
    .B2(_06829_),
    .ZN(_01801_));
 MUX2_X1 _24930_ (.A(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .B(net484),
    .S(_06919_),
    .Z(_01802_));
 NAND2_X1 _24931_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .A2(_06922_),
    .ZN(_06933_));
 OAI21_X1 _24932_ (.A(_06933_),
    .B1(_06923_),
    .B2(_06834_),
    .ZN(_01803_));
 NAND2_X1 _24933_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .A2(_06922_),
    .ZN(_06934_));
 OAI21_X1 _24934_ (.A(_06934_),
    .B1(_06923_),
    .B2(_06836_),
    .ZN(_01804_));
 MUX2_X1 _24935_ (.A(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .B(_06423_),
    .S(_06919_),
    .Z(_01805_));
 NAND2_X1 _24936_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .A2(_06922_),
    .ZN(_06935_));
 OAI21_X2 _24937_ (.A(_06935_),
    .B1(_06923_),
    .B2(_06838_),
    .ZN(_01806_));
 NAND2_X1 _24938_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .A2(_06922_),
    .ZN(_06936_));
 NAND2_X1 _24939_ (.A1(_06623_),
    .A2(_06920_),
    .ZN(_06937_));
 OAI21_X4 _24940_ (.A(_06936_),
    .B1(net358),
    .B2(_06937_),
    .ZN(_01807_));
 NAND2_X4 _24941_ (.A1(_06647_),
    .A2(_06879_),
    .ZN(_06938_));
 BUF_X4 _24942_ (.A(_06938_),
    .Z(_06939_));
 MUX2_X1 _24943_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S(_06939_),
    .Z(_01808_));
 MUX2_X1 _24944_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .S(_06939_),
    .Z(_01809_));
 MUX2_X1 _24945_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S(_06939_),
    .Z(_01810_));
 MUX2_X1 _24946_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .S(_06939_),
    .Z(_01811_));
 NAND2_X1 _24947_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .A2(_06813_),
    .ZN(_06940_));
 OAI21_X2 _24948_ (.A(_06940_),
    .B1(_06814_),
    .B2(_06831_),
    .ZN(_01812_));
 MUX2_X1 _24949_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S(_06939_),
    .Z(_01813_));
 MUX2_X1 _24950_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S(_06939_),
    .Z(_01814_));
 BUF_X4 _24951_ (.A(_06938_),
    .Z(_06941_));
 NAND2_X1 _24952_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .A2(_06941_),
    .ZN(_06942_));
 OAI21_X1 _24953_ (.A(_06942_),
    .B1(_06941_),
    .B2(_06816_),
    .ZN(_01815_));
 NAND2_X4 _24954_ (.A1(_06657_),
    .A2(_06879_),
    .ZN(_06943_));
 MUX2_X1 _24955_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S(_06943_),
    .Z(_01816_));
 MUX2_X1 _24956_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S(_06939_),
    .Z(_01817_));
 MUX2_X1 _24957_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S(_06939_),
    .Z(_01818_));
 BUF_X4 _24958_ (.A(_06943_),
    .Z(_06944_));
 NAND2_X1 _24959_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .A2(_06944_),
    .ZN(_06945_));
 OAI21_X1 _24960_ (.A(_06945_),
    .B1(_06944_),
    .B2(_06905_),
    .ZN(_01819_));
 MUX2_X1 _24961_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S(_06939_),
    .Z(_01820_));
 MUX2_X1 _24962_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S(_06943_),
    .Z(_01821_));
 MUX2_X1 _24963_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S(_06938_),
    .Z(_01822_));
 MUX2_X1 _24964_ (.A(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .B(_06675_),
    .S(_06755_),
    .Z(_01823_));
 MUX2_X1 _24965_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S(_06938_),
    .Z(_01824_));
 MUX2_X1 _24966_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S(_06938_),
    .Z(_01825_));
 MUX2_X1 _24967_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S(_06943_),
    .Z(_01826_));
 NAND2_X1 _24968_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .A2(_06941_),
    .ZN(_06946_));
 OAI21_X1 _24969_ (.A(_06946_),
    .B1(_06944_),
    .B2(_06823_),
    .ZN(_01827_));
 MUX2_X1 _24970_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S(_06943_),
    .Z(_01828_));
 MUX2_X1 _24971_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S(_06943_),
    .Z(_01829_));
 MUX2_X1 _24972_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S(_06943_),
    .Z(_01830_));
 NAND2_X1 _24973_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .A2(_06941_),
    .ZN(_06947_));
 OAI21_X1 _24974_ (.A(_06947_),
    .B1(_06944_),
    .B2(_06825_),
    .ZN(_01831_));
 NAND2_X1 _24975_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .A2(_06941_),
    .ZN(_06948_));
 OAI21_X1 _24976_ (.A(_06948_),
    .B1(_06944_),
    .B2(_06827_),
    .ZN(_01832_));
 MUX2_X1 _24977_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S(_06938_),
    .Z(_01833_));
 NAND2_X1 _24978_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .A2(_06813_),
    .ZN(_06949_));
 OAI21_X1 _24979_ (.A(_06949_),
    .B1(_06814_),
    .B2(_06834_),
    .ZN(_01834_));
 MUX2_X1 _24980_ (.A(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .B(_06654_),
    .S(_06659_),
    .Z(_01835_));
 NAND2_X1 _24981_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .A2(_06941_),
    .ZN(_06950_));
 OAI21_X1 _24982_ (.A(_06950_),
    .B1(_06944_),
    .B2(_06829_),
    .ZN(_01836_));
 NAND2_X1 _24983_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .A2(_06941_),
    .ZN(_06951_));
 OAI21_X2 _24984_ (.A(_06951_),
    .B1(_06944_),
    .B2(net487),
    .ZN(_01837_));
 MUX2_X1 _24985_ (.A(net483),
    .B(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S(_06938_),
    .Z(_01838_));
 NAND2_X1 _24986_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .A2(_06941_),
    .ZN(_06952_));
 OAI21_X1 _24987_ (.A(_06952_),
    .B1(_06944_),
    .B2(_06834_),
    .ZN(_01839_));
 NAND2_X1 _24988_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .A2(_06941_),
    .ZN(_06953_));
 OAI21_X1 _24989_ (.A(_06953_),
    .B1(_06944_),
    .B2(_06836_),
    .ZN(_01840_));
 MUX2_X1 _24990_ (.A(net599),
    .B(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S(_06938_),
    .Z(_01841_));
 NAND2_X1 _24991_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .A2(_06941_),
    .ZN(_06954_));
 OAI21_X2 _24992_ (.A(_06954_),
    .B1(_06944_),
    .B2(net459),
    .ZN(_01842_));
 NAND2_X1 _24993_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .A2(_06939_),
    .ZN(_06955_));
 NAND3_X1 _24994_ (.A1(_06747_),
    .A2(_06682_),
    .A3(_06879_),
    .ZN(_06956_));
 OAI21_X4 _24995_ (.A(_06955_),
    .B1(net358),
    .B2(_06956_),
    .ZN(_01843_));
 NOR2_X4 _24996_ (.A1(_06878_),
    .A2(_05493_),
    .ZN(_06957_));
 NAND2_X4 _24997_ (.A1(_05495_),
    .A2(_06957_),
    .ZN(_06958_));
 BUF_X4 _24998_ (.A(_06958_),
    .Z(_06959_));
 MUX2_X1 _24999_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .S(_06959_),
    .Z(_01844_));
 MUX2_X1 _25000_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .S(_06959_),
    .Z(_01845_));
 NAND2_X1 _25001_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .A2(_06813_),
    .ZN(_06960_));
 OAI21_X1 _25002_ (.A(_06960_),
    .B1(_06814_),
    .B2(_06836_),
    .ZN(_01846_));
 MUX2_X1 _25003_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .S(_06959_),
    .Z(_01847_));
 MUX2_X1 _25004_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .S(_06959_),
    .Z(_01848_));
 MUX2_X1 _25005_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .S(_06959_),
    .Z(_01849_));
 MUX2_X1 _25006_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .S(_06959_),
    .Z(_01850_));
 BUF_X4 _25007_ (.A(_06958_),
    .Z(_06961_));
 NAND2_X1 _25008_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .A2(_06961_),
    .ZN(_06962_));
 OAI21_X1 _25009_ (.A(_06962_),
    .B1(_06961_),
    .B2(_06816_),
    .ZN(_01851_));
 NAND2_X4 _25010_ (.A1(_05737_),
    .A2(_06957_),
    .ZN(_06963_));
 MUX2_X1 _25011_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .S(_06963_),
    .Z(_01852_));
 MUX2_X1 _25012_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .S(_06959_),
    .Z(_01853_));
 MUX2_X1 _25013_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .S(_06959_),
    .Z(_01854_));
 BUF_X4 _25014_ (.A(_06963_),
    .Z(_06964_));
 NAND2_X1 _25015_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .A2(_06964_),
    .ZN(_06965_));
 OAI21_X1 _25016_ (.A(_06965_),
    .B1(_06964_),
    .B2(_06905_),
    .ZN(_01855_));
 MUX2_X1 _25017_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .S(_06959_),
    .Z(_01856_));
 MUX2_X1 _25018_ (.A(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .B(net450),
    .S(_06755_),
    .Z(_01857_));
 MUX2_X1 _25019_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .S(_06963_),
    .Z(_01858_));
 MUX2_X1 _25020_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .S(_06958_),
    .Z(_01859_));
 MUX2_X1 _25021_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .S(_06958_),
    .Z(_01860_));
 MUX2_X1 _25022_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .S(_06958_),
    .Z(_01861_));
 MUX2_X1 _25023_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .S(_06963_),
    .Z(_01862_));
 NAND2_X1 _25024_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .A2(_06961_),
    .ZN(_06966_));
 OAI21_X1 _25025_ (.A(_06966_),
    .B1(_06964_),
    .B2(_06823_),
    .ZN(_01863_));
 MUX2_X1 _25026_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .S(_06963_),
    .Z(_01864_));
 MUX2_X1 _25027_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .S(_06963_),
    .Z(_01865_));
 MUX2_X1 _25028_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .S(_06963_),
    .Z(_01866_));
 NAND2_X1 _25029_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .A2(_06961_),
    .ZN(_06967_));
 OAI21_X1 _25030_ (.A(_06967_),
    .B1(_06964_),
    .B2(_06825_),
    .ZN(_01867_));
 NAND2_X1 _25031_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .A2(_06813_),
    .ZN(_06968_));
 OAI21_X4 _25032_ (.A(_06968_),
    .B1(net459),
    .B2(_06814_),
    .ZN(_01868_));
 NAND2_X1 _25033_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .A2(_06961_),
    .ZN(_06969_));
 OAI21_X1 _25034_ (.A(_06969_),
    .B1(_06964_),
    .B2(_06827_),
    .ZN(_01869_));
 MUX2_X1 _25035_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .S(_06958_),
    .Z(_01870_));
 NAND2_X1 _25036_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .A2(_06961_),
    .ZN(_06970_));
 OAI21_X1 _25037_ (.A(_06970_),
    .B1(_06964_),
    .B2(_06829_),
    .ZN(_01871_));
 NAND2_X1 _25038_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .A2(_06961_),
    .ZN(_06971_));
 OAI21_X2 _25039_ (.A(_06971_),
    .B1(_06964_),
    .B2(net487),
    .ZN(_01872_));
 MUX2_X1 _25040_ (.A(net483),
    .B(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .S(_06958_),
    .Z(_01873_));
 NAND2_X1 _25041_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .A2(_06961_),
    .ZN(_06972_));
 OAI21_X1 _25042_ (.A(_06972_),
    .B1(_06964_),
    .B2(_06834_),
    .ZN(_01874_));
 NAND2_X1 _25043_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .A2(_06961_),
    .ZN(_06973_));
 OAI21_X1 _25044_ (.A(_06973_),
    .B1(_06964_),
    .B2(_06836_),
    .ZN(_01875_));
 MUX2_X1 _25045_ (.A(_06806_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .S(_06958_),
    .Z(_01876_));
 NAND2_X1 _25046_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .A2(_06961_),
    .ZN(_06974_));
 OAI21_X2 _25047_ (.A(_06974_),
    .B1(_06964_),
    .B2(_06838_),
    .ZN(_01877_));
 NAND2_X1 _25048_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A2(_06959_),
    .ZN(_06975_));
 NAND3_X1 _25049_ (.A1(_05591_),
    .A2(_06483_),
    .A3(_06957_),
    .ZN(_06976_));
 OAI21_X4 _25050_ (.A(_06975_),
    .B1(net358),
    .B2(_06976_),
    .ZN(_01878_));
 NAND2_X1 _25051_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A2(_06813_),
    .ZN(_06977_));
 NAND2_X1 _25052_ (.A1(_06623_),
    .A2(_06756_),
    .ZN(_06978_));
 OAI21_X4 _25053_ (.A(_06977_),
    .B1(net358),
    .B2(_06978_),
    .ZN(_01879_));
 AND2_X2 _25054_ (.A1(_05976_),
    .A2(_06957_),
    .ZN(_06979_));
 BUF_X4 _25055_ (.A(_06979_),
    .Z(_06980_));
 MUX2_X1 _25056_ (.A(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .B(_06646_),
    .S(_06980_),
    .Z(_01880_));
 MUX2_X1 _25057_ (.A(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .B(_06650_),
    .S(_06980_),
    .Z(_01881_));
 MUX2_X1 _25058_ (.A(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .B(_06651_),
    .S(_06980_),
    .Z(_01882_));
 MUX2_X1 _25059_ (.A(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .B(_06652_),
    .S(_06980_),
    .Z(_01883_));
 MUX2_X1 _25060_ (.A(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .B(_06653_),
    .S(_06980_),
    .Z(_01884_));
 MUX2_X1 _25061_ (.A(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .B(_06654_),
    .S(_06980_),
    .Z(_01885_));
 NAND2_X2 _25062_ (.A1(_05976_),
    .A2(_06957_),
    .ZN(_06981_));
 BUF_X4 _25063_ (.A(_06981_),
    .Z(_06982_));
 NAND2_X1 _25064_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .A2(_06982_),
    .ZN(_06983_));
 BUF_X4 _25065_ (.A(_06981_),
    .Z(_06984_));
 OAI21_X1 _25066_ (.A(_06983_),
    .B1(_06984_),
    .B2(_06816_),
    .ZN(_01886_));
 MUX2_X1 _25067_ (.A(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .B(_06607_),
    .S(_06980_),
    .Z(_01887_));
 MUX2_X1 _25068_ (.A(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .B(_06660_),
    .S(_06980_),
    .Z(_01888_));
 MUX2_X1 _25069_ (.A(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .B(_06661_),
    .S(_06980_),
    .Z(_01889_));
 NAND2_X4 _25070_ (.A1(_11311_),
    .A2(_06647_),
    .ZN(_06985_));
 BUF_X4 _25071_ (.A(_06985_),
    .Z(_06986_));
 MUX2_X1 _25072_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(_06986_),
    .Z(_01890_));
 NAND2_X1 _25073_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .A2(_06982_),
    .ZN(_06987_));
 OAI21_X1 _25074_ (.A(_06987_),
    .B1(_06984_),
    .B2(_06905_),
    .ZN(_01891_));
 BUF_X4 _25075_ (.A(_06979_),
    .Z(_06988_));
 MUX2_X1 _25076_ (.A(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .B(_06665_),
    .S(_06988_),
    .Z(_01892_));
 MUX2_X1 _25077_ (.A(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .B(_05941_),
    .S(_06988_),
    .Z(_01893_));
 MUX2_X1 _25078_ (.A(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .B(_06666_),
    .S(_06988_),
    .Z(_01894_));
 MUX2_X1 _25079_ (.A(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .B(_06667_),
    .S(_06988_),
    .Z(_01895_));
 MUX2_X1 _25080_ (.A(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .B(_06668_),
    .S(_06988_),
    .Z(_01896_));
 MUX2_X1 _25081_ (.A(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .B(_06088_),
    .S(_06988_),
    .Z(_01897_));
 NAND2_X1 _25082_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .A2(_06982_),
    .ZN(_06989_));
 OAI21_X1 _25083_ (.A(_06989_),
    .B1(_06984_),
    .B2(_06823_),
    .ZN(_01898_));
 MUX2_X1 _25084_ (.A(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .B(_06132_),
    .S(_06988_),
    .Z(_01899_));
 MUX2_X1 _25085_ (.A(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .B(_06156_),
    .S(_06988_),
    .Z(_01900_));
 MUX2_X1 _25086_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(_06986_),
    .Z(_01901_));
 MUX2_X1 _25087_ (.A(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .B(_06178_),
    .S(_06988_),
    .Z(_01902_));
 NAND2_X1 _25088_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .A2(_06982_),
    .ZN(_06990_));
 OAI21_X1 _25089_ (.A(_06990_),
    .B1(_06984_),
    .B2(_06825_),
    .ZN(_01903_));
 NAND2_X1 _25090_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .A2(_06982_),
    .ZN(_06991_));
 OAI21_X1 _25091_ (.A(_06991_),
    .B1(_06984_),
    .B2(_06827_),
    .ZN(_01904_));
 MUX2_X1 _25092_ (.A(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .B(net460),
    .S(_06988_),
    .Z(_01905_));
 NAND2_X1 _25093_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .A2(_06982_),
    .ZN(_06992_));
 OAI21_X1 _25094_ (.A(_06992_),
    .B1(_06984_),
    .B2(_06829_),
    .ZN(_01906_));
 NAND2_X1 _25095_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .A2(_06982_),
    .ZN(_06993_));
 OAI21_X2 _25096_ (.A(_06993_),
    .B1(_06984_),
    .B2(net487),
    .ZN(_01907_));
 MUX2_X1 _25097_ (.A(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .B(net485),
    .S(_06979_),
    .Z(_01908_));
 NAND2_X1 _25098_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .A2(_06982_),
    .ZN(_06994_));
 OAI21_X1 _25099_ (.A(_06994_),
    .B1(_06984_),
    .B2(_06834_),
    .ZN(_01909_));
 NAND2_X1 _25100_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .A2(_06982_),
    .ZN(_06995_));
 OAI21_X1 _25101_ (.A(_06995_),
    .B1(_06984_),
    .B2(_06836_),
    .ZN(_01910_));
 MUX2_X1 _25102_ (.A(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .B(_06679_),
    .S(_06979_),
    .Z(_01911_));
 MUX2_X1 _25103_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(_06986_),
    .Z(_01912_));
 NAND2_X1 _25104_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .A2(_06982_),
    .ZN(_06996_));
 OAI21_X2 _25105_ (.A(_06996_),
    .B1(_06984_),
    .B2(_06838_),
    .ZN(_01913_));
 NAND2_X1 _25106_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .A2(_06981_),
    .ZN(_06997_));
 NAND2_X1 _25107_ (.A1(_06623_),
    .A2(_06980_),
    .ZN(_06998_));
 OAI21_X4 _25108_ (.A(_06997_),
    .B1(_06841_),
    .B2(_06998_),
    .ZN(_01914_));
 AND2_X2 _25109_ (.A1(_06629_),
    .A2(_06957_),
    .ZN(_06999_));
 BUF_X4 _25110_ (.A(_06999_),
    .Z(_07000_));
 MUX2_X1 _25111_ (.A(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .B(_06646_),
    .S(_07000_),
    .Z(_01915_));
 MUX2_X1 _25112_ (.A(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .B(_06650_),
    .S(_07000_),
    .Z(_01916_));
 MUX2_X1 _25113_ (.A(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .B(_06651_),
    .S(_07000_),
    .Z(_01917_));
 MUX2_X1 _25114_ (.A(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .B(_06652_),
    .S(_07000_),
    .Z(_01918_));
 MUX2_X1 _25115_ (.A(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .B(_06653_),
    .S(_07000_),
    .Z(_01919_));
 MUX2_X1 _25116_ (.A(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .B(_06654_),
    .S(_07000_),
    .Z(_01920_));
 NAND2_X2 _25117_ (.A1(_06629_),
    .A2(_06957_),
    .ZN(_07001_));
 BUF_X4 _25118_ (.A(_07001_),
    .Z(_07002_));
 NAND2_X1 _25119_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .A2(_07002_),
    .ZN(_07003_));
 BUF_X4 _25120_ (.A(_07001_),
    .Z(_07004_));
 CLKBUF_X3 _25121_ (.A(_05662_),
    .Z(_07005_));
 OAI21_X1 _25122_ (.A(_07003_),
    .B1(_07004_),
    .B2(_07005_),
    .ZN(_01921_));
 MUX2_X1 _25123_ (.A(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .B(_05736_),
    .S(_07000_),
    .Z(_01922_));
 MUX2_X1 _25124_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(_06986_),
    .Z(_01923_));
 MUX2_X1 _25125_ (.A(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .B(_06660_),
    .S(_07000_),
    .Z(_01924_));
 MUX2_X1 _25126_ (.A(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .B(_06661_),
    .S(_07000_),
    .Z(_01925_));
 NAND2_X1 _25127_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .A2(_07002_),
    .ZN(_07006_));
 OAI21_X1 _25128_ (.A(_07006_),
    .B1(_07004_),
    .B2(_06905_),
    .ZN(_01926_));
 BUF_X4 _25129_ (.A(_06999_),
    .Z(_07007_));
 MUX2_X1 _25130_ (.A(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .B(_06665_),
    .S(_07007_),
    .Z(_01927_));
 MUX2_X1 _25131_ (.A(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .B(_05941_),
    .S(_07007_),
    .Z(_01928_));
 MUX2_X1 _25132_ (.A(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .B(_06666_),
    .S(_07007_),
    .Z(_01929_));
 MUX2_X1 _25133_ (.A(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .B(_06667_),
    .S(_07007_),
    .Z(_01930_));
 MUX2_X1 _25134_ (.A(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .B(_06668_),
    .S(_07007_),
    .Z(_01931_));
 MUX2_X1 _25135_ (.A(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .B(_06088_),
    .S(_07007_),
    .Z(_01932_));
 NAND2_X1 _25136_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .A2(_07002_),
    .ZN(_07008_));
 CLKBUF_X3 _25137_ (.A(_06108_),
    .Z(_07009_));
 OAI21_X1 _25138_ (.A(_07008_),
    .B1(_07004_),
    .B2(_07009_),
    .ZN(_01933_));
 MUX2_X1 _25139_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(_06986_),
    .Z(_01934_));
 MUX2_X1 _25140_ (.A(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .B(_06132_),
    .S(_07007_),
    .Z(_01935_));
 MUX2_X1 _25141_ (.A(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .B(_06156_),
    .S(_07007_),
    .Z(_01936_));
 MUX2_X1 _25142_ (.A(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .B(_06178_),
    .S(_07007_),
    .Z(_01937_));
 NAND2_X1 _25143_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .A2(_07002_),
    .ZN(_07010_));
 CLKBUF_X3 _25144_ (.A(_06202_),
    .Z(_07011_));
 OAI21_X1 _25145_ (.A(_07010_),
    .B1(_07004_),
    .B2(_07011_),
    .ZN(_01938_));
 NAND2_X1 _25146_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .A2(_07002_),
    .ZN(_07012_));
 BUF_X4 _25147_ (.A(_06230_),
    .Z(_07013_));
 OAI21_X1 _25148_ (.A(_07012_),
    .B1(_07004_),
    .B2(_07013_),
    .ZN(_01939_));
 MUX2_X1 _25149_ (.A(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .B(net460),
    .S(_07007_),
    .Z(_01940_));
 NAND2_X1 _25150_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .A2(_07002_),
    .ZN(_07014_));
 CLKBUF_X3 _25151_ (.A(_06283_),
    .Z(_07015_));
 OAI21_X1 _25152_ (.A(_07014_),
    .B1(_07004_),
    .B2(_07015_),
    .ZN(_01941_));
 NAND2_X1 _25153_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .A2(_07002_),
    .ZN(_07016_));
 BUF_X8 _25154_ (.A(_06309_),
    .Z(_07017_));
 OAI21_X1 _25155_ (.A(_07016_),
    .B1(_07004_),
    .B2(_07017_),
    .ZN(_01942_));
 MUX2_X1 _25156_ (.A(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .B(_06675_),
    .S(_06999_),
    .Z(_01943_));
 NAND2_X1 _25157_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .A2(_07002_),
    .ZN(_07018_));
 BUF_X4 _25158_ (.A(_06360_),
    .Z(_07019_));
 OAI21_X1 _25159_ (.A(_07018_),
    .B1(_07004_),
    .B2(_07019_),
    .ZN(_01944_));
 MUX2_X1 _25160_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(_06986_),
    .Z(_01945_));
 NAND2_X1 _25161_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .A2(_05977_),
    .ZN(_07020_));
 OAI21_X1 _25162_ (.A(_07020_),
    .B1(_05663_),
    .B2(_05980_),
    .ZN(_01946_));
 NAND2_X1 _25163_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .A2(_07002_),
    .ZN(_07021_));
 BUF_X4 _25164_ (.A(_06391_),
    .Z(_07022_));
 OAI21_X1 _25165_ (.A(_07021_),
    .B1(_07004_),
    .B2(_07022_),
    .ZN(_01947_));
 MUX2_X1 _25166_ (.A(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .B(net450),
    .S(_06999_),
    .Z(_01948_));
 NAND2_X1 _25167_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .A2(_07002_),
    .ZN(_07023_));
 BUF_X8 _25168_ (.A(_06456_),
    .Z(_07024_));
 OAI21_X4 _25169_ (.A(_07023_),
    .B1(_07024_),
    .B2(_07004_),
    .ZN(_01949_));
 NAND2_X1 _25170_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .A2(_07001_),
    .ZN(_07025_));
 NAND2_X1 _25171_ (.A1(_06747_),
    .A2(_07000_),
    .ZN(_07026_));
 BUF_X16 _25172_ (.A(net372),
    .Z(_07027_));
 OAI21_X4 _25173_ (.A(_07025_),
    .B1(_07027_),
    .B2(_07026_),
    .ZN(_01950_));
 NAND2_X4 _25174_ (.A1(_06647_),
    .A2(_06957_),
    .ZN(_07028_));
 BUF_X4 _25175_ (.A(_07028_),
    .Z(_07029_));
 MUX2_X1 _25176_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S(_07029_),
    .Z(_01951_));
 MUX2_X1 _25177_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S(_07029_),
    .Z(_01952_));
 MUX2_X1 _25178_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S(_07029_),
    .Z(_01953_));
 MUX2_X1 _25179_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S(_07029_),
    .Z(_01954_));
 MUX2_X1 _25180_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S(_07029_),
    .Z(_01955_));
 MUX2_X1 _25181_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S(_07029_),
    .Z(_01956_));
 CLKBUF_X3 _25182_ (.A(_06985_),
    .Z(_07030_));
 NAND2_X1 _25183_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .A2(_07030_),
    .ZN(_07031_));
 OAI21_X1 _25184_ (.A(_07031_),
    .B1(_07030_),
    .B2(_07005_),
    .ZN(_01957_));
 BUF_X4 _25185_ (.A(_07028_),
    .Z(_07032_));
 NAND2_X1 _25186_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .A2(_07032_),
    .ZN(_07033_));
 OAI21_X1 _25187_ (.A(_07033_),
    .B1(_07032_),
    .B2(_07005_),
    .ZN(_01958_));
 NAND2_X4 _25188_ (.A1(_06657_),
    .A2(_06957_),
    .ZN(_07034_));
 MUX2_X1 _25189_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S(_07034_),
    .Z(_01959_));
 MUX2_X1 _25190_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S(_07029_),
    .Z(_01960_));
 MUX2_X1 _25191_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S(_07029_),
    .Z(_01961_));
 BUF_X4 _25192_ (.A(_07034_),
    .Z(_07035_));
 NAND2_X1 _25193_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .A2(_07035_),
    .ZN(_07036_));
 OAI21_X1 _25194_ (.A(_07036_),
    .B1(_07035_),
    .B2(_06905_),
    .ZN(_01962_));
 MUX2_X1 _25195_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S(_07029_),
    .Z(_01963_));
 MUX2_X1 _25196_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S(_07034_),
    .Z(_01964_));
 MUX2_X1 _25197_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S(_07028_),
    .Z(_01965_));
 MUX2_X1 _25198_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S(_07028_),
    .Z(_01966_));
 MUX2_X1 _25199_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S(_07028_),
    .Z(_01967_));
 NAND2_X4 _25200_ (.A1(_11311_),
    .A2(_06657_),
    .ZN(_07037_));
 MUX2_X1 _25201_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(_07037_),
    .Z(_01968_));
 MUX2_X1 _25202_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S(_07034_),
    .Z(_01969_));
 NAND2_X1 _25203_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .A2(_07032_),
    .ZN(_07038_));
 OAI21_X1 _25204_ (.A(_07038_),
    .B1(_07035_),
    .B2(_07009_),
    .ZN(_01970_));
 MUX2_X1 _25205_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S(_07034_),
    .Z(_01971_));
 MUX2_X1 _25206_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S(_07034_),
    .Z(_01972_));
 MUX2_X1 _25207_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S(_07034_),
    .Z(_01973_));
 NAND2_X1 _25208_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .A2(_07032_),
    .ZN(_07039_));
 OAI21_X1 _25209_ (.A(_07039_),
    .B1(_07035_),
    .B2(_07011_),
    .ZN(_01974_));
 NAND2_X1 _25210_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .A2(_07032_),
    .ZN(_07040_));
 OAI21_X1 _25211_ (.A(_07040_),
    .B1(_07035_),
    .B2(_07013_),
    .ZN(_01975_));
 MUX2_X1 _25212_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S(_07028_),
    .Z(_01976_));
 NAND2_X1 _25213_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .A2(_07032_),
    .ZN(_07041_));
 OAI21_X1 _25214_ (.A(_07041_),
    .B1(_07035_),
    .B2(_07015_),
    .ZN(_01977_));
 NAND2_X1 _25215_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .A2(_07032_),
    .ZN(_07042_));
 OAI21_X1 _25216_ (.A(_07042_),
    .B1(_07035_),
    .B2(_07017_),
    .ZN(_01978_));
 MUX2_X1 _25217_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(_06986_),
    .Z(_01979_));
 MUX2_X1 _25218_ (.A(net483),
    .B(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S(_07028_),
    .Z(_01980_));
 NAND2_X1 _25219_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .A2(_07032_),
    .ZN(_07043_));
 OAI21_X1 _25220_ (.A(_07043_),
    .B1(_07035_),
    .B2(_07019_),
    .ZN(_01981_));
 NAND2_X1 _25221_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .A2(_07032_),
    .ZN(_07044_));
 OAI21_X1 _25222_ (.A(_07044_),
    .B1(_07035_),
    .B2(_07022_),
    .ZN(_01982_));
 MUX2_X1 _25223_ (.A(_06806_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S(_07028_),
    .Z(_01983_));
 NAND2_X1 _25224_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .A2(_07032_),
    .ZN(_07045_));
 OAI21_X2 _25225_ (.A(_07045_),
    .B1(_07035_),
    .B2(_07024_),
    .ZN(_01984_));
 NAND2_X1 _25226_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .A2(_07029_),
    .ZN(_07046_));
 NAND3_X1 _25227_ (.A1(_06747_),
    .A2(_06682_),
    .A3(_06957_),
    .ZN(_07047_));
 OAI21_X4 _25228_ (.A(_07046_),
    .B1(net371),
    .B2(_07047_),
    .ZN(_01985_));
 NOR2_X1 _25229_ (.A1(_06878_),
    .A2(_06684_),
    .ZN(_07048_));
 BUF_X4 _25230_ (.A(_07048_),
    .Z(_07049_));
 NAND2_X4 _25231_ (.A1(_05495_),
    .A2(_07049_),
    .ZN(_07050_));
 BUF_X4 _25232_ (.A(_07050_),
    .Z(_07051_));
 MUX2_X1 _25233_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .S(_07051_),
    .Z(_01986_));
 MUX2_X1 _25234_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .S(_07051_),
    .Z(_01987_));
 MUX2_X1 _25235_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .S(_07051_),
    .Z(_01988_));
 MUX2_X1 _25236_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .S(_07051_),
    .Z(_01989_));
 MUX2_X1 _25237_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(_06986_),
    .Z(_01990_));
 MUX2_X1 _25238_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .S(_07051_),
    .Z(_01991_));
 MUX2_X1 _25239_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .S(_07051_),
    .Z(_01992_));
 BUF_X4 _25240_ (.A(_07050_),
    .Z(_07052_));
 NAND2_X1 _25241_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .A2(_07052_),
    .ZN(_07053_));
 OAI21_X1 _25242_ (.A(_07053_),
    .B1(_07052_),
    .B2(_07005_),
    .ZN(_01993_));
 NAND2_X4 _25243_ (.A1(_05737_),
    .A2(_07049_),
    .ZN(_07054_));
 MUX2_X1 _25244_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .S(_07054_),
    .Z(_01994_));
 MUX2_X1 _25245_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .S(_07051_),
    .Z(_01995_));
 MUX2_X1 _25246_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .S(_07051_),
    .Z(_01996_));
 BUF_X4 _25247_ (.A(_07054_),
    .Z(_07055_));
 NAND2_X1 _25248_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .A2(_07055_),
    .ZN(_07056_));
 OAI21_X1 _25249_ (.A(_07056_),
    .B1(_07055_),
    .B2(_06905_),
    .ZN(_01997_));
 MUX2_X1 _25250_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .S(_07051_),
    .Z(_01998_));
 MUX2_X1 _25251_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .S(_07054_),
    .Z(_01999_));
 MUX2_X1 _25252_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .S(_07050_),
    .Z(_02000_));
 CLKBUF_X3 _25253_ (.A(_07037_),
    .Z(_07057_));
 NAND2_X1 _25254_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .A2(_07057_),
    .ZN(_07058_));
 OAI21_X1 _25255_ (.A(_07058_),
    .B1(_07057_),
    .B2(_06905_),
    .ZN(_02001_));
 MUX2_X1 _25256_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .S(_07050_),
    .Z(_02002_));
 MUX2_X1 _25257_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .S(_07050_),
    .Z(_02003_));
 MUX2_X1 _25258_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .S(_07054_),
    .Z(_02004_));
 NAND2_X1 _25259_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .A2(_07052_),
    .ZN(_07059_));
 OAI21_X1 _25260_ (.A(_07059_),
    .B1(_07055_),
    .B2(_07009_),
    .ZN(_02005_));
 MUX2_X1 _25261_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .S(_07054_),
    .Z(_02006_));
 MUX2_X1 _25262_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .S(_07054_),
    .Z(_02007_));
 MUX2_X1 _25263_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .S(_07054_),
    .Z(_02008_));
 NAND2_X1 _25264_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .A2(_07052_),
    .ZN(_07060_));
 OAI21_X1 _25265_ (.A(_07060_),
    .B1(_07055_),
    .B2(_07011_),
    .ZN(_02009_));
 NAND2_X1 _25266_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .A2(_07052_),
    .ZN(_07061_));
 OAI21_X1 _25267_ (.A(_07061_),
    .B1(_07055_),
    .B2(_07013_),
    .ZN(_02010_));
 MUX2_X1 _25268_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .S(_07050_),
    .Z(_02011_));
 MUX2_X1 _25269_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(_06986_),
    .Z(_02012_));
 NAND2_X1 _25270_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .A2(_07052_),
    .ZN(_07062_));
 OAI21_X1 _25271_ (.A(_07062_),
    .B1(_07055_),
    .B2(_07015_),
    .ZN(_02013_));
 NAND2_X1 _25272_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .A2(_07052_),
    .ZN(_07063_));
 OAI21_X1 _25273_ (.A(_07063_),
    .B1(_07055_),
    .B2(_07017_),
    .ZN(_02014_));
 MUX2_X1 _25274_ (.A(_06803_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .S(_07050_),
    .Z(_02015_));
 NAND2_X1 _25275_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .A2(_07052_),
    .ZN(_07064_));
 OAI21_X1 _25276_ (.A(_07064_),
    .B1(_07055_),
    .B2(_07019_),
    .ZN(_02016_));
 NAND2_X1 _25277_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .A2(_07052_),
    .ZN(_07065_));
 OAI21_X1 _25278_ (.A(_07065_),
    .B1(_07055_),
    .B2(_07022_),
    .ZN(_02017_));
 MUX2_X1 _25279_ (.A(net599),
    .B(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .S(_07050_),
    .Z(_02018_));
 NAND2_X1 _25280_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .A2(_07052_),
    .ZN(_07066_));
 OAI21_X4 _25281_ (.A(_07066_),
    .B1(_07024_),
    .B2(_07055_),
    .ZN(_02019_));
 NAND2_X1 _25282_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A2(_07051_),
    .ZN(_07067_));
 NAND3_X1 _25283_ (.A1(_05591_),
    .A2(_06483_),
    .A3(_07049_),
    .ZN(_07068_));
 OAI21_X4 _25284_ (.A(_07067_),
    .B1(_07027_),
    .B2(_07068_),
    .ZN(_02020_));
 AND2_X1 _25285_ (.A1(_05410_),
    .A2(_07049_),
    .ZN(_07069_));
 BUF_X4 _25286_ (.A(_07069_),
    .Z(_07070_));
 BUF_X4 _25287_ (.A(_07070_),
    .Z(_07071_));
 MUX2_X1 _25288_ (.A(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .B(_06646_),
    .S(_07071_),
    .Z(_02021_));
 MUX2_X1 _25289_ (.A(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .B(_06650_),
    .S(_07071_),
    .Z(_02022_));
 MUX2_X1 _25290_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(_07037_),
    .Z(_02023_));
 MUX2_X1 _25291_ (.A(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .B(_06651_),
    .S(_07071_),
    .Z(_02024_));
 MUX2_X1 _25292_ (.A(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .B(_06652_),
    .S(_07071_),
    .Z(_02025_));
 MUX2_X1 _25293_ (.A(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .B(_06653_),
    .S(_07071_),
    .Z(_02026_));
 MUX2_X1 _25294_ (.A(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .B(_06654_),
    .S(_07071_),
    .Z(_02027_));
 NAND2_X4 _25295_ (.A1(_05976_),
    .A2(_07049_),
    .ZN(_07072_));
 CLKBUF_X3 _25296_ (.A(_07072_),
    .Z(_07073_));
 NAND2_X1 _25297_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .A2(_07073_),
    .ZN(_07074_));
 OAI21_X1 _25298_ (.A(_07074_),
    .B1(_07073_),
    .B2(_07005_),
    .ZN(_02028_));
 MUX2_X1 _25299_ (.A(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .B(_05736_),
    .S(_07071_),
    .Z(_02029_));
 BUF_X4 _25300_ (.A(_07070_),
    .Z(_07075_));
 MUX2_X1 _25301_ (.A(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .B(_06660_),
    .S(_07075_),
    .Z(_02030_));
 MUX2_X1 _25302_ (.A(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .B(_06661_),
    .S(_07075_),
    .Z(_02031_));
 NOR2_X1 _25303_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .A2(_07071_),
    .ZN(_07076_));
 AOI21_X1 _25304_ (.A(_07076_),
    .B1(_07071_),
    .B2(_06664_),
    .ZN(_02032_));
 MUX2_X1 _25305_ (.A(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .B(_06665_),
    .S(_07075_),
    .Z(_02033_));
 MUX2_X1 _25306_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(_06985_),
    .Z(_02034_));
 MUX2_X1 _25307_ (.A(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .B(_05941_),
    .S(_07075_),
    .Z(_02035_));
 MUX2_X1 _25308_ (.A(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .B(_06666_),
    .S(_07075_),
    .Z(_02036_));
 MUX2_X1 _25309_ (.A(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .B(_06667_),
    .S(_07075_),
    .Z(_02037_));
 MUX2_X1 _25310_ (.A(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .B(_06668_),
    .S(_07075_),
    .Z(_02038_));
 MUX2_X1 _25311_ (.A(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .B(_06088_),
    .S(_07075_),
    .Z(_02039_));
 NAND2_X1 _25312_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .A2(_07072_),
    .ZN(_07077_));
 OAI21_X1 _25313_ (.A(_07077_),
    .B1(_07073_),
    .B2(_07009_),
    .ZN(_02040_));
 MUX2_X1 _25314_ (.A(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .B(_06132_),
    .S(_07075_),
    .Z(_02041_));
 MUX2_X1 _25315_ (.A(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .B(_06156_),
    .S(_07075_),
    .Z(_02042_));
 MUX2_X1 _25316_ (.A(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .B(_06178_),
    .S(_07070_),
    .Z(_02043_));
 NAND2_X1 _25317_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .A2(_07072_),
    .ZN(_07078_));
 OAI21_X1 _25318_ (.A(_07078_),
    .B1(_07073_),
    .B2(_07011_),
    .ZN(_02044_));
 MUX2_X1 _25319_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(_06985_),
    .Z(_02045_));
 NAND2_X1 _25320_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .A2(_07072_),
    .ZN(_07079_));
 OAI21_X1 _25321_ (.A(_07079_),
    .B1(_07073_),
    .B2(_07013_),
    .ZN(_02046_));
 MUX2_X1 _25322_ (.A(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .B(net460),
    .S(_07070_),
    .Z(_02047_));
 NAND2_X1 _25323_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .A2(_07072_),
    .ZN(_07080_));
 OAI21_X1 _25324_ (.A(_07080_),
    .B1(_07073_),
    .B2(_07015_),
    .ZN(_02048_));
 NAND2_X1 _25325_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .A2(_07072_),
    .ZN(_07081_));
 OAI21_X1 _25326_ (.A(_07081_),
    .B1(_07073_),
    .B2(_07017_),
    .ZN(_02049_));
 MUX2_X1 _25327_ (.A(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .B(net485),
    .S(_07070_),
    .Z(_02050_));
 NAND2_X1 _25328_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .A2(_07072_),
    .ZN(_07082_));
 OAI21_X1 _25329_ (.A(_07082_),
    .B1(_07073_),
    .B2(_07019_),
    .ZN(_02051_));
 NAND2_X1 _25330_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .A2(_07072_),
    .ZN(_07083_));
 OAI21_X1 _25331_ (.A(_07083_),
    .B1(_07073_),
    .B2(_07022_),
    .ZN(_02052_));
 MUX2_X1 _25332_ (.A(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .B(_06679_),
    .S(_07070_),
    .Z(_02053_));
 NAND2_X1 _25333_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A2(_07072_),
    .ZN(_07084_));
 OAI21_X4 _25334_ (.A(_07084_),
    .B1(net456),
    .B2(_07073_),
    .ZN(_02054_));
 NAND2_X1 _25335_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A2(_07072_),
    .ZN(_07085_));
 NAND2_X1 _25336_ (.A1(_06747_),
    .A2(_07071_),
    .ZN(_07086_));
 OAI21_X4 _25337_ (.A(_07085_),
    .B1(_07027_),
    .B2(_07086_),
    .ZN(_02055_));
 MUX2_X1 _25338_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(_06985_),
    .Z(_02056_));
 MUX2_X1 _25339_ (.A(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .B(_05736_),
    .S(_06659_),
    .Z(_02057_));
 AND2_X1 _25340_ (.A1(_06625_),
    .A2(_07049_),
    .ZN(_07087_));
 BUF_X4 _25341_ (.A(_07087_),
    .Z(_07088_));
 BUF_X4 _25342_ (.A(_07088_),
    .Z(_07089_));
 MUX2_X1 _25343_ (.A(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .B(_06646_),
    .S(_07089_),
    .Z(_02058_));
 MUX2_X1 _25344_ (.A(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .B(_06650_),
    .S(_07089_),
    .Z(_02059_));
 MUX2_X1 _25345_ (.A(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .B(_06651_),
    .S(_07089_),
    .Z(_02060_));
 MUX2_X1 _25346_ (.A(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .B(_06652_),
    .S(_07089_),
    .Z(_02061_));
 MUX2_X1 _25347_ (.A(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .B(_06653_),
    .S(_07089_),
    .Z(_02062_));
 MUX2_X1 _25348_ (.A(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .B(_06654_),
    .S(_07089_),
    .Z(_02063_));
 NAND2_X4 _25349_ (.A1(_06629_),
    .A2(_07049_),
    .ZN(_07090_));
 CLKBUF_X3 _25350_ (.A(_07090_),
    .Z(_07091_));
 NAND2_X1 _25351_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .A2(_07091_),
    .ZN(_07092_));
 OAI21_X1 _25352_ (.A(_07092_),
    .B1(_07091_),
    .B2(_07005_),
    .ZN(_02064_));
 MUX2_X1 _25353_ (.A(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .B(_05736_),
    .S(_07089_),
    .Z(_02065_));
 BUF_X4 _25354_ (.A(_07088_),
    .Z(_07093_));
 MUX2_X1 _25355_ (.A(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .B(_06660_),
    .S(_07093_),
    .Z(_02066_));
 MUX2_X1 _25356_ (.A(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .B(_06661_),
    .S(_07093_),
    .Z(_02067_));
 MUX2_X1 _25357_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(_07037_),
    .Z(_02068_));
 NOR2_X1 _25358_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .A2(_07089_),
    .ZN(_07094_));
 AOI21_X1 _25359_ (.A(_07094_),
    .B1(_07089_),
    .B2(_06664_),
    .ZN(_02069_));
 MUX2_X1 _25360_ (.A(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .B(_06665_),
    .S(_07093_),
    .Z(_02070_));
 MUX2_X1 _25361_ (.A(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .B(_05941_),
    .S(_07093_),
    .Z(_02071_));
 MUX2_X1 _25362_ (.A(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .B(_06666_),
    .S(_07093_),
    .Z(_02072_));
 MUX2_X1 _25363_ (.A(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .B(_06667_),
    .S(_07093_),
    .Z(_02073_));
 MUX2_X1 _25364_ (.A(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .B(_06668_),
    .S(_07093_),
    .Z(_02074_));
 MUX2_X1 _25365_ (.A(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .B(_06088_),
    .S(_07093_),
    .Z(_02075_));
 NAND2_X1 _25366_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .A2(_07090_),
    .ZN(_07095_));
 OAI21_X1 _25367_ (.A(_07095_),
    .B1(_07091_),
    .B2(_07009_),
    .ZN(_02076_));
 MUX2_X1 _25368_ (.A(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .B(_06132_),
    .S(_07093_),
    .Z(_02077_));
 MUX2_X1 _25369_ (.A(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .B(_06156_),
    .S(_07093_),
    .Z(_02078_));
 NAND2_X1 _25370_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .A2(_07030_),
    .ZN(_07096_));
 OAI21_X1 _25371_ (.A(_07096_),
    .B1(_07057_),
    .B2(_07009_),
    .ZN(_02079_));
 MUX2_X1 _25372_ (.A(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .B(_06178_),
    .S(_07088_),
    .Z(_02080_));
 NAND2_X1 _25373_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .A2(_07090_),
    .ZN(_07097_));
 OAI21_X1 _25374_ (.A(_07097_),
    .B1(_07091_),
    .B2(_07011_),
    .ZN(_02081_));
 NAND2_X1 _25375_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .A2(_07090_),
    .ZN(_07098_));
 OAI21_X1 _25376_ (.A(_07098_),
    .B1(_07091_),
    .B2(_07013_),
    .ZN(_02082_));
 MUX2_X1 _25377_ (.A(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .B(_06672_),
    .S(_07088_),
    .Z(_02083_));
 NAND2_X1 _25378_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .A2(_07090_),
    .ZN(_07099_));
 OAI21_X1 _25379_ (.A(_07099_),
    .B1(_07091_),
    .B2(_07015_),
    .ZN(_02084_));
 NAND2_X1 _25380_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .A2(_07090_),
    .ZN(_07100_));
 OAI21_X1 _25381_ (.A(_07100_),
    .B1(_07091_),
    .B2(_07017_),
    .ZN(_02085_));
 MUX2_X1 _25382_ (.A(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .B(_06675_),
    .S(_07088_),
    .Z(_02086_));
 NAND2_X1 _25383_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .A2(_07090_),
    .ZN(_07101_));
 OAI21_X1 _25384_ (.A(_07101_),
    .B1(_07091_),
    .B2(_07019_),
    .ZN(_02087_));
 NAND2_X1 _25385_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .A2(_07090_),
    .ZN(_07102_));
 OAI21_X1 _25386_ (.A(_07102_),
    .B1(_07091_),
    .B2(_07022_),
    .ZN(_02088_));
 MUX2_X1 _25387_ (.A(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .B(_06679_),
    .S(_07088_),
    .Z(_02089_));
 MUX2_X1 _25388_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(_07037_),
    .Z(_02090_));
 NAND2_X1 _25389_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .A2(_07090_),
    .ZN(_07103_));
 OAI21_X4 _25390_ (.A(_07103_),
    .B1(net456),
    .B2(_07091_),
    .ZN(_02091_));
 NAND2_X1 _25391_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .A2(_07090_),
    .ZN(_07104_));
 NAND2_X1 _25392_ (.A1(_06747_),
    .A2(_07089_),
    .ZN(_07105_));
 OAI21_X4 _25393_ (.A(_07104_),
    .B1(net371),
    .B2(_07105_),
    .ZN(_02092_));
 NAND2_X4 _25394_ (.A1(_06647_),
    .A2(_07049_),
    .ZN(_07106_));
 BUF_X4 _25395_ (.A(_07106_),
    .Z(_07107_));
 MUX2_X1 _25396_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .S(_07107_),
    .Z(_02093_));
 MUX2_X1 _25397_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .S(_07107_),
    .Z(_02094_));
 MUX2_X1 _25398_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .S(_07107_),
    .Z(_02095_));
 MUX2_X1 _25399_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .S(_07107_),
    .Z(_02096_));
 MUX2_X1 _25400_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S(_07107_),
    .Z(_02097_));
 MUX2_X1 _25401_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .S(_07107_),
    .Z(_02098_));
 BUF_X4 _25402_ (.A(_07106_),
    .Z(_07108_));
 NAND2_X1 _25403_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .A2(_07108_),
    .ZN(_07109_));
 OAI21_X1 _25404_ (.A(_07109_),
    .B1(_07108_),
    .B2(_07005_),
    .ZN(_02099_));
 NAND2_X4 _25405_ (.A1(_06657_),
    .A2(_07049_),
    .ZN(_07110_));
 MUX2_X1 _25406_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .S(_07110_),
    .Z(_02100_));
 MUX2_X1 _25407_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(_07037_),
    .Z(_02101_));
 MUX2_X1 _25408_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .S(_07107_),
    .Z(_02102_));
 MUX2_X1 _25409_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .S(_07107_),
    .Z(_02103_));
 BUF_X4 _25410_ (.A(_07110_),
    .Z(_07111_));
 NAND2_X1 _25411_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .A2(_07111_),
    .ZN(_07112_));
 OAI21_X1 _25412_ (.A(_07112_),
    .B1(_07111_),
    .B2(_06905_),
    .ZN(_02104_));
 MUX2_X1 _25413_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .S(_07107_),
    .Z(_02105_));
 MUX2_X1 _25414_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S(_07110_),
    .Z(_02106_));
 MUX2_X1 _25415_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S(_07106_),
    .Z(_02107_));
 MUX2_X1 _25416_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S(_07106_),
    .Z(_02108_));
 MUX2_X1 _25417_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S(_07106_),
    .Z(_02109_));
 MUX2_X1 _25418_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S(_07110_),
    .Z(_02110_));
 NAND2_X1 _25419_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .A2(_07108_),
    .ZN(_07113_));
 OAI21_X1 _25420_ (.A(_07113_),
    .B1(_07111_),
    .B2(_07009_),
    .ZN(_02111_));
 MUX2_X1 _25421_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(_07037_),
    .Z(_02112_));
 MUX2_X1 _25422_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S(_07110_),
    .Z(_02113_));
 MUX2_X1 _25423_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S(_07110_),
    .Z(_02114_));
 MUX2_X1 _25424_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S(_07110_),
    .Z(_02115_));
 NAND2_X1 _25425_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .A2(_07108_),
    .ZN(_07114_));
 OAI21_X1 _25426_ (.A(_07114_),
    .B1(_07111_),
    .B2(_07011_),
    .ZN(_02116_));
 NAND2_X1 _25427_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .A2(_07108_),
    .ZN(_07115_));
 OAI21_X1 _25428_ (.A(_07115_),
    .B1(_07111_),
    .B2(_07013_),
    .ZN(_02117_));
 MUX2_X1 _25429_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S(_07106_),
    .Z(_02118_));
 NAND2_X1 _25430_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .A2(_07108_),
    .ZN(_07116_));
 OAI21_X1 _25431_ (.A(_07116_),
    .B1(_07111_),
    .B2(_07015_),
    .ZN(_02119_));
 NAND2_X1 _25432_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .A2(_07108_),
    .ZN(_07117_));
 OAI21_X1 _25433_ (.A(_07117_),
    .B1(_07111_),
    .B2(_07017_),
    .ZN(_02120_));
 MUX2_X1 _25434_ (.A(net483),
    .B(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S(_07106_),
    .Z(_02121_));
 NAND2_X1 _25435_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .A2(_07108_),
    .ZN(_07118_));
 OAI21_X1 _25436_ (.A(_07118_),
    .B1(_07111_),
    .B2(_07019_),
    .ZN(_02122_));
 NAND2_X1 _25437_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .A2(_07030_),
    .ZN(_07119_));
 OAI21_X1 _25438_ (.A(_07119_),
    .B1(_07057_),
    .B2(_07011_),
    .ZN(_02123_));
 NAND2_X1 _25439_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .A2(_07108_),
    .ZN(_07120_));
 OAI21_X1 _25440_ (.A(_07120_),
    .B1(_07111_),
    .B2(_07022_),
    .ZN(_02124_));
 MUX2_X1 _25441_ (.A(_06806_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S(_07106_),
    .Z(_02125_));
 NAND2_X1 _25442_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .A2(_07108_),
    .ZN(_07121_));
 OAI21_X4 _25443_ (.A(_07121_),
    .B1(net456),
    .B2(_07111_),
    .ZN(_02126_));
 NAND2_X1 _25444_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .A2(_07107_),
    .ZN(_07122_));
 NAND3_X1 _25445_ (.A1(_06483_),
    .A2(_06682_),
    .A3(_07049_),
    .ZN(_07123_));
 OAI21_X4 _25446_ (.A(_07122_),
    .B1(net371),
    .B2(_07123_),
    .ZN(_02127_));
 NOR2_X4 _25447_ (.A1(_06878_),
    .A2(_06770_),
    .ZN(_07124_));
 NAND2_X4 _25448_ (.A1(_05495_),
    .A2(_07124_),
    .ZN(_07125_));
 BUF_X4 _25449_ (.A(_07125_),
    .Z(_07126_));
 MUX2_X1 _25450_ (.A(_06769_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .S(_07126_),
    .Z(_02128_));
 MUX2_X1 _25451_ (.A(_06775_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .S(_07126_),
    .Z(_02129_));
 MUX2_X1 _25452_ (.A(_06776_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .S(_07126_),
    .Z(_02130_));
 MUX2_X1 _25453_ (.A(_06777_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .S(_07126_),
    .Z(_02131_));
 MUX2_X1 _25454_ (.A(_06778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .S(_07126_),
    .Z(_02132_));
 MUX2_X1 _25455_ (.A(_06779_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .S(_07126_),
    .Z(_02133_));
 NAND2_X1 _25456_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .A2(_07030_),
    .ZN(_07127_));
 OAI21_X1 _25457_ (.A(_07127_),
    .B1(_07057_),
    .B2(_07013_),
    .ZN(_02134_));
 BUF_X4 _25458_ (.A(_07125_),
    .Z(_07128_));
 NAND2_X1 _25459_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .A2(_07128_),
    .ZN(_07129_));
 OAI21_X1 _25460_ (.A(_07129_),
    .B1(_07128_),
    .B2(_07005_),
    .ZN(_02135_));
 NAND2_X4 _25461_ (.A1(_05737_),
    .A2(_07124_),
    .ZN(_07130_));
 MUX2_X1 _25462_ (.A(_06782_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .S(_07130_),
    .Z(_02136_));
 MUX2_X1 _25463_ (.A(_06784_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .S(_07126_),
    .Z(_02137_));
 MUX2_X1 _25464_ (.A(_06785_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .S(_07126_),
    .Z(_02138_));
 BUF_X4 _25465_ (.A(_07130_),
    .Z(_07131_));
 NAND2_X1 _25466_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .A2(_07131_),
    .ZN(_07132_));
 OAI21_X1 _25467_ (.A(_07132_),
    .B1(_07131_),
    .B2(_06905_),
    .ZN(_02139_));
 MUX2_X1 _25468_ (.A(_06788_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .S(_07126_),
    .Z(_02140_));
 MUX2_X1 _25469_ (.A(_06789_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .S(_07130_),
    .Z(_02141_));
 MUX2_X1 _25470_ (.A(_06790_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .S(_07125_),
    .Z(_02142_));
 MUX2_X1 _25471_ (.A(_06791_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .S(_07125_),
    .Z(_02143_));
 MUX2_X1 _25472_ (.A(_06792_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .S(_07125_),
    .Z(_02144_));
 MUX2_X1 _25473_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(_06985_),
    .Z(_02145_));
 MUX2_X1 _25474_ (.A(_06793_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .S(_07130_),
    .Z(_02146_));
 NAND2_X1 _25475_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .A2(_07128_),
    .ZN(_07133_));
 OAI21_X1 _25476_ (.A(_07133_),
    .B1(_07131_),
    .B2(_07009_),
    .ZN(_02147_));
 MUX2_X1 _25477_ (.A(_06795_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .S(_07130_),
    .Z(_02148_));
 MUX2_X1 _25478_ (.A(_06796_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .S(_07130_),
    .Z(_02149_));
 MUX2_X1 _25479_ (.A(_06797_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .S(_07130_),
    .Z(_02150_));
 NAND2_X1 _25480_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .A2(_07128_),
    .ZN(_07134_));
 OAI21_X1 _25481_ (.A(_07134_),
    .B1(_07131_),
    .B2(_07011_),
    .ZN(_02151_));
 NAND2_X1 _25482_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .A2(_07128_),
    .ZN(_07135_));
 OAI21_X1 _25483_ (.A(_07135_),
    .B1(_07131_),
    .B2(_07013_),
    .ZN(_02152_));
 MUX2_X1 _25484_ (.A(_06800_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .S(_07125_),
    .Z(_02153_));
 NAND2_X1 _25485_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .A2(_07128_),
    .ZN(_07136_));
 OAI21_X1 _25486_ (.A(_07136_),
    .B1(_07131_),
    .B2(_07015_),
    .ZN(_02154_));
 NAND2_X1 _25487_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .A2(_07128_),
    .ZN(_07137_));
 OAI21_X1 _25488_ (.A(_07137_),
    .B1(_07131_),
    .B2(_07017_),
    .ZN(_02155_));
 NAND2_X1 _25489_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .A2(_07030_),
    .ZN(_07138_));
 OAI21_X1 _25490_ (.A(_07138_),
    .B1(_07057_),
    .B2(_07015_),
    .ZN(_02156_));
 MUX2_X1 _25491_ (.A(_06803_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .S(_07125_),
    .Z(_02157_));
 NAND2_X1 _25492_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .A2(_07128_),
    .ZN(_07139_));
 OAI21_X1 _25493_ (.A(_07139_),
    .B1(_07131_),
    .B2(_07019_),
    .ZN(_02158_));
 NAND2_X1 _25494_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .A2(_07128_),
    .ZN(_07140_));
 OAI21_X1 _25495_ (.A(_07140_),
    .B1(_07131_),
    .B2(_07022_),
    .ZN(_02159_));
 MUX2_X1 _25496_ (.A(_06806_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .S(_07125_),
    .Z(_02160_));
 NAND2_X1 _25497_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .A2(_07128_),
    .ZN(_07141_));
 OAI21_X4 _25498_ (.A(_07141_),
    .B1(_07024_),
    .B2(_07131_),
    .ZN(_02161_));
 NAND2_X1 _25499_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A2(_07126_),
    .ZN(_07142_));
 NAND3_X1 _25500_ (.A1(_05591_),
    .A2(_06483_),
    .A3(_07124_),
    .ZN(_07143_));
 OAI21_X4 _25501_ (.A(_07142_),
    .B1(_07027_),
    .B2(_07143_),
    .ZN(_02162_));
 AND2_X1 _25502_ (.A1(_05410_),
    .A2(_07124_),
    .ZN(_07144_));
 BUF_X4 _25503_ (.A(_07144_),
    .Z(_07145_));
 BUF_X4 _25504_ (.A(_07145_),
    .Z(_07146_));
 MUX2_X1 _25505_ (.A(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .B(_06646_),
    .S(_07146_),
    .Z(_02163_));
 MUX2_X1 _25506_ (.A(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .B(_06650_),
    .S(_07146_),
    .Z(_02164_));
 MUX2_X1 _25507_ (.A(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .B(_06651_),
    .S(_07146_),
    .Z(_02165_));
 MUX2_X1 _25508_ (.A(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .B(_06652_),
    .S(_07146_),
    .Z(_02166_));
 NAND2_X1 _25509_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .A2(_07030_),
    .ZN(_07147_));
 OAI21_X1 _25510_ (.A(_07147_),
    .B1(_07057_),
    .B2(_07017_),
    .ZN(_02167_));
 MUX2_X1 _25511_ (.A(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .B(_06660_),
    .S(_05411_),
    .Z(_02168_));
 MUX2_X1 _25512_ (.A(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .B(_06653_),
    .S(_07146_),
    .Z(_02169_));
 MUX2_X1 _25513_ (.A(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .B(_06654_),
    .S(_07146_),
    .Z(_02170_));
 NAND2_X4 _25514_ (.A1(_05976_),
    .A2(_07124_),
    .ZN(_07148_));
 BUF_X4 _25515_ (.A(_07148_),
    .Z(_07149_));
 NAND2_X1 _25516_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .A2(_07149_),
    .ZN(_07150_));
 OAI21_X1 _25517_ (.A(_07150_),
    .B1(_07149_),
    .B2(_07005_),
    .ZN(_02171_));
 MUX2_X1 _25518_ (.A(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .B(_05736_),
    .S(_07146_),
    .Z(_02172_));
 BUF_X4 _25519_ (.A(_07145_),
    .Z(_07151_));
 MUX2_X1 _25520_ (.A(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .B(_06660_),
    .S(_07151_),
    .Z(_02173_));
 MUX2_X1 _25521_ (.A(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .B(_06661_),
    .S(_07151_),
    .Z(_02174_));
 NOR2_X1 _25522_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .A2(_07146_),
    .ZN(_07152_));
 AOI21_X1 _25523_ (.A(_07152_),
    .B1(_07146_),
    .B2(_06664_),
    .ZN(_02175_));
 MUX2_X1 _25524_ (.A(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .B(_06665_),
    .S(_07151_),
    .Z(_02176_));
 MUX2_X1 _25525_ (.A(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .B(_05941_),
    .S(_07151_),
    .Z(_02177_));
 MUX2_X1 _25526_ (.A(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .B(_06666_),
    .S(_07151_),
    .Z(_02178_));
 MUX2_X1 _25527_ (.A(_06803_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(_06985_),
    .Z(_02179_));
 MUX2_X1 _25528_ (.A(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .B(_06667_),
    .S(_07151_),
    .Z(_02180_));
 MUX2_X1 _25529_ (.A(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .B(_06668_),
    .S(_07151_),
    .Z(_02181_));
 MUX2_X1 _25530_ (.A(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .B(_06088_),
    .S(_07151_),
    .Z(_02182_));
 NAND2_X1 _25531_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .A2(_07148_),
    .ZN(_07153_));
 OAI21_X1 _25532_ (.A(_07153_),
    .B1(_07149_),
    .B2(_07009_),
    .ZN(_02183_));
 MUX2_X1 _25533_ (.A(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .B(_06132_),
    .S(_07151_),
    .Z(_02184_));
 MUX2_X1 _25534_ (.A(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .B(_06156_),
    .S(_07151_),
    .Z(_02185_));
 MUX2_X1 _25535_ (.A(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .B(_06178_),
    .S(_07145_),
    .Z(_02186_));
 NAND2_X1 _25536_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .A2(_07148_),
    .ZN(_07154_));
 OAI21_X1 _25537_ (.A(_07154_),
    .B1(_07149_),
    .B2(_07011_),
    .ZN(_02187_));
 NAND2_X1 _25538_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .A2(_07148_),
    .ZN(_07155_));
 OAI21_X1 _25539_ (.A(_07155_),
    .B1(_07149_),
    .B2(_07013_),
    .ZN(_02188_));
 MUX2_X1 _25540_ (.A(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .B(net460),
    .S(_07145_),
    .Z(_02189_));
 NAND2_X1 _25541_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .A2(_07030_),
    .ZN(_07156_));
 OAI21_X1 _25542_ (.A(_07156_),
    .B1(_07057_),
    .B2(_07019_),
    .ZN(_02190_));
 NAND2_X1 _25543_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .A2(_07148_),
    .ZN(_07157_));
 OAI21_X1 _25544_ (.A(_07157_),
    .B1(_07149_),
    .B2(_07015_),
    .ZN(_02191_));
 NAND2_X1 _25545_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .A2(_07148_),
    .ZN(_07158_));
 OAI21_X1 _25546_ (.A(_07158_),
    .B1(_07149_),
    .B2(_07017_),
    .ZN(_02192_));
 MUX2_X1 _25547_ (.A(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .B(net485),
    .S(_07145_),
    .Z(_02193_));
 NAND2_X1 _25548_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .A2(_07148_),
    .ZN(_07159_));
 OAI21_X1 _25549_ (.A(_07159_),
    .B1(_07149_),
    .B2(_07019_),
    .ZN(_02194_));
 NAND2_X1 _25550_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .A2(_07148_),
    .ZN(_07160_));
 OAI21_X1 _25551_ (.A(_07160_),
    .B1(_07149_),
    .B2(_07022_),
    .ZN(_02195_));
 MUX2_X1 _25552_ (.A(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .B(_06679_),
    .S(_07145_),
    .Z(_02196_));
 NAND2_X1 _25553_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .A2(_07148_),
    .ZN(_07161_));
 OAI21_X4 _25554_ (.A(_07161_),
    .B1(net456),
    .B2(_07149_),
    .ZN(_02197_));
 NAND2_X1 _25555_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A2(_07148_),
    .ZN(_07162_));
 NAND2_X1 _25556_ (.A1(_06747_),
    .A2(_07146_),
    .ZN(_07163_));
 OAI21_X4 _25557_ (.A(_07162_),
    .B1(net371),
    .B2(_07163_),
    .ZN(_02198_));
 AND2_X1 _25558_ (.A1(_06625_),
    .A2(_07124_),
    .ZN(_07164_));
 BUF_X4 _25559_ (.A(_07164_),
    .Z(_07165_));
 BUF_X4 _25560_ (.A(_07165_),
    .Z(_07166_));
 MUX2_X1 _25561_ (.A(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .B(_06646_),
    .S(_07166_),
    .Z(_02199_));
 MUX2_X1 _25562_ (.A(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .B(_06650_),
    .S(_07166_),
    .Z(_02200_));
 NAND2_X1 _25563_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .A2(_07030_),
    .ZN(_07167_));
 OAI21_X1 _25564_ (.A(_07167_),
    .B1(_07057_),
    .B2(_07022_),
    .ZN(_02201_));
 MUX2_X1 _25565_ (.A(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .B(_06651_),
    .S(_07166_),
    .Z(_02202_));
 MUX2_X1 _25566_ (.A(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .B(_06652_),
    .S(_07166_),
    .Z(_02203_));
 MUX2_X1 _25567_ (.A(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .B(_06653_),
    .S(_07166_),
    .Z(_02204_));
 MUX2_X1 _25568_ (.A(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .B(_06654_),
    .S(_07166_),
    .Z(_02205_));
 NAND2_X4 _25569_ (.A1(_06629_),
    .A2(_07124_),
    .ZN(_07168_));
 BUF_X4 _25570_ (.A(_07168_),
    .Z(_07169_));
 NAND2_X1 _25571_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .A2(_07169_),
    .ZN(_07170_));
 OAI21_X1 _25572_ (.A(_07170_),
    .B1(_07169_),
    .B2(_07005_),
    .ZN(_02206_));
 MUX2_X1 _25573_ (.A(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .B(_05736_),
    .S(_07166_),
    .Z(_02207_));
 BUF_X4 _25574_ (.A(_07165_),
    .Z(_07171_));
 MUX2_X1 _25575_ (.A(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .B(_06660_),
    .S(_07171_),
    .Z(_02208_));
 MUX2_X1 _25576_ (.A(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .B(_06661_),
    .S(_07171_),
    .Z(_02209_));
 NOR2_X1 _25577_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .A2(_07166_),
    .ZN(_07172_));
 AOI21_X1 _25578_ (.A(_07172_),
    .B1(_07166_),
    .B2(_06664_),
    .ZN(_02210_));
 MUX2_X1 _25579_ (.A(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .B(_06665_),
    .S(_07171_),
    .Z(_02211_));
 MUX2_X1 _25580_ (.A(net599),
    .B(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(_06985_),
    .Z(_02212_));
 MUX2_X1 _25581_ (.A(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .B(_05941_),
    .S(_07171_),
    .Z(_02213_));
 MUX2_X1 _25582_ (.A(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .B(_06666_),
    .S(_07171_),
    .Z(_02214_));
 MUX2_X1 _25583_ (.A(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .B(_06667_),
    .S(_07171_),
    .Z(_02215_));
 MUX2_X1 _25584_ (.A(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .B(_06668_),
    .S(_07171_),
    .Z(_02216_));
 MUX2_X1 _25585_ (.A(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .B(_06088_),
    .S(_07171_),
    .Z(_02217_));
 NAND2_X1 _25586_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .A2(_07168_),
    .ZN(_07173_));
 OAI21_X1 _25587_ (.A(_07173_),
    .B1(_07169_),
    .B2(_07009_),
    .ZN(_02218_));
 MUX2_X1 _25588_ (.A(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .B(_06132_),
    .S(_07171_),
    .Z(_02219_));
 MUX2_X1 _25589_ (.A(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .B(_06156_),
    .S(_07171_),
    .Z(_02220_));
 MUX2_X1 _25590_ (.A(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .B(_06178_),
    .S(_07165_),
    .Z(_02221_));
 NAND2_X1 _25591_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .A2(_07168_),
    .ZN(_07174_));
 OAI21_X1 _25592_ (.A(_07174_),
    .B1(_07169_),
    .B2(_07011_),
    .ZN(_02222_));
 NAND2_X1 _25593_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .A2(_07030_),
    .ZN(_07175_));
 OAI21_X4 _25594_ (.A(_07175_),
    .B1(_07024_),
    .B2(_07057_),
    .ZN(_02223_));
 NAND2_X1 _25595_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .A2(_07168_),
    .ZN(_07176_));
 OAI21_X1 _25596_ (.A(_07176_),
    .B1(_07169_),
    .B2(_07013_),
    .ZN(_02224_));
 MUX2_X1 _25597_ (.A(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .B(_06672_),
    .S(_07165_),
    .Z(_02225_));
 NAND2_X1 _25598_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .A2(_07168_),
    .ZN(_07177_));
 OAI21_X1 _25599_ (.A(_07177_),
    .B1(_07169_),
    .B2(_07015_),
    .ZN(_02226_));
 NAND2_X1 _25600_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .A2(_07168_),
    .ZN(_07178_));
 OAI21_X1 _25601_ (.A(_07178_),
    .B1(_07169_),
    .B2(_07017_),
    .ZN(_02227_));
 MUX2_X1 _25602_ (.A(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .B(net485),
    .S(_07165_),
    .Z(_02228_));
 NAND2_X1 _25603_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .A2(_07168_),
    .ZN(_07179_));
 OAI21_X1 _25604_ (.A(_07179_),
    .B1(_07169_),
    .B2(_07019_),
    .ZN(_02229_));
 NAND2_X1 _25605_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .A2(_07168_),
    .ZN(_07180_));
 OAI21_X1 _25606_ (.A(_07180_),
    .B1(_07169_),
    .B2(_07022_),
    .ZN(_02230_));
 MUX2_X1 _25607_ (.A(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .B(net450),
    .S(_07165_),
    .Z(_02231_));
 NAND2_X1 _25608_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .A2(_07168_),
    .ZN(_07181_));
 OAI21_X4 _25609_ (.A(_07181_),
    .B1(net456),
    .B2(_07169_),
    .ZN(_02232_));
 NAND2_X1 _25610_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .A2(_07168_),
    .ZN(_07182_));
 NAND2_X1 _25611_ (.A1(_06747_),
    .A2(_07166_),
    .ZN(_07183_));
 OAI21_X4 _25612_ (.A(_07182_),
    .B1(_07027_),
    .B2(_07183_),
    .ZN(_02233_));
 NAND2_X1 _25613_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .A2(_06986_),
    .ZN(_07184_));
 NAND3_X1 _25614_ (.A1(_11311_),
    .A2(_06482_),
    .A3(_06682_),
    .ZN(_07185_));
 OAI21_X4 _25615_ (.A(_07184_),
    .B1(net371),
    .B2(_07185_),
    .ZN(_02234_));
 NOR2_X4 _25616_ (.A1(_11471_),
    .A2(_06770_),
    .ZN(_07186_));
 NAND2_X4 _25617_ (.A1(_06647_),
    .A2(_07186_),
    .ZN(_07187_));
 BUF_X4 _25618_ (.A(_07187_),
    .Z(_07188_));
 MUX2_X1 _25619_ (.A(_05402_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S(_07188_),
    .Z(_02235_));
 MUX2_X1 _25620_ (.A(_06525_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S(_07188_),
    .Z(_02236_));
 MUX2_X1 _25621_ (.A(_06565_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S(_07188_),
    .Z(_02237_));
 MUX2_X1 _25622_ (.A(_06602_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S(_07188_),
    .Z(_02238_));
 MUX2_X1 _25623_ (.A(_05491_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S(_07188_),
    .Z(_02239_));
 MUX2_X1 _25624_ (.A(_05589_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S(_07188_),
    .Z(_02240_));
 CLKBUF_X3 _25625_ (.A(_07187_),
    .Z(_07189_));
 NAND2_X1 _25626_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .A2(_07189_),
    .ZN(_07190_));
 OAI21_X1 _25627_ (.A(_07190_),
    .B1(_07189_),
    .B2(_05662_),
    .ZN(_02241_));
 NAND2_X4 _25628_ (.A1(_06657_),
    .A2(_07186_),
    .ZN(_07191_));
 MUX2_X1 _25629_ (.A(_05735_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S(_07191_),
    .Z(_02242_));
 MUX2_X1 _25630_ (.A(_05778_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S(_07188_),
    .Z(_02243_));
 MUX2_X1 _25631_ (.A(_05815_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S(_07188_),
    .Z(_02244_));
 MUX2_X1 _25632_ (.A(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .B(_06646_),
    .S(_05497_),
    .Z(_02245_));
 CLKBUF_X3 _25633_ (.A(_07191_),
    .Z(_07192_));
 NAND2_X1 _25634_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .A2(_07192_),
    .ZN(_07193_));
 OAI21_X1 _25635_ (.A(_07193_),
    .B1(_07192_),
    .B2(_05868_),
    .ZN(_02246_));
 MUX2_X1 _25636_ (.A(_05908_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S(_07188_),
    .Z(_02247_));
 MUX2_X1 _25637_ (.A(_05940_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S(_07191_),
    .Z(_02248_));
 MUX2_X1 _25638_ (.A(_05974_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S(_07187_),
    .Z(_02249_));
 MUX2_X1 _25639_ (.A(_06026_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S(_07187_),
    .Z(_02250_));
 MUX2_X1 _25640_ (.A(_06054_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S(_07187_),
    .Z(_02251_));
 MUX2_X1 _25641_ (.A(_06087_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S(_07191_),
    .Z(_02252_));
 NAND2_X1 _25642_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .A2(_07189_),
    .ZN(_07194_));
 OAI21_X1 _25643_ (.A(_07194_),
    .B1(_07192_),
    .B2(_06108_),
    .ZN(_02253_));
 MUX2_X1 _25644_ (.A(_06131_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S(_07191_),
    .Z(_02254_));
 MUX2_X1 _25645_ (.A(_06155_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S(_07191_),
    .Z(_02255_));
 MUX2_X1 _25646_ (.A(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .B(_06650_),
    .S(_05497_),
    .Z(_02256_));
 MUX2_X1 _25647_ (.A(_06177_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S(_07191_),
    .Z(_02257_));
 NAND2_X1 _25648_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .A2(_07189_),
    .ZN(_07195_));
 OAI21_X1 _25649_ (.A(_07195_),
    .B1(_07192_),
    .B2(_06202_),
    .ZN(_02258_));
 NAND2_X1 _25650_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .A2(_07189_),
    .ZN(_07196_));
 OAI21_X1 _25651_ (.A(_07196_),
    .B1(_07192_),
    .B2(_06230_),
    .ZN(_02259_));
 MUX2_X1 _25652_ (.A(net461),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S(_07187_),
    .Z(_02260_));
 NAND2_X1 _25653_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .A2(_07189_),
    .ZN(_07197_));
 OAI21_X1 _25654_ (.A(_07197_),
    .B1(_07192_),
    .B2(_06283_),
    .ZN(_02261_));
 NAND2_X1 _25655_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .A2(_07189_),
    .ZN(_07198_));
 OAI21_X1 _25656_ (.A(_07198_),
    .B1(_07192_),
    .B2(_06309_),
    .ZN(_02262_));
 MUX2_X1 _25657_ (.A(_06328_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S(_07187_),
    .Z(_02263_));
 NAND2_X1 _25658_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .A2(_07189_),
    .ZN(_07199_));
 OAI21_X1 _25659_ (.A(_07199_),
    .B1(_07192_),
    .B2(_06360_),
    .ZN(_02264_));
 NAND2_X1 _25660_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .A2(_07189_),
    .ZN(_07200_));
 OAI21_X2 _25661_ (.A(_07200_),
    .B1(_06391_),
    .B2(_07192_),
    .ZN(_02265_));
 MUX2_X1 _25662_ (.A(_06422_),
    .B(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S(_07187_),
    .Z(_02266_));
 MUX2_X1 _25663_ (.A(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .B(_06651_),
    .S(_05497_),
    .Z(_02267_));
 NAND2_X1 _25664_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .A2(_07189_),
    .ZN(_07201_));
 OAI21_X2 _25665_ (.A(_07201_),
    .B1(_06456_),
    .B2(_07192_),
    .ZN(_02268_));
 NAND2_X1 _25666_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .A2(_07188_),
    .ZN(_07202_));
 NAND3_X1 _25667_ (.A1(_06483_),
    .A2(_06682_),
    .A3(_07186_),
    .ZN(_07203_));
 OAI21_X4 _25668_ (.A(_07202_),
    .B1(net372),
    .B2(_07203_),
    .ZN(_02269_));
 MUX2_X1 _25669_ (.A(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .B(_06652_),
    .S(_05497_),
    .Z(_02270_));
 MUX2_X1 _25670_ (.A(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .B(_06661_),
    .S(_05411_),
    .Z(_02271_));
 NAND2_X4 _25671_ (.A1(_10820_),
    .A2(_11293_),
    .ZN(_07204_));
 AOI21_X1 _25672_ (.A(_07204_),
    .B1(_05408_),
    .B2(_10795_),
    .ZN(_07205_));
 NAND2_X1 _25673_ (.A1(_10794_),
    .A2(_07205_),
    .ZN(_07206_));
 AOI21_X1 _25674_ (.A(_05393_),
    .B1(_04006_),
    .B2(_03528_),
    .ZN(_07207_));
 AND3_X1 _25675_ (.A1(_10942_),
    .A2(_11865_),
    .A3(_04005_),
    .ZN(_07208_));
 OAI21_X1 _25676_ (.A(_10795_),
    .B1(_07207_),
    .B2(_07208_),
    .ZN(_07209_));
 NAND2_X1 _25677_ (.A1(_04005_),
    .A2(_05394_),
    .ZN(_07210_));
 NAND3_X2 _25678_ (.A1(_03687_),
    .A2(_07209_),
    .A3(_07210_),
    .ZN(_07211_));
 AOI21_X4 _25679_ (.A(_03537_),
    .B1(_07206_),
    .B2(_07211_),
    .ZN(_07212_));
 OR4_X1 _25680_ (.A1(\alu_adder_result_ex[14] ),
    .A2(\alu_adder_result_ex[22] ),
    .A3(\alu_adder_result_ex[27] ),
    .A4(\alu_adder_result_ex[29] ),
    .ZN(_07213_));
 NOR3_X1 _25681_ (.A1(\alu_adder_result_ex[26] ),
    .A2(\alu_adder_result_ex[30] ),
    .A3(_07213_),
    .ZN(_07214_));
 OR3_X1 _25682_ (.A1(\alu_adder_result_ex[16] ),
    .A2(\alu_adder_result_ex[18] ),
    .A3(\alu_adder_result_ex[4] ),
    .ZN(_07215_));
 NOR4_X1 _25683_ (.A1(\alu_adder_result_ex[10] ),
    .A2(\alu_adder_result_ex[12] ),
    .A3(\alu_adder_result_ex[25] ),
    .A4(\alu_adder_result_ex[2] ),
    .ZN(_07216_));
 NAND3_X1 _25684_ (.A1(_12271_),
    .A2(_12881_),
    .A3(_03709_),
    .ZN(_07217_));
 NOR4_X1 _25685_ (.A1(\alu_adder_result_ex[15] ),
    .A2(\alu_adder_result_ex[21] ),
    .A3(\alu_adder_result_ex[23] ),
    .A4(_07217_),
    .ZN(_07218_));
 NOR2_X1 _25686_ (.A1(\alu_adder_result_ex[6] ),
    .A2(\alu_adder_result_ex[19] ),
    .ZN(_07219_));
 NAND4_X1 _25687_ (.A1(_12286_),
    .A2(_07216_),
    .A3(_07218_),
    .A4(_07219_),
    .ZN(_07220_));
 NOR4_X1 _25688_ (.A1(\alu_adder_result_ex[24] ),
    .A2(\alu_adder_result_ex[28] ),
    .A3(_07215_),
    .A4(_07220_),
    .ZN(_07221_));
 NOR2_X1 _25689_ (.A1(\alu_adder_result_ex[20] ),
    .A2(net313),
    .ZN(_07222_));
 AND4_X1 _25690_ (.A1(_07214_),
    .A2(_07221_),
    .A3(_07222_),
    .A4(_05200_),
    .ZN(_07223_));
 AOI211_X2 _25691_ (.A(_05198_),
    .B(_07223_),
    .C1(_05199_),
    .C2(_03732_),
    .ZN(_07224_));
 NAND2_X2 _25692_ (.A1(_10796_),
    .A2(_03739_),
    .ZN(_07225_));
 OR4_X4 _25693_ (.A1(_10942_),
    .A2(_04006_),
    .A3(_07224_),
    .A4(_07225_),
    .ZN(_07226_));
 INV_X4 _25694_ (.A(_07226_),
    .ZN(\id_stage_i.branch_set_d ));
 NOR2_X1 _25695_ (.A1(_07212_),
    .A2(\id_stage_i.branch_set_d ),
    .ZN(_07227_));
 NOR3_X4 _25696_ (.A1(_03564_),
    .A2(_03978_),
    .A3(_03994_),
    .ZN(_07228_));
 AOI21_X1 _25697_ (.A(_03998_),
    .B1(_03997_),
    .B2(_10794_),
    .ZN(_07229_));
 OR2_X1 _25698_ (.A1(_04086_),
    .A2(_07229_),
    .ZN(_07230_));
 NAND2_X1 _25699_ (.A1(_03532_),
    .A2(_07230_),
    .ZN(_07231_));
 OR3_X1 _25700_ (.A1(_04009_),
    .A2(_07228_),
    .A3(_07231_),
    .ZN(_07232_));
 OAI21_X1 _25701_ (.A(_03533_),
    .B1(_07227_),
    .B2(_07232_),
    .ZN(_07233_));
 CLKBUF_X3 _25702_ (.A(_04083_),
    .Z(_07234_));
 NOR2_X1 _25703_ (.A1(_11304_),
    .A2(_03668_),
    .ZN(_07235_));
 OR2_X1 _25704_ (.A1(\id_stage_i.controller_i.load_err_d ),
    .A2(\id_stage_i.controller_i.store_err_d ),
    .ZN(_07236_));
 NOR3_X1 _25705_ (.A1(_10711_),
    .A2(_15927_),
    .A3(_03674_),
    .ZN(_07237_));
 NOR3_X1 _25706_ (.A1(_03646_),
    .A2(_11322_),
    .A3(_03669_),
    .ZN(_07238_));
 AOI21_X1 _25707_ (.A(_07237_),
    .B1(_07238_),
    .B2(_15927_),
    .ZN(_07239_));
 OR4_X1 _25708_ (.A1(_10810_),
    .A2(_11323_),
    .A3(_04473_),
    .A4(_07239_),
    .ZN(_07240_));
 INV_X1 _25709_ (.A(_07240_),
    .ZN(_07241_));
 OR4_X2 _25710_ (.A1(_03665_),
    .A2(_07235_),
    .A3(_07236_),
    .A4(_07241_),
    .ZN(_07242_));
 NOR2_X1 _25711_ (.A1(\id_stage_i.controller_i.exc_req_d ),
    .A2(_07242_),
    .ZN(_07243_));
 NOR2_X2 _25712_ (.A1(_04006_),
    .A2(_07225_),
    .ZN(_07244_));
 NAND2_X2 _25713_ (.A1(net333),
    .A2(_07244_),
    .ZN(_07245_));
 NOR2_X2 _25714_ (.A1(_07224_),
    .A2(_07245_),
    .ZN(_07246_));
 OR3_X1 _25715_ (.A1(_07212_),
    .A2(_07230_),
    .A3(_07246_),
    .ZN(_07247_));
 NAND3_X1 _25716_ (.A1(_07234_),
    .A2(_07243_),
    .A3(_07247_),
    .ZN(_07248_));
 NOR3_X2 _25717_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_03678_),
    .A3(_04011_),
    .ZN(_07249_));
 AOI21_X1 _25718_ (.A(_07230_),
    .B1(_07249_),
    .B2(_04018_),
    .ZN(_07250_));
 OR2_X1 _25719_ (.A1(_04014_),
    .A2(_07250_),
    .ZN(_07251_));
 NOR2_X1 _25720_ (.A1(_04015_),
    .A2(_04029_),
    .ZN(_07252_));
 AOI21_X2 _25721_ (.A(_07251_),
    .B1(_07252_),
    .B2(_03665_),
    .ZN(_07253_));
 NOR2_X1 _25722_ (.A1(_03997_),
    .A2(_03998_),
    .ZN(_07254_));
 NAND2_X1 _25723_ (.A1(_03994_),
    .A2(_07254_),
    .ZN(_07255_));
 NOR4_X2 _25724_ (.A1(_03534_),
    .A2(_03976_),
    .A3(_03979_),
    .A4(_07255_),
    .ZN(_07256_));
 NOR2_X1 _25725_ (.A1(_04009_),
    .A2(_03649_),
    .ZN(_07257_));
 NAND2_X1 _25726_ (.A1(_03531_),
    .A2(_03534_),
    .ZN(_07258_));
 AOI221_X1 _25727_ (.A(_04000_),
    .B1(_07231_),
    .B2(_07257_),
    .C1(_07258_),
    .C2(_04009_),
    .ZN(_07259_));
 NOR4_X1 _25728_ (.A1(_04035_),
    .A2(_07253_),
    .A3(_07256_),
    .A4(_07259_),
    .ZN(_07260_));
 AOI22_X1 _25729_ (.A1(_03996_),
    .A2(_07233_),
    .B1(_07248_),
    .B2(_07260_),
    .ZN(_02272_));
 NOR2_X1 _25730_ (.A1(_03649_),
    .A2(_07231_),
    .ZN(_07261_));
 AOI22_X1 _25731_ (.A1(_03531_),
    .A2(_03649_),
    .B1(_07228_),
    .B2(_07261_),
    .ZN(_07262_));
 NOR3_X1 _25732_ (.A1(_04009_),
    .A2(_04000_),
    .A3(_07262_),
    .ZN(_07263_));
 NOR4_X2 _25733_ (.A1(_10875_),
    .A2(_01161_),
    .A3(_11317_),
    .A4(_03674_),
    .ZN(_07264_));
 AOI22_X2 _25734_ (.A1(_03663_),
    .A2(_07264_),
    .B1(_07228_),
    .B2(_07241_),
    .ZN(_07265_));
 NOR3_X1 _25735_ (.A1(_04030_),
    .A2(_07251_),
    .A3(_07265_),
    .ZN(_07266_));
 OR2_X1 _25736_ (.A1(_03656_),
    .A2(_03658_),
    .ZN(_07267_));
 NOR3_X2 _25737_ (.A1(_03672_),
    .A2(_03681_),
    .A3(_07242_),
    .ZN(_07268_));
 AOI21_X4 _25738_ (.A(_04073_),
    .B1(_07267_),
    .B2(_07268_),
    .ZN(_07269_));
 NOR4_X1 _25739_ (.A1(_07256_),
    .A2(_07263_),
    .A3(_07266_),
    .A4(_07269_),
    .ZN(_07270_));
 AOI21_X1 _25740_ (.A(_03531_),
    .B1(_07227_),
    .B2(_07228_),
    .ZN(_07271_));
 NAND2_X1 _25741_ (.A1(_07234_),
    .A2(_07247_),
    .ZN(_07272_));
 OAI21_X1 _25742_ (.A(_07270_),
    .B1(_07271_),
    .B2(_07272_),
    .ZN(_02273_));
 INV_X1 _25743_ (.A(_04026_),
    .ZN(_07273_));
 NAND3_X1 _25744_ (.A1(_03534_),
    .A2(_04310_),
    .A3(_07230_),
    .ZN(_07274_));
 OAI21_X1 _25745_ (.A(_07274_),
    .B1(_03534_),
    .B2(_03533_),
    .ZN(_07275_));
 NAND2_X1 _25746_ (.A1(_03979_),
    .A2(_03996_),
    .ZN(_07276_));
 AOI222_X2 _25747_ (.A1(_07273_),
    .A2(_07253_),
    .B1(_07275_),
    .B2(_03532_),
    .C1(_04009_),
    .C2(_07276_),
    .ZN(_07277_));
 OR2_X1 _25748_ (.A1(\id_stage_i.controller_i.exc_req_d ),
    .A2(_07242_),
    .ZN(_07278_));
 OAI21_X1 _25749_ (.A(_07234_),
    .B1(_07278_),
    .B2(_07247_),
    .ZN(_07279_));
 AOI221_X1 _25750_ (.A(_07256_),
    .B1(_07277_),
    .B2(_07279_),
    .C1(_03996_),
    .C2(_04000_),
    .ZN(_02274_));
 OAI21_X1 _25751_ (.A(_03536_),
    .B1(_04026_),
    .B2(_07250_),
    .ZN(_07280_));
 NOR2_X1 _25752_ (.A1(_04086_),
    .A2(_07229_),
    .ZN(_07281_));
 NAND2_X1 _25753_ (.A1(_03650_),
    .A2(_07281_),
    .ZN(_07282_));
 AOI21_X1 _25754_ (.A(_04013_),
    .B1(_07227_),
    .B2(_07243_),
    .ZN(_07283_));
 OAI21_X1 _25755_ (.A(_07280_),
    .B1(_07282_),
    .B2(_07283_),
    .ZN(_02275_));
 OR3_X4 _25756_ (.A1(_03669_),
    .A2(_03668_),
    .A3(_04065_),
    .ZN(_07284_));
 NAND3_X4 _25757_ (.A1(_03532_),
    .A2(_04000_),
    .A3(_03649_),
    .ZN(_07285_));
 OAI21_X1 _25758_ (.A(_03975_),
    .B1(_03999_),
    .B2(_07285_),
    .ZN(_07286_));
 AND2_X1 _25759_ (.A1(_07284_),
    .A2(_07286_),
    .ZN(_02276_));
 NAND4_X4 _25760_ (.A1(_10971_),
    .A2(_11324_),
    .A3(_03667_),
    .A4(_04033_),
    .ZN(_07287_));
 NOR2_X4 _25761_ (.A1(_04037_),
    .A2(_07287_),
    .ZN(_07288_));
 BUF_X4 _25762_ (.A(_07288_),
    .Z(_07289_));
 OAI22_X1 _25763_ (.A1(_04060_),
    .A2(_03980_),
    .B1(_07289_),
    .B2(_03977_),
    .ZN(_02277_));
 NOR2_X1 _25764_ (.A1(_10942_),
    .A2(_07224_),
    .ZN(_07290_));
 NOR3_X1 _25765_ (.A1(_04006_),
    .A2(_07210_),
    .A3(_07290_),
    .ZN(_07291_));
 NOR3_X1 _25766_ (.A1(_03537_),
    .A2(_05408_),
    .A3(_07204_),
    .ZN(_07292_));
 NOR3_X1 _25767_ (.A1(_03653_),
    .A2(_05393_),
    .A3(_07292_),
    .ZN(_07293_));
 OAI22_X1 _25768_ (.A1(_07225_),
    .A2(_07291_),
    .B1(_07293_),
    .B2(_10796_),
    .ZN(_02278_));
 MUX2_X1 _25769_ (.A(_03786_),
    .B(net276),
    .S(_03925_),
    .Z(_07294_));
 CLKBUF_X3 _25770_ (.A(_03691_),
    .Z(_07295_));
 MUX2_X1 _25771_ (.A(_07294_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .S(_07295_),
    .Z(_02279_));
 CLKBUF_X3 _25772_ (.A(_03766_),
    .Z(_07296_));
 MUX2_X1 _25773_ (.A(\alu_adder_result_ex[10] ),
    .B(_11724_),
    .S(_07296_),
    .Z(_07297_));
 MUX2_X1 _25774_ (.A(_07297_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .S(_07295_),
    .Z(_02280_));
 MUX2_X1 _25775_ (.A(net486),
    .B(_11769_),
    .S(_07296_),
    .Z(_07298_));
 MUX2_X1 _25776_ (.A(_07298_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .S(_07295_),
    .Z(_02281_));
 MUX2_X1 _25777_ (.A(\alu_adder_result_ex[12] ),
    .B(_12420_),
    .S(_07296_),
    .Z(_07299_));
 MUX2_X1 _25778_ (.A(_07299_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .S(_07295_),
    .Z(_02282_));
 MUX2_X1 _25779_ (.A(\alu_adder_result_ex[13] ),
    .B(_12473_),
    .S(_07296_),
    .Z(_07300_));
 MUX2_X1 _25780_ (.A(_07300_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .S(_07295_),
    .Z(_02283_));
 MUX2_X1 _25781_ (.A(net7),
    .B(_12580_),
    .S(_07296_),
    .Z(_07301_));
 MUX2_X1 _25782_ (.A(_07301_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .S(_07295_),
    .Z(_02284_));
 MUX2_X1 _25783_ (.A(net439),
    .B(_12656_),
    .S(_07296_),
    .Z(_07302_));
 MUX2_X1 _25784_ (.A(_07302_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .S(_07295_),
    .Z(_02285_));
 MUX2_X1 _25785_ (.A(\alu_adder_result_ex[16] ),
    .B(net281),
    .S(_07296_),
    .Z(_07303_));
 MUX2_X1 _25786_ (.A(_07303_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .S(_07295_),
    .Z(_02286_));
 NAND2_X1 _25787_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .A2(_03692_),
    .ZN(_07304_));
 MUX2_X1 _25788_ (.A(_12881_),
    .B(_12825_),
    .S(_03925_),
    .Z(_07305_));
 OAI21_X1 _25789_ (.A(_07304_),
    .B1(_07305_),
    .B2(_03692_),
    .ZN(_02287_));
 MUX2_X1 _25790_ (.A(\alu_adder_result_ex[18] ),
    .B(net286),
    .S(_07296_),
    .Z(_07306_));
 MUX2_X1 _25791_ (.A(_07306_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .S(_07295_),
    .Z(_02288_));
 MUX2_X1 _25792_ (.A(\alu_adder_result_ex[19] ),
    .B(net283),
    .S(_07296_),
    .Z(_07307_));
 CLKBUF_X3 _25793_ (.A(_03690_),
    .Z(_07308_));
 MUX2_X1 _25794_ (.A(_07307_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .S(_07308_),
    .Z(_02289_));
 MUX2_X1 _25795_ (.A(_16491_),
    .B(net301),
    .S(_03766_),
    .Z(_07309_));
 NOR2_X1 _25796_ (.A1(_04172_),
    .A2(_07309_),
    .ZN(_07310_));
 MUX2_X1 _25797_ (.A(_07310_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .S(_07308_),
    .Z(_02290_));
 MUX2_X1 _25798_ (.A(\alu_adder_result_ex[20] ),
    .B(net368),
    .S(_07296_),
    .Z(_07311_));
 MUX2_X1 _25799_ (.A(_07311_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .S(_07308_),
    .Z(_02291_));
 CLKBUF_X3 _25800_ (.A(_03766_),
    .Z(_07312_));
 MUX2_X1 _25801_ (.A(\alu_adder_result_ex[21] ),
    .B(_13198_),
    .S(_07312_),
    .Z(_07313_));
 MUX2_X1 _25802_ (.A(_07313_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .S(_07308_),
    .Z(_02292_));
 MUX2_X1 _25803_ (.A(\alu_adder_result_ex[22] ),
    .B(net323),
    .S(_07312_),
    .Z(_07314_));
 MUX2_X1 _25804_ (.A(_07314_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .S(_07308_),
    .Z(_02293_));
 MUX2_X1 _25805_ (.A(net357),
    .B(net319),
    .S(_07312_),
    .Z(_07315_));
 MUX2_X1 _25806_ (.A(_07315_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .S(_07308_),
    .Z(_02294_));
 MUX2_X1 _25807_ (.A(\alu_adder_result_ex[24] ),
    .B(_13480_),
    .S(_07312_),
    .Z(_07316_));
 MUX2_X1 _25808_ (.A(_07316_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .S(_07308_),
    .Z(_02295_));
 MUX2_X1 _25809_ (.A(net389),
    .B(_13555_),
    .S(_07312_),
    .Z(_07317_));
 MUX2_X1 _25810_ (.A(_07317_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .S(_07308_),
    .Z(_02296_));
 NAND2_X1 _25811_ (.A1(_13648_),
    .A2(_03925_),
    .ZN(_07318_));
 OAI21_X1 _25812_ (.A(_07318_),
    .B1(_03925_),
    .B2(net392),
    .ZN(_07319_));
 MUX2_X1 _25813_ (.A(_07319_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .S(_07308_),
    .Z(_02297_));
 MUX2_X1 _25814_ (.A(\alu_adder_result_ex[27] ),
    .B(_03104_),
    .S(_07312_),
    .Z(_07320_));
 MUX2_X1 _25815_ (.A(_07320_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .S(_07308_),
    .Z(_02298_));
 MUX2_X1 _25816_ (.A(net386),
    .B(_03198_),
    .S(_07312_),
    .Z(_07321_));
 MUX2_X1 _25817_ (.A(_07321_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .S(_03691_),
    .Z(_02299_));
 MUX2_X1 _25818_ (.A(net411),
    .B(_03276_),
    .S(_07312_),
    .Z(_07322_));
 MUX2_X1 _25819_ (.A(_07322_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .S(_03691_),
    .Z(_02300_));
 MUX2_X1 _25820_ (.A(\alu_adder_result_ex[2] ),
    .B(net364),
    .S(_07312_),
    .Z(_07323_));
 MUX2_X1 _25821_ (.A(_07323_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .S(_03691_),
    .Z(_02301_));
 MUX2_X1 _25822_ (.A(net345),
    .B(_03372_),
    .S(_07312_),
    .Z(_07324_));
 MUX2_X1 _25823_ (.A(_07324_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .S(_03691_),
    .Z(_02302_));
 NAND2_X1 _25824_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .A2(_03692_),
    .ZN(_07325_));
 INV_X1 _25825_ (.A(_03765_),
    .ZN(_07326_));
 OAI21_X1 _25826_ (.A(_03452_),
    .B1(net289),
    .B2(_07326_),
    .ZN(_07327_));
 OAI21_X1 _25827_ (.A(_07325_),
    .B1(_07327_),
    .B2(_03692_),
    .ZN(_02303_));
 AND3_X1 _25828_ (.A1(_04176_),
    .A2(_03739_),
    .A3(_03773_),
    .ZN(_07328_));
 AND3_X1 _25829_ (.A1(_03686_),
    .A2(_07328_),
    .A3(_05152_),
    .ZN(_07329_));
 NOR2_X4 _25830_ (.A1(_03685_),
    .A2(_03774_),
    .ZN(_07330_));
 NOR4_X4 _25831_ (.A1(_03492_),
    .A2(_03493_),
    .A3(_03742_),
    .A4(_03683_),
    .ZN(_07331_));
 INV_X2 _25832_ (.A(_03490_),
    .ZN(_07332_));
 AOI221_X1 _25833_ (.A(_07331_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B2(_03683_),
    .C1(_07332_),
    .C2(_03786_),
    .ZN(_07333_));
 MUX2_X1 _25834_ (.A(_00118_),
    .B(_00116_),
    .S(_04967_),
    .Z(_07334_));
 MUX2_X1 _25835_ (.A(_00119_),
    .B(_00117_),
    .S(_04967_),
    .Z(_07335_));
 MUX2_X1 _25836_ (.A(_07334_),
    .B(_07335_),
    .S(_04964_),
    .Z(_07336_));
 MUX2_X1 _25837_ (.A(_00126_),
    .B(_00124_),
    .S(_04967_),
    .Z(_07337_));
 MUX2_X1 _25838_ (.A(_00127_),
    .B(_00125_),
    .S(_04967_),
    .Z(_07338_));
 MUX2_X1 _25839_ (.A(_07337_),
    .B(_07338_),
    .S(_04964_),
    .Z(_07339_));
 MUX2_X1 _25840_ (.A(_07336_),
    .B(_07339_),
    .S(_04978_),
    .Z(_07340_));
 MUX2_X1 _25841_ (.A(_00122_),
    .B(_00120_),
    .S(_04967_),
    .Z(_07341_));
 MUX2_X1 _25842_ (.A(_00123_),
    .B(_00121_),
    .S(_04968_),
    .Z(_07342_));
 MUX2_X1 _25843_ (.A(_07341_),
    .B(_07342_),
    .S(_04964_),
    .Z(_07343_));
 MUX2_X1 _25844_ (.A(_00130_),
    .B(_00128_),
    .S(_04967_),
    .Z(_07344_));
 MUX2_X1 _25845_ (.A(_00131_),
    .B(_00129_),
    .S(_04968_),
    .Z(_07345_));
 MUX2_X1 _25846_ (.A(_07344_),
    .B(_07345_),
    .S(_04964_),
    .Z(_07346_));
 MUX2_X1 _25847_ (.A(_07343_),
    .B(_07346_),
    .S(_04978_),
    .Z(_07347_));
 MUX2_X1 _25848_ (.A(_07340_),
    .B(_07347_),
    .S(_04973_),
    .Z(_07348_));
 MUX2_X1 _25849_ (.A(_00102_),
    .B(_00100_),
    .S(_04967_),
    .Z(_07349_));
 MUX2_X1 _25850_ (.A(_00103_),
    .B(_00101_),
    .S(_04968_),
    .Z(_07350_));
 MUX2_X1 _25851_ (.A(_07349_),
    .B(_07350_),
    .S(_04964_),
    .Z(_07351_));
 MUX2_X1 _25852_ (.A(_00110_),
    .B(_00108_),
    .S(_04968_),
    .Z(_07352_));
 MUX2_X1 _25853_ (.A(_00111_),
    .B(_00109_),
    .S(_04968_),
    .Z(_07353_));
 MUX2_X1 _25854_ (.A(_07352_),
    .B(_07353_),
    .S(_04964_),
    .Z(_07354_));
 MUX2_X1 _25855_ (.A(_07351_),
    .B(_07354_),
    .S(_04978_),
    .Z(_07355_));
 MUX2_X1 _25856_ (.A(_00106_),
    .B(_00104_),
    .S(_04968_),
    .Z(_07356_));
 MUX2_X1 _25857_ (.A(_00107_),
    .B(_00105_),
    .S(_04968_),
    .Z(_07357_));
 MUX2_X1 _25858_ (.A(_07356_),
    .B(_07357_),
    .S(_04964_),
    .Z(_07358_));
 MUX2_X1 _25859_ (.A(_00114_),
    .B(_00112_),
    .S(_04968_),
    .Z(_07359_));
 MUX2_X1 _25860_ (.A(_00115_),
    .B(_00113_),
    .S(_04968_),
    .Z(_07360_));
 MUX2_X1 _25861_ (.A(_07359_),
    .B(_07360_),
    .S(_04964_),
    .Z(_07361_));
 MUX2_X1 _25862_ (.A(_07358_),
    .B(_07361_),
    .S(_04978_),
    .Z(_07362_));
 MUX2_X1 _25863_ (.A(_07355_),
    .B(_07362_),
    .S(_04973_),
    .Z(_07363_));
 MUX2_X1 _25864_ (.A(_07348_),
    .B(_07363_),
    .S(_04981_),
    .Z(_07364_));
 OAI21_X1 _25865_ (.A(_07333_),
    .B1(_07364_),
    .B2(_03699_),
    .ZN(_07365_));
 NAND2_X2 _25866_ (.A1(_07331_),
    .A2(_03761_),
    .ZN(_07366_));
 OAI21_X1 _25867_ (.A(_07365_),
    .B1(_07366_),
    .B2(_03796_),
    .ZN(_07367_));
 INV_X1 _25868_ (.A(_07367_),
    .ZN(_07368_));
 CLKBUF_X3 _25869_ (.A(_03774_),
    .Z(_07369_));
 AOI221_X2 _25870_ (.A(_07329_),
    .B1(_07330_),
    .B2(_07368_),
    .C1(_07369_),
    .C2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .ZN(_07370_));
 INV_X1 _25871_ (.A(_03492_),
    .ZN(_07371_));
 OAI21_X1 _25872_ (.A(_07330_),
    .B1(_07366_),
    .B2(_11967_),
    .ZN(_07372_));
 OR2_X1 _25873_ (.A1(_07371_),
    .A2(_07372_),
    .ZN(_07373_));
 CLKBUF_X3 _25874_ (.A(_07373_),
    .Z(_07374_));
 MUX2_X1 _25875_ (.A(_00217_),
    .B(_16502_),
    .S(_05033_),
    .Z(_07375_));
 CLKBUF_X3 _25876_ (.A(_03761_),
    .Z(_07376_));
 MUX2_X1 _25877_ (.A(_05036_),
    .B(_07375_),
    .S(_07376_),
    .Z(_07377_));
 OAI21_X1 _25878_ (.A(_07370_),
    .B1(_07374_),
    .B2(_07377_),
    .ZN(_02304_));
 BUF_X4 _25879_ (.A(_07331_),
    .Z(_07378_));
 AOI21_X1 _25880_ (.A(_07378_),
    .B1(\alu_adder_result_ex[1] ),
    .B2(_07332_),
    .ZN(_07379_));
 MUX2_X1 _25881_ (.A(_00185_),
    .B(_16491_),
    .S(_05033_),
    .Z(_07380_));
 MUX2_X1 _25882_ (.A(_05080_),
    .B(_07380_),
    .S(_03761_),
    .Z(_07381_));
 OAI221_X2 _25883_ (.A(_07379_),
    .B1(_07381_),
    .B2(_07371_),
    .C1(_03699_),
    .C2(_07375_),
    .ZN(_07382_));
 CLKBUF_X3 _25884_ (.A(_07366_),
    .Z(_07383_));
 OAI21_X1 _25885_ (.A(_07382_),
    .B1(_07383_),
    .B2(_03811_),
    .ZN(_07384_));
 CLKBUF_X3 _25886_ (.A(_03738_),
    .Z(_07385_));
 AOI21_X1 _25887_ (.A(_06490_),
    .B1(_07384_),
    .B2(_07385_),
    .ZN(_07386_));
 CLKBUF_X3 _25888_ (.A(_07328_),
    .Z(_07387_));
 CLKBUF_X3 _25889_ (.A(_07387_),
    .Z(_07388_));
 MUX2_X1 _25890_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .B(_07386_),
    .S(_07388_),
    .Z(_02305_));
 CLKBUF_X3 _25891_ (.A(_03686_),
    .Z(_07389_));
 AND3_X1 _25892_ (.A1(_07389_),
    .A2(_07387_),
    .A3(_06535_),
    .ZN(_07390_));
 CLKBUF_X3 _25893_ (.A(_07369_),
    .Z(_07391_));
 AOI21_X1 _25894_ (.A(_07390_),
    .B1(_07391_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .ZN(_07392_));
 NOR2_X1 _25895_ (.A1(_03700_),
    .A2(_07380_),
    .ZN(_07393_));
 OAI21_X1 _25896_ (.A(_03771_),
    .B1(_04072_),
    .B2(_03490_),
    .ZN(_07394_));
 NOR2_X1 _25897_ (.A1(_07393_),
    .A2(_07394_),
    .ZN(_07395_));
 CLKBUF_X3 _25898_ (.A(_07330_),
    .Z(_07396_));
 CLKBUF_X3 _25899_ (.A(_07366_),
    .Z(_07397_));
 OAI21_X1 _25900_ (.A(_07396_),
    .B1(_07397_),
    .B2(_03820_),
    .ZN(_07398_));
 MUX2_X1 _25901_ (.A(_00558_),
    .B(_04072_),
    .S(_05033_),
    .Z(_07399_));
 MUX2_X1 _25902_ (.A(_05120_),
    .B(_07399_),
    .S(_07376_),
    .Z(_07400_));
 OAI221_X1 _25903_ (.A(_07392_),
    .B1(_07395_),
    .B2(_07398_),
    .C1(_07400_),
    .C2(_07374_),
    .ZN(_02306_));
 BUF_X2 _25904_ (.A(_07369_),
    .Z(_07401_));
 OR3_X1 _25905_ (.A1(_07385_),
    .A2(_07401_),
    .A3(_06583_),
    .ZN(_07402_));
 AOI21_X1 _25906_ (.A(_07378_),
    .B1(\alu_adder_result_ex[3] ),
    .B2(_07332_),
    .ZN(_07403_));
 OAI21_X1 _25907_ (.A(_07403_),
    .B1(_07399_),
    .B2(_03700_),
    .ZN(_07404_));
 NOR2_X2 _25908_ (.A1(_10882_),
    .A2(_03686_),
    .ZN(_07405_));
 CLKBUF_X3 _25909_ (.A(_07405_),
    .Z(_07406_));
 BUF_X4 _25910_ (.A(_07406_),
    .Z(_07407_));
 BUF_X4 _25911_ (.A(_05110_),
    .Z(_07408_));
 NOR2_X1 _25912_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_07408_),
    .ZN(_07409_));
 BUF_X4 _25913_ (.A(_07408_),
    .Z(_07410_));
 AOI21_X2 _25914_ (.A(_07409_),
    .B1(_07410_),
    .B2(_00559_),
    .ZN(_07411_));
 NOR2_X1 _25915_ (.A1(_07407_),
    .A2(_07411_),
    .ZN(_07412_));
 AOI21_X1 _25916_ (.A(_07412_),
    .B1(_05130_),
    .B2(_07407_),
    .ZN(_07413_));
 AOI21_X1 _25917_ (.A(_07404_),
    .B1(_07413_),
    .B2(_03781_),
    .ZN(_07414_));
 CLKBUF_X3 _25918_ (.A(_07387_),
    .Z(_07415_));
 OAI221_X1 _25919_ (.A(_07402_),
    .B1(_07414_),
    .B2(_07372_),
    .C1(_07415_),
    .C2(_06584_),
    .ZN(_02307_));
 AND3_X1 _25920_ (.A1(_07389_),
    .A2(_07328_),
    .A3(_05431_),
    .ZN(_07416_));
 AOI21_X1 _25921_ (.A(_07416_),
    .B1(_07391_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .ZN(_07417_));
 BUF_X4 _25922_ (.A(_07378_),
    .Z(_07418_));
 AOI221_X2 _25923_ (.A(_07418_),
    .B1(_07411_),
    .B2(_03784_),
    .C1(_07332_),
    .C2(\alu_adder_result_ex[4] ),
    .ZN(_07419_));
 OAI21_X1 _25924_ (.A(_07396_),
    .B1(_07397_),
    .B2(_12008_),
    .ZN(_07420_));
 MUX2_X1 _25925_ (.A(_00560_),
    .B(_03725_),
    .S(_05033_),
    .Z(_07421_));
 MUX2_X1 _25926_ (.A(_05134_),
    .B(_07421_),
    .S(_07376_),
    .Z(_07422_));
 OAI221_X1 _25927_ (.A(_07417_),
    .B1(_07419_),
    .B2(_07420_),
    .C1(_07422_),
    .C2(_07374_),
    .ZN(_02308_));
 NAND3_X1 _25928_ (.A1(_07389_),
    .A2(_07388_),
    .A3(_05510_),
    .ZN(_07423_));
 AOI21_X1 _25929_ (.A(_07378_),
    .B1(\alu_adder_result_ex[5] ),
    .B2(_07332_),
    .ZN(_07424_));
 OAI21_X1 _25930_ (.A(_07424_),
    .B1(_07421_),
    .B2(_03700_),
    .ZN(_07425_));
 CLKBUF_X3 _25931_ (.A(_05110_),
    .Z(_07426_));
 CLKBUF_X3 _25932_ (.A(_07426_),
    .Z(_07427_));
 NAND2_X1 _25933_ (.A1(_00561_),
    .A2(_07427_),
    .ZN(_07428_));
 OAI21_X1 _25934_ (.A(_07428_),
    .B1(_07410_),
    .B2(\alu_adder_result_ex[5] ),
    .ZN(_07429_));
 OR2_X1 _25935_ (.A1(_07406_),
    .A2(_07429_),
    .ZN(_07430_));
 OAI21_X1 _25936_ (.A(_07430_),
    .B1(_05137_),
    .B2(_07376_),
    .ZN(_07431_));
 AOI21_X1 _25937_ (.A(_07425_),
    .B1(_07431_),
    .B2(_03780_),
    .ZN(_07432_));
 CLKBUF_X3 _25938_ (.A(_07330_),
    .Z(_07433_));
 OAI21_X1 _25939_ (.A(_07433_),
    .B1(_07397_),
    .B2(_12051_),
    .ZN(_07434_));
 INV_X1 _25940_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .ZN(_07435_));
 OAI221_X1 _25941_ (.A(_07423_),
    .B1(_07432_),
    .B2(_07434_),
    .C1(_07415_),
    .C2(_07435_),
    .ZN(_02309_));
 NAND2_X1 _25942_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .A2(_03692_),
    .ZN(_07436_));
 MUX2_X1 _25943_ (.A(\alu_adder_result_ex[3] ),
    .B(_11427_),
    .S(_03925_),
    .Z(_07437_));
 NAND2_X1 _25944_ (.A1(_04179_),
    .A2(_07437_),
    .ZN(_07438_));
 OAI21_X1 _25945_ (.A(_07436_),
    .B1(_07438_),
    .B2(_03692_),
    .ZN(_02310_));
 OR3_X1 _25946_ (.A1(_07385_),
    .A2(_07401_),
    .A3(_05598_),
    .ZN(_07439_));
 AOI21_X1 _25947_ (.A(_07378_),
    .B1(net8),
    .B2(_07332_),
    .ZN(_07440_));
 OAI21_X1 _25948_ (.A(_07440_),
    .B1(_07429_),
    .B2(_03700_),
    .ZN(_07441_));
 NAND2_X1 _25949_ (.A1(_00562_),
    .A2(_07427_),
    .ZN(_07442_));
 OAI21_X1 _25950_ (.A(_07442_),
    .B1(_07410_),
    .B2(net8),
    .ZN(_07443_));
 OR2_X1 _25951_ (.A1(_07406_),
    .A2(_07443_),
    .ZN(_07444_));
 OAI21_X1 _25952_ (.A(_07444_),
    .B1(_05140_),
    .B2(_07376_),
    .ZN(_07445_));
 AOI21_X1 _25953_ (.A(_07441_),
    .B1(_07445_),
    .B2(_03780_),
    .ZN(_07446_));
 OAI21_X1 _25954_ (.A(_07433_),
    .B1(_07397_),
    .B2(_03854_),
    .ZN(_07447_));
 OAI221_X1 _25955_ (.A(_07439_),
    .B1(_07446_),
    .B2(_07447_),
    .C1(_07415_),
    .C2(_05599_),
    .ZN(_02311_));
 NOR2_X1 _25956_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .A2(_07415_),
    .ZN(_07448_));
 AOI21_X1 _25957_ (.A(_07391_),
    .B1(_05688_),
    .B2(_07389_),
    .ZN(_07449_));
 AOI21_X1 _25958_ (.A(_07418_),
    .B1(\alu_adder_result_ex[7] ),
    .B2(_03744_),
    .ZN(_07450_));
 OAI21_X1 _25959_ (.A(_07450_),
    .B1(_07443_),
    .B2(_03700_),
    .ZN(_07451_));
 NOR2_X1 _25960_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_05110_),
    .ZN(_07452_));
 AOI21_X1 _25961_ (.A(_07452_),
    .B1(_07426_),
    .B2(_00563_),
    .ZN(_07453_));
 NAND2_X1 _25962_ (.A1(_07376_),
    .A2(_07453_),
    .ZN(_07454_));
 BUF_X4 _25963_ (.A(_03761_),
    .Z(_07455_));
 OAI21_X1 _25964_ (.A(_07454_),
    .B1(_05143_),
    .B2(_07455_),
    .ZN(_07456_));
 AOI21_X1 _25965_ (.A(_07451_),
    .B1(_07456_),
    .B2(_03781_),
    .ZN(_07457_));
 OAI21_X1 _25966_ (.A(_07396_),
    .B1(_07397_),
    .B2(_03861_),
    .ZN(_07458_));
 OAI22_X1 _25967_ (.A1(_07448_),
    .A2(_07449_),
    .B1(_07457_),
    .B2(_07458_),
    .ZN(_02312_));
 OR3_X1 _25968_ (.A1(_07385_),
    .A2(_07401_),
    .A3(_05755_),
    .ZN(_07459_));
 OAI21_X1 _25969_ (.A(_07396_),
    .B1(_07397_),
    .B2(_03872_),
    .ZN(_07460_));
 AOI221_X1 _25970_ (.A(_07331_),
    .B1(_07453_),
    .B2(_03493_),
    .C1(_03742_),
    .C2(\alu_adder_result_ex[8] ),
    .ZN(_07461_));
 INV_X1 _25971_ (.A(_07461_),
    .ZN(_07462_));
 NOR2_X1 _25972_ (.A1(\alu_adder_result_ex[8] ),
    .A2(_07408_),
    .ZN(_07463_));
 AOI21_X2 _25973_ (.A(_07463_),
    .B1(_07427_),
    .B2(_00564_),
    .ZN(_07464_));
 NOR2_X1 _25974_ (.A1(_07406_),
    .A2(_07464_),
    .ZN(_07465_));
 AOI21_X1 _25975_ (.A(_07465_),
    .B1(_05146_),
    .B2(_07407_),
    .ZN(_07466_));
 AOI21_X1 _25976_ (.A(_07462_),
    .B1(_07466_),
    .B2(_03780_),
    .ZN(_07467_));
 OAI221_X1 _25977_ (.A(_07459_),
    .B1(_07460_),
    .B2(_07467_),
    .C1(_07415_),
    .C2(_05756_),
    .ZN(_02313_));
 OAI21_X1 _25978_ (.A(_07387_),
    .B1(_05785_),
    .B2(_07385_),
    .ZN(_07468_));
 OAI21_X1 _25979_ (.A(_07468_),
    .B1(_07388_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .ZN(_07469_));
 AOI221_X2 _25980_ (.A(_07418_),
    .B1(_07464_),
    .B2(_03784_),
    .C1(_03744_),
    .C2(\alu_adder_result_ex[9] ),
    .ZN(_07470_));
 OAI21_X1 _25981_ (.A(_07433_),
    .B1(_07383_),
    .B2(_03880_),
    .ZN(_07471_));
 MUX2_X1 _25982_ (.A(_00565_),
    .B(_12271_),
    .S(_05033_),
    .Z(_07472_));
 MUX2_X1 _25983_ (.A(_05149_),
    .B(_07472_),
    .S(_07376_),
    .Z(_07473_));
 OAI221_X1 _25984_ (.A(_07469_),
    .B1(_07470_),
    .B2(_07471_),
    .C1(_07473_),
    .C2(_07374_),
    .ZN(_02314_));
 NOR2_X1 _25985_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .A2(_07415_),
    .ZN(_07474_));
 AOI21_X1 _25986_ (.A(_07391_),
    .B1(_05860_),
    .B2(_07389_),
    .ZN(_07475_));
 AOI21_X1 _25987_ (.A(_07418_),
    .B1(\alu_adder_result_ex[10] ),
    .B2(_03743_),
    .ZN(_07476_));
 OAI21_X1 _25988_ (.A(_07476_),
    .B1(_07472_),
    .B2(_03700_),
    .ZN(_07477_));
 NAND2_X1 _25989_ (.A1(_00566_),
    .A2(_07427_),
    .ZN(_07478_));
 OAI21_X1 _25990_ (.A(_07478_),
    .B1(_07410_),
    .B2(\alu_adder_result_ex[10] ),
    .ZN(_07479_));
 OR2_X1 _25991_ (.A1(_07406_),
    .A2(_07479_),
    .ZN(_07480_));
 OAI21_X1 _25992_ (.A(_07480_),
    .B1(_05044_),
    .B2(_07455_),
    .ZN(_07481_));
 AOI21_X1 _25993_ (.A(_07477_),
    .B1(_07481_),
    .B2(_03781_),
    .ZN(_07482_));
 OAI21_X1 _25994_ (.A(_07396_),
    .B1(_07397_),
    .B2(_03889_),
    .ZN(_07483_));
 OAI22_X1 _25995_ (.A1(_07474_),
    .A2(_07475_),
    .B1(_07482_),
    .B2(_07483_),
    .ZN(_02315_));
 NOR2_X1 _25996_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .A2(_07415_),
    .ZN(_07484_));
 AOI21_X1 _25997_ (.A(_07391_),
    .B1(_05893_),
    .B2(_07389_),
    .ZN(_07485_));
 AOI21_X1 _25998_ (.A(_07418_),
    .B1(net486),
    .B2(_03743_),
    .ZN(_07486_));
 OAI21_X1 _25999_ (.A(_07486_),
    .B1(_07479_),
    .B2(_03700_),
    .ZN(_07487_));
 NOR2_X1 _26000_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_07408_),
    .ZN(_07488_));
 AOI21_X2 _26001_ (.A(_07488_),
    .B1(_07410_),
    .B2(_00567_),
    .ZN(_07489_));
 NAND2_X1 _26002_ (.A1(_07376_),
    .A2(_07489_),
    .ZN(_07490_));
 OAI21_X1 _26003_ (.A(_07490_),
    .B1(_05048_),
    .B2(_07455_),
    .ZN(_07491_));
 AOI21_X1 _26004_ (.A(_07487_),
    .B1(_07491_),
    .B2(_03781_),
    .ZN(_07492_));
 OAI21_X1 _26005_ (.A(_07396_),
    .B1(_07397_),
    .B2(_03896_),
    .ZN(_07493_));
 OAI22_X1 _26006_ (.A1(_07484_),
    .A2(_07485_),
    .B1(_07492_),
    .B2(_07493_),
    .ZN(_02316_));
 OAI21_X1 _26007_ (.A(_07387_),
    .B1(_05915_),
    .B2(_03738_),
    .ZN(_07494_));
 OAI21_X1 _26008_ (.A(_07494_),
    .B1(_07388_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .ZN(_07495_));
 AOI221_X2 _26009_ (.A(_07418_),
    .B1(_07489_),
    .B2(_03784_),
    .C1(_03744_),
    .C2(\alu_adder_result_ex[12] ),
    .ZN(_07496_));
 OAI21_X1 _26010_ (.A(_07433_),
    .B1(_07383_),
    .B2(_03905_),
    .ZN(_07497_));
 NOR2_X1 _26011_ (.A1(_07455_),
    .A2(_05052_),
    .ZN(_07498_));
 NOR2_X1 _26012_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_07408_),
    .ZN(_07499_));
 AOI21_X2 _26013_ (.A(_07499_),
    .B1(_07410_),
    .B2(_00568_),
    .ZN(_07500_));
 CLKBUF_X3 _26014_ (.A(_03761_),
    .Z(_07501_));
 AOI21_X1 _26015_ (.A(_07498_),
    .B1(_07500_),
    .B2(_07501_),
    .ZN(_07502_));
 OAI221_X1 _26016_ (.A(_07495_),
    .B1(_07496_),
    .B2(_07497_),
    .C1(_07502_),
    .C2(_07374_),
    .ZN(_02317_));
 MUX2_X1 _26017_ (.A(_04163_),
    .B(_05961_),
    .S(_06144_),
    .Z(_07503_));
 NOR3_X1 _26018_ (.A1(_03738_),
    .A2(_07369_),
    .A3(_07503_),
    .ZN(_07504_));
 AOI21_X1 _26019_ (.A(_07504_),
    .B1(_07391_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .ZN(_07505_));
 AOI221_X2 _26020_ (.A(_07418_),
    .B1(_07500_),
    .B2(_03784_),
    .C1(_03744_),
    .C2(\alu_adder_result_ex[13] ),
    .ZN(_07506_));
 OAI21_X1 _26021_ (.A(_07433_),
    .B1(_07383_),
    .B2(_03914_),
    .ZN(_07507_));
 NOR2_X1 _26022_ (.A1(_07455_),
    .A2(_05055_),
    .ZN(_07508_));
 NOR2_X1 _26023_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_07408_),
    .ZN(_07509_));
 AOI21_X2 _26024_ (.A(_07509_),
    .B1(_07410_),
    .B2(_04163_),
    .ZN(_07510_));
 AOI21_X1 _26025_ (.A(_07508_),
    .B1(_07510_),
    .B2(_07501_),
    .ZN(_07511_));
 OAI221_X1 _26026_ (.A(_07505_),
    .B1(_07506_),
    .B2(_07507_),
    .C1(_07511_),
    .C2(_07374_),
    .ZN(_02318_));
 MUX2_X1 _26027_ (.A(_00630_),
    .B(_05989_),
    .S(_06144_),
    .Z(_07512_));
 NOR3_X1 _26028_ (.A1(_03738_),
    .A2(_07369_),
    .A3(_07512_),
    .ZN(_07513_));
 AOI21_X1 _26029_ (.A(_07513_),
    .B1(_07391_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .ZN(_07514_));
 AOI221_X2 _26030_ (.A(_07418_),
    .B1(_07510_),
    .B2(_03783_),
    .C1(_03744_),
    .C2(net7),
    .ZN(_07515_));
 OAI21_X1 _26031_ (.A(_07433_),
    .B1(_07383_),
    .B2(_03921_),
    .ZN(_07516_));
 NOR2_X1 _26032_ (.A1(_07455_),
    .A2(_05058_),
    .ZN(_07517_));
 NOR2_X1 _26033_ (.A1(net7),
    .A2(_07408_),
    .ZN(_07518_));
 AOI21_X2 _26034_ (.A(_07518_),
    .B1(_07410_),
    .B2(_00630_),
    .ZN(_07519_));
 AOI21_X1 _26035_ (.A(_07517_),
    .B1(_07519_),
    .B2(_07501_),
    .ZN(_07520_));
 OAI221_X1 _26036_ (.A(_07514_),
    .B1(_07515_),
    .B2(_07516_),
    .C1(_07520_),
    .C2(_07374_),
    .ZN(_02319_));
 OR2_X1 _26037_ (.A1(_00661_),
    .A2(_06144_),
    .ZN(_07521_));
 OAI21_X1 _26038_ (.A(_07521_),
    .B1(_06049_),
    .B2(_05884_),
    .ZN(_07522_));
 AOI22_X1 _26039_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .A2(_07391_),
    .B1(_03775_),
    .B2(_07522_),
    .ZN(_07523_));
 AOI221_X2 _26040_ (.A(_07418_),
    .B1(_07519_),
    .B2(_03783_),
    .C1(_03744_),
    .C2(net438),
    .ZN(_07524_));
 OAI21_X1 _26041_ (.A(_07433_),
    .B1(_07383_),
    .B2(_03928_),
    .ZN(_07525_));
 INV_X1 _26042_ (.A(\alu_adder_result_ex[15] ),
    .ZN(_07526_));
 MUX2_X1 _26043_ (.A(_00661_),
    .B(_07526_),
    .S(_05033_),
    .Z(_07527_));
 MUX2_X1 _26044_ (.A(_05061_),
    .B(_07527_),
    .S(_07376_),
    .Z(_07528_));
 OAI221_X1 _26045_ (.A(_07523_),
    .B1(_07524_),
    .B2(_07525_),
    .C1(_07528_),
    .C2(_07373_),
    .ZN(_02320_));
 NAND2_X1 _26046_ (.A1(net330),
    .A2(_03925_),
    .ZN(_07529_));
 OAI21_X1 _26047_ (.A(_07529_),
    .B1(_03925_),
    .B2(_03725_),
    .ZN(_07530_));
 MUX2_X1 _26048_ (.A(_07530_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .S(_03691_),
    .Z(_02321_));
 NAND3_X1 _26049_ (.A1(_07389_),
    .A2(_07388_),
    .A3(_06083_),
    .ZN(_07531_));
 OAI21_X1 _26050_ (.A(_07396_),
    .B1(_07397_),
    .B2(_04344_),
    .ZN(_07532_));
 AOI21_X1 _26051_ (.A(_07378_),
    .B1(\alu_adder_result_ex[16] ),
    .B2(_03743_),
    .ZN(_07533_));
 OAI21_X1 _26052_ (.A(_07533_),
    .B1(_07527_),
    .B2(_03700_),
    .ZN(_07534_));
 NOR2_X1 _26053_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_05110_),
    .ZN(_07535_));
 AOI21_X2 _26054_ (.A(_07535_),
    .B1(_07408_),
    .B2(_03800_),
    .ZN(_07536_));
 NAND2_X1 _26055_ (.A1(_03761_),
    .A2(_07536_),
    .ZN(_07537_));
 OAI21_X1 _26056_ (.A(_07537_),
    .B1(_05066_),
    .B2(_07376_),
    .ZN(_07538_));
 AOI21_X2 _26057_ (.A(_07534_),
    .B1(_07538_),
    .B2(_03780_),
    .ZN(_07539_));
 INV_X1 _26058_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .ZN(_07540_));
 OAI221_X1 _26059_ (.A(_07531_),
    .B1(_07532_),
    .B2(_07539_),
    .C1(_07415_),
    .C2(_07540_),
    .ZN(_02322_));
 AND2_X1 _26060_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A2(_07401_),
    .ZN(_07541_));
 NOR3_X1 _26061_ (.A1(_07385_),
    .A2(_07401_),
    .A3(_06104_),
    .ZN(_07542_));
 OAI21_X1 _26062_ (.A(_07433_),
    .B1(_07383_),
    .B2(_03812_),
    .ZN(_07543_));
 AOI221_X2 _26063_ (.A(_07378_),
    .B1(_07536_),
    .B2(_03783_),
    .C1(_03743_),
    .C2(\alu_adder_result_ex[17] ),
    .ZN(_07544_));
 NOR2_X1 _26064_ (.A1(_07543_),
    .A2(_07544_),
    .ZN(_07545_));
 NOR3_X1 _26065_ (.A1(_07541_),
    .A2(_07542_),
    .A3(_07545_),
    .ZN(_07546_));
 NOR2_X1 _26066_ (.A1(_07501_),
    .A2(_05069_),
    .ZN(_07547_));
 NOR2_X1 _26067_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_07426_),
    .ZN(_07548_));
 AOI21_X2 _26068_ (.A(_07548_),
    .B1(_07408_),
    .B2(_03940_),
    .ZN(_07549_));
 AOI21_X1 _26069_ (.A(_07547_),
    .B1(_07549_),
    .B2(_07501_),
    .ZN(_07550_));
 OAI21_X1 _26070_ (.A(_07546_),
    .B1(_07550_),
    .B2(_07374_),
    .ZN(_02323_));
 AND2_X1 _26071_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A2(_07401_),
    .ZN(_07551_));
 NOR3_X1 _26072_ (.A1(_07385_),
    .A2(_07401_),
    .A3(_06120_),
    .ZN(_07552_));
 OAI21_X1 _26073_ (.A(_07433_),
    .B1(_07383_),
    .B2(_03822_),
    .ZN(_07553_));
 AOI221_X2 _26074_ (.A(_07331_),
    .B1(_07549_),
    .B2(_03783_),
    .C1(_03742_),
    .C2(\alu_adder_result_ex[18] ),
    .ZN(_07554_));
 NOR2_X1 _26075_ (.A1(_07553_),
    .A2(_07554_),
    .ZN(_07555_));
 NOR3_X1 _26076_ (.A1(_07551_),
    .A2(_07552_),
    .A3(_07555_),
    .ZN(_07556_));
 NOR2_X1 _26077_ (.A1(_07501_),
    .A2(_05072_),
    .ZN(_07557_));
 NOR2_X1 _26078_ (.A1(\alu_adder_result_ex[18] ),
    .A2(_05110_),
    .ZN(_07558_));
 AOI21_X2 _26079_ (.A(_07558_),
    .B1(_05110_),
    .B2(_03944_),
    .ZN(_07559_));
 AOI21_X1 _26080_ (.A(_07557_),
    .B1(_07559_),
    .B2(_07501_),
    .ZN(_07560_));
 OAI21_X1 _26081_ (.A(_07556_),
    .B1(_07560_),
    .B2(_07374_),
    .ZN(_02324_));
 OAI21_X1 _26082_ (.A(_07330_),
    .B1(_07366_),
    .B2(_03828_),
    .ZN(_07561_));
 AOI221_X2 _26083_ (.A(_07331_),
    .B1(_07559_),
    .B2(_03493_),
    .C1(_03742_),
    .C2(\alu_adder_result_ex[19] ),
    .ZN(_07562_));
 NOR2_X1 _26084_ (.A1(_07561_),
    .A2(_07562_),
    .ZN(_07563_));
 AOI221_X2 _26085_ (.A(_07563_),
    .B1(_06145_),
    .B2(_03775_),
    .C1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .C2(_07369_),
    .ZN(_07564_));
 NOR2_X1 _26086_ (.A1(_07501_),
    .A2(_05075_),
    .ZN(_07565_));
 NOR2_X1 _26087_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_07426_),
    .ZN(_07566_));
 AOI21_X2 _26088_ (.A(_07566_),
    .B1(_07408_),
    .B2(_03946_),
    .ZN(_07567_));
 AOI21_X1 _26089_ (.A(_07565_),
    .B1(_07567_),
    .B2(_07501_),
    .ZN(_07568_));
 OAI21_X1 _26090_ (.A(_07564_),
    .B1(_07568_),
    .B2(_07374_),
    .ZN(_02325_));
 AOI22_X1 _26091_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_07391_),
    .B1(_03775_),
    .B2(_06167_),
    .ZN(_07569_));
 AOI221_X2 _26092_ (.A(_07378_),
    .B1(_07567_),
    .B2(_03783_),
    .C1(_03743_),
    .C2(\alu_adder_result_ex[20] ),
    .ZN(_07570_));
 INV_X1 _26093_ (.A(_07570_),
    .ZN(_07571_));
 NOR2_X1 _26094_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_07427_),
    .ZN(_07572_));
 AOI21_X2 _26095_ (.A(_07572_),
    .B1(_07410_),
    .B2(_03948_),
    .ZN(_07573_));
 OAI21_X1 _26096_ (.A(_03780_),
    .B1(_07406_),
    .B2(_07573_),
    .ZN(_07574_));
 AOI21_X1 _26097_ (.A(_07574_),
    .B1(_05084_),
    .B2(_04962_),
    .ZN(_07575_));
 OAI221_X1 _26098_ (.A(_07396_),
    .B1(_07571_),
    .B2(_07575_),
    .C1(_07397_),
    .C2(_03836_),
    .ZN(_07576_));
 NAND2_X1 _26099_ (.A1(_07569_),
    .A2(_07576_),
    .ZN(_02326_));
 OR3_X1 _26100_ (.A1(_10924_),
    .A2(_07369_),
    .A3(_06191_),
    .ZN(_07577_));
 NOR2_X2 _26101_ (.A1(_03771_),
    .A2(_07405_),
    .ZN(_07578_));
 NAND2_X2 _26102_ (.A1(_07330_),
    .A2(_07578_),
    .ZN(_07579_));
 OAI221_X1 _26103_ (.A(_07577_),
    .B1(_07579_),
    .B2(_03846_),
    .C1(_07387_),
    .C2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .ZN(_07580_));
 NOR2_X1 _26104_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_05110_),
    .ZN(_07581_));
 AOI21_X2 _26105_ (.A(_07581_),
    .B1(_07426_),
    .B2(_03950_),
    .ZN(_07582_));
 NOR2_X1 _26106_ (.A1(_07407_),
    .A2(_07582_),
    .ZN(_07583_));
 AOI21_X1 _26107_ (.A(_07583_),
    .B1(_05087_),
    .B2(_07407_),
    .ZN(_07584_));
 NAND2_X1 _26108_ (.A1(_03781_),
    .A2(_07584_),
    .ZN(_07585_));
 NAND2_X4 _26109_ (.A1(_03771_),
    .A2(_07330_),
    .ZN(_07586_));
 AOI221_X2 _26110_ (.A(_07586_),
    .B1(\alu_adder_result_ex[21] ),
    .B2(_03743_),
    .C1(_03784_),
    .C2(_07573_),
    .ZN(_07587_));
 AOI21_X1 _26111_ (.A(_07580_),
    .B1(_07585_),
    .B2(_07587_),
    .ZN(_02327_));
 OAI22_X1 _26112_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_07328_),
    .B1(_07579_),
    .B2(_03855_),
    .ZN(_07588_));
 AOI221_X2 _26113_ (.A(_07586_),
    .B1(_07582_),
    .B2(_03783_),
    .C1(_03742_),
    .C2(\alu_adder_result_ex[22] ),
    .ZN(_07589_));
 MUX2_X1 _26114_ (.A(_03953_),
    .B(\alu_adder_result_ex[22] ),
    .S(_05032_),
    .Z(_07590_));
 NOR2_X1 _26115_ (.A1(_07406_),
    .A2(_07590_),
    .ZN(_07591_));
 AOI21_X1 _26116_ (.A(_07591_),
    .B1(_05090_),
    .B2(_07406_),
    .ZN(_07592_));
 NAND2_X1 _26117_ (.A1(_03780_),
    .A2(_07592_),
    .ZN(_07593_));
 AOI221_X1 _26118_ (.A(_07588_),
    .B1(_07589_),
    .B2(_07593_),
    .C1(_06227_),
    .C2(_07387_),
    .ZN(_02328_));
 NOR2_X1 _26119_ (.A1(_07369_),
    .A2(_06251_),
    .ZN(_07594_));
 NOR2_X1 _26120_ (.A1(net356),
    .A2(_05110_),
    .ZN(_07595_));
 AOI21_X2 _26121_ (.A(_07595_),
    .B1(_07426_),
    .B2(_03955_),
    .ZN(_07596_));
 OAI21_X1 _26122_ (.A(_03492_),
    .B1(_07406_),
    .B2(_07596_),
    .ZN(_07597_));
 AOI21_X1 _26123_ (.A(_07597_),
    .B1(_05093_),
    .B2(_04962_),
    .ZN(_07598_));
 AOI221_X2 _26124_ (.A(_07331_),
    .B1(_07590_),
    .B2(_03493_),
    .C1(_03742_),
    .C2(net356),
    .ZN(_07599_));
 AOI21_X1 _26125_ (.A(_07599_),
    .B1(_07578_),
    .B2(_13422_),
    .ZN(_07600_));
 NOR2_X1 _26126_ (.A1(_07598_),
    .A2(_07600_),
    .ZN(_07601_));
 INV_X1 _26127_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .ZN(_07602_));
 AOI221_X2 _26128_ (.A(_07594_),
    .B1(_07601_),
    .B2(_07433_),
    .C1(_07401_),
    .C2(_07602_),
    .ZN(_02329_));
 NOR2_X1 _26129_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_07426_),
    .ZN(_07603_));
 AOI21_X1 _26130_ (.A(_07603_),
    .B1(_07427_),
    .B2(_03957_),
    .ZN(_07604_));
 OAI21_X1 _26131_ (.A(_03780_),
    .B1(_07407_),
    .B2(_07604_),
    .ZN(_07605_));
 AOI21_X1 _26132_ (.A(_07605_),
    .B1(_05097_),
    .B2(_04962_),
    .ZN(_07606_));
 AOI221_X2 _26133_ (.A(_07331_),
    .B1(_07596_),
    .B2(_03493_),
    .C1(_03742_),
    .C2(\alu_adder_result_ex[24] ),
    .ZN(_07607_));
 AOI21_X1 _26134_ (.A(_07607_),
    .B1(_07578_),
    .B2(_13518_),
    .ZN(_07608_));
 OAI21_X1 _26135_ (.A(_07396_),
    .B1(_07606_),
    .B2(_07608_),
    .ZN(_07609_));
 INV_X1 _26136_ (.A(_03775_),
    .ZN(_07610_));
 INV_X1 _26137_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .ZN(_07611_));
 OAI221_X1 _26138_ (.A(_07609_),
    .B1(_06272_),
    .B2(_07610_),
    .C1(_07611_),
    .C2(_07415_),
    .ZN(_02330_));
 AOI221_X1 _26139_ (.A(_07586_),
    .B1(_07604_),
    .B2(_03783_),
    .C1(_03743_),
    .C2(net388),
    .ZN(_07612_));
 INV_X1 _26140_ (.A(_07612_),
    .ZN(_07613_));
 NOR2_X1 _26141_ (.A1(net388),
    .A2(_07427_),
    .ZN(_07614_));
 AOI21_X2 _26142_ (.A(_07614_),
    .B1(_07410_),
    .B2(_03959_),
    .ZN(_07615_));
 NAND2_X1 _26143_ (.A1(_07455_),
    .A2(_07615_),
    .ZN(_07616_));
 OAI21_X1 _26144_ (.A(_07616_),
    .B1(_05100_),
    .B2(_07501_),
    .ZN(_07617_));
 AOI21_X1 _26145_ (.A(_07613_),
    .B1(_07617_),
    .B2(_03781_),
    .ZN(_07618_));
 NAND2_X1 _26146_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(_07369_),
    .ZN(_07619_));
 OAI21_X1 _26147_ (.A(_07619_),
    .B1(_06306_),
    .B2(_07401_),
    .ZN(_07620_));
 OAI21_X1 _26148_ (.A(_07620_),
    .B1(_07579_),
    .B2(_03881_),
    .ZN(_07621_));
 NOR2_X1 _26149_ (.A1(_07618_),
    .A2(_07621_),
    .ZN(_02331_));
 NAND2_X1 _26150_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .A2(_03692_),
    .ZN(_07622_));
 MUX2_X1 _26151_ (.A(\alu_adder_result_ex[5] ),
    .B(_03831_),
    .S(_03925_),
    .Z(_07623_));
 NAND2_X1 _26152_ (.A1(_04179_),
    .A2(_07623_),
    .ZN(_07624_));
 OAI21_X1 _26153_ (.A(_07622_),
    .B1(_07624_),
    .B2(_03692_),
    .ZN(_02332_));
 NAND2_X1 _26154_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A2(_07369_),
    .ZN(_07625_));
 NOR2_X1 _26155_ (.A1(_10924_),
    .A2(_06318_),
    .ZN(_07626_));
 OAI21_X1 _26156_ (.A(_07625_),
    .B1(_07626_),
    .B2(_07401_),
    .ZN(_07627_));
 OAI21_X1 _26157_ (.A(_07627_),
    .B1(_07579_),
    .B2(_13686_),
    .ZN(_07628_));
 MUX2_X1 _26158_ (.A(_03961_),
    .B(\alu_adder_result_ex[26] ),
    .S(_05033_),
    .Z(_07629_));
 NOR2_X1 _26159_ (.A1(_07407_),
    .A2(_07629_),
    .ZN(_07630_));
 AOI21_X1 _26160_ (.A(_07630_),
    .B1(_05103_),
    .B2(_07407_),
    .ZN(_07631_));
 NAND2_X1 _26161_ (.A1(_03781_),
    .A2(_07631_),
    .ZN(_07632_));
 AOI221_X2 _26162_ (.A(_07586_),
    .B1(_07615_),
    .B2(_03784_),
    .C1(_03744_),
    .C2(\alu_adder_result_ex[26] ),
    .ZN(_07633_));
 AOI21_X1 _26163_ (.A(_07628_),
    .B1(_07632_),
    .B2(_07633_),
    .ZN(_02333_));
 OAI22_X1 _26164_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A2(_07328_),
    .B1(_07579_),
    .B2(_03139_),
    .ZN(_07634_));
 NAND2_X1 _26165_ (.A1(_01033_),
    .A2(_07426_),
    .ZN(_07635_));
 OAI21_X1 _26166_ (.A(_07635_),
    .B1(_07426_),
    .B2(\alu_adder_result_ex[27] ),
    .ZN(_07636_));
 MUX2_X1 _26167_ (.A(_05106_),
    .B(_07636_),
    .S(_03761_),
    .Z(_07637_));
 OR2_X1 _26168_ (.A1(_07371_),
    .A2(_07637_),
    .ZN(_07638_));
 AOI221_X2 _26169_ (.A(_07586_),
    .B1(_07629_),
    .B2(_03493_),
    .C1(_03742_),
    .C2(\alu_adder_result_ex[27] ),
    .ZN(_07639_));
 INV_X1 _26170_ (.A(_06351_),
    .ZN(_07640_));
 AOI221_X1 _26171_ (.A(_07634_),
    .B1(_07638_),
    .B2(_07639_),
    .C1(_07387_),
    .C2(_07640_),
    .ZN(_02334_));
 NAND2_X1 _26172_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A2(_07391_),
    .ZN(_07641_));
 NAND3_X1 _26173_ (.A1(_03237_),
    .A2(_07385_),
    .A3(_07578_),
    .ZN(_07642_));
 NAND3_X1 _26174_ (.A1(_07388_),
    .A2(_06379_),
    .A3(_07642_),
    .ZN(_07643_));
 NAND2_X1 _26175_ (.A1(_07407_),
    .A2(_05112_),
    .ZN(_07644_));
 NAND2_X1 _26176_ (.A1(_03967_),
    .A2(_07427_),
    .ZN(_07645_));
 OAI21_X1 _26177_ (.A(_07645_),
    .B1(_07427_),
    .B2(net386),
    .ZN(_07646_));
 NAND2_X1 _26178_ (.A1(_07455_),
    .A2(_07646_),
    .ZN(_07647_));
 NAND3_X1 _26179_ (.A1(_03781_),
    .A2(_07644_),
    .A3(_07647_),
    .ZN(_07648_));
 INV_X1 _26180_ (.A(_07636_),
    .ZN(_07649_));
 AOI221_X2 _26181_ (.A(_07586_),
    .B1(_07649_),
    .B2(_03784_),
    .C1(_03744_),
    .C2(net386),
    .ZN(_07650_));
 AOI22_X1 _26182_ (.A1(_07641_),
    .A2(_07643_),
    .B1(_07648_),
    .B2(_07650_),
    .ZN(_02335_));
 OAI21_X1 _26183_ (.A(_03738_),
    .B1(_07366_),
    .B2(_03915_),
    .ZN(_07651_));
 AOI21_X1 _26184_ (.A(_07331_),
    .B1(net411),
    .B2(_03742_),
    .ZN(_07652_));
 OAI21_X1 _26185_ (.A(_07652_),
    .B1(_07646_),
    .B2(_03699_),
    .ZN(_07653_));
 MUX2_X1 _26186_ (.A(_03969_),
    .B(net411),
    .S(_05033_),
    .Z(_07654_));
 NOR2_X1 _26187_ (.A1(_07405_),
    .A2(_07654_),
    .ZN(_07655_));
 AOI21_X1 _26188_ (.A(_07655_),
    .B1(_05117_),
    .B2(_07406_),
    .ZN(_07656_));
 AOI21_X2 _26189_ (.A(_07653_),
    .B1(_07656_),
    .B2(_03780_),
    .ZN(_07657_));
 OAI22_X1 _26190_ (.A1(_07385_),
    .A2(_06411_),
    .B1(_07651_),
    .B2(_07657_),
    .ZN(_07658_));
 MUX2_X1 _26191_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .B(_07658_),
    .S(_07388_),
    .Z(_02336_));
 AOI221_X2 _26192_ (.A(_07378_),
    .B1(_07654_),
    .B2(_03783_),
    .C1(_03743_),
    .C2(net345),
    .ZN(_07659_));
 NOR2_X1 _26193_ (.A1(_03922_),
    .A2(_07383_),
    .ZN(_07660_));
 NOR2_X1 _26194_ (.A1(_03761_),
    .A2(_05123_),
    .ZN(_07661_));
 NOR2_X1 _26195_ (.A1(net345),
    .A2(_07426_),
    .ZN(_07662_));
 AOI21_X1 _26196_ (.A(_07662_),
    .B1(_07427_),
    .B2(_03971_),
    .ZN(_07663_));
 AOI21_X1 _26197_ (.A(_07661_),
    .B1(_07663_),
    .B2(_07455_),
    .ZN(_07664_));
 OAI221_X2 _26198_ (.A(_07396_),
    .B1(_07659_),
    .B2(_07660_),
    .C1(_07664_),
    .C2(_07371_),
    .ZN(_07665_));
 NOR2_X1 _26199_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(_07387_),
    .ZN(_07666_));
 AOI21_X1 _26200_ (.A(_07666_),
    .B1(_06430_),
    .B2(_07388_),
    .ZN(_07667_));
 AND2_X1 _26201_ (.A1(_07665_),
    .A2(_07667_),
    .ZN(_02337_));
 OAI21_X1 _26202_ (.A(_03738_),
    .B1(_07383_),
    .B2(_03488_),
    .ZN(_07668_));
 AND2_X1 _26203_ (.A1(_03499_),
    .A2(net289),
    .ZN(_07669_));
 NAND2_X1 _26204_ (.A1(_00099_),
    .A2(_04962_),
    .ZN(_07670_));
 OAI221_X2 _26205_ (.A(_03780_),
    .B1(_04962_),
    .B2(_07669_),
    .C1(_07670_),
    .C2(_05126_),
    .ZN(_07671_));
 AOI221_X1 _26206_ (.A(_07378_),
    .B1(_07663_),
    .B2(_03783_),
    .C1(_03743_),
    .C2(net289),
    .ZN(_07672_));
 AOI21_X1 _26207_ (.A(_07668_),
    .B1(_07671_),
    .B2(_07672_),
    .ZN(_07673_));
 OAI21_X1 _26208_ (.A(_07387_),
    .B1(_06466_),
    .B2(_07385_),
    .ZN(_07674_));
 OAI22_X1 _26209_ (.A1(_03499_),
    .A2(_07415_),
    .B1(_07673_),
    .B2(_07674_),
    .ZN(_07675_));
 INV_X1 _26210_ (.A(_07675_),
    .ZN(_02338_));
 OAI21_X1 _26211_ (.A(_06463_),
    .B1(_06428_),
    .B2(_06462_),
    .ZN(_07676_));
 AOI21_X1 _26212_ (.A(_16224_),
    .B1(_07676_),
    .B2(_16225_),
    .ZN(_07677_));
 XNOR2_X1 _26213_ (.A(_16231_),
    .B(_07677_),
    .ZN(_07678_));
 NAND3_X1 _26214_ (.A1(_07389_),
    .A2(_06144_),
    .A3(_07678_),
    .ZN(_07679_));
 AOI22_X4 _26215_ (.A1(_07418_),
    .A2(_07407_),
    .B1(_07669_),
    .B2(_03784_),
    .ZN(_07680_));
 OAI21_X1 _26216_ (.A(_07679_),
    .B1(_07680_),
    .B2(_07389_),
    .ZN(_07681_));
 MUX2_X1 _26217_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B(_07681_),
    .S(_07388_),
    .Z(_02339_));
 NAND2_X1 _26218_ (.A1(_07389_),
    .A2(_06144_),
    .ZN(_07682_));
 XNOR2_X1 _26219_ (.A(_15745_),
    .B(_16134_),
    .ZN(_07683_));
 XNOR2_X1 _26220_ (.A(_15741_),
    .B(_07683_),
    .ZN(_07684_));
 XOR2_X1 _26221_ (.A(_15732_),
    .B(_15702_),
    .Z(_07685_));
 XNOR2_X1 _26222_ (.A(_16227_),
    .B(_15749_),
    .ZN(_07686_));
 XNOR2_X1 _26223_ (.A(_07685_),
    .B(_07686_),
    .ZN(_07687_));
 XNOR2_X1 _26224_ (.A(_15660_),
    .B(_15214_),
    .ZN(_07688_));
 XNOR2_X1 _26225_ (.A(_07687_),
    .B(_07688_),
    .ZN(_07689_));
 XOR2_X1 _26226_ (.A(_15736_),
    .B(_15739_),
    .Z(_07690_));
 XNOR2_X1 _26227_ (.A(_15701_),
    .B(_15728_),
    .ZN(_07691_));
 XNOR2_X1 _26228_ (.A(_07690_),
    .B(_07691_),
    .ZN(_07692_));
 XNOR2_X1 _26229_ (.A(_15752_),
    .B(_15725_),
    .ZN(_07693_));
 XNOR2_X1 _26230_ (.A(_15724_),
    .B(_15619_),
    .ZN(_07694_));
 XNOR2_X1 _26231_ (.A(_07693_),
    .B(_07694_),
    .ZN(_07695_));
 XNOR2_X2 _26232_ (.A(_07692_),
    .B(_07695_),
    .ZN(_07696_));
 XNOR2_X2 _26233_ (.A(_07689_),
    .B(_07696_),
    .ZN(_07697_));
 XNOR2_X2 _26234_ (.A(_07684_),
    .B(_07697_),
    .ZN(_07698_));
 OAI21_X1 _26235_ (.A(_03933_),
    .B1(_03757_),
    .B2(_01163_),
    .ZN(_07699_));
 INV_X1 _26236_ (.A(_07699_),
    .ZN(_07700_));
 NOR3_X1 _26237_ (.A1(_00132_),
    .A2(_03843_),
    .A3(_07700_),
    .ZN(_07701_));
 XNOR2_X1 _26238_ (.A(_07698_),
    .B(_07701_),
    .ZN(_07702_));
 AOI21_X1 _26239_ (.A(_16224_),
    .B1(_06464_),
    .B2(_16225_),
    .ZN(_07703_));
 INV_X1 _26240_ (.A(_07703_),
    .ZN(_07704_));
 AOI21_X1 _26241_ (.A(_16230_),
    .B1(_07704_),
    .B2(_16231_),
    .ZN(_07705_));
 XNOR2_X1 _26242_ (.A(_07702_),
    .B(_07705_),
    .ZN(_07706_));
 OAI22_X1 _26243_ (.A1(_03771_),
    .A2(_07455_),
    .B1(_07682_),
    .B2(_07706_),
    .ZN(_07707_));
 MUX2_X1 _26244_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .B(_07707_),
    .S(_07388_),
    .Z(_02340_));
 MUX2_X1 _26245_ (.A(net8),
    .B(net361),
    .S(_03766_),
    .Z(_07708_));
 MUX2_X1 _26246_ (.A(_07708_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .S(_03691_),
    .Z(_02341_));
 NAND2_X1 _26247_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .A2(_07295_),
    .ZN(_07709_));
 MUX2_X1 _26248_ (.A(\alu_adder_result_ex[7] ),
    .B(_03849_),
    .S(_03925_),
    .Z(_07710_));
 NAND2_X1 _26249_ (.A1(_04179_),
    .A2(_07710_),
    .ZN(_07711_));
 OAI21_X1 _26250_ (.A(_07709_),
    .B1(_07711_),
    .B2(_03692_),
    .ZN(_02342_));
 MUX2_X1 _26251_ (.A(\alu_adder_result_ex[8] ),
    .B(_11648_),
    .S(_03766_),
    .Z(_07712_));
 MUX2_X1 _26252_ (.A(_07712_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .S(_03691_),
    .Z(_02343_));
 MUX2_X1 _26253_ (.A(\alu_adder_result_ex[9] ),
    .B(_03867_),
    .S(_03766_),
    .Z(_07713_));
 MUX2_X1 _26254_ (.A(_07713_),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .S(_03691_),
    .Z(_02344_));
 NAND2_X1 _26255_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .A2(_04100_),
    .ZN(_07714_));
 NAND2_X4 _26256_ (.A1(_04034_),
    .A2(_04040_),
    .ZN(_07715_));
 OAI21_X1 _26257_ (.A(_04078_),
    .B1(_07715_),
    .B2(net1),
    .ZN(_07716_));
 AOI221_X2 _26258_ (.A(_04042_),
    .B1(_04066_),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .C1(_04068_),
    .C2(\cs_registers_i.csr_mepc_o[10] ),
    .ZN(_07717_));
 INV_X1 _26259_ (.A(_04034_),
    .ZN(_07718_));
 OAI33_X1 _26260_ (.A1(_04013_),
    .A2(_04000_),
    .A3(_03649_),
    .B1(_04086_),
    .B2(_07718_),
    .B3(_04040_),
    .ZN(_07719_));
 NAND2_X4 _26261_ (.A1(_03531_),
    .A2(_07719_),
    .ZN(_07720_));
 OAI21_X1 _26262_ (.A(_07717_),
    .B1(_07720_),
    .B2(_01171_),
    .ZN(_07721_));
 AOI21_X2 _26263_ (.A(_07721_),
    .B1(_04083_),
    .B2(\alu_adder_result_ex[10] ),
    .ZN(_07722_));
 OAI21_X2 _26264_ (.A(_07714_),
    .B1(_07716_),
    .B2(_07722_),
    .ZN(_07723_));
 BUF_X4 _26265_ (.A(_04042_),
    .Z(_07724_));
 NOR2_X1 _26266_ (.A1(_03990_),
    .A2(_04061_),
    .ZN(_07725_));
 NAND2_X1 _26267_ (.A1(net125),
    .A2(\cs_registers_i.mie_q[15] ),
    .ZN(_07726_));
 OAI21_X1 _26268_ (.A(_07725_),
    .B1(_07726_),
    .B2(_03985_),
    .ZN(_07727_));
 NAND2_X1 _26269_ (.A1(_03995_),
    .A2(_07727_),
    .ZN(_07728_));
 OAI21_X1 _26270_ (.A(_07728_),
    .B1(_07284_),
    .B2(_01167_),
    .ZN(_07729_));
 AOI221_X1 _26271_ (.A(_07729_),
    .B1(\alu_adder_result_ex[5] ),
    .B2(_03652_),
    .C1(\cs_registers_i.csr_mepc_o[5] ),
    .C2(_07288_),
    .ZN(_07730_));
 OR3_X1 _26272_ (.A1(_04032_),
    .A2(_07724_),
    .A3(_07730_),
    .ZN(_07731_));
 INV_X1 _26273_ (.A(_07731_),
    .ZN(_07732_));
 AOI21_X2 _26274_ (.A(_07732_),
    .B1(_04100_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .ZN(_07733_));
 NAND2_X1 _26275_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .A2(_04100_),
    .ZN(_07734_));
 NAND2_X1 _26276_ (.A1(_03981_),
    .A2(_03982_),
    .ZN(_07735_));
 NAND3_X1 _26277_ (.A1(_07735_),
    .A2(_03986_),
    .A3(_03987_),
    .ZN(_07736_));
 NAND4_X1 _26278_ (.A1(_03988_),
    .A2(_03989_),
    .A3(_04089_),
    .A4(_07736_),
    .ZN(_07737_));
 AOI21_X1 _26279_ (.A(_07737_),
    .B1(_03993_),
    .B2(_03991_),
    .ZN(_07738_));
 OR2_X1 _26280_ (.A1(_04044_),
    .A2(_07738_),
    .ZN(_07739_));
 OAI21_X1 _26281_ (.A(_07739_),
    .B1(_07284_),
    .B2(_01166_),
    .ZN(_07740_));
 AOI21_X2 _26282_ (.A(_07740_),
    .B1(_04070_),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .ZN(_07741_));
 OAI21_X1 _26283_ (.A(_07741_),
    .B1(_03725_),
    .B2(_04073_),
    .ZN(_07742_));
 NAND2_X2 _26284_ (.A1(_04043_),
    .A2(_07742_),
    .ZN(_07743_));
 AOI21_X2 _26285_ (.A(_07733_),
    .B1(_07734_),
    .B2(_07743_),
    .ZN(_07744_));
 NOR2_X1 _26286_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .A2(_04078_),
    .ZN(_07745_));
 OAI21_X1 _26287_ (.A(_03995_),
    .B1(_04061_),
    .B2(_04088_),
    .ZN(_07746_));
 OAI21_X2 _26288_ (.A(_07746_),
    .B1(_07284_),
    .B2(_01168_),
    .ZN(_07747_));
 AOI221_X2 _26289_ (.A(_07747_),
    .B1(_04083_),
    .B2(\alu_adder_result_ex[6] ),
    .C1(\cs_registers_i.csr_mepc_o[6] ),
    .C2(_07288_),
    .ZN(_07748_));
 AOI21_X2 _26290_ (.A(_07745_),
    .B1(_07748_),
    .B2(_04078_),
    .ZN(_07749_));
 NAND2_X1 _26291_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_04083_),
    .ZN(_07750_));
 NOR2_X4 _26292_ (.A1(_03669_),
    .A2(_07287_),
    .ZN(_07751_));
 AOI22_X2 _26293_ (.A1(\cs_registers_i.csr_mepc_o[7] ),
    .A2(_07288_),
    .B1(_07751_),
    .B2(\cs_registers_i.csr_depc_o[7] ),
    .ZN(_07752_));
 AND3_X1 _26294_ (.A1(_04043_),
    .A2(_07750_),
    .A3(_07752_),
    .ZN(_07753_));
 INV_X1 _26295_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .ZN(_07754_));
 AOI21_X2 _26296_ (.A(_07753_),
    .B1(_04100_),
    .B2(_07754_),
    .ZN(_07755_));
 AND2_X1 _26297_ (.A1(_07749_),
    .A2(_07755_),
    .ZN(_07756_));
 AND3_X1 _26298_ (.A1(_16513_),
    .A2(_07744_),
    .A3(_07756_),
    .ZN(_07757_));
 NOR2_X1 _26299_ (.A1(net32),
    .A2(_07715_),
    .ZN(_07758_));
 AOI22_X1 _26300_ (.A1(\cs_registers_i.csr_mepc_o[9] ),
    .A2(_07288_),
    .B1(_07751_),
    .B2(\cs_registers_i.csr_depc_o[9] ),
    .ZN(_07759_));
 INV_X1 _26301_ (.A(_01170_),
    .ZN(_07760_));
 NAND3_X1 _26302_ (.A1(_03531_),
    .A2(_07760_),
    .A3(_07719_),
    .ZN(_07761_));
 NAND2_X1 _26303_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_03652_),
    .ZN(_07762_));
 AND4_X1 _26304_ (.A1(_07715_),
    .A2(_07759_),
    .A3(_07761_),
    .A4(_07762_),
    .ZN(_07763_));
 NOR3_X2 _26305_ (.A1(_04032_),
    .A2(_07758_),
    .A3(_07763_),
    .ZN(_07764_));
 AOI21_X2 _26306_ (.A(_07764_),
    .B1(_04032_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .ZN(_07765_));
 NAND2_X1 _26307_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .A2(_04100_),
    .ZN(_07766_));
 NOR4_X4 _26308_ (.A1(_12275_),
    .A2(_12282_),
    .A3(_12285_),
    .A4(_04010_),
    .ZN(_07767_));
 AOI221_X2 _26309_ (.A(_04042_),
    .B1(_04066_),
    .B2(\cs_registers_i.csr_depc_o[8] ),
    .C1(_04068_),
    .C2(\cs_registers_i.csr_mepc_o[8] ),
    .ZN(_07768_));
 OAI21_X2 _26310_ (.A(_07768_),
    .B1(_07720_),
    .B2(_01169_),
    .ZN(_07769_));
 OAI221_X2 _26311_ (.A(_04078_),
    .B1(_07767_),
    .B2(_07769_),
    .C1(_07715_),
    .C2(net31),
    .ZN(_07770_));
 AOI21_X1 _26312_ (.A(_07765_),
    .B1(_07766_),
    .B2(_07770_),
    .ZN(_07771_));
 NAND2_X1 _26313_ (.A1(_07757_),
    .A2(_07771_),
    .ZN(_07772_));
 XNOR2_X1 _26314_ (.A(_07723_),
    .B(_07772_),
    .ZN(_07773_));
 NAND2_X4 _26315_ (.A1(_04304_),
    .A2(_04313_),
    .ZN(_07774_));
 BUF_X4 _26316_ (.A(_07774_),
    .Z(_07775_));
 MUX2_X1 _26317_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .B(_07773_),
    .S(_07775_),
    .Z(_02345_));
 NOR2_X1 _26318_ (.A1(net2),
    .A2(_07715_),
    .ZN(_07776_));
 NOR2_X4 _26319_ (.A1(_07718_),
    .A2(_04040_),
    .ZN(_07777_));
 NAND3_X1 _26320_ (.A1(_00551_),
    .A2(_04085_),
    .A3(_04084_),
    .ZN(_07778_));
 NAND2_X1 _26321_ (.A1(_03536_),
    .A2(_04015_),
    .ZN(_07779_));
 NAND3_X1 _26322_ (.A1(_04495_),
    .A2(_07285_),
    .A3(_07779_),
    .ZN(_07780_));
 NAND3_X1 _26323_ (.A1(_07777_),
    .A2(_07778_),
    .A3(_07780_),
    .ZN(_07781_));
 AOI22_X1 _26324_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_07288_),
    .B1(_07751_),
    .B2(\cs_registers_i.csr_depc_o[11] ),
    .ZN(_07782_));
 NAND2_X1 _26325_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_03652_),
    .ZN(_07783_));
 AND4_X1 _26326_ (.A1(_07715_),
    .A2(_07781_),
    .A3(_07782_),
    .A4(_07783_),
    .ZN(_07784_));
 OR3_X1 _26327_ (.A1(_04032_),
    .A2(_07776_),
    .A3(_07784_),
    .ZN(_07785_));
 INV_X1 _26328_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .ZN(_07786_));
 OAI21_X1 _26329_ (.A(_07785_),
    .B1(_04078_),
    .B2(_07786_),
    .ZN(_07787_));
 AND3_X2 _26330_ (.A1(_16511_),
    .A2(_16512_),
    .A3(_07744_),
    .ZN(_07788_));
 AND4_X1 _26331_ (.A1(_07723_),
    .A2(_07756_),
    .A3(_07771_),
    .A4(_07788_),
    .ZN(_07789_));
 XOR2_X1 _26332_ (.A(_07787_),
    .B(_07789_),
    .Z(_07790_));
 MUX2_X1 _26333_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .B(_07790_),
    .S(_07775_),
    .Z(_02346_));
 NOR2_X1 _26334_ (.A1(_04081_),
    .A2(_16509_),
    .ZN(_07791_));
 AOI221_X2 _26335_ (.A(_04042_),
    .B1(_04066_),
    .B2(\cs_registers_i.csr_depc_o[12] ),
    .C1(_04068_),
    .C2(\cs_registers_i.csr_mepc_o[12] ),
    .ZN(_07792_));
 OAI21_X1 _26336_ (.A(_07792_),
    .B1(_07720_),
    .B2(_00550_),
    .ZN(_07793_));
 AOI21_X2 _26337_ (.A(_07793_),
    .B1(_04083_),
    .B2(\alu_adder_result_ex[12] ),
    .ZN(_07794_));
 OAI21_X2 _26338_ (.A(_04078_),
    .B1(_07715_),
    .B2(net3),
    .ZN(_07795_));
 NOR2_X1 _26339_ (.A1(_07794_),
    .A2(_07795_),
    .ZN(_07796_));
 AND3_X1 _26340_ (.A1(_07723_),
    .A2(_07771_),
    .A3(_07787_),
    .ZN(_07797_));
 AND2_X1 _26341_ (.A1(_07757_),
    .A2(_07797_),
    .ZN(_07798_));
 NOR2_X1 _26342_ (.A1(_07796_),
    .A2(_07798_),
    .ZN(_07799_));
 NAND2_X1 _26343_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .A2(_04032_),
    .ZN(_07800_));
 OAI21_X2 _26344_ (.A(_07800_),
    .B1(_07795_),
    .B2(_07794_),
    .ZN(_07801_));
 AOI22_X1 _26345_ (.A1(_04081_),
    .A2(_07799_),
    .B1(_07801_),
    .B2(_07798_),
    .ZN(_07802_));
 NOR2_X1 _26346_ (.A1(_07791_),
    .A2(_07799_),
    .ZN(_07803_));
 OAI22_X1 _26347_ (.A1(_07791_),
    .A2(_07802_),
    .B1(_07803_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .ZN(_07804_));
 INV_X1 _26348_ (.A(_07804_),
    .ZN(_02347_));
 AOI22_X1 _26349_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_04066_),
    .B1(_04068_),
    .B2(\cs_registers_i.csr_mepc_o[13] ),
    .ZN(_07805_));
 INV_X1 _26350_ (.A(_07805_),
    .ZN(_07806_));
 AOI221_X1 _26351_ (.A(_07806_),
    .B1(_03652_),
    .B2(\alu_adder_result_ex[13] ),
    .C1(net4),
    .C2(_04042_),
    .ZN(_07807_));
 OAI21_X1 _26352_ (.A(_07807_),
    .B1(_07720_),
    .B2(_01172_),
    .ZN(_07808_));
 NOR2_X2 _26353_ (.A1(_04032_),
    .A2(_07808_),
    .ZN(_07809_));
 INV_X1 _26354_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .ZN(_07810_));
 AOI21_X2 _26355_ (.A(_07809_),
    .B1(_04100_),
    .B2(_07810_),
    .ZN(_07811_));
 NAND4_X1 _26356_ (.A1(_07756_),
    .A2(_07788_),
    .A3(_07797_),
    .A4(_07801_),
    .ZN(_07812_));
 XNOR2_X1 _26357_ (.A(_07811_),
    .B(_07812_),
    .ZN(_07813_));
 MUX2_X1 _26358_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .B(_07813_),
    .S(_07775_),
    .Z(_02348_));
 AND2_X1 _26359_ (.A1(\alu_adder_result_ex[14] ),
    .A2(_04083_),
    .ZN(_07814_));
 AOI221_X2 _26360_ (.A(_04042_),
    .B1(_07288_),
    .B2(\cs_registers_i.csr_mepc_o[14] ),
    .C1(_07751_),
    .C2(\cs_registers_i.csr_depc_o[14] ),
    .ZN(_07815_));
 OAI21_X1 _26361_ (.A(_07815_),
    .B1(_07720_),
    .B2(_01173_),
    .ZN(_07816_));
 BUF_X4 _26362_ (.A(_07715_),
    .Z(_07817_));
 OAI221_X2 _26363_ (.A(_04078_),
    .B1(_07814_),
    .B2(_07816_),
    .C1(_07817_),
    .C2(net5),
    .ZN(_07818_));
 INV_X1 _26364_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .ZN(_07819_));
 OAI21_X2 _26365_ (.A(_07818_),
    .B1(_04079_),
    .B2(_07819_),
    .ZN(_07820_));
 AND4_X1 _26366_ (.A1(_07749_),
    .A2(_07755_),
    .A3(_07801_),
    .A4(_07811_),
    .ZN(_07821_));
 NAND4_X1 _26367_ (.A1(_16513_),
    .A2(_07744_),
    .A3(_07797_),
    .A4(_07821_),
    .ZN(_07822_));
 XNOR2_X1 _26368_ (.A(_07820_),
    .B(_07822_),
    .ZN(_07823_));
 MUX2_X1 _26369_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .B(_07823_),
    .S(_07775_),
    .Z(_02349_));
 INV_X1 _26370_ (.A(\cs_registers_i.csr_depc_o[15] ),
    .ZN(_07824_));
 NOR3_X1 _26371_ (.A1(_07824_),
    .A2(_03669_),
    .A3(_07287_),
    .ZN(_07825_));
 AOI221_X2 _26372_ (.A(_07825_),
    .B1(_04042_),
    .B2(net6),
    .C1(\cs_registers_i.csr_mepc_o[15] ),
    .C2(_07288_),
    .ZN(_07826_));
 CLKBUF_X3 _26373_ (.A(_07720_),
    .Z(_07827_));
 OAI221_X2 _26374_ (.A(_07826_),
    .B1(_04073_),
    .B2(_07526_),
    .C1(_01174_),
    .C2(_07827_),
    .ZN(_07828_));
 NAND2_X1 _26375_ (.A1(_04079_),
    .A2(_07828_),
    .ZN(_07829_));
 INV_X1 _26376_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .ZN(_07830_));
 OAI21_X2 _26377_ (.A(_07829_),
    .B1(_04079_),
    .B2(_07830_),
    .ZN(_07831_));
 NAND4_X1 _26378_ (.A1(_07788_),
    .A2(_07797_),
    .A3(_07820_),
    .A4(_07821_),
    .ZN(_07832_));
 XNOR2_X1 _26379_ (.A(_07831_),
    .B(_07832_),
    .ZN(_07833_));
 MUX2_X1 _26380_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .B(_07833_),
    .S(_07775_),
    .Z(_02350_));
 NAND3_X1 _26381_ (.A1(_04085_),
    .A2(_01175_),
    .A3(_04084_),
    .ZN(_07834_));
 BUF_X4 _26382_ (.A(_07779_),
    .Z(_07835_));
 NAND3_X1 _26383_ (.A1(_04646_),
    .A2(_07285_),
    .A3(_07835_),
    .ZN(_07836_));
 NAND3_X1 _26384_ (.A1(_07777_),
    .A2(_07834_),
    .A3(_07836_),
    .ZN(_07837_));
 AOI22_X2 _26385_ (.A1(\cs_registers_i.csr_mepc_o[16] ),
    .A2(_07289_),
    .B1(_07751_),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .ZN(_07838_));
 NAND3_X1 _26386_ (.A1(_07817_),
    .A2(_07837_),
    .A3(_07838_),
    .ZN(_07839_));
 AOI21_X2 _26387_ (.A(_04073_),
    .B1(_12896_),
    .B2(_12889_),
    .ZN(_07840_));
 OAI221_X2 _26388_ (.A(_04079_),
    .B1(_07840_),
    .B2(_07839_),
    .C1(_07817_),
    .C2(net15),
    .ZN(_07841_));
 NAND2_X1 _26389_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .A2(_04303_),
    .ZN(_07842_));
 AND2_X1 _26390_ (.A1(_07841_),
    .A2(_07842_),
    .ZN(_07843_));
 NAND2_X1 _26391_ (.A1(_16513_),
    .A2(_07744_),
    .ZN(_07844_));
 NAND4_X1 _26392_ (.A1(_07797_),
    .A2(_07820_),
    .A3(_07821_),
    .A4(_07831_),
    .ZN(_07845_));
 NOR2_X1 _26393_ (.A1(_07844_),
    .A2(_07845_),
    .ZN(_07846_));
 XNOR2_X1 _26394_ (.A(_07843_),
    .B(_07846_),
    .ZN(_07847_));
 MUX2_X1 _26395_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .B(_07847_),
    .S(_07775_),
    .Z(_02351_));
 NOR2_X1 _26396_ (.A1(_12881_),
    .A2(_04073_),
    .ZN(_07848_));
 AOI221_X2 _26397_ (.A(_07724_),
    .B1(_04066_),
    .B2(\cs_registers_i.csr_depc_o[17] ),
    .C1(_04069_),
    .C2(\cs_registers_i.csr_mepc_o[17] ),
    .ZN(_07849_));
 OAI21_X1 _26398_ (.A(_07849_),
    .B1(_07827_),
    .B2(_01176_),
    .ZN(_07850_));
 OAI221_X2 _26399_ (.A(_04079_),
    .B1(_07848_),
    .B2(_07850_),
    .C1(_07817_),
    .C2(net16),
    .ZN(_07851_));
 NAND2_X1 _26400_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .A2(_04303_),
    .ZN(_07852_));
 NAND2_X1 _26401_ (.A1(_07851_),
    .A2(_07852_),
    .ZN(_07853_));
 NAND2_X1 _26402_ (.A1(_07841_),
    .A2(_07842_),
    .ZN(_07854_));
 AND4_X1 _26403_ (.A1(_07797_),
    .A2(_07820_),
    .A3(_07821_),
    .A4(_07831_),
    .ZN(_07855_));
 NAND3_X1 _26404_ (.A1(_07788_),
    .A2(_07854_),
    .A3(_07855_),
    .ZN(_07856_));
 XNOR2_X1 _26405_ (.A(_07853_),
    .B(_07856_),
    .ZN(_07857_));
 MUX2_X1 _26406_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .B(_07857_),
    .S(_07775_),
    .Z(_02352_));
 BUF_X4 _26407_ (.A(_04304_),
    .Z(_07858_));
 AND2_X1 _26408_ (.A1(_07851_),
    .A2(_07852_),
    .ZN(_07859_));
 OR4_X2 _26409_ (.A1(_07844_),
    .A2(_07843_),
    .A3(_07845_),
    .A4(_07859_),
    .ZN(_07860_));
 INV_X1 _26410_ (.A(_07860_),
    .ZN(_07861_));
 NAND3_X1 _26411_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .A2(_16509_),
    .A3(_07861_),
    .ZN(_07862_));
 OAI21_X1 _26412_ (.A(_07862_),
    .B1(_16509_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .ZN(_07863_));
 NAND2_X1 _26413_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .A2(_04303_),
    .ZN(_07864_));
 NOR4_X4 _26414_ (.A1(_13065_),
    .A2(_13067_),
    .A3(_13070_),
    .A4(_04073_),
    .ZN(_07865_));
 AOI221_X2 _26415_ (.A(_07724_),
    .B1(_04066_),
    .B2(\cs_registers_i.csr_depc_o[18] ),
    .C1(_04069_),
    .C2(\cs_registers_i.csr_mepc_o[18] ),
    .ZN(_07866_));
 OAI21_X1 _26416_ (.A(_07866_),
    .B1(_07827_),
    .B2(_01177_),
    .ZN(_07867_));
 BUF_X4 _26417_ (.A(_07817_),
    .Z(_07868_));
 OAI221_X2 _26418_ (.A(_04079_),
    .B1(_07865_),
    .B2(_07867_),
    .C1(_07868_),
    .C2(net17),
    .ZN(_07869_));
 XNOR2_X1 _26419_ (.A(_07860_),
    .B(_07869_),
    .ZN(_07870_));
 AOI22_X1 _26420_ (.A1(_07858_),
    .A2(_07863_),
    .B1(_07864_),
    .B2(_07870_),
    .ZN(_02353_));
 AOI22_X2 _26421_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_04067_),
    .B1(_04069_),
    .B2(\cs_registers_i.csr_mepc_o[19] ),
    .ZN(_07871_));
 INV_X1 _26422_ (.A(net18),
    .ZN(_07872_));
 OAI221_X2 _26423_ (.A(_07871_),
    .B1(_07817_),
    .B2(_07872_),
    .C1(_01178_),
    .C2(_07827_),
    .ZN(_07873_));
 AOI21_X1 _26424_ (.A(_07873_),
    .B1(_07234_),
    .B2(\alu_adder_result_ex[19] ),
    .ZN(_07874_));
 OR2_X2 _26425_ (.A1(_04303_),
    .A2(_07874_),
    .ZN(_07875_));
 INV_X1 _26426_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .ZN(_07876_));
 OAI21_X1 _26427_ (.A(_07875_),
    .B1(_04080_),
    .B2(_07876_),
    .ZN(_07877_));
 NAND2_X2 _26428_ (.A1(_07864_),
    .A2(_07869_),
    .ZN(_07878_));
 AND4_X1 _26429_ (.A1(_07788_),
    .A2(_07854_),
    .A3(_07855_),
    .A4(_07853_),
    .ZN(_07879_));
 NAND2_X1 _26430_ (.A1(_07878_),
    .A2(_07879_),
    .ZN(_07880_));
 XNOR2_X1 _26431_ (.A(_07877_),
    .B(_07880_),
    .ZN(_07881_));
 MUX2_X1 _26432_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .B(_07881_),
    .S(_07775_),
    .Z(_02354_));
 NAND3_X1 _26433_ (.A1(_04085_),
    .A2(_01179_),
    .A3(_04084_),
    .ZN(_07882_));
 NAND3_X1 _26434_ (.A1(_04722_),
    .A2(_07285_),
    .A3(_07835_),
    .ZN(_07883_));
 NAND3_X1 _26435_ (.A1(_07777_),
    .A2(_07882_),
    .A3(_07883_),
    .ZN(_07884_));
 AOI221_X2 _26436_ (.A(_07724_),
    .B1(_04067_),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .C1(_04070_),
    .C2(\cs_registers_i.csr_mepc_o[20] ),
    .ZN(_07885_));
 AND2_X1 _26437_ (.A1(_07884_),
    .A2(_07885_),
    .ZN(_07886_));
 OAI21_X2 _26438_ (.A(_07886_),
    .B1(_04073_),
    .B2(_13266_),
    .ZN(_07887_));
 INV_X1 _26439_ (.A(net19),
    .ZN(_07888_));
 AOI21_X4 _26440_ (.A(_04303_),
    .B1(_07724_),
    .B2(_07888_),
    .ZN(_07889_));
 AOI22_X4 _26441_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .A2(_04303_),
    .B1(_07887_),
    .B2(_07889_),
    .ZN(_07890_));
 NAND2_X1 _26442_ (.A1(_07878_),
    .A2(_07877_),
    .ZN(_07891_));
 NOR2_X1 _26443_ (.A1(_07860_),
    .A2(_07891_),
    .ZN(_07892_));
 XNOR2_X1 _26444_ (.A(_07890_),
    .B(_07892_),
    .ZN(_07893_));
 MUX2_X1 _26445_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .B(_07893_),
    .S(_07775_),
    .Z(_02355_));
 NOR2_X1 _26446_ (.A1(net20),
    .A2(_07817_),
    .ZN(_07894_));
 AOI22_X1 _26447_ (.A1(\cs_registers_i.csr_mepc_o[21] ),
    .A2(_07289_),
    .B1(_07751_),
    .B2(\cs_registers_i.csr_depc_o[21] ),
    .ZN(_07895_));
 OAI21_X1 _26448_ (.A(_07895_),
    .B1(_07720_),
    .B2(_01180_),
    .ZN(_07896_));
 AOI21_X1 _26449_ (.A(_07896_),
    .B1(_07234_),
    .B2(\alu_adder_result_ex[21] ),
    .ZN(_07897_));
 AOI21_X1 _26450_ (.A(_07894_),
    .B1(_07897_),
    .B2(_07817_),
    .ZN(_07898_));
 NAND2_X2 _26451_ (.A1(_04079_),
    .A2(_07898_),
    .ZN(_07899_));
 INV_X1 _26452_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .ZN(_07900_));
 OAI21_X2 _26453_ (.A(_07899_),
    .B1(_04080_),
    .B2(_07900_),
    .ZN(_07901_));
 NOR2_X2 _26454_ (.A1(_07890_),
    .A2(_07891_),
    .ZN(_07902_));
 NAND2_X2 _26455_ (.A1(_07879_),
    .A2(_07902_),
    .ZN(_07903_));
 XNOR2_X1 _26456_ (.A(_07901_),
    .B(_07903_),
    .ZN(_07904_));
 MUX2_X1 _26457_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .B(_07904_),
    .S(_07775_),
    .Z(_02356_));
 NAND2_X1 _26458_ (.A1(net21),
    .A2(_04370_),
    .ZN(_07905_));
 AOI22_X1 _26459_ (.A1(\cs_registers_i.csr_mepc_o[22] ),
    .A2(_07289_),
    .B1(_07751_),
    .B2(\cs_registers_i.csr_depc_o[22] ),
    .ZN(_07906_));
 OAI21_X1 _26460_ (.A(_07906_),
    .B1(_07827_),
    .B2(_01181_),
    .ZN(_07907_));
 NOR3_X1 _26461_ (.A1(_13441_),
    .A2(_13443_),
    .A3(_04073_),
    .ZN(_07908_));
 OAI21_X1 _26462_ (.A(_04043_),
    .B1(_07907_),
    .B2(_07908_),
    .ZN(_07909_));
 NAND2_X1 _26463_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .A2(_04303_),
    .ZN(_07910_));
 NAND3_X2 _26464_ (.A1(_07905_),
    .A2(_07909_),
    .A3(_07910_),
    .ZN(_07911_));
 NAND3_X1 _26465_ (.A1(_07861_),
    .A2(_07902_),
    .A3(_07901_),
    .ZN(_07912_));
 XNOR2_X1 _26466_ (.A(_07911_),
    .B(_07912_),
    .ZN(_07913_));
 BUF_X4 _26467_ (.A(_07774_),
    .Z(_07914_));
 MUX2_X1 _26468_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .B(_07913_),
    .S(_07914_),
    .Z(_02357_));
 AND2_X2 _26469_ (.A1(_04083_),
    .A2(\alu_adder_result_ex[23] ),
    .ZN(_07915_));
 AOI221_X2 _26470_ (.A(_07724_),
    .B1(_04066_),
    .B2(\cs_registers_i.csr_depc_o[23] ),
    .C1(_04069_),
    .C2(\cs_registers_i.csr_mepc_o[23] ),
    .ZN(_07916_));
 OAI21_X1 _26471_ (.A(_07916_),
    .B1(_07827_),
    .B2(_01182_),
    .ZN(_07917_));
 OAI221_X2 _26472_ (.A(_04079_),
    .B1(_07917_),
    .B2(_07915_),
    .C1(_07868_),
    .C2(net22),
    .ZN(_07918_));
 INV_X1 _26473_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .ZN(_07919_));
 OAI21_X4 _26474_ (.A(_07918_),
    .B1(_04080_),
    .B2(_07919_),
    .ZN(_07920_));
 NAND4_X1 _26475_ (.A1(_07879_),
    .A2(_07902_),
    .A3(_07901_),
    .A4(_07911_),
    .ZN(_07921_));
 XNOR2_X1 _26476_ (.A(_07920_),
    .B(_07921_),
    .ZN(_07922_));
 MUX2_X1 _26477_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .B(_07922_),
    .S(_07914_),
    .Z(_02358_));
 OR2_X1 _26478_ (.A1(_07890_),
    .A2(_07891_),
    .ZN(_07923_));
 NAND3_X1 _26479_ (.A1(_07901_),
    .A2(_07911_),
    .A3(_07920_),
    .ZN(_07924_));
 NOR3_X1 _26480_ (.A1(_07860_),
    .A2(_07923_),
    .A3(_07924_),
    .ZN(_07925_));
 NAND3_X1 _26481_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .A2(_16509_),
    .A3(_07925_),
    .ZN(_07926_));
 OAI21_X1 _26482_ (.A(_07926_),
    .B1(_16509_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .ZN(_07927_));
 NAND2_X1 _26483_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .A2(_04303_),
    .ZN(_07928_));
 AOI221_X2 _26484_ (.A(_07724_),
    .B1(_04067_),
    .B2(\cs_registers_i.csr_depc_o[24] ),
    .C1(_04069_),
    .C2(\cs_registers_i.csr_mepc_o[24] ),
    .ZN(_07929_));
 OAI21_X1 _26485_ (.A(_07929_),
    .B1(_07827_),
    .B2(_01183_),
    .ZN(_07930_));
 AOI21_X1 _26486_ (.A(_07930_),
    .B1(_07234_),
    .B2(\alu_adder_result_ex[24] ),
    .ZN(_07931_));
 OAI21_X1 _26487_ (.A(_04080_),
    .B1(_07868_),
    .B2(net23),
    .ZN(_07932_));
 OR2_X1 _26488_ (.A1(_07931_),
    .A2(_07932_),
    .ZN(_07933_));
 XOR2_X1 _26489_ (.A(_07925_),
    .B(_07933_),
    .Z(_07934_));
 AOI22_X1 _26490_ (.A1(_07858_),
    .A2(_07927_),
    .B1(_07928_),
    .B2(_07934_),
    .ZN(_02359_));
 NAND3_X1 _26491_ (.A1(_04085_),
    .A2(_01184_),
    .A3(_04084_),
    .ZN(_07935_));
 NAND3_X1 _26492_ (.A1(_04823_),
    .A2(_07285_),
    .A3(_07835_),
    .ZN(_07936_));
 NAND3_X1 _26493_ (.A1(_07777_),
    .A2(_07935_),
    .A3(_07936_),
    .ZN(_07937_));
 AOI22_X2 _26494_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(_04067_),
    .B1(_04070_),
    .B2(\cs_registers_i.csr_mepc_o[25] ),
    .ZN(_07938_));
 NAND3_X1 _26495_ (.A1(_07817_),
    .A2(_07937_),
    .A3(_07938_),
    .ZN(_07939_));
 AND2_X1 _26496_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_04083_),
    .ZN(_07940_));
 OAI221_X2 _26497_ (.A(_04079_),
    .B1(_07939_),
    .B2(_07940_),
    .C1(_07868_),
    .C2(net24),
    .ZN(_07941_));
 INV_X1 _26498_ (.A(_07941_),
    .ZN(_07942_));
 AOI21_X2 _26499_ (.A(_07942_),
    .B1(_04304_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .ZN(_07943_));
 OAI21_X1 _26500_ (.A(_07928_),
    .B1(_07931_),
    .B2(_07932_),
    .ZN(_07944_));
 NAND4_X1 _26501_ (.A1(_07901_),
    .A2(_07911_),
    .A3(_07920_),
    .A4(_07944_),
    .ZN(_07945_));
 NOR2_X1 _26502_ (.A1(_07903_),
    .A2(_07945_),
    .ZN(_07946_));
 XNOR2_X1 _26503_ (.A(_07943_),
    .B(_07946_),
    .ZN(_07947_));
 MUX2_X1 _26504_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .B(_07947_),
    .S(_07914_),
    .Z(_02360_));
 AOI22_X4 _26505_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(_04066_),
    .B1(_04069_),
    .B2(\cs_registers_i.csr_mepc_o[26] ),
    .ZN(_07948_));
 OAI221_X2 _26506_ (.A(_07948_),
    .B1(_04010_),
    .B2(_03162_),
    .C1(_01185_),
    .C2(_07720_),
    .ZN(_07949_));
 AOI222_X2 _26507_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .A2(_04100_),
    .B1(_04043_),
    .B2(_07949_),
    .C1(_04370_),
    .C2(net25),
    .ZN(_07950_));
 OR2_X2 _26508_ (.A1(_07943_),
    .A2(_07945_),
    .ZN(_07951_));
 NOR3_X2 _26509_ (.A1(_07860_),
    .A2(_07923_),
    .A3(_07951_),
    .ZN(_07952_));
 XNOR2_X1 _26510_ (.A(_07950_),
    .B(_07952_),
    .ZN(_07953_));
 MUX2_X1 _26511_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .B(_07953_),
    .S(_07914_),
    .Z(_02361_));
 NAND3_X1 _26512_ (.A1(_04085_),
    .A2(_00007_),
    .A3(_04084_),
    .ZN(_07954_));
 NAND3_X1 _26513_ (.A1(_04854_),
    .A2(_07285_),
    .A3(_07835_),
    .ZN(_07955_));
 NAND3_X1 _26514_ (.A1(_07777_),
    .A2(_07954_),
    .A3(_07955_),
    .ZN(_07956_));
 AOI22_X1 _26515_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(_04067_),
    .B1(_04069_),
    .B2(\cs_registers_i.csr_mepc_o[27] ),
    .ZN(_07957_));
 NAND3_X1 _26516_ (.A1(_07715_),
    .A2(_07956_),
    .A3(_07957_),
    .ZN(_07958_));
 AND2_X2 _26517_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_04083_),
    .ZN(_07959_));
 OAI221_X2 _26518_ (.A(_04078_),
    .B1(_07958_),
    .B2(_07959_),
    .C1(_07817_),
    .C2(net26),
    .ZN(_07960_));
 NAND2_X1 _26519_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .A2(_04100_),
    .ZN(_07961_));
 AND2_X4 _26520_ (.A1(_07960_),
    .A2(_07961_),
    .ZN(_07962_));
 NOR3_X1 _26521_ (.A1(_07903_),
    .A2(_07950_),
    .A3(_07951_),
    .ZN(_07963_));
 XNOR2_X1 _26522_ (.A(_07962_),
    .B(_07963_),
    .ZN(_07964_));
 MUX2_X1 _26523_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .B(_07964_),
    .S(_07914_),
    .Z(_02362_));
 NAND2_X2 _26524_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .A2(_04304_),
    .ZN(_07965_));
 NOR2_X1 _26525_ (.A1(_07950_),
    .A2(_07962_),
    .ZN(_07966_));
 NAND2_X1 _26526_ (.A1(_07952_),
    .A2(_07966_),
    .ZN(_07967_));
 NOR2_X1 _26527_ (.A1(_04313_),
    .A2(_07967_),
    .ZN(_07968_));
 NAND3_X1 _26528_ (.A1(_04085_),
    .A2(_00008_),
    .A3(_04084_),
    .ZN(_07969_));
 NAND3_X1 _26529_ (.A1(_04869_),
    .A2(_07285_),
    .A3(_07835_),
    .ZN(_07970_));
 NAND3_X1 _26530_ (.A1(_07777_),
    .A2(_07969_),
    .A3(_07970_),
    .ZN(_07971_));
 AOI22_X2 _26531_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(_04067_),
    .B1(_04070_),
    .B2(\cs_registers_i.csr_mepc_o[28] ),
    .ZN(_07972_));
 NAND3_X1 _26532_ (.A1(_07868_),
    .A2(_07971_),
    .A3(_07972_),
    .ZN(_07973_));
 AND2_X2 _26533_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_07234_),
    .ZN(_07974_));
 OAI221_X2 _26534_ (.A(_04080_),
    .B1(_07974_),
    .B2(_07973_),
    .C1(_07868_),
    .C2(net27),
    .ZN(_07975_));
 AOI21_X1 _26535_ (.A(_07967_),
    .B1(_07975_),
    .B2(_07965_),
    .ZN(_07976_));
 INV_X1 _26536_ (.A(_07975_),
    .ZN(_07977_));
 AOI21_X1 _26537_ (.A(_07977_),
    .B1(_07966_),
    .B2(_07952_),
    .ZN(_07978_));
 OR2_X1 _26538_ (.A1(_07791_),
    .A2(_07978_),
    .ZN(_07979_));
 OAI22_X1 _26539_ (.A1(_07965_),
    .A2(_07968_),
    .B1(_07976_),
    .B2(_07979_),
    .ZN(_02363_));
 NAND2_X2 _26540_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .A2(_04303_),
    .ZN(_07980_));
 NAND2_X2 _26541_ (.A1(_07975_),
    .A2(_07965_),
    .ZN(_07981_));
 NAND2_X1 _26542_ (.A1(_07966_),
    .A2(_07981_),
    .ZN(_07982_));
 OR3_X1 _26543_ (.A1(_07903_),
    .A2(_07951_),
    .A3(_07982_),
    .ZN(_07983_));
 NOR2_X1 _26544_ (.A1(_04313_),
    .A2(_07983_),
    .ZN(_07984_));
 AND2_X4 _26545_ (.A1(_07234_),
    .A2(\alu_adder_result_ex[29] ),
    .ZN(_07985_));
 AOI221_X2 _26546_ (.A(_07724_),
    .B1(_04066_),
    .B2(\cs_registers_i.csr_depc_o[29] ),
    .C1(_04069_),
    .C2(\cs_registers_i.csr_mepc_o[29] ),
    .ZN(_07986_));
 OAI21_X1 _26547_ (.A(_07986_),
    .B1(_07827_),
    .B2(_00009_),
    .ZN(_07987_));
 OAI221_X2 _26548_ (.A(_04080_),
    .B1(_07987_),
    .B2(_07985_),
    .C1(_07868_),
    .C2(net28),
    .ZN(_07988_));
 AOI21_X1 _26549_ (.A(_07983_),
    .B1(_07988_),
    .B2(_07980_),
    .ZN(_07989_));
 NOR3_X1 _26550_ (.A1(_07903_),
    .A2(_07951_),
    .A3(_07982_),
    .ZN(_07990_));
 INV_X1 _26551_ (.A(_07988_),
    .ZN(_07991_));
 OAI21_X1 _26552_ (.A(_07774_),
    .B1(_07990_),
    .B2(_07991_),
    .ZN(_07992_));
 OAI22_X1 _26553_ (.A1(_07980_),
    .A2(_07984_),
    .B1(_07989_),
    .B2(_07992_),
    .ZN(_02364_));
 MUX2_X1 _26554_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ),
    .S(_07914_),
    .Z(_02365_));
 AND2_X2 _26555_ (.A1(_07234_),
    .A2(\alu_adder_result_ex[30] ),
    .ZN(_07993_));
 AOI221_X2 _26556_ (.A(_07724_),
    .B1(_04067_),
    .B2(\cs_registers_i.csr_depc_o[30] ),
    .C1(_04070_),
    .C2(\cs_registers_i.csr_mepc_o[30] ),
    .ZN(_07994_));
 OAI21_X1 _26557_ (.A(_07994_),
    .B1(_07827_),
    .B2(_00010_),
    .ZN(_07995_));
 OAI221_X2 _26558_ (.A(_04080_),
    .B1(_07995_),
    .B2(_07993_),
    .C1(_07868_),
    .C2(net29),
    .ZN(_07996_));
 INV_X1 _26559_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .ZN(_07997_));
 OAI21_X2 _26560_ (.A(_07996_),
    .B1(_04080_),
    .B2(_07997_),
    .ZN(_07998_));
 OR2_X1 _26561_ (.A1(_07950_),
    .A2(_07962_),
    .ZN(_07999_));
 AOI221_X2 _26562_ (.A(_07999_),
    .B1(_07980_),
    .B2(_07988_),
    .C1(_07975_),
    .C2(_07965_),
    .ZN(_08000_));
 NAND2_X1 _26563_ (.A1(_07952_),
    .A2(_08000_),
    .ZN(_08001_));
 XNOR2_X1 _26564_ (.A(_07998_),
    .B(_08001_),
    .ZN(_08002_));
 MUX2_X1 _26565_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .B(_08002_),
    .S(_07914_),
    .Z(_02366_));
 AND2_X2 _26566_ (.A1(_07234_),
    .A2(_03517_),
    .ZN(_08003_));
 AOI221_X2 _26567_ (.A(_07724_),
    .B1(_04067_),
    .B2(\cs_registers_i.csr_depc_o[31] ),
    .C1(_04070_),
    .C2(\cs_registers_i.csr_mepc_o[31] ),
    .ZN(_08004_));
 OAI21_X1 _26568_ (.A(_08004_),
    .B1(_07827_),
    .B2(_00011_),
    .ZN(_08005_));
 OAI221_X2 _26569_ (.A(_04080_),
    .B1(_08003_),
    .B2(_08005_),
    .C1(_07868_),
    .C2(net30),
    .ZN(_08006_));
 INV_X1 _26570_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .ZN(_08007_));
 OAI21_X2 _26571_ (.A(_08006_),
    .B1(_04081_),
    .B2(_08007_),
    .ZN(_08008_));
 NAND2_X1 _26572_ (.A1(_07998_),
    .A2(_08000_),
    .ZN(_08009_));
 NOR3_X1 _26573_ (.A1(_07903_),
    .A2(_07951_),
    .A3(_08009_),
    .ZN(_08010_));
 XOR2_X1 _26574_ (.A(_08008_),
    .B(_08010_),
    .Z(_08011_));
 MUX2_X1 _26575_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .B(_08011_),
    .S(_07914_),
    .Z(_02367_));
 MUX2_X1 _26576_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ),
    .S(_07914_),
    .Z(_02368_));
 NAND2_X1 _26577_ (.A1(_07743_),
    .A2(_07734_),
    .ZN(_08012_));
 XOR2_X1 _26578_ (.A(_16513_),
    .B(_08012_),
    .Z(_08013_));
 MUX2_X1 _26579_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .B(_08013_),
    .S(_07914_),
    .Z(_02369_));
 NAND3_X1 _26580_ (.A1(_16511_),
    .A2(_16512_),
    .A3(_08012_),
    .ZN(_08014_));
 XOR2_X1 _26581_ (.A(_07733_),
    .B(_08014_),
    .Z(_08015_));
 MUX2_X1 _26582_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .B(_08015_),
    .S(_07774_),
    .Z(_02370_));
 XNOR2_X1 _26583_ (.A(_07844_),
    .B(_07749_),
    .ZN(_08016_));
 MUX2_X1 _26584_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .B(_08016_),
    .S(_07774_),
    .Z(_02371_));
 NAND2_X1 _26585_ (.A1(_07749_),
    .A2(_07788_),
    .ZN(_08017_));
 XNOR2_X1 _26586_ (.A(_07755_),
    .B(_08017_),
    .ZN(_08018_));
 MUX2_X1 _26587_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .B(_08018_),
    .S(_07774_),
    .Z(_02372_));
 NAND3_X1 _26588_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .A2(_16509_),
    .A3(_07757_),
    .ZN(_08019_));
 OAI21_X1 _26589_ (.A(_08019_),
    .B1(_16509_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .ZN(_08020_));
 NOR2_X1 _26590_ (.A1(_07767_),
    .A2(_07769_),
    .ZN(_08021_));
 OAI21_X1 _26591_ (.A(_04081_),
    .B1(_07868_),
    .B2(net31),
    .ZN(_08022_));
 NOR2_X2 _26592_ (.A1(_08021_),
    .A2(_08022_),
    .ZN(_08023_));
 XNOR2_X1 _26593_ (.A(_07757_),
    .B(_08023_),
    .ZN(_08024_));
 AOI22_X1 _26594_ (.A1(_07858_),
    .A2(_08020_),
    .B1(_08024_),
    .B2(_07766_),
    .ZN(_02373_));
 AND2_X1 _26595_ (.A1(_07766_),
    .A2(_07770_),
    .ZN(_08025_));
 NAND2_X1 _26596_ (.A1(_07756_),
    .A2(_07788_),
    .ZN(_08026_));
 NOR2_X1 _26597_ (.A1(_08025_),
    .A2(_08026_),
    .ZN(_08027_));
 XNOR2_X1 _26598_ (.A(_07765_),
    .B(_08027_),
    .ZN(_08028_));
 MUX2_X1 _26599_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .B(_08028_),
    .S(_07774_),
    .Z(_02374_));
 CLKBUF_X3 _26600_ (.A(_04308_),
    .Z(_08029_));
 CLKBUF_X3 _26601_ (.A(_08029_),
    .Z(_08030_));
 MUX2_X1 _26602_ (.A(_04108_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .S(_08030_),
    .Z(_08031_));
 INV_X1 _26603_ (.A(_00135_),
    .ZN(_08032_));
 BUF_X4 _26604_ (.A(_04107_),
    .Z(_08033_));
 INV_X1 _26605_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .ZN(_08034_));
 NAND2_X1 _26606_ (.A1(_04305_),
    .A2(net124),
    .ZN(_08035_));
 INV_X1 _26607_ (.A(_08035_),
    .ZN(_08036_));
 NAND2_X2 _26608_ (.A1(_08034_),
    .A2(_08036_),
    .ZN(_08037_));
 NOR3_X1 _26609_ (.A1(_08033_),
    .A2(_04308_),
    .A3(_08037_),
    .ZN(_08038_));
 OR2_X1 _26610_ (.A1(_08032_),
    .A2(_08038_),
    .ZN(_08039_));
 BUF_X4 _26611_ (.A(_04121_),
    .Z(_08040_));
 NOR2_X1 _26612_ (.A1(_08040_),
    .A2(_08037_),
    .ZN(_08041_));
 OR2_X1 _26613_ (.A1(_07224_),
    .A2(_07245_),
    .ZN(_08042_));
 BUF_X4 _26614_ (.A(_08042_),
    .Z(_08043_));
 NAND2_X1 _26615_ (.A1(_00137_),
    .A2(_04122_),
    .ZN(_08044_));
 NOR2_X2 _26616_ (.A1(_03534_),
    .A2(_03979_),
    .ZN(_08045_));
 OAI21_X1 _26617_ (.A(_03650_),
    .B1(_07228_),
    .B2(_07281_),
    .ZN(_08046_));
 INV_X1 _26618_ (.A(_08046_),
    .ZN(_08047_));
 NOR3_X2 _26619_ (.A1(_03536_),
    .A2(_08045_),
    .A3(_08047_),
    .ZN(_08048_));
 OAI21_X1 _26620_ (.A(_00135_),
    .B1(_08037_),
    .B2(_00136_),
    .ZN(_08049_));
 NAND2_X1 _26621_ (.A1(_00136_),
    .A2(_08037_),
    .ZN(_08050_));
 MUX2_X1 _26622_ (.A(_08049_),
    .B(_08050_),
    .S(_04116_),
    .Z(_08051_));
 NAND2_X2 _26623_ (.A1(_08048_),
    .A2(_08051_),
    .ZN(_08052_));
 NOR3_X4 _26624_ (.A1(_07212_),
    .A2(_07269_),
    .A3(_08052_),
    .ZN(_08053_));
 NAND3_X2 _26625_ (.A1(_08043_),
    .A2(_08044_),
    .A3(_08053_),
    .ZN(_08054_));
 MUX2_X1 _26626_ (.A(_08039_),
    .B(_08041_),
    .S(_08054_),
    .Z(_08055_));
 CLKBUF_X3 _26627_ (.A(_08055_),
    .Z(_08056_));
 BUF_X4 _26628_ (.A(_08056_),
    .Z(_08057_));
 MUX2_X1 _26629_ (.A(_04113_),
    .B(_08031_),
    .S(_08057_),
    .Z(_02375_));
 BUF_X4 _26630_ (.A(_04306_),
    .Z(_08058_));
 MUX2_X1 _26631_ (.A(_04108_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .S(_08058_),
    .Z(_08059_));
 INV_X1 _26632_ (.A(_04306_),
    .ZN(_08060_));
 INV_X1 _26633_ (.A(_04308_),
    .ZN(_08061_));
 OAI21_X1 _26634_ (.A(_08060_),
    .B1(_08037_),
    .B2(_08061_),
    .ZN(_08062_));
 MUX2_X1 _26635_ (.A(_08062_),
    .B(_08038_),
    .S(_08054_),
    .Z(_08063_));
 CLKBUF_X3 _26636_ (.A(_08063_),
    .Z(_08064_));
 BUF_X4 _26637_ (.A(_08064_),
    .Z(_08065_));
 MUX2_X1 _26638_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B(_08059_),
    .S(_08065_),
    .Z(_02376_));
 NOR3_X4 _26639_ (.A1(_08061_),
    .A2(_04306_),
    .A3(_08037_),
    .ZN(_08066_));
 BUF_X4 _26640_ (.A(_08066_),
    .Z(_08067_));
 MUX2_X1 _26641_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .B(_04108_),
    .S(_08067_),
    .Z(_02377_));
 BUF_X4 _26642_ (.A(_04081_),
    .Z(_08068_));
 INV_X1 _26643_ (.A(_00555_),
    .ZN(_08069_));
 AOI22_X2 _26644_ (.A1(\cs_registers_i.csr_mepc_o[1] ),
    .A2(_07289_),
    .B1(_07751_),
    .B2(_08069_),
    .ZN(_08070_));
 OAI21_X2 _26645_ (.A(_08070_),
    .B1(_04073_),
    .B2(_16491_),
    .ZN(_08071_));
 NAND2_X1 _26646_ (.A1(_08068_),
    .A2(_08071_),
    .ZN(_08072_));
 INV_X2 _26647_ (.A(_04104_),
    .ZN(_08073_));
 BUF_X4 _26648_ (.A(_08073_),
    .Z(_08074_));
 NAND3_X1 _26649_ (.A1(_08074_),
    .A2(_04304_),
    .A3(_04122_),
    .ZN(_08075_));
 NAND2_X4 _26650_ (.A1(_08043_),
    .A2(_08053_),
    .ZN(_08076_));
 BUF_X4 _26651_ (.A(_08076_),
    .Z(_08077_));
 CLKBUF_X3 _26652_ (.A(_07246_),
    .Z(_08078_));
 OR3_X1 _26653_ (.A1(_07212_),
    .A2(_08078_),
    .A3(_07269_),
    .ZN(_08079_));
 INV_X1 _26654_ (.A(_04115_),
    .ZN(_08080_));
 NAND3_X1 _26655_ (.A1(_08080_),
    .A2(_08048_),
    .A3(_08050_),
    .ZN(_08081_));
 OAI21_X1 _26656_ (.A(_04123_),
    .B1(_08079_),
    .B2(_08081_),
    .ZN(_08082_));
 OAI221_X2 _26657_ (.A(_08072_),
    .B1(_08075_),
    .B2(_08077_),
    .C1(_08082_),
    .C2(_08068_),
    .ZN(_02378_));
 BUF_X1 _26658_ (.A(\cs_registers_i.pc_if_i[11] ),
    .Z(_08083_));
 OR3_X1 _26659_ (.A1(_07212_),
    .A2(_07269_),
    .A3(_08052_),
    .ZN(_08084_));
 CLKBUF_X3 _26660_ (.A(_08084_),
    .Z(_08085_));
 CLKBUF_X2 _26661_ (.A(\cs_registers_i.pc_if_i[9] ),
    .Z(_08086_));
 NAND2_X1 _26662_ (.A1(_08086_),
    .A2(\cs_registers_i.pc_if_i[10] ),
    .ZN(_08087_));
 INV_X1 _26663_ (.A(\cs_registers_i.pc_if_i[5] ),
    .ZN(_08088_));
 INV_X1 _26664_ (.A(\cs_registers_i.pc_if_i[3] ),
    .ZN(_08089_));
 INV_X1 _26665_ (.A(\cs_registers_i.pc_if_i[4] ),
    .ZN(_08090_));
 OR3_X1 _26666_ (.A1(_08089_),
    .A2(_08090_),
    .A3(_15757_),
    .ZN(_08091_));
 OR2_X1 _26667_ (.A1(_08088_),
    .A2(_08091_),
    .ZN(_08092_));
 CLKBUF_X2 _26668_ (.A(\cs_registers_i.pc_if_i[7] ),
    .Z(_08093_));
 NAND3_X2 _26669_ (.A1(\cs_registers_i.pc_if_i[6] ),
    .A2(_08093_),
    .A3(\cs_registers_i.pc_if_i[8] ),
    .ZN(_08094_));
 NOR2_X1 _26670_ (.A1(_08092_),
    .A2(_08094_),
    .ZN(_08095_));
 INV_X1 _26671_ (.A(_08095_),
    .ZN(_08096_));
 NOR4_X1 _26672_ (.A1(_08078_),
    .A2(_08085_),
    .A3(_08087_),
    .A4(_08096_),
    .ZN(_08097_));
 XNOR2_X1 _26673_ (.A(_08083_),
    .B(_08097_),
    .ZN(_08098_));
 OAI21_X1 _26674_ (.A(_07785_),
    .B1(_08098_),
    .B2(_08068_),
    .ZN(_02379_));
 OAI21_X1 _26675_ (.A(_04304_),
    .B1(_08078_),
    .B2(_08085_),
    .ZN(_08099_));
 CLKBUF_X3 _26676_ (.A(_08099_),
    .Z(_08100_));
 OR2_X1 _26677_ (.A1(_07794_),
    .A2(_07795_),
    .ZN(_08101_));
 AND2_X1 _26678_ (.A1(_08086_),
    .A2(\cs_registers_i.pc_if_i[10] ),
    .ZN(_08102_));
 AOI21_X1 _26679_ (.A(_16233_),
    .B1(_04169_),
    .B2(_16234_),
    .ZN(_08103_));
 NOR3_X1 _26680_ (.A1(_08089_),
    .A2(_08090_),
    .A3(_08103_),
    .ZN(_08104_));
 INV_X1 _26681_ (.A(_08104_),
    .ZN(_08105_));
 NOR3_X4 _26682_ (.A1(_08088_),
    .A2(_08094_),
    .A3(_08105_),
    .ZN(_08106_));
 NAND3_X1 _26683_ (.A1(_08083_),
    .A2(_08102_),
    .A3(_08106_),
    .ZN(_08107_));
 NAND2_X1 _26684_ (.A1(_08101_),
    .A2(_08107_),
    .ZN(_08108_));
 AOI21_X1 _26685_ (.A(\cs_registers_i.pc_if_i[12] ),
    .B1(_08100_),
    .B2(_08108_),
    .ZN(_08109_));
 CLKBUF_X3 _26686_ (.A(_04304_),
    .Z(_08110_));
 NAND3_X1 _26687_ (.A1(_08083_),
    .A2(\cs_registers_i.pc_if_i[12] ),
    .A3(_08102_),
    .ZN(_08111_));
 NAND3_X2 _26688_ (.A1(_08043_),
    .A2(_08053_),
    .A3(_08106_),
    .ZN(_08112_));
 OAI21_X1 _26689_ (.A(_08110_),
    .B1(_08111_),
    .B2(_08112_),
    .ZN(_08113_));
 AOI21_X1 _26690_ (.A(_08109_),
    .B1(_08113_),
    .B2(_08101_),
    .ZN(_02380_));
 NOR4_X1 _26691_ (.A1(_08078_),
    .A2(_08085_),
    .A3(_08096_),
    .A4(_08111_),
    .ZN(_08114_));
 XNOR2_X1 _26692_ (.A(\cs_registers_i.pc_if_i[13] ),
    .B(_08114_),
    .ZN(_08115_));
 AOI21_X1 _26693_ (.A(_07809_),
    .B1(_08115_),
    .B2(_07858_),
    .ZN(_02381_));
 INV_X1 _26694_ (.A(\cs_registers_i.pc_if_i[13] ),
    .ZN(_08116_));
 NOR2_X1 _26695_ (.A1(_08116_),
    .A2(_08111_),
    .ZN(_08117_));
 NAND2_X1 _26696_ (.A1(_08106_),
    .A2(_08117_),
    .ZN(_08118_));
 NAND2_X1 _26697_ (.A1(_07818_),
    .A2(_08118_),
    .ZN(_08119_));
 AOI21_X1 _26698_ (.A(\cs_registers_i.pc_if_i[14] ),
    .B1(_08100_),
    .B2(_08119_),
    .ZN(_08120_));
 NAND2_X1 _26699_ (.A1(\cs_registers_i.pc_if_i[14] ),
    .A2(_08117_),
    .ZN(_08121_));
 OAI21_X1 _26700_ (.A(_08110_),
    .B1(_08112_),
    .B2(_08121_),
    .ZN(_08122_));
 AOI21_X1 _26701_ (.A(_08120_),
    .B1(_08122_),
    .B2(_07818_),
    .ZN(_02382_));
 CLKBUF_X2 _26702_ (.A(\cs_registers_i.pc_if_i[15] ),
    .Z(_08123_));
 OAI21_X1 _26703_ (.A(_07829_),
    .B1(_08096_),
    .B2(_08121_),
    .ZN(_08124_));
 AOI21_X1 _26704_ (.A(_08123_),
    .B1(_08100_),
    .B2(_08124_),
    .ZN(_08125_));
 NOR2_X1 _26705_ (.A1(_08096_),
    .A2(_08121_),
    .ZN(_08126_));
 NAND2_X1 _26706_ (.A1(_08123_),
    .A2(_08126_),
    .ZN(_08127_));
 OAI21_X1 _26707_ (.A(_08110_),
    .B1(_08077_),
    .B2(_08127_),
    .ZN(_08128_));
 AOI21_X1 _26708_ (.A(_08125_),
    .B1(_08128_),
    .B2(_07829_),
    .ZN(_02383_));
 INV_X1 _26709_ (.A(_08106_),
    .ZN(_08129_));
 NOR2_X1 _26710_ (.A1(_08129_),
    .A2(_08121_),
    .ZN(_08130_));
 NAND2_X1 _26711_ (.A1(_08123_),
    .A2(_08130_),
    .ZN(_08131_));
 NAND2_X1 _26712_ (.A1(_07841_),
    .A2(_08131_),
    .ZN(_08132_));
 AOI21_X1 _26713_ (.A(\cs_registers_i.pc_if_i[16] ),
    .B1(_08100_),
    .B2(_08132_),
    .ZN(_08133_));
 AND3_X1 _26714_ (.A1(_08123_),
    .A2(\cs_registers_i.pc_if_i[16] ),
    .A3(_08130_),
    .ZN(_08134_));
 INV_X1 _26715_ (.A(_08134_),
    .ZN(_08135_));
 OAI21_X1 _26716_ (.A(_08110_),
    .B1(_08077_),
    .B2(_08135_),
    .ZN(_08136_));
 AOI21_X1 _26717_ (.A(_08133_),
    .B1(_08136_),
    .B2(_07841_),
    .ZN(_02384_));
 CLKBUF_X3 _26718_ (.A(_04304_),
    .Z(_08137_));
 BUF_X1 _26719_ (.A(\cs_registers_i.pc_if_i[17] ),
    .Z(_08138_));
 AND3_X1 _26720_ (.A1(_08123_),
    .A2(\cs_registers_i.pc_if_i[16] ),
    .A3(_08126_),
    .ZN(_08139_));
 NAND2_X1 _26721_ (.A1(_08138_),
    .A2(_08139_),
    .ZN(_08140_));
 OAI21_X1 _26722_ (.A(_08137_),
    .B1(_08077_),
    .B2(_08140_),
    .ZN(_08141_));
 CLKBUF_X3 _26723_ (.A(_08099_),
    .Z(_08142_));
 INV_X1 _26724_ (.A(_07851_),
    .ZN(_08143_));
 OAI21_X1 _26725_ (.A(_08142_),
    .B1(_08139_),
    .B2(_08143_),
    .ZN(_08144_));
 INV_X1 _26726_ (.A(_08138_),
    .ZN(_08145_));
 AOI22_X1 _26727_ (.A1(_07851_),
    .A2(_08141_),
    .B1(_08144_),
    .B2(_08145_),
    .ZN(_02385_));
 OAI21_X1 _26728_ (.A(_07869_),
    .B1(_08135_),
    .B2(_08145_),
    .ZN(_08146_));
 AOI21_X1 _26729_ (.A(\cs_registers_i.pc_if_i[18] ),
    .B1(_08100_),
    .B2(_08146_),
    .ZN(_08147_));
 AND3_X1 _26730_ (.A1(_08138_),
    .A2(\cs_registers_i.pc_if_i[18] ),
    .A3(_08134_),
    .ZN(_08148_));
 NAND3_X1 _26731_ (.A1(_08043_),
    .A2(_08053_),
    .A3(_08148_),
    .ZN(_08149_));
 NAND2_X1 _26732_ (.A1(_08110_),
    .A2(_08149_),
    .ZN(_08150_));
 AOI21_X1 _26733_ (.A(_08147_),
    .B1(_08150_),
    .B2(_07869_),
    .ZN(_02386_));
 CLKBUF_X2 _26734_ (.A(\cs_registers_i.pc_if_i[19] ),
    .Z(_08151_));
 NOR2_X2 _26735_ (.A1(_07246_),
    .A2(_08085_),
    .ZN(_08152_));
 BUF_X8 _26736_ (.A(_08152_),
    .Z(_08153_));
 AND3_X1 _26737_ (.A1(_08138_),
    .A2(\cs_registers_i.pc_if_i[18] ),
    .A3(_08139_),
    .ZN(_08154_));
 AND4_X1 _26738_ (.A1(_08151_),
    .A2(_07875_),
    .A3(_08153_),
    .A4(_08154_),
    .ZN(_08155_));
 NOR3_X1 _26739_ (.A1(_08151_),
    .A2(_08068_),
    .A3(_08153_),
    .ZN(_08156_));
 NOR2_X1 _26740_ (.A1(_08151_),
    .A2(_08154_),
    .ZN(_08157_));
 OAI21_X1 _26741_ (.A(_07875_),
    .B1(_08157_),
    .B2(_04081_),
    .ZN(_08158_));
 INV_X1 _26742_ (.A(_08158_),
    .ZN(_08159_));
 NOR3_X1 _26743_ (.A1(_08155_),
    .A2(_08156_),
    .A3(_08159_),
    .ZN(_02387_));
 NAND2_X1 _26744_ (.A1(_07887_),
    .A2(_07889_),
    .ZN(_08160_));
 NAND2_X1 _26745_ (.A1(_08151_),
    .A2(_08148_),
    .ZN(_08161_));
 NAND2_X1 _26746_ (.A1(_08160_),
    .A2(_08161_),
    .ZN(_08162_));
 AOI21_X1 _26747_ (.A(\cs_registers_i.pc_if_i[20] ),
    .B1(_08100_),
    .B2(_08162_),
    .ZN(_08163_));
 NAND2_X1 _26748_ (.A1(_08151_),
    .A2(\cs_registers_i.pc_if_i[20] ),
    .ZN(_08164_));
 OAI21_X1 _26749_ (.A(_08110_),
    .B1(_08149_),
    .B2(_08164_),
    .ZN(_08165_));
 AOI21_X1 _26750_ (.A(_08163_),
    .B1(_08165_),
    .B2(_08160_),
    .ZN(_02388_));
 NOR3_X1 _26751_ (.A1(_15758_),
    .A2(_08078_),
    .A3(_08085_),
    .ZN(_08166_));
 AOI21_X1 _26752_ (.A(_08166_),
    .B1(_08077_),
    .B2(\cs_registers_i.pc_if_i[2] ),
    .ZN(_08167_));
 OAI21_X1 _26753_ (.A(_04075_),
    .B1(_08167_),
    .B2(_08068_),
    .ZN(_02389_));
 BUF_X1 _26754_ (.A(\cs_registers_i.pc_if_i[21] ),
    .Z(_08168_));
 AND2_X1 _26755_ (.A1(_08151_),
    .A2(\cs_registers_i.pc_if_i[20] ),
    .ZN(_08169_));
 NAND4_X1 _26756_ (.A1(_08043_),
    .A2(_08053_),
    .A3(_08154_),
    .A4(_08169_),
    .ZN(_08170_));
 XOR2_X1 _26757_ (.A(_08168_),
    .B(_08170_),
    .Z(_08171_));
 OAI21_X1 _26758_ (.A(_07899_),
    .B1(_08171_),
    .B2(_08068_),
    .ZN(_02390_));
 AND2_X1 _26759_ (.A1(_07905_),
    .A2(_07909_),
    .ZN(_08172_));
 NAND3_X1 _26760_ (.A1(_08168_),
    .A2(_08148_),
    .A3(_08169_),
    .ZN(_08173_));
 NAND2_X1 _26761_ (.A1(_08172_),
    .A2(_08173_),
    .ZN(_08174_));
 AOI21_X1 _26762_ (.A(\cs_registers_i.pc_if_i[22] ),
    .B1(_08100_),
    .B2(_08174_),
    .ZN(_08175_));
 AND3_X1 _26763_ (.A1(_08168_),
    .A2(\cs_registers_i.pc_if_i[22] ),
    .A3(_08169_),
    .ZN(_08176_));
 NAND2_X2 _26764_ (.A1(_08148_),
    .A2(_08176_),
    .ZN(_08177_));
 OR3_X2 _26765_ (.A1(_08078_),
    .A2(_08085_),
    .A3(_08177_),
    .ZN(_08178_));
 NAND2_X1 _26766_ (.A1(_08110_),
    .A2(_08178_),
    .ZN(_08179_));
 AOI21_X1 _26767_ (.A(_08175_),
    .B1(_08179_),
    .B2(_08172_),
    .ZN(_02391_));
 AND2_X1 _26768_ (.A1(_08068_),
    .A2(_07918_),
    .ZN(_08180_));
 INV_X1 _26769_ (.A(\cs_registers_i.pc_if_i[23] ),
    .ZN(_08181_));
 NAND2_X2 _26770_ (.A1(_08154_),
    .A2(_08176_),
    .ZN(_08182_));
 OR3_X2 _26771_ (.A1(_08078_),
    .A2(_08085_),
    .A3(_08182_),
    .ZN(_08183_));
 XNOR2_X1 _26772_ (.A(_08181_),
    .B(_08183_),
    .ZN(_08184_));
 AOI21_X1 _26773_ (.A(_08180_),
    .B1(_08184_),
    .B2(_07858_),
    .ZN(_02392_));
 OAI21_X1 _26774_ (.A(_07933_),
    .B1(_08177_),
    .B2(_08181_),
    .ZN(_08185_));
 AOI21_X1 _26775_ (.A(\cs_registers_i.pc_if_i[24] ),
    .B1(_08100_),
    .B2(_08185_),
    .ZN(_08186_));
 NAND2_X1 _26776_ (.A1(\cs_registers_i.pc_if_i[23] ),
    .A2(\cs_registers_i.pc_if_i[24] ),
    .ZN(_08187_));
 OAI21_X1 _26777_ (.A(_08110_),
    .B1(_08178_),
    .B2(_08187_),
    .ZN(_08188_));
 AOI21_X1 _26778_ (.A(_08186_),
    .B1(_08188_),
    .B2(_07933_),
    .ZN(_02393_));
 OAI21_X1 _26779_ (.A(_07941_),
    .B1(_08182_),
    .B2(_08187_),
    .ZN(_08189_));
 AOI21_X1 _26780_ (.A(\cs_registers_i.pc_if_i[25] ),
    .B1(_08100_),
    .B2(_08189_),
    .ZN(_08190_));
 AND3_X1 _26781_ (.A1(\cs_registers_i.pc_if_i[23] ),
    .A2(\cs_registers_i.pc_if_i[24] ),
    .A3(\cs_registers_i.pc_if_i[25] ),
    .ZN(_08191_));
 INV_X1 _26782_ (.A(_08191_),
    .ZN(_08192_));
 OAI21_X1 _26783_ (.A(_08110_),
    .B1(_08183_),
    .B2(_08192_),
    .ZN(_08193_));
 AOI21_X1 _26784_ (.A(_08190_),
    .B1(_08193_),
    .B2(_07941_),
    .ZN(_02394_));
 CLKBUF_X2 _26785_ (.A(\cs_registers_i.pc_if_i[26] ),
    .Z(_08194_));
 AOI22_X2 _26786_ (.A1(net25),
    .A2(_04370_),
    .B1(_07949_),
    .B2(_04043_),
    .ZN(_08195_));
 OAI21_X1 _26787_ (.A(_08195_),
    .B1(_08177_),
    .B2(_08192_),
    .ZN(_08196_));
 AOI21_X1 _26788_ (.A(_08194_),
    .B1(_08142_),
    .B2(_08196_),
    .ZN(_08197_));
 NAND2_X1 _26789_ (.A1(_08194_),
    .A2(_08191_),
    .ZN(_08198_));
 OAI21_X1 _26790_ (.A(_08110_),
    .B1(_08178_),
    .B2(_08198_),
    .ZN(_08199_));
 AOI21_X1 _26791_ (.A(_08197_),
    .B1(_08199_),
    .B2(_08195_),
    .ZN(_02395_));
 OAI21_X1 _26792_ (.A(_07960_),
    .B1(_08182_),
    .B2(_08198_),
    .ZN(_08200_));
 AOI21_X1 _26793_ (.A(\cs_registers_i.pc_if_i[27] ),
    .B1(_08142_),
    .B2(_08200_),
    .ZN(_08201_));
 NAND3_X1 _26794_ (.A1(_08194_),
    .A2(\cs_registers_i.pc_if_i[27] ),
    .A3(_08191_),
    .ZN(_08202_));
 OAI21_X1 _26795_ (.A(_08137_),
    .B1(_08183_),
    .B2(_08202_),
    .ZN(_08203_));
 AOI21_X1 _26796_ (.A(_08201_),
    .B1(_08203_),
    .B2(_07960_),
    .ZN(_02396_));
 OAI21_X1 _26797_ (.A(_07975_),
    .B1(_08177_),
    .B2(_08202_),
    .ZN(_08204_));
 AOI21_X1 _26798_ (.A(\cs_registers_i.pc_if_i[28] ),
    .B1(_08142_),
    .B2(_08204_),
    .ZN(_08205_));
 AND3_X1 _26799_ (.A1(_08194_),
    .A2(\cs_registers_i.pc_if_i[27] ),
    .A3(_08191_),
    .ZN(_08206_));
 NAND2_X1 _26800_ (.A1(\cs_registers_i.pc_if_i[28] ),
    .A2(_08206_),
    .ZN(_08207_));
 OAI21_X1 _26801_ (.A(_08137_),
    .B1(_08178_),
    .B2(_08207_),
    .ZN(_08208_));
 AOI21_X1 _26802_ (.A(_08205_),
    .B1(_08208_),
    .B2(_07975_),
    .ZN(_02397_));
 BUF_X1 _26803_ (.A(\cs_registers_i.pc_if_i[29] ),
    .Z(_08209_));
 OAI21_X1 _26804_ (.A(_07988_),
    .B1(_08182_),
    .B2(_08207_),
    .ZN(_08210_));
 AOI21_X1 _26805_ (.A(_08209_),
    .B1(_08142_),
    .B2(_08210_),
    .ZN(_08211_));
 AND2_X1 _26806_ (.A1(\cs_registers_i.pc_if_i[28] ),
    .A2(_08206_),
    .ZN(_08212_));
 NAND2_X1 _26807_ (.A1(_08209_),
    .A2(_08212_),
    .ZN(_08213_));
 OAI21_X1 _26808_ (.A(_08137_),
    .B1(_08183_),
    .B2(_08213_),
    .ZN(_08214_));
 AOI21_X1 _26809_ (.A(_08211_),
    .B1(_08214_),
    .B2(_07988_),
    .ZN(_02398_));
 OAI21_X1 _26810_ (.A(_07996_),
    .B1(_08177_),
    .B2(_08213_),
    .ZN(_08215_));
 AOI21_X1 _26811_ (.A(\cs_registers_i.pc_if_i[30] ),
    .B1(_08142_),
    .B2(_08215_),
    .ZN(_08216_));
 NAND3_X1 _26812_ (.A1(_08209_),
    .A2(\cs_registers_i.pc_if_i[30] ),
    .A3(_08212_),
    .ZN(_08217_));
 OAI21_X1 _26813_ (.A(_08137_),
    .B1(_08178_),
    .B2(_08217_),
    .ZN(_08218_));
 AOI21_X1 _26814_ (.A(_08216_),
    .B1(_08218_),
    .B2(_07996_),
    .ZN(_02399_));
 NOR3_X1 _26815_ (.A1(_15757_),
    .A2(_08078_),
    .A3(_08085_),
    .ZN(_08219_));
 XNOR2_X1 _26816_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(_08219_),
    .ZN(_08220_));
 AOI21_X1 _26817_ (.A(_04099_),
    .B1(_08220_),
    .B2(_07858_),
    .ZN(_02400_));
 OAI21_X1 _26818_ (.A(_08006_),
    .B1(_08182_),
    .B2(_08217_),
    .ZN(_08221_));
 AOI21_X1 _26819_ (.A(\cs_registers_i.pc_if_i[31] ),
    .B1(_08142_),
    .B2(_08221_),
    .ZN(_08222_));
 NOR2_X1 _26820_ (.A1(_08182_),
    .A2(_08217_),
    .ZN(_08223_));
 NAND2_X1 _26821_ (.A1(\cs_registers_i.pc_if_i[31] ),
    .A2(_08223_),
    .ZN(_08224_));
 OAI21_X1 _26822_ (.A(_08137_),
    .B1(_08077_),
    .B2(_08224_),
    .ZN(_08225_));
 AOI21_X1 _26823_ (.A(_08222_),
    .B1(_08225_),
    .B2(_08006_),
    .ZN(_02401_));
 OAI21_X1 _26824_ (.A(_07743_),
    .B1(_08103_),
    .B2(_08089_),
    .ZN(_08226_));
 AOI21_X1 _26825_ (.A(\cs_registers_i.pc_if_i[4] ),
    .B1(_08142_),
    .B2(_08226_),
    .ZN(_08227_));
 OAI21_X1 _26826_ (.A(_08137_),
    .B1(_08077_),
    .B2(_08105_),
    .ZN(_08228_));
 AOI21_X1 _26827_ (.A(_08227_),
    .B1(_08228_),
    .B2(_07743_),
    .ZN(_02402_));
 NAND2_X1 _26828_ (.A1(_07731_),
    .A2(_08091_),
    .ZN(_08229_));
 AOI21_X1 _26829_ (.A(\cs_registers_i.pc_if_i[5] ),
    .B1(_08142_),
    .B2(_08229_),
    .ZN(_08230_));
 OAI21_X1 _26830_ (.A(_08137_),
    .B1(_08077_),
    .B2(_08092_),
    .ZN(_08231_));
 AOI21_X1 _26831_ (.A(_08230_),
    .B1(_08231_),
    .B2(_07731_),
    .ZN(_02403_));
 OR2_X1 _26832_ (.A1(_04304_),
    .A2(_07748_),
    .ZN(_08232_));
 INV_X1 _26833_ (.A(\cs_registers_i.pc_if_i[6] ),
    .ZN(_08233_));
 NOR2_X1 _26834_ (.A1(_08088_),
    .A2(_08105_),
    .ZN(_08234_));
 NAND3_X1 _26835_ (.A1(_08043_),
    .A2(_08053_),
    .A3(_08234_),
    .ZN(_08235_));
 XNOR2_X1 _26836_ (.A(_08233_),
    .B(_08235_),
    .ZN(_08236_));
 OAI21_X1 _26837_ (.A(_08232_),
    .B1(_08236_),
    .B2(_08068_),
    .ZN(_02404_));
 NOR4_X1 _26838_ (.A1(_08233_),
    .A2(_08078_),
    .A3(_08085_),
    .A4(_08092_),
    .ZN(_08237_));
 XNOR2_X1 _26839_ (.A(_08093_),
    .B(_08237_),
    .ZN(_08238_));
 AOI21_X1 _26840_ (.A(_07753_),
    .B1(_08238_),
    .B2(_07858_),
    .ZN(_02405_));
 AOI21_X1 _26841_ (.A(_08023_),
    .B1(_08112_),
    .B2(_08137_),
    .ZN(_08239_));
 AND3_X1 _26842_ (.A1(\cs_registers_i.pc_if_i[6] ),
    .A2(_08093_),
    .A3(_08234_),
    .ZN(_08240_));
 OAI21_X1 _26843_ (.A(_08100_),
    .B1(_08240_),
    .B2(_08023_),
    .ZN(_08241_));
 INV_X1 _26844_ (.A(\cs_registers_i.pc_if_i[8] ),
    .ZN(_08242_));
 AOI21_X1 _26845_ (.A(_08239_),
    .B1(_08241_),
    .B2(_08242_),
    .ZN(_02406_));
 INV_X1 _26846_ (.A(_07764_),
    .ZN(_08243_));
 NOR3_X1 _26847_ (.A1(_08078_),
    .A2(_08085_),
    .A3(_08096_),
    .ZN(_08244_));
 XNOR2_X1 _26848_ (.A(_08086_),
    .B(_08244_),
    .ZN(_08245_));
 OAI21_X1 _26849_ (.A(_08243_),
    .B1(_08245_),
    .B2(_08068_),
    .ZN(_02407_));
 OR2_X1 _26850_ (.A1(_07722_),
    .A2(_07716_),
    .ZN(_08246_));
 INV_X1 _26851_ (.A(_08086_),
    .ZN(_08247_));
 OAI21_X1 _26852_ (.A(_08246_),
    .B1(_08129_),
    .B2(_08247_),
    .ZN(_08248_));
 AOI21_X1 _26853_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B1(_08142_),
    .B2(_08248_),
    .ZN(_08249_));
 OAI21_X1 _26854_ (.A(_08137_),
    .B1(_08087_),
    .B2(_08112_),
    .ZN(_08250_));
 AOI21_X1 _26855_ (.A(_08249_),
    .B1(_08250_),
    .B2(_08246_),
    .ZN(_02408_));
 MUX2_X1 _26856_ (.A(net94),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_08251_));
 MUX2_X1 _26857_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .B(_08251_),
    .S(_08057_),
    .Z(_02409_));
 MUX2_X1 _26858_ (.A(net95),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(_04307_),
    .Z(_08252_));
 MUX2_X1 _26859_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .B(_08252_),
    .S(_08057_),
    .Z(_02410_));
 MUX2_X1 _26860_ (.A(net96),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_08253_));
 MUX2_X1 _26861_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .B(_08253_),
    .S(_08057_),
    .Z(_02411_));
 MUX2_X1 _26862_ (.A(net97),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(_04308_),
    .Z(_08254_));
 MUX2_X1 _26863_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .B(_08254_),
    .S(_08057_),
    .Z(_02412_));
 MUX2_X1 _26864_ (.A(net98),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(_04308_),
    .Z(_08255_));
 MUX2_X1 _26865_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .B(_08255_),
    .S(_08057_),
    .Z(_02413_));
 MUX2_X1 _26866_ (.A(net99),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(_04307_),
    .Z(_08256_));
 MUX2_X1 _26867_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .B(_08256_),
    .S(_08057_),
    .Z(_02414_));
 MUX2_X1 _26868_ (.A(net100),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(_04308_),
    .Z(_08257_));
 MUX2_X1 _26869_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .B(_08257_),
    .S(_08057_),
    .Z(_02415_));
 MUX2_X1 _26870_ (.A(_04110_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .S(_08030_),
    .Z(_08258_));
 MUX2_X1 _26871_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .B(_08258_),
    .S(_08057_),
    .Z(_02416_));
 MUX2_X1 _26872_ (.A(_04109_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .S(_08030_),
    .Z(_08259_));
 MUX2_X1 _26873_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .B(_08259_),
    .S(_08057_),
    .Z(_02417_));
 MUX2_X1 _26874_ (.A(net101),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .S(_08030_),
    .Z(_08260_));
 BUF_X4 _26875_ (.A(_08056_),
    .Z(_08261_));
 MUX2_X1 _26876_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .B(_08260_),
    .S(_08261_),
    .Z(_02418_));
 MUX2_X1 _26877_ (.A(net102),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .S(_08030_),
    .Z(_08262_));
 MUX2_X1 _26878_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .B(_08262_),
    .S(_08261_),
    .Z(_02419_));
 MUX2_X1 _26879_ (.A(net103),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(_04307_),
    .Z(_08263_));
 MUX2_X1 _26880_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B(_08263_),
    .S(_08261_),
    .Z(_02420_));
 MUX2_X1 _26881_ (.A(net104),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .S(_08030_),
    .Z(_08264_));
 MUX2_X1 _26882_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .B(_08264_),
    .S(_08261_),
    .Z(_02421_));
 MUX2_X1 _26883_ (.A(net105),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .S(_08030_),
    .Z(_08265_));
 MUX2_X1 _26884_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .B(_08265_),
    .S(_08261_),
    .Z(_02422_));
 MUX2_X1 _26885_ (.A(net106),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .S(_08030_),
    .Z(_08266_));
 MUX2_X1 _26886_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .B(_08266_),
    .S(_08261_),
    .Z(_02423_));
 MUX2_X1 _26887_ (.A(net107),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .S(_08030_),
    .Z(_08267_));
 MUX2_X1 _26888_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .B(_08267_),
    .S(_08261_),
    .Z(_02424_));
 MUX2_X1 _26889_ (.A(net108),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .S(_08030_),
    .Z(_08268_));
 MUX2_X1 _26890_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .B(_08268_),
    .S(_08261_),
    .Z(_02425_));
 MUX2_X1 _26891_ (.A(net109),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .S(_08029_),
    .Z(_08269_));
 MUX2_X1 _26892_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .B(_08269_),
    .S(_08261_),
    .Z(_02426_));
 MUX2_X1 _26893_ (.A(net110),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .S(_08029_),
    .Z(_08270_));
 MUX2_X1 _26894_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .B(_08270_),
    .S(_08261_),
    .Z(_02427_));
 MUX2_X1 _26895_ (.A(net111),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .S(_08029_),
    .Z(_08271_));
 BUF_X4 _26896_ (.A(_08056_),
    .Z(_08272_));
 MUX2_X1 _26897_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .B(_08271_),
    .S(_08272_),
    .Z(_02428_));
 MUX2_X1 _26898_ (.A(net112),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .S(_08029_),
    .Z(_08273_));
 MUX2_X1 _26899_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .B(_08273_),
    .S(_08272_),
    .Z(_02429_));
 MUX2_X1 _26900_ (.A(net113),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .S(_08029_),
    .Z(_08274_));
 MUX2_X1 _26901_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .B(_08274_),
    .S(_08272_),
    .Z(_02430_));
 MUX2_X1 _26902_ (.A(net114),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(_04307_),
    .Z(_08275_));
 MUX2_X1 _26903_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .B(_08275_),
    .S(_08272_),
    .Z(_02431_));
 MUX2_X1 _26904_ (.A(net115),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .S(_08029_),
    .Z(_08276_));
 MUX2_X1 _26905_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .B(_08276_),
    .S(_08272_),
    .Z(_02432_));
 MUX2_X1 _26906_ (.A(net116),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .S(_08029_),
    .Z(_08277_));
 MUX2_X1 _26907_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .B(_08277_),
    .S(_08272_),
    .Z(_02433_));
 MUX2_X1 _26908_ (.A(net94),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(_08058_),
    .Z(_08278_));
 MUX2_X1 _26909_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .B(_08278_),
    .S(_08065_),
    .Z(_02434_));
 MUX2_X1 _26910_ (.A(net103),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(_08058_),
    .Z(_08279_));
 MUX2_X1 _26911_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .B(_08279_),
    .S(_08065_),
    .Z(_02435_));
 MUX2_X1 _26912_ (.A(net114),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(_08058_),
    .Z(_08280_));
 MUX2_X1 _26913_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .B(_08280_),
    .S(_08065_),
    .Z(_02436_));
 MUX2_X1 _26914_ (.A(net117),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(_08058_),
    .Z(_08281_));
 MUX2_X1 _26915_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .B(_08281_),
    .S(_08065_),
    .Z(_02437_));
 MUX2_X1 _26916_ (.A(net118),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(_08058_),
    .Z(_08282_));
 MUX2_X1 _26917_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .B(_08282_),
    .S(_08065_),
    .Z(_02438_));
 MUX2_X1 _26918_ (.A(net119),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(_08058_),
    .Z(_08283_));
 MUX2_X1 _26919_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .B(_08283_),
    .S(_08065_),
    .Z(_02439_));
 MUX2_X1 _26920_ (.A(net120),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(_08058_),
    .Z(_08284_));
 MUX2_X1 _26921_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .B(_08284_),
    .S(_08065_),
    .Z(_02440_));
 MUX2_X1 _26922_ (.A(net121),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(_08058_),
    .Z(_08285_));
 MUX2_X1 _26923_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .B(_08285_),
    .S(_08065_),
    .Z(_02441_));
 MUX2_X1 _26924_ (.A(net117),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(_04308_),
    .Z(_08286_));
 MUX2_X1 _26925_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .B(_08286_),
    .S(_08272_),
    .Z(_02442_));
 MUX2_X1 _26926_ (.A(net122),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(_08058_),
    .Z(_08287_));
 MUX2_X1 _26927_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .B(_08287_),
    .S(_08065_),
    .Z(_02443_));
 CLKBUF_X3 _26928_ (.A(_04306_),
    .Z(_08288_));
 MUX2_X1 _26929_ (.A(net123),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(_08288_),
    .Z(_08289_));
 BUF_X4 _26930_ (.A(_08064_),
    .Z(_08290_));
 MUX2_X1 _26931_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .B(_08289_),
    .S(_08290_),
    .Z(_02444_));
 MUX2_X1 _26932_ (.A(net95),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(_08288_),
    .Z(_08291_));
 MUX2_X1 _26933_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .B(_08291_),
    .S(_08290_),
    .Z(_02445_));
 MUX2_X1 _26934_ (.A(net96),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(_08288_),
    .Z(_08292_));
 MUX2_X1 _26935_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .B(_08292_),
    .S(_08290_),
    .Z(_02446_));
 MUX2_X1 _26936_ (.A(net97),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(_08288_),
    .Z(_08293_));
 MUX2_X1 _26937_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .B(_08293_),
    .S(_08290_),
    .Z(_02447_));
 MUX2_X1 _26938_ (.A(net98),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(_08288_),
    .Z(_08294_));
 MUX2_X1 _26939_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .B(_08294_),
    .S(_08290_),
    .Z(_02448_));
 MUX2_X1 _26940_ (.A(net99),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(_08288_),
    .Z(_08295_));
 MUX2_X1 _26941_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .B(_08295_),
    .S(_08290_),
    .Z(_02449_));
 MUX2_X1 _26942_ (.A(net100),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(_08288_),
    .Z(_08296_));
 MUX2_X1 _26943_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .B(_08296_),
    .S(_08290_),
    .Z(_02450_));
 MUX2_X1 _26944_ (.A(_04110_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(_08288_),
    .Z(_08297_));
 MUX2_X1 _26945_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .B(_08297_),
    .S(_08290_),
    .Z(_02451_));
 MUX2_X1 _26946_ (.A(_04109_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(_08288_),
    .Z(_08298_));
 MUX2_X1 _26947_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .B(_08298_),
    .S(_08290_),
    .Z(_02452_));
 MUX2_X1 _26948_ (.A(net118),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(_04307_),
    .Z(_08299_));
 MUX2_X1 _26949_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .B(_08299_),
    .S(_08272_),
    .Z(_02453_));
 MUX2_X1 _26950_ (.A(net101),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(_08288_),
    .Z(_08300_));
 MUX2_X1 _26951_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .B(_08300_),
    .S(_08290_),
    .Z(_02454_));
 CLKBUF_X3 _26952_ (.A(_04306_),
    .Z(_08301_));
 MUX2_X1 _26953_ (.A(net102),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(_08301_),
    .Z(_08302_));
 BUF_X4 _26954_ (.A(_08064_),
    .Z(_08303_));
 MUX2_X1 _26955_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .B(_08302_),
    .S(_08303_),
    .Z(_02455_));
 MUX2_X1 _26956_ (.A(net104),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(_08301_),
    .Z(_08304_));
 MUX2_X1 _26957_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .B(_08304_),
    .S(_08303_),
    .Z(_02456_));
 MUX2_X1 _26958_ (.A(net105),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(_08301_),
    .Z(_08305_));
 MUX2_X1 _26959_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .B(_08305_),
    .S(_08303_),
    .Z(_02457_));
 MUX2_X1 _26960_ (.A(net106),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(_08301_),
    .Z(_08306_));
 MUX2_X1 _26961_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .B(_08306_),
    .S(_08303_),
    .Z(_02458_));
 MUX2_X1 _26962_ (.A(net107),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(_08301_),
    .Z(_08307_));
 MUX2_X1 _26963_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .B(_08307_),
    .S(_08303_),
    .Z(_02459_));
 MUX2_X1 _26964_ (.A(net108),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(_08301_),
    .Z(_08308_));
 MUX2_X1 _26965_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .B(_08308_),
    .S(_08303_),
    .Z(_02460_));
 MUX2_X1 _26966_ (.A(net109),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(_08301_),
    .Z(_08309_));
 MUX2_X1 _26967_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .B(_08309_),
    .S(_08303_),
    .Z(_02461_));
 MUX2_X1 _26968_ (.A(net110),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(_08301_),
    .Z(_08310_));
 MUX2_X1 _26969_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .B(_08310_),
    .S(_08303_),
    .Z(_02462_));
 MUX2_X1 _26970_ (.A(net111),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(_08301_),
    .Z(_08311_));
 MUX2_X1 _26971_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .B(_08311_),
    .S(_08303_),
    .Z(_02463_));
 MUX2_X1 _26972_ (.A(net119),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(_04307_),
    .Z(_08312_));
 MUX2_X1 _26973_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .B(_08312_),
    .S(_08272_),
    .Z(_02464_));
 MUX2_X1 _26974_ (.A(net112),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(_08301_),
    .Z(_08313_));
 MUX2_X1 _26975_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .B(_08313_),
    .S(_08303_),
    .Z(_02465_));
 MUX2_X1 _26976_ (.A(net113),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(_04306_),
    .Z(_08314_));
 MUX2_X1 _26977_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .B(_08314_),
    .S(_08064_),
    .Z(_02466_));
 MUX2_X1 _26978_ (.A(net115),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(_04306_),
    .Z(_08315_));
 MUX2_X1 _26979_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .B(_08315_),
    .S(_08064_),
    .Z(_02467_));
 MUX2_X1 _26980_ (.A(net116),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(_04306_),
    .Z(_08316_));
 MUX2_X1 _26981_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .B(_08316_),
    .S(_08064_),
    .Z(_02468_));
 MUX2_X1 _26982_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .B(net94),
    .S(_08067_),
    .Z(_02469_));
 MUX2_X1 _26983_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .B(net103),
    .S(_08067_),
    .Z(_02470_));
 MUX2_X1 _26984_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .B(net114),
    .S(_08067_),
    .Z(_02471_));
 MUX2_X1 _26985_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .B(net117),
    .S(_08067_),
    .Z(_02472_));
 MUX2_X1 _26986_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .B(net118),
    .S(_08067_),
    .Z(_02473_));
 MUX2_X1 _26987_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .B(net119),
    .S(_08067_),
    .Z(_02474_));
 MUX2_X1 _26988_ (.A(net120),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(_04308_),
    .Z(_08317_));
 MUX2_X1 _26989_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .B(_08317_),
    .S(_08272_),
    .Z(_02475_));
 MUX2_X1 _26990_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .B(net120),
    .S(_08067_),
    .Z(_02476_));
 MUX2_X1 _26991_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .B(net121),
    .S(_08067_),
    .Z(_02477_));
 MUX2_X1 _26992_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .B(net122),
    .S(_08067_),
    .Z(_02478_));
 CLKBUF_X3 _26993_ (.A(_08066_),
    .Z(_08318_));
 MUX2_X1 _26994_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .B(net123),
    .S(_08318_),
    .Z(_02479_));
 MUX2_X1 _26995_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .B(net95),
    .S(_08318_),
    .Z(_02480_));
 MUX2_X1 _26996_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .B(net96),
    .S(_08318_),
    .Z(_02481_));
 MUX2_X1 _26997_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .B(net97),
    .S(_08318_),
    .Z(_02482_));
 MUX2_X1 _26998_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .B(net98),
    .S(_08318_),
    .Z(_02483_));
 MUX2_X1 _26999_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .B(net99),
    .S(_08318_),
    .Z(_02484_));
 MUX2_X1 _27000_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .B(net100),
    .S(_08318_),
    .Z(_02485_));
 MUX2_X1 _27001_ (.A(net121),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(_04307_),
    .Z(_08319_));
 MUX2_X1 _27002_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .B(_08319_),
    .S(_08056_),
    .Z(_02486_));
 MUX2_X1 _27003_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .B(_04110_),
    .S(_08318_),
    .Z(_02487_));
 MUX2_X1 _27004_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .B(_04109_),
    .S(_08318_),
    .Z(_02488_));
 MUX2_X1 _27005_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .B(net101),
    .S(_08318_),
    .Z(_02489_));
 CLKBUF_X3 _27006_ (.A(_08066_),
    .Z(_08320_));
 MUX2_X1 _27007_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .B(net102),
    .S(_08320_),
    .Z(_02490_));
 MUX2_X1 _27008_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .B(net104),
    .S(_08320_),
    .Z(_02491_));
 MUX2_X1 _27009_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .B(net105),
    .S(_08320_),
    .Z(_02492_));
 MUX2_X1 _27010_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .B(net106),
    .S(_08320_),
    .Z(_02493_));
 MUX2_X1 _27011_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .B(net107),
    .S(_08320_),
    .Z(_02494_));
 MUX2_X1 _27012_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .B(net108),
    .S(_08320_),
    .Z(_02495_));
 MUX2_X1 _27013_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .B(net109),
    .S(_08320_),
    .Z(_02496_));
 MUX2_X1 _27014_ (.A(net122),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(_04307_),
    .Z(_08321_));
 MUX2_X1 _27015_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .B(_08321_),
    .S(_08056_),
    .Z(_02497_));
 MUX2_X1 _27016_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .B(net110),
    .S(_08320_),
    .Z(_02498_));
 MUX2_X1 _27017_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .B(net111),
    .S(_08320_),
    .Z(_02499_));
 MUX2_X1 _27018_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .B(net112),
    .S(_08320_),
    .Z(_02500_));
 MUX2_X1 _27019_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .B(net113),
    .S(_08066_),
    .Z(_02501_));
 MUX2_X1 _27020_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .B(net115),
    .S(_08066_),
    .Z(_02502_));
 MUX2_X1 _27021_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .B(net116),
    .S(_08066_),
    .Z(_02503_));
 MUX2_X1 _27022_ (.A(net123),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(_04307_),
    .Z(_08322_));
 MUX2_X1 _27023_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .B(_08322_),
    .S(_08056_),
    .Z(_02504_));
 INV_X4 _27024_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .ZN(_08323_));
 CLKBUF_X3 _27025_ (.A(_08323_),
    .Z(_08324_));
 MUX2_X1 _27026_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .B(_07723_),
    .S(_08324_),
    .Z(net215));
 NOR2_X2 _27027_ (.A1(net93),
    .A2(_04313_),
    .ZN(_08325_));
 CLKBUF_X3 _27028_ (.A(_08325_),
    .Z(_08326_));
 MUX2_X1 _27029_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .B(net215),
    .S(_08326_),
    .Z(_02505_));
 MUX2_X1 _27030_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .B(_07787_),
    .S(_08324_),
    .Z(net216));
 MUX2_X1 _27031_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .B(net216),
    .S(_08326_),
    .Z(_02506_));
 MUX2_X1 _27032_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .B(_07801_),
    .S(_08324_),
    .Z(net217));
 MUX2_X1 _27033_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .B(net217),
    .S(_08326_),
    .Z(_02507_));
 MUX2_X1 _27034_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .B(_07811_),
    .S(_08324_),
    .Z(net218));
 MUX2_X1 _27035_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .B(net218),
    .S(_08326_),
    .Z(_02508_));
 MUX2_X1 _27036_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .B(_07820_),
    .S(_08324_),
    .Z(net219));
 MUX2_X1 _27037_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .B(net219),
    .S(_08326_),
    .Z(_02509_));
 MUX2_X1 _27038_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .B(_07831_),
    .S(_08324_),
    .Z(net220));
 MUX2_X1 _27039_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .B(net220),
    .S(_08326_),
    .Z(_02510_));
 CLKBUF_X3 _27040_ (.A(_08323_),
    .Z(_08327_));
 MUX2_X1 _27041_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .B(_07854_),
    .S(_08327_),
    .Z(net221));
 MUX2_X1 _27042_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .B(net221),
    .S(_08326_),
    .Z(_02511_));
 MUX2_X1 _27043_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .B(_07853_),
    .S(_08327_),
    .Z(net222));
 MUX2_X1 _27044_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .B(net222),
    .S(_08326_),
    .Z(_02512_));
 MUX2_X1 _27045_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .B(_07878_),
    .S(_08327_),
    .Z(net223));
 MUX2_X1 _27046_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .B(net223),
    .S(_08326_),
    .Z(_02513_));
 MUX2_X1 _27047_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .B(_07877_),
    .S(_08327_),
    .Z(net224));
 MUX2_X1 _27048_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .B(net224),
    .S(_08326_),
    .Z(_02514_));
 CLKBUF_X3 _27049_ (.A(_08323_),
    .Z(_08328_));
 NOR2_X1 _27050_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .A2(_08328_),
    .ZN(_08329_));
 AOI21_X1 _27051_ (.A(_08329_),
    .B1(_07890_),
    .B2(_08328_),
    .ZN(net225));
 CLKBUF_X3 _27052_ (.A(_08325_),
    .Z(_08330_));
 MUX2_X1 _27053_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .B(net225),
    .S(_08330_),
    .Z(_02515_));
 MUX2_X1 _27054_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .B(_07901_),
    .S(_08327_),
    .Z(net226));
 MUX2_X1 _27055_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .B(net226),
    .S(_08330_),
    .Z(_02516_));
 MUX2_X1 _27056_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .B(_07911_),
    .S(_08327_),
    .Z(net227));
 MUX2_X1 _27057_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .B(net227),
    .S(_08330_),
    .Z(_02517_));
 MUX2_X1 _27058_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .B(_07920_),
    .S(_08327_),
    .Z(net228));
 MUX2_X1 _27059_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .B(net228),
    .S(_08330_),
    .Z(_02518_));
 MUX2_X1 _27060_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .B(_07944_),
    .S(_08327_),
    .Z(net229));
 MUX2_X1 _27061_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .B(net229),
    .S(_08330_),
    .Z(_02519_));
 NOR2_X1 _27062_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .A2(_08328_),
    .ZN(_08331_));
 AOI21_X1 _27063_ (.A(_08331_),
    .B1(_07943_),
    .B2(_08328_),
    .ZN(net230));
 MUX2_X1 _27064_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .B(net230),
    .S(_08330_),
    .Z(_02520_));
 NOR2_X1 _27065_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .A2(_08328_),
    .ZN(_08332_));
 AOI21_X1 _27066_ (.A(_08332_),
    .B1(_07950_),
    .B2(_08328_),
    .ZN(net231));
 MUX2_X1 _27067_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .B(net231),
    .S(_08330_),
    .Z(_02521_));
 NOR2_X1 _27068_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .A2(_08324_),
    .ZN(_08333_));
 AOI21_X2 _27069_ (.A(_08333_),
    .B1(_07962_),
    .B2(_08328_),
    .ZN(net232));
 MUX2_X1 _27070_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .B(net232),
    .S(_08330_),
    .Z(_02522_));
 MUX2_X1 _27071_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .B(_07981_),
    .S(_08327_),
    .Z(net233));
 MUX2_X1 _27072_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .B(net233),
    .S(_08330_),
    .Z(_02523_));
 NAND2_X1 _27073_ (.A1(_07988_),
    .A2(_07980_),
    .ZN(_08334_));
 MUX2_X1 _27074_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .B(_08334_),
    .S(_08327_),
    .Z(net234));
 MUX2_X1 _27075_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .B(net234),
    .S(_08330_),
    .Z(_02524_));
 MUX2_X1 _27076_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .B(_16510_),
    .S(_08323_),
    .Z(net235));
 CLKBUF_X3 _27077_ (.A(_08325_),
    .Z(_08335_));
 MUX2_X1 _27078_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .B(net235),
    .S(_08335_),
    .Z(_02525_));
 MUX2_X1 _27079_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .B(_07998_),
    .S(_08323_),
    .Z(net236));
 MUX2_X1 _27080_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .B(net236),
    .S(_08335_),
    .Z(_02526_));
 MUX2_X1 _27081_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .B(_08008_),
    .S(_08323_),
    .Z(net237));
 MUX2_X1 _27082_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .B(net237),
    .S(_08335_),
    .Z(_02527_));
 MUX2_X1 _27083_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .B(_16512_),
    .S(_08323_),
    .Z(net238));
 MUX2_X1 _27084_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .B(net238),
    .S(_08335_),
    .Z(_02528_));
 MUX2_X1 _27085_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .B(_08012_),
    .S(_08323_),
    .Z(net239));
 MUX2_X1 _27086_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .B(net239),
    .S(_08335_),
    .Z(_02529_));
 NOR2_X1 _27087_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .A2(_08324_),
    .ZN(_08336_));
 AOI21_X1 _27088_ (.A(_08336_),
    .B1(_07733_),
    .B2(_08328_),
    .ZN(net240));
 MUX2_X1 _27089_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .B(net240),
    .S(_08335_),
    .Z(_02530_));
 MUX2_X1 _27090_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .B(_07749_),
    .S(_08323_),
    .Z(net241));
 MUX2_X1 _27091_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .B(net241),
    .S(_08335_),
    .Z(_02531_));
 MUX2_X1 _27092_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .B(_07755_),
    .S(_08323_),
    .Z(net242));
 MUX2_X1 _27093_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .B(net242),
    .S(_08335_),
    .Z(_02532_));
 NOR2_X1 _27094_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .A2(_08324_),
    .ZN(_08337_));
 AOI21_X1 _27095_ (.A(_08337_),
    .B1(_08025_),
    .B2(_08328_),
    .ZN(net243));
 MUX2_X1 _27096_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .B(net243),
    .S(_08335_),
    .Z(_02533_));
 NOR2_X1 _27097_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .A2(_08324_),
    .ZN(_08338_));
 AOI21_X1 _27098_ (.A(_08338_),
    .B1(_07765_),
    .B2(_08328_),
    .ZN(net244));
 MUX2_X1 _27099_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .B(net244),
    .S(_08335_),
    .Z(_02534_));
 NOR2_X2 _27100_ (.A1(_10771_),
    .A2(_05407_),
    .ZN(_08339_));
 NAND2_X1 _27101_ (.A1(_10770_),
    .A2(_08339_),
    .ZN(_08340_));
 NOR2_X2 _27102_ (.A1(net33),
    .A2(_08340_),
    .ZN(_08341_));
 NAND3_X2 _27103_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_03525_),
    .A3(_08341_),
    .ZN(_08342_));
 NAND3_X4 _27104_ (.A1(_10796_),
    .A2(_03739_),
    .A3(_04006_),
    .ZN(_08343_));
 NOR2_X2 _27105_ (.A1(_03524_),
    .A2(_08343_),
    .ZN(_08344_));
 AOI21_X1 _27106_ (.A(_10772_),
    .B1(_03524_),
    .B2(\load_store_unit_i.lsu_err_q ),
    .ZN(_08345_));
 NOR2_X1 _27107_ (.A1(_08344_),
    .A2(_08345_),
    .ZN(_08346_));
 INV_X1 _27108_ (.A(_08346_),
    .ZN(_08347_));
 AOI21_X2 _27109_ (.A(_08341_),
    .B1(_08347_),
    .B2(_10768_),
    .ZN(_08348_));
 BUF_X2 _27110_ (.A(data_gnt_i),
    .Z(_08349_));
 INV_X1 _27111_ (.A(_08349_),
    .ZN(_08350_));
 OAI21_X4 _27112_ (.A(_08342_),
    .B1(_08348_),
    .B2(_08350_),
    .ZN(_08351_));
 CLKBUF_X3 _27113_ (.A(_08351_),
    .Z(_08352_));
 MUX2_X1 _27114_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .B(_03786_),
    .S(_08352_),
    .Z(_02618_));
 MUX2_X1 _27115_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .B(\alu_adder_result_ex[10] ),
    .S(_08352_),
    .Z(_02619_));
 MUX2_X1 _27116_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .B(net486),
    .S(_08352_),
    .Z(_02620_));
 MUX2_X1 _27117_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .B(\alu_adder_result_ex[12] ),
    .S(_08352_),
    .Z(_02621_));
 MUX2_X1 _27118_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .B(\alu_adder_result_ex[13] ),
    .S(_08352_),
    .Z(_02622_));
 MUX2_X1 _27119_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .B(\alu_adder_result_ex[14] ),
    .S(_08352_),
    .Z(_02623_));
 MUX2_X1 _27120_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .B(\alu_adder_result_ex[15] ),
    .S(_08352_),
    .Z(_02624_));
 MUX2_X1 _27121_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .B(\alu_adder_result_ex[16] ),
    .S(_08352_),
    .Z(_02625_));
 MUX2_X1 _27122_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .B(\alu_adder_result_ex[17] ),
    .S(_08352_),
    .Z(_02626_));
 MUX2_X1 _27123_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .B(\alu_adder_result_ex[18] ),
    .S(_08352_),
    .Z(_02627_));
 CLKBUF_X3 _27124_ (.A(_08351_),
    .Z(_08353_));
 MUX2_X1 _27125_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .B(\alu_adder_result_ex[19] ),
    .S(_08353_),
    .Z(_02628_));
 MUX2_X1 _27126_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .B(\alu_adder_result_ex[1] ),
    .S(_08353_),
    .Z(_02629_));
 MUX2_X1 _27127_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .B(\alu_adder_result_ex[20] ),
    .S(_08353_),
    .Z(_02630_));
 MUX2_X1 _27128_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .B(\alu_adder_result_ex[21] ),
    .S(_08353_),
    .Z(_02631_));
 MUX2_X1 _27129_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .B(\alu_adder_result_ex[22] ),
    .S(_08353_),
    .Z(_02632_));
 MUX2_X1 _27130_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .B(\alu_adder_result_ex[23] ),
    .S(_08353_),
    .Z(_02633_));
 MUX2_X1 _27131_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .B(\alu_adder_result_ex[24] ),
    .S(_08353_),
    .Z(_02634_));
 MUX2_X1 _27132_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .B(net390),
    .S(_08353_),
    .Z(_02635_));
 MUX2_X1 _27133_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .B(\alu_adder_result_ex[26] ),
    .S(_08353_),
    .Z(_02636_));
 MUX2_X1 _27134_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .B(\alu_adder_result_ex[27] ),
    .S(_08353_),
    .Z(_02637_));
 CLKBUF_X3 _27135_ (.A(_08351_),
    .Z(_08354_));
 MUX2_X1 _27136_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .B(net386),
    .S(_08354_),
    .Z(_02638_));
 MUX2_X1 _27137_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .B(net411),
    .S(_08354_),
    .Z(_02639_));
 MUX2_X1 _27138_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .B(\alu_adder_result_ex[2] ),
    .S(_08354_),
    .Z(_02640_));
 MUX2_X1 _27139_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .B(\alu_adder_result_ex[30] ),
    .S(_08354_),
    .Z(_02641_));
 MUX2_X1 _27140_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .B(net289),
    .S(_08354_),
    .Z(_02642_));
 MUX2_X1 _27141_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .B(\alu_adder_result_ex[3] ),
    .S(_08354_),
    .Z(_02643_));
 MUX2_X1 _27142_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .B(\alu_adder_result_ex[4] ),
    .S(_08354_),
    .Z(_02644_));
 MUX2_X1 _27143_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .B(\alu_adder_result_ex[5] ),
    .S(_08354_),
    .Z(_02645_));
 MUX2_X1 _27144_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .B(\alu_adder_result_ex[6] ),
    .S(_08354_),
    .Z(_02646_));
 MUX2_X1 _27145_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .B(\alu_adder_result_ex[7] ),
    .S(_08354_),
    .Z(_02647_));
 MUX2_X1 _27146_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .B(\alu_adder_result_ex[8] ),
    .S(_08351_),
    .Z(_02648_));
 MUX2_X1 _27147_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .B(\alu_adder_result_ex[9] ),
    .S(_08351_),
    .Z(_02649_));
 NOR3_X1 _27148_ (.A1(_10785_),
    .A2(_10924_),
    .A3(_07204_),
    .ZN(_08355_));
 NOR2_X1 _27149_ (.A1(_03523_),
    .A2(_08350_),
    .ZN(_08356_));
 OAI21_X4 _27150_ (.A(_08356_),
    .B1(_08344_),
    .B2(_10771_),
    .ZN(_08357_));
 MUX2_X1 _27151_ (.A(_08355_),
    .B(\load_store_unit_i.data_sign_ext_q ),
    .S(_08357_),
    .Z(_02650_));
 NOR2_X4 _27152_ (.A1(_10821_),
    .A2(_03537_),
    .ZN(net214));
 MUX2_X1 _27153_ (.A(net214),
    .B(\load_store_unit_i.data_we_q ),
    .S(_08357_),
    .Z(_02651_));
 CLKBUF_X2 _27154_ (.A(_16496_),
    .Z(_08358_));
 NOR2_X4 _27155_ (.A1(_10882_),
    .A2(_07204_),
    .ZN(_08359_));
 NAND3_X1 _27156_ (.A1(_10828_),
    .A2(_08358_),
    .A3(_08359_),
    .ZN(_08360_));
 OAI21_X2 _27157_ (.A(_08360_),
    .B1(_08359_),
    .B2(_03704_),
    .ZN(_08361_));
 AOI21_X1 _27158_ (.A(_08361_),
    .B1(_03526_),
    .B2(_10768_),
    .ZN(_08362_));
 AOI21_X1 _27159_ (.A(_10816_),
    .B1(_08339_),
    .B2(_08350_),
    .ZN(_08363_));
 NOR2_X1 _27160_ (.A1(_08362_),
    .A2(_08363_),
    .ZN(_08364_));
 NOR2_X2 _27161_ (.A1(_07204_),
    .A2(_07225_),
    .ZN(_08365_));
 OAI21_X1 _27162_ (.A(_08349_),
    .B1(_08365_),
    .B2(_10771_),
    .ZN(_08366_));
 OAI21_X1 _27163_ (.A(_03524_),
    .B1(_08349_),
    .B2(_08339_),
    .ZN(_08367_));
 AOI21_X1 _27164_ (.A(_03523_),
    .B1(_08366_),
    .B2(_08367_),
    .ZN(_08368_));
 MUX2_X1 _27165_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B(_08364_),
    .S(_08368_),
    .Z(_02652_));
 NAND2_X1 _27166_ (.A1(_03524_),
    .A2(_05407_),
    .ZN(_08369_));
 INV_X1 _27167_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .ZN(_08370_));
 AOI21_X1 _27168_ (.A(_10771_),
    .B1(_03524_),
    .B2(_05407_),
    .ZN(_08371_));
 OAI33_X1 _27169_ (.A1(_08370_),
    .A2(net59),
    .A3(_03526_),
    .B1(_08371_),
    .B2(_08349_),
    .B3(_03523_),
    .ZN(_08372_));
 AOI21_X2 _27170_ (.A(_08372_),
    .B1(_08343_),
    .B2(_03527_),
    .ZN(_08373_));
 AOI21_X1 _27171_ (.A(_10771_),
    .B1(_08369_),
    .B2(_08373_),
    .ZN(_08374_));
 NOR3_X1 _27172_ (.A1(_03523_),
    .A2(_08349_),
    .A3(_08374_),
    .ZN(_02653_));
 AOI21_X1 _27173_ (.A(_10771_),
    .B1(_08349_),
    .B2(_08361_),
    .ZN(_08375_));
 NOR2_X1 _27174_ (.A1(_03524_),
    .A2(_08361_),
    .ZN(_08376_));
 AOI21_X1 _27175_ (.A(_08376_),
    .B1(_08339_),
    .B2(_03524_),
    .ZN(_08377_));
 OAI22_X1 _27176_ (.A1(_03524_),
    .A2(_08375_),
    .B1(_08377_),
    .B2(_08349_),
    .ZN(_08378_));
 NAND3_X1 _27177_ (.A1(_10768_),
    .A2(_08373_),
    .A3(_08378_),
    .ZN(_08379_));
 INV_X1 _27178_ (.A(_03524_),
    .ZN(_08380_));
 OAI21_X1 _27179_ (.A(_08379_),
    .B1(_08373_),
    .B2(_08380_),
    .ZN(_02654_));
 NOR3_X1 _27180_ (.A1(_10771_),
    .A2(net59),
    .A3(_10816_),
    .ZN(_08381_));
 MUX2_X1 _27181_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(_08381_),
    .S(_08373_),
    .Z(_02655_));
 NAND2_X1 _27182_ (.A1(_03527_),
    .A2(_08343_),
    .ZN(_08382_));
 AOI21_X1 _27183_ (.A(\load_store_unit_i.lsu_err_q ),
    .B1(_03527_),
    .B2(_08370_),
    .ZN(_08383_));
 NAND3_X1 _27184_ (.A1(_10772_),
    .A2(net33),
    .A3(_10770_),
    .ZN(_08384_));
 NAND3_X1 _27185_ (.A1(_08370_),
    .A2(_08384_),
    .A3(_08365_),
    .ZN(_08385_));
 OAI21_X1 _27186_ (.A(_08385_),
    .B1(_08365_),
    .B2(\load_store_unit_i.lsu_err_q ),
    .ZN(_08386_));
 AOI222_X2 _27187_ (.A1(_08341_),
    .A2(_08382_),
    .B1(_08383_),
    .B2(_08340_),
    .C1(_03527_),
    .C2(_08386_),
    .ZN(_02656_));
 MUX2_X1 _27188_ (.A(_03786_),
    .B(_05361_),
    .S(_08357_),
    .Z(_02657_));
 MUX2_X1 _27189_ (.A(\alu_adder_result_ex[1] ),
    .B(_05387_),
    .S(_08357_),
    .Z(_02658_));
 OR2_X1 _27190_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_08340_),
    .ZN(_08387_));
 CLKBUF_X3 _27191_ (.A(_08387_),
    .Z(_08388_));
 BUF_X4 _27192_ (.A(_08388_),
    .Z(_08389_));
 MUX2_X1 _27193_ (.A(_05374_),
    .B(\load_store_unit_i.rdata_q[8] ),
    .S(_08389_),
    .Z(_02659_));
 MUX2_X1 _27194_ (.A(net38),
    .B(\load_store_unit_i.rdata_q[18] ),
    .S(_08389_),
    .Z(_02660_));
 MUX2_X1 _27195_ (.A(net39),
    .B(\load_store_unit_i.rdata_q[19] ),
    .S(_08389_),
    .Z(_02661_));
 MUX2_X1 _27196_ (.A(net41),
    .B(\load_store_unit_i.rdata_q[20] ),
    .S(_08389_),
    .Z(_02662_));
 MUX2_X1 _27197_ (.A(net42),
    .B(\load_store_unit_i.rdata_q[21] ),
    .S(_08389_),
    .Z(_02663_));
 MUX2_X1 _27198_ (.A(net43),
    .B(\load_store_unit_i.rdata_q[22] ),
    .S(_08389_),
    .Z(_02664_));
 MUX2_X1 _27199_ (.A(net44),
    .B(\load_store_unit_i.rdata_q[23] ),
    .S(_08389_),
    .Z(_02665_));
 MUX2_X1 _27200_ (.A(net45),
    .B(\load_store_unit_i.rdata_q[24] ),
    .S(_08389_),
    .Z(_02666_));
 MUX2_X1 _27201_ (.A(net46),
    .B(\load_store_unit_i.rdata_q[25] ),
    .S(_08389_),
    .Z(_02667_));
 MUX2_X1 _27202_ (.A(net47),
    .B(\load_store_unit_i.rdata_q[26] ),
    .S(_08389_),
    .Z(_02668_));
 BUF_X4 _27203_ (.A(_08388_),
    .Z(_08390_));
 MUX2_X1 _27204_ (.A(net48),
    .B(\load_store_unit_i.rdata_q[27] ),
    .S(_08390_),
    .Z(_02669_));
 MUX2_X1 _27205_ (.A(_05808_),
    .B(\load_store_unit_i.rdata_q[9] ),
    .S(_08390_),
    .Z(_02670_));
 MUX2_X1 _27206_ (.A(net49),
    .B(\load_store_unit_i.rdata_q[28] ),
    .S(_08390_),
    .Z(_02671_));
 MUX2_X1 _27207_ (.A(net50),
    .B(\load_store_unit_i.rdata_q[29] ),
    .S(_08390_),
    .Z(_02672_));
 MUX2_X1 _27208_ (.A(net52),
    .B(\load_store_unit_i.rdata_q[30] ),
    .S(_08390_),
    .Z(_02673_));
 MUX2_X1 _27209_ (.A(net53),
    .B(\load_store_unit_i.rdata_q[31] ),
    .S(_08390_),
    .Z(_02674_));
 MUX2_X1 _27210_ (.A(_05821_),
    .B(\load_store_unit_i.rdata_q[10] ),
    .S(_08390_),
    .Z(_02675_));
 MUX2_X1 _27211_ (.A(_05900_),
    .B(\load_store_unit_i.rdata_q[11] ),
    .S(_08390_),
    .Z(_02676_));
 MUX2_X1 _27212_ (.A(_05419_),
    .B(\load_store_unit_i.rdata_q[12] ),
    .S(_08390_),
    .Z(_02677_));
 MUX2_X1 _27213_ (.A(_05500_),
    .B(\load_store_unit_i.rdata_q[13] ),
    .S(_08390_),
    .Z(_02678_));
 MUX2_X1 _27214_ (.A(net35),
    .B(\load_store_unit_i.rdata_q[14] ),
    .S(_08388_),
    .Z(_02679_));
 MUX2_X1 _27215_ (.A(_05674_),
    .B(\load_store_unit_i.rdata_q[15] ),
    .S(_08388_),
    .Z(_02680_));
 MUX2_X1 _27216_ (.A(net36),
    .B(\load_store_unit_i.rdata_q[16] ),
    .S(_08388_),
    .Z(_02681_));
 MUX2_X1 _27217_ (.A(net37),
    .B(\load_store_unit_i.rdata_q[17] ),
    .S(_08388_),
    .Z(_02682_));
 MUX2_X1 _27218_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .S(_03775_),
    .Z(_02683_));
 MUX2_X1 _27219_ (.A(_03752_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .S(_03775_),
    .Z(_02684_));
 MUX2_X1 _27220_ (.A(_03744_),
    .B(_03781_),
    .S(_03702_),
    .Z(_02685_));
 MUX2_X1 _27221_ (.A(_03683_),
    .B(_03734_),
    .S(_03689_),
    .Z(_02686_));
 MUX2_X1 _27222_ (.A(_03701_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .S(_03689_),
    .Z(_02687_));
 NOR2_X1 _27223_ (.A1(_10939_),
    .A2(_07204_),
    .ZN(_08391_));
 MUX2_X1 _27224_ (.A(_08391_),
    .B(_05363_),
    .S(_08357_),
    .Z(_02688_));
 NAND2_X1 _27225_ (.A1(_05379_),
    .A2(_08357_),
    .ZN(_08392_));
 NAND2_X1 _27226_ (.A1(_10967_),
    .A2(_04006_),
    .ZN(_08393_));
 OAI21_X1 _27227_ (.A(_08392_),
    .B1(_08393_),
    .B2(_08357_),
    .ZN(_02689_));
 MUX2_X1 _27228_ (.A(_11772_),
    .B(_04465_),
    .S(_16239_),
    .Z(_08394_));
 NOR2_X1 _27229_ (.A1(_04469_),
    .A2(_08394_),
    .ZN(_08395_));
 AOI21_X4 _27230_ (.A(_08395_),
    .B1(_05356_),
    .B2(_16239_),
    .ZN(_08396_));
 NAND3_X1 _27231_ (.A1(_16274_),
    .A2(_15908_),
    .A3(_04455_),
    .ZN(_08397_));
 NOR2_X1 _27232_ (.A1(_08397_),
    .A2(_04542_),
    .ZN(_08398_));
 MUX2_X1 _27233_ (.A(\cs_registers_i.mcountinhibit[0] ),
    .B(_08396_),
    .S(_08398_),
    .Z(_02690_));
 MUX2_X1 _27234_ (.A(_04465_),
    .B(_11772_),
    .S(_16254_),
    .Z(_08399_));
 NOR2_X1 _27235_ (.A1(_04469_),
    .A2(_08399_),
    .ZN(_08400_));
 AOI21_X4 _27236_ (.A(_08400_),
    .B1(_06563_),
    .B2(_16258_),
    .ZN(_08401_));
 BUF_X4 _27237_ (.A(_08401_),
    .Z(_08402_));
 MUX2_X1 _27238_ (.A(\cs_registers_i.mcountinhibit[2] ),
    .B(_08402_),
    .S(_08398_),
    .Z(_02691_));
 NAND2_X1 _27239_ (.A1(_04380_),
    .A2(_04608_),
    .ZN(_08403_));
 NOR2_X2 _27240_ (.A1(_03631_),
    .A2(_03603_),
    .ZN(_08404_));
 XNOR2_X1 _27241_ (.A(_03576_),
    .B(_08404_),
    .ZN(_08405_));
 AND4_X1 _27242_ (.A1(_15911_),
    .A2(_15915_),
    .A3(_15919_),
    .A4(_08405_),
    .ZN(_08406_));
 NAND3_X1 _27243_ (.A1(_16266_),
    .A2(_16274_),
    .A3(_05216_),
    .ZN(_08407_));
 NAND2_X1 _27244_ (.A1(_11329_),
    .A2(_08407_),
    .ZN(_08408_));
 AND2_X1 _27245_ (.A1(_08406_),
    .A2(_08408_),
    .ZN(_08409_));
 NAND3_X1 _27246_ (.A1(_08403_),
    .A2(_04490_),
    .A3(_08409_),
    .ZN(_08410_));
 CLKBUF_X3 _27247_ (.A(_08410_),
    .Z(_08411_));
 INV_X2 _27248_ (.A(_08411_),
    .ZN(_08412_));
 MUX2_X1 _27249_ (.A(_00552_),
    .B(_08396_),
    .S(_08412_),
    .Z(_08413_));
 MUX2_X1 _27250_ (.A(_04756_),
    .B(_00554_),
    .S(_08411_),
    .Z(_08414_));
 BUF_X2 _27251_ (.A(_08414_),
    .Z(_08415_));
 CLKBUF_X3 _27252_ (.A(_08415_),
    .Z(_08416_));
 MUX2_X1 _27253_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(_08413_),
    .S(_08416_),
    .Z(_02692_));
 CLKBUF_X3 _27254_ (.A(_08415_),
    .Z(_08417_));
 CLKBUF_X3 _27255_ (.A(_08411_),
    .Z(_08418_));
 NAND2_X2 _27256_ (.A1(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .A2(_15936_),
    .ZN(_08419_));
 NAND3_X2 _27257_ (.A1(_06595_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .ZN(_08420_));
 NOR2_X1 _27258_ (.A1(_08419_),
    .A2(_08420_),
    .ZN(_08421_));
 NAND3_X1 _27259_ (.A1(_05606_),
    .A2(_05693_),
    .A3(_08421_),
    .ZN(_08422_));
 NAND2_X1 _27260_ (.A1(_04931_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .ZN(_08423_));
 OAI21_X1 _27261_ (.A(_08418_),
    .B1(_08422_),
    .B2(_08423_),
    .ZN(_08424_));
 AOI21_X1 _27262_ (.A(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .B1(_08417_),
    .B2(_08424_),
    .ZN(_08425_));
 AND3_X1 _27263_ (.A1(_04931_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .ZN(_08426_));
 AND3_X2 _27264_ (.A1(_04373_),
    .A2(_04378_),
    .A3(_03584_),
    .ZN(_08427_));
 NOR2_X2 _27265_ (.A1(_08427_),
    .A2(_06500_),
    .ZN(_08428_));
 NAND2_X1 _27266_ (.A1(_08406_),
    .A2(_08408_),
    .ZN(_08429_));
 NOR3_X4 _27267_ (.A1(_08428_),
    .A2(_04542_),
    .A3(_08429_),
    .ZN(_08430_));
 BUF_X2 _27268_ (.A(_08430_),
    .Z(_08431_));
 NOR2_X1 _27269_ (.A1(_08431_),
    .A2(_08422_),
    .ZN(_08432_));
 NAND2_X1 _27270_ (.A1(_08426_),
    .A2(_08432_),
    .ZN(_08433_));
 CLKBUF_X3 _27271_ (.A(_08430_),
    .Z(_08434_));
 NAND2_X1 _27272_ (.A1(_16321_),
    .A2(_05840_),
    .ZN(_08435_));
 MUX2_X1 _27273_ (.A(_04642_),
    .B(_04643_),
    .S(_16317_),
    .Z(_08436_));
 OAI21_X4 _27274_ (.A(_08435_),
    .B1(_08436_),
    .B2(_04600_),
    .ZN(_08437_));
 NAND2_X1 _27275_ (.A1(_08434_),
    .A2(_08437_),
    .ZN(_08438_));
 NAND2_X1 _27276_ (.A1(_08433_),
    .A2(_08438_),
    .ZN(_08439_));
 CLKBUF_X3 _27277_ (.A(_08415_),
    .Z(_08440_));
 AOI21_X1 _27278_ (.A(_08425_),
    .B1(_08439_),
    .B2(_08440_),
    .ZN(_02693_));
 INV_X1 _27279_ (.A(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .ZN(_08441_));
 INV_X1 _27280_ (.A(_05606_),
    .ZN(_08442_));
 INV_X1 _27281_ (.A(_05693_),
    .ZN(_08443_));
 NAND3_X2 _27282_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .ZN(_08444_));
 OR2_X1 _27283_ (.A1(_08420_),
    .A2(_08444_),
    .ZN(_08445_));
 NOR3_X2 _27284_ (.A1(_08442_),
    .A2(_08443_),
    .A3(_08445_),
    .ZN(_08446_));
 AND2_X1 _27285_ (.A1(_08426_),
    .A2(_08446_),
    .ZN(_08447_));
 OAI21_X1 _27286_ (.A(_08417_),
    .B1(_08447_),
    .B2(_08412_),
    .ZN(_08448_));
 NAND2_X1 _27287_ (.A1(_04472_),
    .A2(_08431_),
    .ZN(_08449_));
 AND2_X1 _27288_ (.A1(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .A2(_08447_),
    .ZN(_08450_));
 INV_X1 _27289_ (.A(_08450_),
    .ZN(_08451_));
 CLKBUF_X3 _27290_ (.A(_08431_),
    .Z(_08452_));
 OAI21_X1 _27291_ (.A(_08449_),
    .B1(_08451_),
    .B2(_08452_),
    .ZN(_08453_));
 CLKBUF_X3 _27292_ (.A(_08415_),
    .Z(_08454_));
 AOI22_X1 _27293_ (.A1(_08441_),
    .A2(_08448_),
    .B1(_08453_),
    .B2(_08454_),
    .ZN(_02694_));
 INV_X1 _27294_ (.A(_04503_),
    .ZN(_08455_));
 NAND4_X2 _27295_ (.A1(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .A2(_05606_),
    .A3(_05693_),
    .A4(_08426_),
    .ZN(_08456_));
 NOR3_X4 _27296_ (.A1(_08419_),
    .A2(_08420_),
    .A3(_08456_),
    .ZN(_08457_));
 OAI21_X1 _27297_ (.A(_08417_),
    .B1(_08457_),
    .B2(_08412_),
    .ZN(_08458_));
 CLKBUF_X3 _27298_ (.A(_08411_),
    .Z(_08459_));
 NAND3_X1 _27299_ (.A1(_04503_),
    .A2(_08459_),
    .A3(_08457_),
    .ZN(_08460_));
 BUF_X2 _27300_ (.A(_08430_),
    .Z(_08461_));
 NAND2_X1 _27301_ (.A1(_04528_),
    .A2(_08461_),
    .ZN(_08462_));
 NAND2_X1 _27302_ (.A1(_08460_),
    .A2(_08462_),
    .ZN(_08463_));
 AOI22_X1 _27303_ (.A1(_08455_),
    .A2(_08458_),
    .B1(_08463_),
    .B2(_08454_),
    .ZN(_02695_));
 OAI21_X1 _27304_ (.A(_08418_),
    .B1(_08451_),
    .B2(_08455_),
    .ZN(_08464_));
 AOI21_X1 _27305_ (.A(_04549_),
    .B1(_08417_),
    .B2(_08464_),
    .ZN(_08465_));
 NAND2_X1 _27306_ (.A1(_04562_),
    .A2(_08434_),
    .ZN(_08466_));
 NAND3_X1 _27307_ (.A1(_04503_),
    .A2(_04549_),
    .A3(_08450_),
    .ZN(_08467_));
 OAI21_X1 _27308_ (.A(_08466_),
    .B1(_08467_),
    .B2(_08452_),
    .ZN(_08468_));
 AOI21_X1 _27309_ (.A(_08465_),
    .B1(_08468_),
    .B2(_08440_),
    .ZN(_02696_));
 CLKBUF_X3 _27310_ (.A(_08411_),
    .Z(_08469_));
 NAND3_X1 _27311_ (.A1(_04503_),
    .A2(_04549_),
    .A3(_08457_),
    .ZN(_08470_));
 NAND2_X1 _27312_ (.A1(_08469_),
    .A2(_08470_),
    .ZN(_08471_));
 AOI21_X1 _27313_ (.A(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .B1(_08417_),
    .B2(_08471_),
    .ZN(_08472_));
 NAND2_X1 _27314_ (.A1(_04597_),
    .A2(_08434_),
    .ZN(_08473_));
 NAND2_X1 _27315_ (.A1(_04549_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .ZN(_08474_));
 OAI21_X1 _27316_ (.A(_08473_),
    .B1(_08474_),
    .B2(_08460_),
    .ZN(_08475_));
 AOI21_X1 _27317_ (.A(_08472_),
    .B1(_08475_),
    .B2(_08440_),
    .ZN(_02697_));
 INV_X1 _27318_ (.A(_04605_),
    .ZN(_08476_));
 NOR2_X1 _27319_ (.A1(_08455_),
    .A2(_08474_),
    .ZN(_08477_));
 NOR2_X1 _27320_ (.A1(_08445_),
    .A2(_08456_),
    .ZN(_08478_));
 AND2_X1 _27321_ (.A1(_08477_),
    .A2(_08478_),
    .ZN(_08479_));
 OAI21_X1 _27322_ (.A(_08417_),
    .B1(_08479_),
    .B2(_08412_),
    .ZN(_08480_));
 OR3_X2 _27323_ (.A1(_08428_),
    .A2(_04542_),
    .A3(_08429_),
    .ZN(_08481_));
 CLKBUF_X3 _27324_ (.A(_08481_),
    .Z(_08482_));
 NAND3_X1 _27325_ (.A1(_04605_),
    .A2(_08482_),
    .A3(_08479_),
    .ZN(_08483_));
 NAND2_X1 _27326_ (.A1(_04620_),
    .A2(_08431_),
    .ZN(_08484_));
 NAND2_X1 _27327_ (.A1(_08483_),
    .A2(_08484_),
    .ZN(_08485_));
 AOI22_X1 _27328_ (.A1(_08476_),
    .A2(_08480_),
    .B1(_08485_),
    .B2(_08454_),
    .ZN(_02698_));
 NAND3_X2 _27329_ (.A1(_04605_),
    .A2(_08457_),
    .A3(_08477_),
    .ZN(_08486_));
 NAND2_X1 _27330_ (.A1(_08469_),
    .A2(_08486_),
    .ZN(_08487_));
 AOI21_X1 _27331_ (.A(_04626_),
    .B1(_08417_),
    .B2(_08487_),
    .ZN(_08488_));
 INV_X1 _27332_ (.A(_04626_),
    .ZN(_08489_));
 OR3_X1 _27333_ (.A1(_08489_),
    .A2(_08430_),
    .A3(_08486_),
    .ZN(_08490_));
 CLKBUF_X3 _27334_ (.A(_08411_),
    .Z(_08491_));
 NOR2_X1 _27335_ (.A1(_04668_),
    .A2(_04644_),
    .ZN(_08492_));
 AOI21_X4 _27336_ (.A(_08492_),
    .B1(_04640_),
    .B2(_16369_),
    .ZN(_08493_));
 OAI21_X1 _27337_ (.A(_08490_),
    .B1(_08491_),
    .B2(_08493_),
    .ZN(_08494_));
 AOI21_X1 _27338_ (.A(_08488_),
    .B1(_08494_),
    .B2(_08440_),
    .ZN(_02699_));
 NAND3_X1 _27339_ (.A1(_04605_),
    .A2(_04626_),
    .A3(_08479_),
    .ZN(_08495_));
 NAND2_X1 _27340_ (.A1(_08469_),
    .A2(_08495_),
    .ZN(_08496_));
 AOI21_X1 _27341_ (.A(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .B1(_08417_),
    .B2(_08496_),
    .ZN(_08497_));
 NAND2_X1 _27342_ (.A1(_04665_),
    .A2(_08434_),
    .ZN(_08498_));
 NAND2_X2 _27343_ (.A1(_04626_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .ZN(_08499_));
 OAI21_X1 _27344_ (.A(_08498_),
    .B1(_08499_),
    .B2(_08483_),
    .ZN(_08500_));
 AOI21_X1 _27345_ (.A(_08497_),
    .B1(_08500_),
    .B2(_08440_),
    .ZN(_02700_));
 CLKBUF_X3 _27346_ (.A(_08415_),
    .Z(_08501_));
 OAI21_X1 _27347_ (.A(_08418_),
    .B1(_08486_),
    .B2(_08499_),
    .ZN(_08502_));
 AOI21_X1 _27348_ (.A(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .B1(_08501_),
    .B2(_08502_),
    .ZN(_08503_));
 INV_X1 _27349_ (.A(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .ZN(_08504_));
 NOR3_X1 _27350_ (.A1(_08504_),
    .A2(_08486_),
    .A3(_08499_),
    .ZN(_08505_));
 MUX2_X1 _27351_ (.A(_04685_),
    .B(_08505_),
    .S(_08459_),
    .Z(_08506_));
 AOI21_X1 _27352_ (.A(_08503_),
    .B1(_08506_),
    .B2(_08440_),
    .ZN(_02701_));
 NAND2_X1 _27353_ (.A1(_04605_),
    .A2(_08477_),
    .ZN(_08507_));
 NOR3_X2 _27354_ (.A1(_08504_),
    .A2(_08507_),
    .A3(_08499_),
    .ZN(_08508_));
 AND2_X1 _27355_ (.A1(_08478_),
    .A2(_08508_),
    .ZN(_08509_));
 OR2_X1 _27356_ (.A1(_08431_),
    .A2(_08509_),
    .ZN(_08510_));
 AOI21_X1 _27357_ (.A(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .B1(_08501_),
    .B2(_08510_),
    .ZN(_08511_));
 NAND2_X1 _27358_ (.A1(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .A2(_08509_),
    .ZN(_08512_));
 OR2_X1 _27359_ (.A1(_08431_),
    .A2(_08512_),
    .ZN(_08513_));
 NAND2_X1 _27360_ (.A1(_04700_),
    .A2(_08431_),
    .ZN(_08514_));
 NAND2_X1 _27361_ (.A1(_08513_),
    .A2(_08514_),
    .ZN(_08515_));
 AOI21_X1 _27362_ (.A(_08511_),
    .B1(_08515_),
    .B2(_08440_),
    .ZN(_02702_));
 NAND2_X1 _27363_ (.A1(_15937_),
    .A2(_08459_),
    .ZN(_08516_));
 MUX2_X1 _27364_ (.A(_04466_),
    .B(_04467_),
    .S(_16246_),
    .Z(_08517_));
 OAI22_X4 _27365_ (.A1(_16246_),
    .A2(_06507_),
    .B1(_08517_),
    .B2(_04469_),
    .ZN(_08518_));
 BUF_X4 _27366_ (.A(_08518_),
    .Z(_08519_));
 CLKBUF_X3 _27367_ (.A(_08411_),
    .Z(_08520_));
 OAI21_X1 _27368_ (.A(_08516_),
    .B1(_08519_),
    .B2(_08520_),
    .ZN(_08521_));
 MUX2_X1 _27369_ (.A(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .B(_08521_),
    .S(_08415_),
    .Z(_02703_));
 NAND3_X2 _27370_ (.A1(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .A2(_08457_),
    .A3(_08508_),
    .ZN(_08522_));
 NAND2_X1 _27371_ (.A1(_08469_),
    .A2(_08522_),
    .ZN(_08523_));
 AOI21_X1 _27372_ (.A(_04705_),
    .B1(_08501_),
    .B2(_08523_),
    .ZN(_08524_));
 INV_X1 _27373_ (.A(_04705_),
    .ZN(_08525_));
 OR3_X1 _27374_ (.A1(_08525_),
    .A2(_08431_),
    .A3(_08522_),
    .ZN(_08526_));
 NAND2_X1 _27375_ (.A1(_04721_),
    .A2(_08434_),
    .ZN(_08527_));
 NAND2_X1 _27376_ (.A1(_08526_),
    .A2(_08527_),
    .ZN(_08528_));
 AOI21_X1 _27377_ (.A(_08524_),
    .B1(_08528_),
    .B2(_08440_),
    .ZN(_02704_));
 OAI21_X1 _27378_ (.A(_08418_),
    .B1(_08512_),
    .B2(_08525_),
    .ZN(_08529_));
 AOI21_X1 _27379_ (.A(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .B1(_08501_),
    .B2(_08529_),
    .ZN(_08530_));
 NAND2_X1 _27380_ (.A1(_04742_),
    .A2(_08461_),
    .ZN(_08531_));
 NAND2_X1 _27381_ (.A1(_04705_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .ZN(_08532_));
 OAI21_X1 _27382_ (.A(_08531_),
    .B1(_08532_),
    .B2(_08513_),
    .ZN(_08533_));
 AOI21_X1 _27383_ (.A(_08530_),
    .B1(_08533_),
    .B2(_08440_),
    .ZN(_02705_));
 OAI21_X1 _27384_ (.A(_08418_),
    .B1(_08522_),
    .B2(_08532_),
    .ZN(_08534_));
 AOI21_X1 _27385_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .B1(_08501_),
    .B2(_08534_),
    .ZN(_08535_));
 NAND3_X1 _27386_ (.A1(_04705_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .ZN(_08536_));
 NOR2_X1 _27387_ (.A1(_08522_),
    .A2(_08536_),
    .ZN(_08537_));
 MUX2_X1 _27388_ (.A(_04761_),
    .B(_08537_),
    .S(_08459_),
    .Z(_08538_));
 CLKBUF_X3 _27389_ (.A(_08415_),
    .Z(_08539_));
 AOI21_X1 _27390_ (.A(_08535_),
    .B1(_08538_),
    .B2(_08539_),
    .ZN(_02706_));
 INV_X1 _27391_ (.A(_04779_),
    .ZN(_08540_));
 NOR2_X2 _27392_ (.A1(_08512_),
    .A2(_08536_),
    .ZN(_08541_));
 OAI21_X1 _27393_ (.A(_08417_),
    .B1(_08541_),
    .B2(_08412_),
    .ZN(_08542_));
 NAND3_X1 _27394_ (.A1(_04779_),
    .A2(_08482_),
    .A3(_08541_),
    .ZN(_08543_));
 NAND2_X1 _27395_ (.A1(_04783_),
    .A2(_08461_),
    .ZN(_08544_));
 NAND2_X1 _27396_ (.A1(_08543_),
    .A2(_08544_),
    .ZN(_08545_));
 AOI22_X1 _27397_ (.A1(_08540_),
    .A2(_08542_),
    .B1(_08545_),
    .B2(_08454_),
    .ZN(_02707_));
 NAND2_X1 _27398_ (.A1(_04779_),
    .A2(_08537_),
    .ZN(_08546_));
 NAND2_X1 _27399_ (.A1(_08469_),
    .A2(_08546_),
    .ZN(_08547_));
 AOI21_X1 _27400_ (.A(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .B1(_08501_),
    .B2(_08547_),
    .ZN(_08548_));
 AND3_X1 _27401_ (.A1(_04779_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .A3(_08537_),
    .ZN(_08549_));
 NAND2_X1 _27402_ (.A1(_08459_),
    .A2(_08549_),
    .ZN(_08550_));
 NAND2_X1 _27403_ (.A1(_04805_),
    .A2(_08431_),
    .ZN(_08551_));
 NAND2_X1 _27404_ (.A1(_08550_),
    .A2(_08551_),
    .ZN(_08552_));
 AOI21_X1 _27405_ (.A(_08548_),
    .B1(_08552_),
    .B2(_08539_),
    .ZN(_02708_));
 NAND3_X2 _27406_ (.A1(_04779_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .A3(_08541_),
    .ZN(_08553_));
 NAND2_X1 _27407_ (.A1(_08469_),
    .A2(_08553_),
    .ZN(_08554_));
 AOI21_X1 _27408_ (.A(_04815_),
    .B1(_08501_),
    .B2(_08554_),
    .ZN(_08555_));
 NAND2_X1 _27409_ (.A1(_04822_),
    .A2(_08434_),
    .ZN(_08556_));
 OR2_X1 _27410_ (.A1(_08430_),
    .A2(_08553_),
    .ZN(_08557_));
 INV_X1 _27411_ (.A(_04815_),
    .ZN(_08558_));
 OAI21_X1 _27412_ (.A(_08556_),
    .B1(_08557_),
    .B2(_08558_),
    .ZN(_08559_));
 AOI21_X1 _27413_ (.A(_08555_),
    .B1(_08559_),
    .B2(_08539_),
    .ZN(_02709_));
 INV_X2 _27414_ (.A(_08549_),
    .ZN(_08560_));
 OAI21_X1 _27415_ (.A(_08418_),
    .B1(_08560_),
    .B2(_08558_),
    .ZN(_08561_));
 AOI21_X1 _27416_ (.A(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .B1(_08501_),
    .B2(_08561_),
    .ZN(_08562_));
 NAND2_X1 _27417_ (.A1(_04838_),
    .A2(_08434_),
    .ZN(_08563_));
 NAND2_X1 _27418_ (.A1(_04815_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .ZN(_08564_));
 OAI21_X1 _27419_ (.A(_08563_),
    .B1(_08564_),
    .B2(_08550_),
    .ZN(_08565_));
 AOI21_X1 _27420_ (.A(_08562_),
    .B1(_08565_),
    .B2(_08539_),
    .ZN(_02710_));
 OAI21_X1 _27421_ (.A(_08418_),
    .B1(_08553_),
    .B2(_08564_),
    .ZN(_08566_));
 AOI21_X1 _27422_ (.A(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .B1(_08501_),
    .B2(_08566_),
    .ZN(_08567_));
 NAND2_X1 _27423_ (.A1(_04853_),
    .A2(_08461_),
    .ZN(_08568_));
 AND3_X1 _27424_ (.A1(_04815_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .ZN(_08569_));
 INV_X1 _27425_ (.A(_08569_),
    .ZN(_08570_));
 OAI21_X1 _27426_ (.A(_08568_),
    .B1(_08570_),
    .B2(_08557_),
    .ZN(_08571_));
 AOI21_X1 _27427_ (.A(_08567_),
    .B1(_08571_),
    .B2(_08539_),
    .ZN(_02711_));
 OAI21_X1 _27428_ (.A(_08418_),
    .B1(_08560_),
    .B2(_08570_),
    .ZN(_08572_));
 AOI21_X1 _27429_ (.A(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .B1(_08501_),
    .B2(_08572_),
    .ZN(_08573_));
 NAND2_X1 _27430_ (.A1(_04868_),
    .A2(_08461_),
    .ZN(_08574_));
 NAND2_X1 _27431_ (.A1(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .A2(_08569_),
    .ZN(_08575_));
 OAI21_X1 _27432_ (.A(_08574_),
    .B1(_08575_),
    .B2(_08550_),
    .ZN(_08576_));
 AOI21_X1 _27433_ (.A(_08573_),
    .B1(_08576_),
    .B2(_08539_),
    .ZN(_02712_));
 OAI21_X1 _27434_ (.A(_08418_),
    .B1(_08553_),
    .B2(_08575_),
    .ZN(_08577_));
 AOI21_X1 _27435_ (.A(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .B1(_08416_),
    .B2(_08577_),
    .ZN(_08578_));
 NAND2_X1 _27436_ (.A1(_04885_),
    .A2(_08461_),
    .ZN(_08579_));
 AND3_X1 _27437_ (.A1(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .A3(_08569_),
    .ZN(_08580_));
 INV_X1 _27438_ (.A(_08580_),
    .ZN(_08581_));
 OAI21_X1 _27439_ (.A(_08579_),
    .B1(_08581_),
    .B2(_08557_),
    .ZN(_08582_));
 AOI21_X1 _27440_ (.A(_08578_),
    .B1(_08582_),
    .B2(_08539_),
    .ZN(_02713_));
 INV_X1 _27441_ (.A(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .ZN(_08583_));
 OAI21_X1 _27442_ (.A(_08417_),
    .B1(_08452_),
    .B2(_15936_),
    .ZN(_08584_));
 OR2_X1 _27443_ (.A1(_08430_),
    .A2(_08419_),
    .ZN(_08585_));
 OAI21_X1 _27444_ (.A(_08585_),
    .B1(_08491_),
    .B2(_08402_),
    .ZN(_08586_));
 AOI22_X1 _27445_ (.A1(_08583_),
    .A2(_08584_),
    .B1(_08586_),
    .B2(_08454_),
    .ZN(_02714_));
 CLKBUF_X3 _27446_ (.A(_08411_),
    .Z(_08587_));
 OAI21_X1 _27447_ (.A(_08587_),
    .B1(_08560_),
    .B2(_08581_),
    .ZN(_08588_));
 AOI21_X1 _27448_ (.A(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .B1(_08416_),
    .B2(_08588_),
    .ZN(_08589_));
 NAND2_X1 _27449_ (.A1(_04905_),
    .A2(_08461_),
    .ZN(_08590_));
 NAND2_X2 _27450_ (.A1(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .A2(_08580_),
    .ZN(_08591_));
 OAI21_X1 _27451_ (.A(_08590_),
    .B1(_08591_),
    .B2(_08550_),
    .ZN(_08592_));
 AOI21_X1 _27452_ (.A(_08589_),
    .B1(_08592_),
    .B2(_08539_),
    .ZN(_02715_));
 OR2_X2 _27453_ (.A1(_08553_),
    .A2(_08591_),
    .ZN(_08593_));
 NAND2_X1 _27454_ (.A1(_08469_),
    .A2(_08593_),
    .ZN(_08594_));
 AOI21_X1 _27455_ (.A(_04911_),
    .B1(_08416_),
    .B2(_08594_),
    .ZN(_08595_));
 NAND2_X1 _27456_ (.A1(_04924_),
    .A2(_08461_),
    .ZN(_08596_));
 OR2_X1 _27457_ (.A1(_08430_),
    .A2(_08593_),
    .ZN(_08597_));
 INV_X1 _27458_ (.A(_04911_),
    .ZN(_08598_));
 OAI21_X1 _27459_ (.A(_08596_),
    .B1(_08597_),
    .B2(_08598_),
    .ZN(_08599_));
 AOI21_X1 _27460_ (.A(_08595_),
    .B1(_08599_),
    .B2(_08539_),
    .ZN(_02716_));
 NAND2_X1 _27461_ (.A1(_04490_),
    .A2(_08409_),
    .ZN(_08600_));
 OAI21_X1 _27462_ (.A(_00554_),
    .B1(_04629_),
    .B2(_08600_),
    .ZN(_08601_));
 OAI21_X1 _27463_ (.A(_08601_),
    .B1(_08600_),
    .B2(_04756_),
    .ZN(_08602_));
 CLKBUF_X3 _27464_ (.A(_08602_),
    .Z(_08603_));
 CLKBUF_X3 _27465_ (.A(_08603_),
    .Z(_08604_));
 NOR2_X2 _27466_ (.A1(_08560_),
    .A2(_08591_),
    .ZN(_08605_));
 NAND2_X1 _27467_ (.A1(_04911_),
    .A2(_08605_),
    .ZN(_08606_));
 NAND2_X1 _27468_ (.A1(_08469_),
    .A2(_08606_),
    .ZN(_08607_));
 AOI21_X1 _27469_ (.A(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .B1(_08604_),
    .B2(_08607_),
    .ZN(_08608_));
 NAND2_X1 _27470_ (.A1(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .A2(_04911_),
    .ZN(_08609_));
 NAND2_X1 _27471_ (.A1(_08459_),
    .A2(_08605_),
    .ZN(_08610_));
 OAI22_X1 _27472_ (.A1(_08396_),
    .A2(_08491_),
    .B1(_08609_),
    .B2(_08610_),
    .ZN(_08611_));
 CLKBUF_X3 _27473_ (.A(_08603_),
    .Z(_08612_));
 AOI21_X1 _27474_ (.A(_08608_),
    .B1(_08611_),
    .B2(_08612_),
    .ZN(_02717_));
 OAI21_X1 _27475_ (.A(_08587_),
    .B1(_08593_),
    .B2(_08609_),
    .ZN(_08613_));
 AOI21_X1 _27476_ (.A(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .B1(_08604_),
    .B2(_08613_),
    .ZN(_08614_));
 NAND2_X1 _27477_ (.A1(_08452_),
    .A2(_08519_),
    .ZN(_08615_));
 AND3_X1 _27478_ (.A1(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .A3(_04911_),
    .ZN(_08616_));
 INV_X1 _27479_ (.A(_08616_),
    .ZN(_08617_));
 OAI21_X1 _27480_ (.A(_08615_),
    .B1(_08617_),
    .B2(_08597_),
    .ZN(_08618_));
 AOI21_X1 _27481_ (.A(_08614_),
    .B1(_08618_),
    .B2(_08612_),
    .ZN(_02718_));
 CLKBUF_X3 _27482_ (.A(_08603_),
    .Z(_08619_));
 NAND2_X1 _27483_ (.A1(_08605_),
    .A2(_08616_),
    .ZN(_08620_));
 NAND2_X1 _27484_ (.A1(_08469_),
    .A2(_08620_),
    .ZN(_08621_));
 AOI21_X1 _27485_ (.A(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .B1(_08619_),
    .B2(_08621_),
    .ZN(_08622_));
 AND2_X1 _27486_ (.A1(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .A2(_08616_),
    .ZN(_08623_));
 INV_X1 _27487_ (.A(_08623_),
    .ZN(_08624_));
 OAI22_X1 _27488_ (.A1(_08402_),
    .A2(_08491_),
    .B1(_08610_),
    .B2(_08624_),
    .ZN(_08625_));
 AOI21_X1 _27489_ (.A(_08622_),
    .B1(_08625_),
    .B2(_08612_),
    .ZN(_02719_));
 OAI21_X1 _27490_ (.A(_08587_),
    .B1(_08593_),
    .B2(_08624_),
    .ZN(_08626_));
 AOI21_X1 _27491_ (.A(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .B1(_08619_),
    .B2(_08626_),
    .ZN(_08627_));
 MUX2_X1 _27492_ (.A(_04466_),
    .B(_04467_),
    .S(_16261_),
    .Z(_08628_));
 OAI22_X4 _27493_ (.A1(_16261_),
    .A2(_06600_),
    .B1(_08628_),
    .B2(_04470_),
    .ZN(_08629_));
 INV_X2 _27494_ (.A(_08629_),
    .ZN(_08630_));
 AND2_X1 _27495_ (.A1(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .A2(_08623_),
    .ZN(_08631_));
 INV_X1 _27496_ (.A(_08631_),
    .ZN(_08632_));
 OAI22_X1 _27497_ (.A1(_08482_),
    .A2(_08630_),
    .B1(_08632_),
    .B2(_08597_),
    .ZN(_08633_));
 AOI21_X1 _27498_ (.A(_08627_),
    .B1(_08633_),
    .B2(_08612_),
    .ZN(_02720_));
 CLKBUF_X3 _27499_ (.A(_08411_),
    .Z(_08634_));
 NAND2_X1 _27500_ (.A1(_08605_),
    .A2(_08631_),
    .ZN(_08635_));
 NAND2_X1 _27501_ (.A1(_08634_),
    .A2(_08635_),
    .ZN(_08636_));
 AOI21_X1 _27502_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .B1(_08619_),
    .B2(_08636_),
    .ZN(_08637_));
 MUX2_X1 _27503_ (.A(_11772_),
    .B(_04465_),
    .S(_16273_),
    .Z(_08638_));
 OAI22_X4 _27504_ (.A1(_16269_),
    .A2(_05488_),
    .B1(_08638_),
    .B2(_04469_),
    .ZN(_08639_));
 NAND2_X1 _27505_ (.A1(_08434_),
    .A2(_08639_),
    .ZN(_08640_));
 NAND2_X1 _27506_ (.A1(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .A2(_08631_),
    .ZN(_08641_));
 OAI21_X1 _27507_ (.A(_08640_),
    .B1(_08641_),
    .B2(_08610_),
    .ZN(_08642_));
 AOI21_X1 _27508_ (.A(_08637_),
    .B1(_08642_),
    .B2(_08612_),
    .ZN(_02721_));
 OAI21_X1 _27509_ (.A(_08587_),
    .B1(_08593_),
    .B2(_08641_),
    .ZN(_08643_));
 AOI21_X1 _27510_ (.A(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .B1(_08619_),
    .B2(_08643_),
    .ZN(_08644_));
 MUX2_X1 _27511_ (.A(_04643_),
    .B(_04601_),
    .S(_16281_),
    .Z(_08645_));
 OAI22_X4 _27512_ (.A1(_16277_),
    .A2(_05523_),
    .B1(_08645_),
    .B2(_04668_),
    .ZN(_08646_));
 NAND2_X1 _27513_ (.A1(_08434_),
    .A2(_08646_),
    .ZN(_08647_));
 NAND3_X2 _27514_ (.A1(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .A3(_08631_),
    .ZN(_08648_));
 OAI21_X1 _27515_ (.A(_08647_),
    .B1(_08648_),
    .B2(_08597_),
    .ZN(_08649_));
 AOI21_X1 _27516_ (.A(_08644_),
    .B1(_08649_),
    .B2(_08612_),
    .ZN(_02722_));
 INV_X1 _27517_ (.A(_05603_),
    .ZN(_08650_));
 NOR3_X4 _27518_ (.A1(_08560_),
    .A2(_08591_),
    .A3(_08648_),
    .ZN(_08651_));
 OAI21_X1 _27519_ (.A(_08604_),
    .B1(_08651_),
    .B2(_08452_),
    .ZN(_08652_));
 NAND3_X1 _27520_ (.A1(_05603_),
    .A2(_08482_),
    .A3(_08651_),
    .ZN(_08653_));
 MUX2_X1 _27521_ (.A(_04601_),
    .B(_15928_),
    .S(_16285_),
    .Z(_08654_));
 OAI22_X4 _27522_ (.A1(_16285_),
    .A2(_05616_),
    .B1(_08654_),
    .B2(_04668_),
    .ZN(_08655_));
 NAND2_X1 _27523_ (.A1(_08461_),
    .A2(_08655_),
    .ZN(_08656_));
 NAND2_X1 _27524_ (.A1(_08653_),
    .A2(_08656_),
    .ZN(_08657_));
 CLKBUF_X3 _27525_ (.A(_08603_),
    .Z(_08658_));
 AOI22_X1 _27526_ (.A1(_08650_),
    .A2(_08652_),
    .B1(_08657_),
    .B2(_08658_),
    .ZN(_02723_));
 NOR2_X2 _27527_ (.A1(_08593_),
    .A2(_08648_),
    .ZN(_08659_));
 NAND2_X1 _27528_ (.A1(_05603_),
    .A2(_08659_),
    .ZN(_08660_));
 NAND2_X1 _27529_ (.A1(_08634_),
    .A2(_08660_),
    .ZN(_08661_));
 AOI21_X1 _27530_ (.A(_05690_),
    .B1(_08619_),
    .B2(_08661_),
    .ZN(_08662_));
 MUX2_X1 _27531_ (.A(_04465_),
    .B(_11772_),
    .S(_16293_),
    .Z(_08663_));
 NOR2_X2 _27532_ (.A1(_04469_),
    .A2(_08663_),
    .ZN(_08664_));
 AOI21_X4 _27533_ (.A(_08664_),
    .B1(_05704_),
    .B2(_16297_),
    .ZN(_08665_));
 BUF_X4 _27534_ (.A(_08665_),
    .Z(_08666_));
 NAND2_X1 _27535_ (.A1(_05603_),
    .A2(_05690_),
    .ZN(_08667_));
 NAND2_X1 _27536_ (.A1(_08482_),
    .A2(_08659_),
    .ZN(_08668_));
 OAI22_X1 _27537_ (.A1(_08482_),
    .A2(_08666_),
    .B1(_08667_),
    .B2(_08668_),
    .ZN(_08669_));
 AOI21_X1 _27538_ (.A(_08662_),
    .B1(_08669_),
    .B2(_08612_),
    .ZN(_02724_));
 NAND2_X1 _27539_ (.A1(_08634_),
    .A2(_08444_),
    .ZN(_08670_));
 AOI21_X1 _27540_ (.A(_06595_),
    .B1(_08416_),
    .B2(_08670_),
    .ZN(_08671_));
 INV_X1 _27541_ (.A(_06595_),
    .ZN(_08672_));
 OR3_X1 _27542_ (.A1(_08672_),
    .A2(_08430_),
    .A3(_08444_),
    .ZN(_08673_));
 OAI21_X1 _27543_ (.A(_08673_),
    .B1(_08630_),
    .B2(_08491_),
    .ZN(_08674_));
 AOI21_X1 _27544_ (.A(_08671_),
    .B1(_08674_),
    .B2(_08539_),
    .ZN(_02725_));
 NAND3_X1 _27545_ (.A1(_05603_),
    .A2(_05690_),
    .A3(_08651_),
    .ZN(_08675_));
 NAND2_X1 _27546_ (.A1(_08634_),
    .A2(_08675_),
    .ZN(_08676_));
 AOI21_X1 _27547_ (.A(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .B1(_08619_),
    .B2(_08676_),
    .ZN(_08677_));
 AND3_X1 _27548_ (.A1(_05603_),
    .A2(_05690_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .ZN(_08678_));
 NAND3_X1 _27549_ (.A1(_08482_),
    .A2(_08651_),
    .A3(_08678_),
    .ZN(_08679_));
 NAND2_X1 _27550_ (.A1(_04942_),
    .A2(_08434_),
    .ZN(_08680_));
 NAND2_X1 _27551_ (.A1(_08679_),
    .A2(_08680_),
    .ZN(_08681_));
 AOI21_X1 _27552_ (.A(_08677_),
    .B1(_08681_),
    .B2(_08612_),
    .ZN(_02726_));
 NAND2_X1 _27553_ (.A1(_08659_),
    .A2(_08678_),
    .ZN(_08682_));
 NAND2_X1 _27554_ (.A1(_08634_),
    .A2(_08682_),
    .ZN(_08683_));
 AOI21_X1 _27555_ (.A(_04945_),
    .B1(_08619_),
    .B2(_08683_),
    .ZN(_08684_));
 NAND2_X1 _27556_ (.A1(_04960_),
    .A2(_08461_),
    .ZN(_08685_));
 NAND2_X1 _27557_ (.A1(_04945_),
    .A2(_08678_),
    .ZN(_08686_));
 OAI21_X1 _27558_ (.A(_08685_),
    .B1(_08686_),
    .B2(_08668_),
    .ZN(_08687_));
 AOI21_X1 _27559_ (.A(_08684_),
    .B1(_08687_),
    .B2(_08612_),
    .ZN(_02727_));
 NAND3_X1 _27560_ (.A1(_04945_),
    .A2(_08651_),
    .A3(_08678_),
    .ZN(_08688_));
 NAND2_X1 _27561_ (.A1(_08634_),
    .A2(_08688_),
    .ZN(_08689_));
 AOI21_X1 _27562_ (.A(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .B1(_08619_),
    .B2(_08689_),
    .ZN(_08690_));
 AND3_X1 _27563_ (.A1(_04945_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .A3(_08678_),
    .ZN(_08691_));
 NAND3_X1 _27564_ (.A1(_08482_),
    .A2(_08651_),
    .A3(_08691_),
    .ZN(_08692_));
 NAND2_X1 _27565_ (.A1(_08438_),
    .A2(_08692_),
    .ZN(_08693_));
 AOI21_X1 _27566_ (.A(_08690_),
    .B1(_08693_),
    .B2(_08612_),
    .ZN(_02728_));
 NAND2_X1 _27567_ (.A1(_08659_),
    .A2(_08691_),
    .ZN(_08694_));
 NAND2_X1 _27568_ (.A1(_08634_),
    .A2(_08694_),
    .ZN(_08695_));
 AOI21_X1 _27569_ (.A(_04382_),
    .B1(_08619_),
    .B2(_08695_),
    .ZN(_08696_));
 NAND2_X1 _27570_ (.A1(_04382_),
    .A2(_08691_),
    .ZN(_08697_));
 OAI21_X1 _27571_ (.A(_08449_),
    .B1(_08668_),
    .B2(_08697_),
    .ZN(_08698_));
 CLKBUF_X3 _27572_ (.A(_08603_),
    .Z(_08699_));
 AOI21_X1 _27573_ (.A(_08696_),
    .B1(_08698_),
    .B2(_08699_),
    .ZN(_02729_));
 NAND3_X1 _27574_ (.A1(_04382_),
    .A2(_08651_),
    .A3(_08691_),
    .ZN(_08700_));
 NAND2_X1 _27575_ (.A1(_08634_),
    .A2(_08700_),
    .ZN(_08701_));
 AOI21_X1 _27576_ (.A(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .B1(_08619_),
    .B2(_08701_),
    .ZN(_08702_));
 AND3_X1 _27577_ (.A1(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .A2(_04382_),
    .A3(_08691_),
    .ZN(_08703_));
 AND2_X1 _27578_ (.A1(_08651_),
    .A2(_08703_),
    .ZN(_08704_));
 NAND2_X1 _27579_ (.A1(_08459_),
    .A2(_08704_),
    .ZN(_08705_));
 NAND2_X1 _27580_ (.A1(_08462_),
    .A2(_08705_),
    .ZN(_08706_));
 AOI21_X1 _27581_ (.A(_08702_),
    .B1(_08706_),
    .B2(_08699_),
    .ZN(_02730_));
 CLKBUF_X3 _27582_ (.A(_08603_),
    .Z(_08707_));
 NAND2_X2 _27583_ (.A1(_08659_),
    .A2(_08703_),
    .ZN(_08708_));
 NAND2_X1 _27584_ (.A1(_08634_),
    .A2(_08708_),
    .ZN(_08709_));
 AOI21_X1 _27585_ (.A(_04546_),
    .B1(_08707_),
    .B2(_08709_),
    .ZN(_08710_));
 OR2_X1 _27586_ (.A1(_08430_),
    .A2(_08708_),
    .ZN(_08711_));
 INV_X1 _27587_ (.A(_04546_),
    .ZN(_08712_));
 OAI21_X1 _27588_ (.A(_08466_),
    .B1(_08711_),
    .B2(_08712_),
    .ZN(_08713_));
 AOI21_X1 _27589_ (.A(_08710_),
    .B1(_08713_),
    .B2(_08699_),
    .ZN(_02731_));
 NAND2_X1 _27590_ (.A1(_04546_),
    .A2(_08704_),
    .ZN(_08714_));
 NAND2_X1 _27591_ (.A1(_08634_),
    .A2(_08714_),
    .ZN(_08715_));
 AOI21_X1 _27592_ (.A(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .B1(_08707_),
    .B2(_08715_),
    .ZN(_08716_));
 NAND2_X1 _27593_ (.A1(_04597_),
    .A2(_08412_),
    .ZN(_08717_));
 NAND2_X1 _27594_ (.A1(_04546_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .ZN(_08718_));
 OAI21_X1 _27595_ (.A(_08717_),
    .B1(_08705_),
    .B2(_08718_),
    .ZN(_08719_));
 AOI21_X1 _27596_ (.A(_08716_),
    .B1(_08719_),
    .B2(_08699_),
    .ZN(_02732_));
 OAI21_X1 _27597_ (.A(_08587_),
    .B1(_08708_),
    .B2(_08718_),
    .ZN(_08720_));
 AOI21_X1 _27598_ (.A(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .B1(_08707_),
    .B2(_08720_),
    .ZN(_08721_));
 AND3_X1 _27599_ (.A1(_04546_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .ZN(_08722_));
 INV_X1 _27600_ (.A(_08722_),
    .ZN(_08723_));
 OAI21_X1 _27601_ (.A(_08484_),
    .B1(_08711_),
    .B2(_08723_),
    .ZN(_08724_));
 AOI21_X1 _27602_ (.A(_08721_),
    .B1(_08724_),
    .B2(_08699_),
    .ZN(_02733_));
 NAND2_X1 _27603_ (.A1(_08704_),
    .A2(_08722_),
    .ZN(_08725_));
 NAND2_X1 _27604_ (.A1(_08520_),
    .A2(_08725_),
    .ZN(_08726_));
 AOI21_X1 _27605_ (.A(_04623_),
    .B1(_08707_),
    .B2(_08726_),
    .ZN(_08727_));
 NAND2_X1 _27606_ (.A1(_04623_),
    .A2(_08722_),
    .ZN(_08728_));
 OAI22_X1 _27607_ (.A1(_08493_),
    .A2(_08491_),
    .B1(_08705_),
    .B2(_08728_),
    .ZN(_08729_));
 AOI21_X1 _27608_ (.A(_08727_),
    .B1(_08729_),
    .B2(_08699_),
    .ZN(_02734_));
 OAI21_X1 _27609_ (.A(_08587_),
    .B1(_08708_),
    .B2(_08728_),
    .ZN(_08730_));
 AOI21_X1 _27610_ (.A(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .B1(_08707_),
    .B2(_08730_),
    .ZN(_08731_));
 NAND3_X2 _27611_ (.A1(_04623_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .A3(_08722_),
    .ZN(_08732_));
 OAI21_X1 _27612_ (.A(_08498_),
    .B1(_08711_),
    .B2(_08732_),
    .ZN(_08733_));
 AOI21_X1 _27613_ (.A(_08731_),
    .B1(_08733_),
    .B2(_08699_),
    .ZN(_02735_));
 OAI21_X1 _27614_ (.A(_08587_),
    .B1(_08419_),
    .B2(_08672_),
    .ZN(_08734_));
 AOI21_X1 _27615_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B1(_08416_),
    .B2(_08734_),
    .ZN(_08735_));
 NAND2_X1 _27616_ (.A1(_06595_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .ZN(_08736_));
 OAI21_X1 _27617_ (.A(_08640_),
    .B1(_08585_),
    .B2(_08736_),
    .ZN(_08737_));
 AOI21_X1 _27618_ (.A(_08735_),
    .B1(_08737_),
    .B2(_08454_),
    .ZN(_02736_));
 INV_X1 _27619_ (.A(_04670_),
    .ZN(_08738_));
 AND3_X1 _27620_ (.A1(_04623_),
    .A2(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .A3(_08722_),
    .ZN(_08739_));
 AND2_X1 _27621_ (.A1(_08704_),
    .A2(_08739_),
    .ZN(_08740_));
 OAI21_X1 _27622_ (.A(_08604_),
    .B1(_08740_),
    .B2(_08452_),
    .ZN(_08741_));
 NAND3_X1 _27623_ (.A1(_04670_),
    .A2(_08459_),
    .A3(_08740_),
    .ZN(_08742_));
 INV_X2 _27624_ (.A(_04685_),
    .ZN(_08743_));
 OAI21_X1 _27625_ (.A(_08742_),
    .B1(_08491_),
    .B2(_08743_),
    .ZN(_08744_));
 AOI22_X1 _27626_ (.A1(_08738_),
    .A2(_08741_),
    .B1(_08744_),
    .B2(_08658_),
    .ZN(_02737_));
 INV_X1 _27627_ (.A(_04696_),
    .ZN(_08745_));
 NOR3_X1 _27628_ (.A1(_08738_),
    .A2(_08708_),
    .A3(_08732_),
    .ZN(_08746_));
 OAI21_X1 _27629_ (.A(_08604_),
    .B1(_08746_),
    .B2(_08452_),
    .ZN(_08747_));
 NAND3_X1 _27630_ (.A1(_04670_),
    .A2(_04696_),
    .A3(_08739_),
    .ZN(_08748_));
 OAI21_X1 _27631_ (.A(_08514_),
    .B1(_08711_),
    .B2(_08748_),
    .ZN(_08749_));
 AOI22_X1 _27632_ (.A1(_08745_),
    .A2(_08747_),
    .B1(_08749_),
    .B2(_08658_),
    .ZN(_02738_));
 NAND3_X1 _27633_ (.A1(_04670_),
    .A2(_04696_),
    .A3(_08740_),
    .ZN(_08750_));
 NAND2_X1 _27634_ (.A1(_08520_),
    .A2(_08750_),
    .ZN(_08751_));
 AOI21_X1 _27635_ (.A(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .B1(_08707_),
    .B2(_08751_),
    .ZN(_08752_));
 AND4_X1 _27636_ (.A1(_04670_),
    .A2(_04696_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .A4(_08740_),
    .ZN(_08753_));
 NAND2_X1 _27637_ (.A1(_08418_),
    .A2(_08753_),
    .ZN(_08754_));
 NAND2_X1 _27638_ (.A1(_08527_),
    .A2(_08754_),
    .ZN(_08755_));
 AOI21_X1 _27639_ (.A(_08752_),
    .B1(_08755_),
    .B2(_08699_),
    .ZN(_02739_));
 INV_X1 _27640_ (.A(_04738_),
    .ZN(_08756_));
 NAND3_X1 _27641_ (.A1(_04670_),
    .A2(_04696_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .ZN(_08757_));
 NOR3_X4 _27642_ (.A1(_08708_),
    .A2(_08732_),
    .A3(_08757_),
    .ZN(_08758_));
 OAI21_X1 _27643_ (.A(_08604_),
    .B1(_08758_),
    .B2(_08452_),
    .ZN(_08759_));
 NAND3_X1 _27644_ (.A1(_04738_),
    .A2(_08482_),
    .A3(_08758_),
    .ZN(_08760_));
 NAND2_X1 _27645_ (.A1(_08531_),
    .A2(_08760_),
    .ZN(_08761_));
 AOI22_X1 _27646_ (.A1(_08756_),
    .A2(_08759_),
    .B1(_08761_),
    .B2(_08658_),
    .ZN(_02740_));
 NAND2_X1 _27647_ (.A1(_04738_),
    .A2(_08753_),
    .ZN(_08762_));
 NAND2_X1 _27648_ (.A1(_08520_),
    .A2(_08762_),
    .ZN(_08763_));
 AOI21_X1 _27649_ (.A(_04757_),
    .B1(_08707_),
    .B2(_08763_),
    .ZN(_08764_));
 INV_X1 _27650_ (.A(_04762_),
    .ZN(_08765_));
 NAND2_X1 _27651_ (.A1(_04738_),
    .A2(_04757_),
    .ZN(_08766_));
 OAI22_X1 _27652_ (.A1(_08765_),
    .A2(_08491_),
    .B1(_08754_),
    .B2(_08766_),
    .ZN(_08767_));
 AOI21_X1 _27653_ (.A(_08764_),
    .B1(_08767_),
    .B2(_08699_),
    .ZN(_02741_));
 NAND3_X1 _27654_ (.A1(_04738_),
    .A2(_04757_),
    .A3(_08758_),
    .ZN(_08768_));
 NAND2_X1 _27655_ (.A1(_08520_),
    .A2(_08768_),
    .ZN(_08769_));
 AOI21_X1 _27656_ (.A(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .B1(_08707_),
    .B2(_08769_),
    .ZN(_08770_));
 NAND4_X2 _27657_ (.A1(_04738_),
    .A2(_04757_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .A4(_08758_),
    .ZN(_08771_));
 OR2_X1 _27658_ (.A1(_08430_),
    .A2(_08771_),
    .ZN(_08772_));
 NAND2_X1 _27659_ (.A1(_08544_),
    .A2(_08772_),
    .ZN(_08773_));
 AOI21_X1 _27660_ (.A(_08770_),
    .B1(_08773_),
    .B2(_08699_),
    .ZN(_02742_));
 INV_X1 _27661_ (.A(_04788_),
    .ZN(_08774_));
 AND4_X1 _27662_ (.A1(_04738_),
    .A2(_04757_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .A4(_08753_),
    .ZN(_08775_));
 OAI21_X1 _27663_ (.A(_08604_),
    .B1(_08775_),
    .B2(_08412_),
    .ZN(_08776_));
 NAND2_X1 _27664_ (.A1(_08481_),
    .A2(_08775_),
    .ZN(_08777_));
 OAI21_X1 _27665_ (.A(_08551_),
    .B1(_08777_),
    .B2(_08774_),
    .ZN(_08778_));
 AOI22_X1 _27666_ (.A1(_08774_),
    .A2(_08776_),
    .B1(_08778_),
    .B2(_08604_),
    .ZN(_02743_));
 OAI21_X1 _27667_ (.A(_08587_),
    .B1(_08771_),
    .B2(_08774_),
    .ZN(_08779_));
 AOI21_X1 _27668_ (.A(_04818_),
    .B1(_08707_),
    .B2(_08779_),
    .ZN(_08780_));
 NAND2_X1 _27669_ (.A1(_04788_),
    .A2(_04818_),
    .ZN(_08781_));
 OAI21_X1 _27670_ (.A(_08556_),
    .B1(_08772_),
    .B2(_08781_),
    .ZN(_08782_));
 AOI21_X1 _27671_ (.A(_08780_),
    .B1(_08782_),
    .B2(_08658_),
    .ZN(_02744_));
 NAND3_X1 _27672_ (.A1(_04788_),
    .A2(_04818_),
    .A3(_08775_),
    .ZN(_08783_));
 NAND2_X1 _27673_ (.A1(_08520_),
    .A2(_08783_),
    .ZN(_08784_));
 AOI21_X1 _27674_ (.A(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .B1(_08707_),
    .B2(_08784_),
    .ZN(_08785_));
 NAND3_X1 _27675_ (.A1(_04788_),
    .A2(_04818_),
    .A3(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .ZN(_08786_));
 OAI21_X1 _27676_ (.A(_08563_),
    .B1(_08777_),
    .B2(_08786_),
    .ZN(_08787_));
 AOI21_X1 _27677_ (.A(_08785_),
    .B1(_08787_),
    .B2(_08658_),
    .ZN(_02745_));
 OAI21_X1 _27678_ (.A(_08587_),
    .B1(_08771_),
    .B2(_08786_),
    .ZN(_08788_));
 AOI21_X1 _27679_ (.A(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .B1(_08603_),
    .B2(_08788_),
    .ZN(_08789_));
 INV_X1 _27680_ (.A(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .ZN(_08790_));
 NOR2_X1 _27681_ (.A1(_08790_),
    .A2(_08786_),
    .ZN(_08791_));
 INV_X1 _27682_ (.A(_08791_),
    .ZN(_08792_));
 OAI21_X1 _27683_ (.A(_08568_),
    .B1(_08772_),
    .B2(_08792_),
    .ZN(_08793_));
 AOI21_X1 _27684_ (.A(_08789_),
    .B1(_08793_),
    .B2(_08658_),
    .ZN(_02746_));
 OAI21_X1 _27685_ (.A(_08587_),
    .B1(_08736_),
    .B2(_08444_),
    .ZN(_08794_));
 AOI21_X1 _27686_ (.A(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .B1(_08416_),
    .B2(_08794_),
    .ZN(_08795_));
 NOR3_X1 _27687_ (.A1(_08431_),
    .A2(_08420_),
    .A3(_08444_),
    .ZN(_08796_));
 AOI21_X1 _27688_ (.A(_08796_),
    .B1(_08646_),
    .B2(_08412_),
    .ZN(_08797_));
 INV_X1 _27689_ (.A(_08797_),
    .ZN(_08798_));
 AOI21_X1 _27690_ (.A(_08795_),
    .B1(_08798_),
    .B2(_08454_),
    .ZN(_02747_));
 NAND2_X1 _27691_ (.A1(_08775_),
    .A2(_08791_),
    .ZN(_08799_));
 NAND2_X1 _27692_ (.A1(_08520_),
    .A2(_08799_),
    .ZN(_08800_));
 AOI21_X1 _27693_ (.A(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .B1(_08603_),
    .B2(_08800_),
    .ZN(_08801_));
 NAND2_X1 _27694_ (.A1(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .A2(_08791_),
    .ZN(_08802_));
 OAI21_X1 _27695_ (.A(_08574_),
    .B1(_08777_),
    .B2(_08802_),
    .ZN(_08803_));
 AOI21_X1 _27696_ (.A(_08801_),
    .B1(_08803_),
    .B2(_08658_),
    .ZN(_02748_));
 OAI21_X1 _27697_ (.A(_08459_),
    .B1(_08771_),
    .B2(_08802_),
    .ZN(_08804_));
 AOI21_X1 _27698_ (.A(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .B1(_08603_),
    .B2(_08804_),
    .ZN(_08805_));
 AND3_X1 _27699_ (.A1(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .A3(_08791_),
    .ZN(_08806_));
 INV_X1 _27700_ (.A(_08806_),
    .ZN(_08807_));
 OAI21_X1 _27701_ (.A(_08579_),
    .B1(_08772_),
    .B2(_08807_),
    .ZN(_08808_));
 AOI21_X1 _27702_ (.A(_08805_),
    .B1(_08808_),
    .B2(_08658_),
    .ZN(_02749_));
 NAND2_X1 _27703_ (.A1(_08775_),
    .A2(_08806_),
    .ZN(_08809_));
 NAND2_X1 _27704_ (.A1(_08520_),
    .A2(_08809_),
    .ZN(_08810_));
 AOI21_X1 _27705_ (.A(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .B1(_08603_),
    .B2(_08810_),
    .ZN(_08811_));
 NAND2_X1 _27706_ (.A1(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .A2(_08806_),
    .ZN(_08812_));
 OAI21_X1 _27707_ (.A(_08590_),
    .B1(_08777_),
    .B2(_08812_),
    .ZN(_08813_));
 AOI21_X1 _27708_ (.A(_08811_),
    .B1(_08813_),
    .B2(_08658_),
    .ZN(_02750_));
 INV_X1 _27709_ (.A(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .ZN(_08814_));
 NOR2_X1 _27710_ (.A1(_08771_),
    .A2(_08812_),
    .ZN(_08815_));
 OAI21_X1 _27711_ (.A(_08604_),
    .B1(_08815_),
    .B2(_08452_),
    .ZN(_08816_));
 NAND3_X1 _27712_ (.A1(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .A2(_08482_),
    .A3(_08815_),
    .ZN(_08817_));
 NAND2_X1 _27713_ (.A1(_08596_),
    .A2(_08817_),
    .ZN(_08818_));
 AOI22_X1 _27714_ (.A1(_08814_),
    .A2(_08816_),
    .B1(_08818_),
    .B2(_08604_),
    .ZN(_02751_));
 NAND3_X1 _27715_ (.A1(_05606_),
    .A2(_08469_),
    .A3(_08421_),
    .ZN(_08819_));
 NAND2_X1 _27716_ (.A1(_08656_),
    .A2(_08819_),
    .ZN(_08820_));
 OAI21_X1 _27717_ (.A(_08415_),
    .B1(_08421_),
    .B2(_08452_),
    .ZN(_08821_));
 AOI22_X1 _27718_ (.A1(_08440_),
    .A2(_08820_),
    .B1(_08821_),
    .B2(_08442_),
    .ZN(_02752_));
 OAI21_X1 _27719_ (.A(_08459_),
    .B1(_08445_),
    .B2(_08442_),
    .ZN(_08822_));
 AOI21_X1 _27720_ (.A(_05693_),
    .B1(_08416_),
    .B2(_08822_),
    .ZN(_08823_));
 NAND2_X1 _27721_ (.A1(_08491_),
    .A2(_08446_),
    .ZN(_08824_));
 OAI21_X1 _27722_ (.A(_08824_),
    .B1(_08666_),
    .B2(_08491_),
    .ZN(_08825_));
 AOI21_X1 _27723_ (.A(_08823_),
    .B1(_08825_),
    .B2(_08454_),
    .ZN(_02753_));
 NAND2_X1 _27724_ (.A1(_08520_),
    .A2(_08422_),
    .ZN(_08826_));
 AOI21_X1 _27725_ (.A(_04931_),
    .B1(_08416_),
    .B2(_08826_),
    .ZN(_08827_));
 NAND2_X1 _27726_ (.A1(_04931_),
    .A2(_08432_),
    .ZN(_08828_));
 NAND2_X1 _27727_ (.A1(_08680_),
    .A2(_08828_),
    .ZN(_08829_));
 AOI21_X1 _27728_ (.A(_08827_),
    .B1(_08829_),
    .B2(_08454_),
    .ZN(_02754_));
 NAND2_X1 _27729_ (.A1(_04931_),
    .A2(_08446_),
    .ZN(_08830_));
 NAND2_X1 _27730_ (.A1(_08520_),
    .A2(_08830_),
    .ZN(_08831_));
 AOI21_X1 _27731_ (.A(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .B1(_08416_),
    .B2(_08831_),
    .ZN(_08832_));
 OAI21_X1 _27732_ (.A(_08685_),
    .B1(_08824_),
    .B2(_08423_),
    .ZN(_08833_));
 AOI21_X1 _27733_ (.A(_08832_),
    .B1(_08833_),
    .B2(_08454_),
    .ZN(_02755_));
 INV_X1 _27734_ (.A(_03645_),
    .ZN(_08834_));
 NOR4_X4 _27735_ (.A1(_08834_),
    .A2(_03565_),
    .A3(_03644_),
    .A4(_03654_),
    .ZN(_08835_));
 XNOR2_X2 _27736_ (.A(_16266_),
    .B(_05216_),
    .ZN(_08836_));
 XNOR2_X2 _27737_ (.A(_11490_),
    .B(_11379_),
    .ZN(_08837_));
 NOR2_X2 _27738_ (.A1(_15911_),
    .A2(_15915_),
    .ZN(_08838_));
 NAND2_X1 _27739_ (.A1(_03571_),
    .A2(_08838_),
    .ZN(_08839_));
 NOR4_X4 _27740_ (.A1(_16242_),
    .A2(_08836_),
    .A3(_08837_),
    .A4(_08839_),
    .ZN(_08840_));
 AND3_X1 _27741_ (.A1(_03594_),
    .A2(_08835_),
    .A3(_08840_),
    .ZN(_08841_));
 BUF_X4 _27742_ (.A(_08841_),
    .Z(_08842_));
 NAND2_X2 _27743_ (.A1(_04588_),
    .A2(_08842_),
    .ZN(_08843_));
 CLKBUF_X3 _27744_ (.A(_08843_),
    .Z(_08844_));
 NAND2_X1 _27745_ (.A1(_03648_),
    .A2(_01158_),
    .ZN(_08845_));
 OR4_X1 _27746_ (.A1(_03679_),
    .A2(_07212_),
    .A3(_07236_),
    .A4(_08845_),
    .ZN(_08846_));
 OR3_X1 _27747_ (.A1(_03688_),
    .A2(_05665_),
    .A3(_08846_),
    .ZN(_08847_));
 OAI33_X1 _27748_ (.A1(_03571_),
    .A2(_03688_),
    .A3(_08846_),
    .B1(_08847_),
    .B2(_03644_),
    .B3(_03565_),
    .ZN(_08848_));
 INV_X2 _27749_ (.A(_08848_),
    .ZN(_08849_));
 AOI21_X2 _27750_ (.A(_08849_),
    .B1(_07244_),
    .B2(net333),
    .ZN(_08850_));
 AOI211_X2 _27751_ (.A(_05198_),
    .B(_08849_),
    .C1(_05200_),
    .C2(_03745_),
    .ZN(_08851_));
 NAND4_X2 _27752_ (.A1(_05166_),
    .A2(_05167_),
    .A3(_03732_),
    .A4(_05187_),
    .ZN(_08852_));
 AOI21_X4 _27753_ (.A(_08850_),
    .B1(_08851_),
    .B2(_08852_),
    .ZN(_08853_));
 BUF_X4 _27754_ (.A(_08853_),
    .Z(_08854_));
 BUF_X4 _27755_ (.A(_08854_),
    .Z(_08855_));
 BUF_X4 _27756_ (.A(_08842_),
    .Z(_08856_));
 BUF_X4 _27757_ (.A(_08856_),
    .Z(_08857_));
 OAI21_X4 _27758_ (.A(_08844_),
    .B1(_08855_),
    .B2(_08857_),
    .ZN(_08858_));
 NOR2_X1 _27759_ (.A1(\cs_registers_i.mhpmcounter[2][0] ),
    .A2(_08858_),
    .ZN(_08859_));
 INV_X1 _27760_ (.A(_08396_),
    .ZN(_08860_));
 NAND3_X2 _27761_ (.A1(_03594_),
    .A2(_08835_),
    .A3(_08840_),
    .ZN(_08861_));
 BUF_X4 _27762_ (.A(_08861_),
    .Z(_08862_));
 NOR2_X1 _27763_ (.A1(_08860_),
    .A2(_08862_),
    .ZN(_08863_));
 CLKBUF_X3 _27764_ (.A(_08862_),
    .Z(_08864_));
 AOI21_X1 _27765_ (.A(_08863_),
    .B1(_08864_),
    .B2(_00553_),
    .ZN(_08865_));
 AOI21_X1 _27766_ (.A(_08859_),
    .B1(_08858_),
    .B2(_08865_),
    .ZN(_02756_));
 NOR2_X1 _27767_ (.A1(_04668_),
    .A2(_08436_),
    .ZN(_08866_));
 AOI21_X4 _27768_ (.A(_08866_),
    .B1(_05840_),
    .B2(_16321_),
    .ZN(_08867_));
 NAND3_X2 _27769_ (.A1(_11173_),
    .A2(_11329_),
    .A3(_08838_),
    .ZN(_08868_));
 NOR4_X4 _27770_ (.A1(_04542_),
    .A2(_08836_),
    .A3(_08837_),
    .A4(_08868_),
    .ZN(_08869_));
 AND2_X1 _27771_ (.A1(_08403_),
    .A2(_08869_),
    .ZN(_08870_));
 BUF_X4 _27772_ (.A(_08870_),
    .Z(_08871_));
 AND2_X1 _27773_ (.A1(_04756_),
    .A2(_08871_),
    .ZN(_08872_));
 OR3_X2 _27774_ (.A1(_03688_),
    .A2(_05399_),
    .A3(_08846_),
    .ZN(_08873_));
 OR2_X2 _27775_ (.A1(_08873_),
    .A2(_08870_),
    .ZN(_08874_));
 NAND2_X1 _27776_ (.A1(_04932_),
    .A2(_04948_),
    .ZN(_08875_));
 CLKBUF_X3 _27777_ (.A(_15934_),
    .Z(_08876_));
 AND4_X1 _27778_ (.A1(_06560_),
    .A2(_06596_),
    .A3(\cs_registers_i.mhpmcounter[2][4] ),
    .A4(_05519_),
    .ZN(_08877_));
 AND2_X1 _27779_ (.A1(\cs_registers_i.mhpmcounter[2][6] ),
    .A2(_08877_),
    .ZN(_08878_));
 AND2_X1 _27780_ (.A1(_05694_),
    .A2(_08878_),
    .ZN(_08879_));
 NAND2_X2 _27781_ (.A1(_08876_),
    .A2(_08879_),
    .ZN(_08880_));
 NOR4_X2 _27782_ (.A1(\id_stage_i.branch_set_d ),
    .A2(_08874_),
    .A3(_08875_),
    .A4(_08880_),
    .ZN(_08881_));
 INV_X1 _27783_ (.A(\cs_registers_i.mhpmcounter[2][10] ),
    .ZN(_08882_));
 AOI22_X1 _27784_ (.A1(_08867_),
    .A2(_08872_),
    .B1(_08881_),
    .B2(_08882_),
    .ZN(_08883_));
 CLKBUF_X3 _27785_ (.A(_08843_),
    .Z(_08884_));
 NAND2_X1 _27786_ (.A1(\cs_registers_i.mhpmcounter[2][10] ),
    .A2(_08884_),
    .ZN(_08885_));
 OAI21_X1 _27787_ (.A(_08883_),
    .B1(_08881_),
    .B2(_08885_),
    .ZN(_02757_));
 BUF_X4 _27788_ (.A(_08857_),
    .Z(_08886_));
 INV_X1 _27789_ (.A(_04948_),
    .ZN(_08887_));
 NAND2_X1 _27790_ (.A1(_05694_),
    .A2(_04932_),
    .ZN(_08888_));
 NOR3_X2 _27791_ (.A1(_08887_),
    .A2(_08882_),
    .A3(_08888_),
    .ZN(_08889_));
 INV_X1 _27792_ (.A(_08889_),
    .ZN(_08890_));
 AND2_X1 _27793_ (.A1(\cs_registers_i.mhpmcounter[2][1] ),
    .A2(\cs_registers_i.mhpmcounter[2][0] ),
    .ZN(_08891_));
 CLKBUF_X3 _27794_ (.A(_08891_),
    .Z(_08892_));
 NAND2_X2 _27795_ (.A1(_08878_),
    .A2(_08892_),
    .ZN(_08893_));
 NOR4_X1 _27796_ (.A1(_04396_),
    .A2(_08886_),
    .A3(_08890_),
    .A4(_08893_),
    .ZN(_08894_));
 BUF_X2 _27797_ (.A(_08861_),
    .Z(_08895_));
 CLKBUF_X3 _27798_ (.A(_08895_),
    .Z(_08896_));
 NOR2_X1 _27799_ (.A1(_04472_),
    .A2(_08896_),
    .ZN(_08897_));
 OAI21_X1 _27800_ (.A(_08858_),
    .B1(_08894_),
    .B2(_08897_),
    .ZN(_08898_));
 OR2_X1 _27801_ (.A1(\id_stage_i.branch_set_d ),
    .A2(_08874_),
    .ZN(_08899_));
 NOR3_X1 _27802_ (.A1(_08899_),
    .A2(_08890_),
    .A3(_08893_),
    .ZN(_08900_));
 NAND2_X1 _27803_ (.A1(_04396_),
    .A2(_08884_),
    .ZN(_08901_));
 OAI21_X1 _27804_ (.A(_08898_),
    .B1(_08900_),
    .B2(_08901_),
    .ZN(_02758_));
 NAND3_X1 _27805_ (.A1(_11173_),
    .A2(_11329_),
    .A3(_08838_),
    .ZN(_08902_));
 NOR3_X1 _27806_ (.A1(_08836_),
    .A2(_08837_),
    .A3(_08902_),
    .ZN(_08903_));
 AND2_X1 _27807_ (.A1(_04490_),
    .A2(_08903_),
    .ZN(_08904_));
 AND2_X1 _27808_ (.A1(_08403_),
    .A2(_08904_),
    .ZN(_08905_));
 NAND2_X1 _27809_ (.A1(_04756_),
    .A2(_08905_),
    .ZN(_08906_));
 CLKBUF_X3 _27810_ (.A(_08906_),
    .Z(_08907_));
 NOR2_X1 _27811_ (.A1(_04528_),
    .A2(_08907_),
    .ZN(_08908_));
 NAND2_X1 _27812_ (.A1(_04504_),
    .A2(_08843_),
    .ZN(_08909_));
 NAND4_X2 _27813_ (.A1(_04396_),
    .A2(_04932_),
    .A3(_04948_),
    .A4(\cs_registers_i.mhpmcounter[2][10] ),
    .ZN(_08910_));
 NOR2_X1 _27814_ (.A1(_08880_),
    .A2(_08910_),
    .ZN(_08911_));
 NOR2_X4 _27815_ (.A1(_08842_),
    .A2(_08853_),
    .ZN(_08912_));
 AOI21_X1 _27816_ (.A(_08909_),
    .B1(_08911_),
    .B2(_08912_),
    .ZN(_08913_));
 NOR2_X2 _27817_ (.A1(_08873_),
    .A2(_08905_),
    .ZN(_08914_));
 NAND2_X2 _27818_ (.A1(_07226_),
    .A2(_08914_),
    .ZN(_08915_));
 NOR4_X1 _27819_ (.A1(_04504_),
    .A2(_08915_),
    .A3(_08880_),
    .A4(_08910_),
    .ZN(_08916_));
 OR3_X1 _27820_ (.A1(_08908_),
    .A2(_08913_),
    .A3(_08916_),
    .ZN(_02759_));
 AND2_X1 _27821_ (.A1(_04550_),
    .A2(_08844_),
    .ZN(_08917_));
 AND4_X2 _27822_ (.A1(_04504_),
    .A2(_04396_),
    .A3(_08878_),
    .A4(_08889_),
    .ZN(_08918_));
 NAND2_X1 _27823_ (.A1(_08892_),
    .A2(_08918_),
    .ZN(_08919_));
 CLKBUF_X3 _27824_ (.A(_08915_),
    .Z(_08920_));
 OAI21_X1 _27825_ (.A(_08917_),
    .B1(_08919_),
    .B2(_08920_),
    .ZN(_08921_));
 NAND2_X4 _27826_ (.A1(_04756_),
    .A2(_08871_),
    .ZN(_08922_));
 NOR2_X4 _27827_ (.A1(\id_stage_i.branch_set_d ),
    .A2(_08874_),
    .ZN(_08923_));
 NAND3_X1 _27828_ (.A1(_08923_),
    .A2(_08892_),
    .A3(_08918_),
    .ZN(_08924_));
 OAI221_X1 _27829_ (.A(_08921_),
    .B1(_08922_),
    .B2(_04562_),
    .C1(_04550_),
    .C2(_08924_),
    .ZN(_02760_));
 OAI22_X1 _27830_ (.A1(_04586_),
    .A2(_08871_),
    .B1(_08844_),
    .B2(_04596_),
    .ZN(_08925_));
 NAND2_X1 _27831_ (.A1(_04586_),
    .A2(_08844_),
    .ZN(_08926_));
 OAI21_X1 _27832_ (.A(_08926_),
    .B1(_08844_),
    .B2(_04597_),
    .ZN(_08927_));
 NAND3_X1 _27833_ (.A1(_04504_),
    .A2(_08876_),
    .A3(_04550_),
    .ZN(_08928_));
 NOR2_X1 _27834_ (.A1(_08910_),
    .A2(_08928_),
    .ZN(_08929_));
 NAND3_X1 _27835_ (.A1(_08912_),
    .A2(_08879_),
    .A3(_08929_),
    .ZN(_08930_));
 MUX2_X1 _27836_ (.A(_08925_),
    .B(_08927_),
    .S(_08930_),
    .Z(_02761_));
 AND3_X1 _27837_ (.A1(_04504_),
    .A2(_04550_),
    .A3(_04586_),
    .ZN(_08931_));
 AND4_X1 _27838_ (.A1(_04396_),
    .A2(_08878_),
    .A3(_08889_),
    .A4(_08931_),
    .ZN(_08932_));
 NAND2_X2 _27839_ (.A1(_08892_),
    .A2(_08932_),
    .ZN(_08933_));
 NOR4_X1 _27840_ (.A1(_04606_),
    .A2(_08857_),
    .A3(_08855_),
    .A4(_08933_),
    .ZN(_08934_));
 AND2_X2 _27841_ (.A1(_04588_),
    .A2(_08856_),
    .ZN(_08935_));
 INV_X1 _27842_ (.A(_04620_),
    .ZN(_08936_));
 AOI21_X1 _27843_ (.A(_08934_),
    .B1(_08935_),
    .B2(_08936_),
    .ZN(_08937_));
 NAND2_X1 _27844_ (.A1(_04606_),
    .A2(_08884_),
    .ZN(_08938_));
 NOR3_X4 _27845_ (.A1(_08856_),
    .A2(_08853_),
    .A3(_08933_),
    .ZN(_08939_));
 OAI21_X1 _27846_ (.A(_08937_),
    .B1(_08938_),
    .B2(_08939_),
    .ZN(_02762_));
 INV_X1 _27847_ (.A(_04606_),
    .ZN(_08940_));
 NAND4_X4 _27848_ (.A1(_08876_),
    .A2(_04550_),
    .A3(_04586_),
    .A4(_08918_),
    .ZN(_08941_));
 NOR4_X2 _27849_ (.A1(_08940_),
    .A2(\id_stage_i.branch_set_d ),
    .A3(_08874_),
    .A4(_08941_),
    .ZN(_08942_));
 INV_X1 _27850_ (.A(_04627_),
    .ZN(_08943_));
 AOI22_X1 _27851_ (.A1(_08493_),
    .A2(_08872_),
    .B1(_08942_),
    .B2(_08943_),
    .ZN(_08944_));
 NAND2_X1 _27852_ (.A1(_04627_),
    .A2(_08884_),
    .ZN(_08945_));
 OAI21_X1 _27853_ (.A(_08944_),
    .B1(_08942_),
    .B2(_08945_),
    .ZN(_02763_));
 INV_X1 _27854_ (.A(\cs_registers_i.mhpmcounter[2][17] ),
    .ZN(_08946_));
 NAND4_X1 _27855_ (.A1(_04606_),
    .A2(_04627_),
    .A3(_08946_),
    .A4(_08939_),
    .ZN(_08947_));
 AND3_X1 _27856_ (.A1(_04606_),
    .A2(_04627_),
    .A3(_08939_),
    .ZN(_08948_));
 NAND2_X1 _27857_ (.A1(\cs_registers_i.mhpmcounter[2][17] ),
    .A2(_08884_),
    .ZN(_08949_));
 OAI221_X1 _27858_ (.A(_08947_),
    .B1(_08948_),
    .B2(_08949_),
    .C1(_04665_),
    .C2(_08922_),
    .ZN(_02764_));
 NAND2_X1 _27859_ (.A1(_04673_),
    .A2(_08907_),
    .ZN(_08950_));
 AND4_X1 _27860_ (.A1(_08876_),
    .A2(_04550_),
    .A3(_04586_),
    .A4(_08918_),
    .ZN(_08951_));
 AND3_X1 _27861_ (.A1(_04606_),
    .A2(_04627_),
    .A3(\cs_registers_i.mhpmcounter[2][17] ),
    .ZN(_08952_));
 AND3_X1 _27862_ (.A1(_08923_),
    .A2(_08951_),
    .A3(_08952_),
    .ZN(_08953_));
 INV_X1 _27863_ (.A(_04673_),
    .ZN(_08954_));
 AND2_X1 _27864_ (.A1(_08954_),
    .A2(_08952_),
    .ZN(_08955_));
 NOR2_X1 _27865_ (.A1(_08871_),
    .A2(_08941_),
    .ZN(_08956_));
 AOI22_X1 _27866_ (.A1(_08743_),
    .A2(_08905_),
    .B1(_08955_),
    .B2(_08956_),
    .ZN(_08957_));
 AND2_X1 _27867_ (.A1(_08915_),
    .A2(_08906_),
    .ZN(_08958_));
 OAI22_X1 _27868_ (.A1(_08950_),
    .A2(_08953_),
    .B1(_08957_),
    .B2(_08958_),
    .ZN(_02765_));
 NOR2_X1 _27869_ (.A1(\cs_registers_i.mhpmcounter[2][19] ),
    .A2(_08935_),
    .ZN(_08959_));
 NAND3_X1 _27870_ (.A1(_04673_),
    .A2(_08939_),
    .A3(_08952_),
    .ZN(_08960_));
 NAND3_X1 _27871_ (.A1(_04673_),
    .A2(\cs_registers_i.mhpmcounter[2][19] ),
    .A3(_08952_),
    .ZN(_08961_));
 NOR2_X1 _27872_ (.A1(_08933_),
    .A2(_08961_),
    .ZN(_08962_));
 MUX2_X1 _27873_ (.A(_04700_),
    .B(_08962_),
    .S(_08862_),
    .Z(_08963_));
 AOI22_X1 _27874_ (.A1(_08959_),
    .A2(_08960_),
    .B1(_08963_),
    .B2(_08858_),
    .ZN(_02766_));
 NOR2_X1 _27875_ (.A1(\cs_registers_i.mhpmcounter[2][1] ),
    .A2(_08858_),
    .ZN(_08964_));
 NOR2_X1 _27876_ (.A1(_08519_),
    .A2(_08862_),
    .ZN(_08965_));
 AOI21_X1 _27877_ (.A(_08965_),
    .B1(_08864_),
    .B2(_15935_),
    .ZN(_08966_));
 AOI21_X1 _27878_ (.A(_08964_),
    .B1(_08966_),
    .B2(_08858_),
    .ZN(_02767_));
 AND3_X1 _27879_ (.A1(_04673_),
    .A2(\cs_registers_i.mhpmcounter[2][19] ),
    .A3(_08952_),
    .ZN(_08967_));
 NAND4_X1 _27880_ (.A1(_07226_),
    .A2(_08914_),
    .A3(_08951_),
    .A4(_08967_),
    .ZN(_08968_));
 NAND3_X1 _27881_ (.A1(_04706_),
    .A2(_08907_),
    .A3(_08968_),
    .ZN(_08969_));
 NAND3_X1 _27882_ (.A1(_08923_),
    .A2(_08951_),
    .A3(_08967_),
    .ZN(_08970_));
 OAI221_X1 _27883_ (.A(_08969_),
    .B1(_08922_),
    .B2(_04721_),
    .C1(_04706_),
    .C2(_08970_),
    .ZN(_02768_));
 INV_X1 _27884_ (.A(_04742_),
    .ZN(_08971_));
 NAND2_X1 _27885_ (.A1(_04706_),
    .A2(_08967_),
    .ZN(_08972_));
 NOR4_X1 _27886_ (.A1(_04736_),
    .A2(_08857_),
    .A3(_08933_),
    .A4(_08972_),
    .ZN(_08973_));
 AOI22_X1 _27887_ (.A1(_08971_),
    .A2(_08935_),
    .B1(_08973_),
    .B2(_08912_),
    .ZN(_08974_));
 NOR3_X1 _27888_ (.A1(_08920_),
    .A2(_08933_),
    .A3(_08972_),
    .ZN(_08975_));
 NAND2_X1 _27889_ (.A1(_04736_),
    .A2(_08884_),
    .ZN(_08976_));
 OAI21_X1 _27890_ (.A(_08974_),
    .B1(_08975_),
    .B2(_08976_),
    .ZN(_02769_));
 AND2_X1 _27891_ (.A1(_04754_),
    .A2(_08844_),
    .ZN(_08977_));
 AND3_X1 _27892_ (.A1(_04706_),
    .A2(_04736_),
    .A3(_08967_),
    .ZN(_08978_));
 NAND2_X1 _27893_ (.A1(_08951_),
    .A2(_08978_),
    .ZN(_08979_));
 OAI21_X1 _27894_ (.A(_08977_),
    .B1(_08979_),
    .B2(_08920_),
    .ZN(_08980_));
 NAND3_X1 _27895_ (.A1(_08923_),
    .A2(_08951_),
    .A3(_08978_),
    .ZN(_08981_));
 OAI221_X1 _27896_ (.A(_08980_),
    .B1(_08922_),
    .B2(_04762_),
    .C1(_04754_),
    .C2(_08981_),
    .ZN(_02770_));
 INV_X1 _27897_ (.A(_04783_),
    .ZN(_08982_));
 INV_X1 _27898_ (.A(\cs_registers_i.mhpmcounter[2][23] ),
    .ZN(_08983_));
 NOR2_X1 _27899_ (.A1(_08983_),
    .A2(_08935_),
    .ZN(_08984_));
 NAND2_X1 _27900_ (.A1(_04754_),
    .A2(_08978_),
    .ZN(_08985_));
 OR4_X1 _27901_ (.A1(_08857_),
    .A2(_08854_),
    .A3(_08933_),
    .A4(_08985_),
    .ZN(_08986_));
 AOI22_X1 _27902_ (.A1(_08982_),
    .A2(_08872_),
    .B1(_08984_),
    .B2(_08986_),
    .ZN(_08987_));
 OAI21_X1 _27903_ (.A(_08987_),
    .B1(_08986_),
    .B2(\cs_registers_i.mhpmcounter[2][23] ),
    .ZN(_02771_));
 NAND3_X1 _27904_ (.A1(_04706_),
    .A2(_04736_),
    .A3(_04754_),
    .ZN(_08988_));
 NAND2_X1 _27905_ (.A1(\cs_registers_i.mhpmcounter[2][23] ),
    .A2(\cs_registers_i.mhpmcounter[2][24] ),
    .ZN(_08989_));
 NOR3_X2 _27906_ (.A1(_08961_),
    .A2(_08988_),
    .A3(_08989_),
    .ZN(_08990_));
 AOI22_X1 _27907_ (.A1(_04804_),
    .A2(_08905_),
    .B1(_08956_),
    .B2(_08990_),
    .ZN(_08991_));
 AOI21_X1 _27908_ (.A(_08991_),
    .B1(_08907_),
    .B2(_08920_),
    .ZN(_08992_));
 NOR2_X1 _27909_ (.A1(\cs_registers_i.mhpmcounter[2][24] ),
    .A2(_08872_),
    .ZN(_08993_));
 OR4_X1 _27910_ (.A1(_08983_),
    .A2(_08915_),
    .A3(_08941_),
    .A4(_08985_),
    .ZN(_08994_));
 AOI21_X1 _27911_ (.A(_08992_),
    .B1(_08993_),
    .B2(_08994_),
    .ZN(_02772_));
 INV_X1 _27912_ (.A(_04816_),
    .ZN(_08995_));
 NAND3_X1 _27913_ (.A1(_08995_),
    .A2(_08939_),
    .A3(_08990_),
    .ZN(_08996_));
 NAND2_X1 _27914_ (.A1(_04816_),
    .A2(_08884_),
    .ZN(_08997_));
 AND2_X1 _27915_ (.A1(_08939_),
    .A2(_08990_),
    .ZN(_08998_));
 OAI221_X1 _27916_ (.A(_08996_),
    .B1(_08997_),
    .B2(_08998_),
    .C1(_08907_),
    .C2(_04822_),
    .ZN(_02773_));
 INV_X1 _27917_ (.A(_04832_),
    .ZN(_08999_));
 CLKBUF_X3 _27918_ (.A(_08857_),
    .Z(_09000_));
 AND4_X1 _27919_ (.A1(_08876_),
    .A2(_04816_),
    .A3(_08932_),
    .A4(_08990_),
    .ZN(_09001_));
 INV_X1 _27920_ (.A(_09001_),
    .ZN(_09002_));
 NOR4_X1 _27921_ (.A1(_08999_),
    .A2(_09000_),
    .A3(_08855_),
    .A4(_09002_),
    .ZN(_09003_));
 NOR2_X1 _27922_ (.A1(_04837_),
    .A2(_08843_),
    .ZN(_09004_));
 AOI221_X2 _27923_ (.A(_09004_),
    .B1(_09001_),
    .B2(_08912_),
    .C1(_04832_),
    .C2(_08843_),
    .ZN(_09005_));
 NOR2_X1 _27924_ (.A1(_09003_),
    .A2(_09005_),
    .ZN(_02774_));
 INV_X1 _27925_ (.A(\cs_registers_i.mhpmcounter[2][27] ),
    .ZN(_09006_));
 NAND2_X1 _27926_ (.A1(_04816_),
    .A2(_08990_),
    .ZN(_09007_));
 OR2_X1 _27927_ (.A1(_08933_),
    .A2(_09007_),
    .ZN(_09008_));
 NOR3_X2 _27928_ (.A1(_08842_),
    .A2(_08853_),
    .A3(_09008_),
    .ZN(_09009_));
 AOI221_X1 _27929_ (.A(_09006_),
    .B1(_04756_),
    .B2(_08871_),
    .C1(_09009_),
    .C2(_04832_),
    .ZN(_09010_));
 NOR2_X1 _27930_ (.A1(_04853_),
    .A2(_08922_),
    .ZN(_09011_));
 AND3_X1 _27931_ (.A1(_04832_),
    .A2(_09006_),
    .A3(_09009_),
    .ZN(_09012_));
 OR3_X1 _27932_ (.A1(_09010_),
    .A2(_09011_),
    .A3(_09012_),
    .ZN(_02775_));
 OR2_X1 _27933_ (.A1(\cs_registers_i.mhpmcounter[2][28] ),
    .A2(_08935_),
    .ZN(_09013_));
 NOR3_X1 _27934_ (.A1(_08999_),
    .A2(_09006_),
    .A3(_09002_),
    .ZN(_09014_));
 AOI21_X1 _27935_ (.A(_09013_),
    .B1(_09014_),
    .B2(_08912_),
    .ZN(_09015_));
 NAND3_X2 _27936_ (.A1(_04832_),
    .A2(\cs_registers_i.mhpmcounter[2][27] ),
    .A3(\cs_registers_i.mhpmcounter[2][28] ),
    .ZN(_09016_));
 NOR3_X2 _27937_ (.A1(_08941_),
    .A2(_09007_),
    .A3(_09016_),
    .ZN(_09017_));
 NAND2_X1 _27938_ (.A1(_08403_),
    .A2(_08904_),
    .ZN(_09018_));
 MUX2_X1 _27939_ (.A(_04867_),
    .B(_09017_),
    .S(_09018_),
    .Z(_09019_));
 NAND2_X1 _27940_ (.A1(_08920_),
    .A2(_08907_),
    .ZN(_09020_));
 AOI21_X1 _27941_ (.A(_09015_),
    .B1(_09019_),
    .B2(_09020_),
    .ZN(_02776_));
 NOR2_X1 _27942_ (.A1(_04885_),
    .A2(_08906_),
    .ZN(_09021_));
 NOR2_X1 _27943_ (.A1(_04880_),
    .A2(_09016_),
    .ZN(_09022_));
 AOI21_X1 _27944_ (.A(_09021_),
    .B1(_09022_),
    .B2(_09009_),
    .ZN(_09023_));
 NOR3_X1 _27945_ (.A1(_08920_),
    .A2(_09008_),
    .A3(_09016_),
    .ZN(_09024_));
 NAND2_X1 _27946_ (.A1(_04880_),
    .A2(_08884_),
    .ZN(_09025_));
 OAI21_X1 _27947_ (.A(_09023_),
    .B1(_09024_),
    .B2(_09025_),
    .ZN(_02777_));
 NAND2_X1 _27948_ (.A1(_06560_),
    .A2(_08844_),
    .ZN(_09026_));
 NAND3_X2 _27949_ (.A1(_08876_),
    .A2(_07226_),
    .A3(_08914_),
    .ZN(_09027_));
 MUX2_X1 _27950_ (.A(_06560_),
    .B(_09026_),
    .S(_09027_),
    .Z(_09028_));
 INV_X2 _27951_ (.A(_08401_),
    .ZN(_09029_));
 OAI21_X1 _27952_ (.A(_09028_),
    .B1(_08907_),
    .B2(_09029_),
    .ZN(_02778_));
 AND2_X1 _27953_ (.A1(\cs_registers_i.mhpmcounter[2][30] ),
    .A2(_08844_),
    .ZN(_09030_));
 NAND2_X1 _27954_ (.A1(_04880_),
    .A2(_09017_),
    .ZN(_09031_));
 OAI21_X1 _27955_ (.A(_09030_),
    .B1(_09031_),
    .B2(_08920_),
    .ZN(_09032_));
 NAND3_X1 _27956_ (.A1(_04880_),
    .A2(_08923_),
    .A3(_09017_),
    .ZN(_09033_));
 OAI221_X1 _27957_ (.A(_09032_),
    .B1(_08922_),
    .B2(_04905_),
    .C1(\cs_registers_i.mhpmcounter[2][30] ),
    .C2(_09033_),
    .ZN(_02779_));
 INV_X1 _27958_ (.A(\cs_registers_i.mhpmcounter[2][31] ),
    .ZN(_09034_));
 NAND2_X1 _27959_ (.A1(_04880_),
    .A2(\cs_registers_i.mhpmcounter[2][30] ),
    .ZN(_09035_));
 NOR2_X1 _27960_ (.A1(_09016_),
    .A2(_09035_),
    .ZN(_09036_));
 AOI221_X1 _27961_ (.A(_09034_),
    .B1(_04756_),
    .B2(_08871_),
    .C1(_09009_),
    .C2(_09036_),
    .ZN(_09037_));
 NOR2_X1 _27962_ (.A1(_04924_),
    .A2(_08922_),
    .ZN(_09038_));
 AND3_X1 _27963_ (.A1(_09034_),
    .A2(_09009_),
    .A3(_09036_),
    .ZN(_09039_));
 OR3_X1 _27964_ (.A1(_09037_),
    .A2(_09038_),
    .A3(_09039_),
    .ZN(_02780_));
 NAND2_X1 _27965_ (.A1(\cs_registers_i.mhpmcounter[2][31] ),
    .A2(_09036_),
    .ZN(_09040_));
 OR3_X2 _27966_ (.A1(_08941_),
    .A2(_09007_),
    .A3(_09040_),
    .ZN(_09041_));
 AND3_X1 _27967_ (.A1(_05347_),
    .A2(_08895_),
    .A3(_09041_),
    .ZN(_09042_));
 INV_X1 _27968_ (.A(_05347_),
    .ZN(_09043_));
 BUF_X4 _27969_ (.A(_08835_),
    .Z(_09044_));
 CLKBUF_X3 _27970_ (.A(_08840_),
    .Z(_09045_));
 AOI21_X1 _27971_ (.A(_09043_),
    .B1(_09044_),
    .B2(_09045_),
    .ZN(_09046_));
 OAI21_X4 _27972_ (.A(_04588_),
    .B1(_08842_),
    .B2(_08849_),
    .ZN(_09047_));
 OAI21_X4 _27973_ (.A(_09047_),
    .B1(_07245_),
    .B2(_07224_),
    .ZN(_09048_));
 CLKBUF_X3 _27974_ (.A(_09048_),
    .Z(_09049_));
 AOI221_X1 _27975_ (.A(_09042_),
    .B1(_09046_),
    .B2(_08855_),
    .C1(_09049_),
    .C2(_05347_),
    .ZN(_09050_));
 NAND2_X1 _27976_ (.A1(_08835_),
    .A2(_08840_),
    .ZN(_09051_));
 BUF_X2 _27977_ (.A(_09051_),
    .Z(_09052_));
 AOI21_X1 _27978_ (.A(_09048_),
    .B1(_09052_),
    .B2(_08854_),
    .ZN(_09053_));
 CLKBUF_X3 _27979_ (.A(_09053_),
    .Z(_09054_));
 CLKBUF_X3 _27980_ (.A(_08857_),
    .Z(_09055_));
 NOR3_X1 _27981_ (.A1(_05347_),
    .A2(_09055_),
    .A3(_09041_),
    .ZN(_09056_));
 OAI21_X1 _27982_ (.A(_09054_),
    .B1(_09056_),
    .B2(_08863_),
    .ZN(_09057_));
 NAND2_X1 _27983_ (.A1(_09050_),
    .A2(_09057_),
    .ZN(_02781_));
 BUF_X2 _27984_ (.A(_09051_),
    .Z(_09058_));
 AND3_X1 _27985_ (.A1(_06493_),
    .A2(_08854_),
    .A3(_09058_),
    .ZN(_09059_));
 OR3_X1 _27986_ (.A1(_09043_),
    .A2(_09008_),
    .A3(_09040_),
    .ZN(_09060_));
 AND2_X1 _27987_ (.A1(_06493_),
    .A2(_09060_),
    .ZN(_09061_));
 CLKBUF_X3 _27988_ (.A(_09048_),
    .Z(_09062_));
 AOI221_X1 _27989_ (.A(_09059_),
    .B1(_09061_),
    .B2(_08862_),
    .C1(_06493_),
    .C2(_09062_),
    .ZN(_09063_));
 NOR3_X1 _27990_ (.A1(_06493_),
    .A2(_09055_),
    .A3(_09060_),
    .ZN(_09064_));
 OAI21_X1 _27991_ (.A(_09054_),
    .B1(_09064_),
    .B2(_08965_),
    .ZN(_09065_));
 NAND2_X1 _27992_ (.A1(_09063_),
    .A2(_09065_),
    .ZN(_02782_));
 BUF_X2 _27993_ (.A(_08861_),
    .Z(_09066_));
 NOR2_X1 _27994_ (.A1(_09043_),
    .A2(_09040_),
    .ZN(_09067_));
 NAND3_X1 _27995_ (.A1(_06493_),
    .A2(_09001_),
    .A3(_09067_),
    .ZN(_09068_));
 AND3_X1 _27996_ (.A1(_06548_),
    .A2(_09066_),
    .A3(_09068_),
    .ZN(_09069_));
 INV_X1 _27997_ (.A(_06548_),
    .ZN(_09070_));
 AOI21_X1 _27998_ (.A(_09070_),
    .B1(_08835_),
    .B2(_09045_),
    .ZN(_09071_));
 BUF_X4 _27999_ (.A(_08854_),
    .Z(_09072_));
 BUF_X4 _28000_ (.A(_09048_),
    .Z(_09073_));
 AOI221_X1 _28001_ (.A(_09069_),
    .B1(_09071_),
    .B2(_09072_),
    .C1(_09073_),
    .C2(_06548_),
    .ZN(_09074_));
 NOR3_X1 _28002_ (.A1(_06548_),
    .A2(_08886_),
    .A3(_09068_),
    .ZN(_09075_));
 AOI21_X1 _28003_ (.A(_09075_),
    .B1(_09000_),
    .B2(_08402_),
    .ZN(_09076_));
 NAND2_X1 _28004_ (.A1(_08855_),
    .A2(_09052_),
    .ZN(_09077_));
 NAND3_X4 _28005_ (.A1(_08043_),
    .A2(_09047_),
    .A3(_09077_),
    .ZN(_09078_));
 OAI21_X1 _28006_ (.A(_09074_),
    .B1(_09076_),
    .B2(_09078_),
    .ZN(_02783_));
 AND3_X1 _28007_ (.A1(_06598_),
    .A2(_08854_),
    .A3(_09058_),
    .ZN(_09079_));
 NAND2_X1 _28008_ (.A1(_06493_),
    .A2(_06548_),
    .ZN(_09080_));
 OR2_X1 _28009_ (.A1(_09060_),
    .A2(_09080_),
    .ZN(_09081_));
 AND2_X1 _28010_ (.A1(_06598_),
    .A2(_09081_),
    .ZN(_09082_));
 AOI221_X1 _28011_ (.A(_09079_),
    .B1(_09082_),
    .B2(_08862_),
    .C1(_06598_),
    .C2(_09062_),
    .ZN(_09083_));
 NOR3_X1 _28012_ (.A1(_06598_),
    .A2(_09055_),
    .A3(_09081_),
    .ZN(_09084_));
 NOR2_X1 _28013_ (.A1(_08629_),
    .A2(_08864_),
    .ZN(_09085_));
 OAI21_X1 _28014_ (.A(_09054_),
    .B1(_09084_),
    .B2(_09085_),
    .ZN(_09086_));
 NAND2_X1 _28015_ (.A1(_09083_),
    .A2(_09086_),
    .ZN(_02784_));
 INV_X1 _28016_ (.A(\cs_registers_i.mhpmcounter[2][36] ),
    .ZN(_09087_));
 NAND2_X1 _28017_ (.A1(_09087_),
    .A2(_09049_),
    .ZN(_09088_));
 NOR2_X1 _28018_ (.A1(_09070_),
    .A2(_09068_),
    .ZN(_09089_));
 AOI21_X1 _28019_ (.A(\cs_registers_i.mhpmcounter[2][36] ),
    .B1(_09089_),
    .B2(_06598_),
    .ZN(_09090_));
 NAND2_X1 _28020_ (.A1(_08896_),
    .A2(_09090_),
    .ZN(_09091_));
 NAND3_X1 _28021_ (.A1(_09087_),
    .A2(_08855_),
    .A3(_09052_),
    .ZN(_09092_));
 NAND3_X1 _28022_ (.A1(_09088_),
    .A2(_09091_),
    .A3(_09092_),
    .ZN(_09093_));
 NAND2_X1 _28023_ (.A1(_06598_),
    .A2(\cs_registers_i.mhpmcounter[2][36] ),
    .ZN(_09094_));
 NOR4_X2 _28024_ (.A1(_09043_),
    .A2(_09041_),
    .A3(_09080_),
    .A4(_09094_),
    .ZN(_09095_));
 MUX2_X1 _28025_ (.A(_08639_),
    .B(_09095_),
    .S(_08862_),
    .Z(_09096_));
 AOI21_X1 _28026_ (.A(_09093_),
    .B1(_09096_),
    .B2(_09054_),
    .ZN(_02785_));
 INV_X1 _28027_ (.A(_05521_),
    .ZN(_09097_));
 NOR2_X2 _28028_ (.A1(_09081_),
    .A2(_09094_),
    .ZN(_09098_));
 NOR3_X1 _28029_ (.A1(_09097_),
    .A2(_08857_),
    .A3(_09098_),
    .ZN(_09099_));
 AOI21_X1 _28030_ (.A(_09097_),
    .B1(_09044_),
    .B2(_09045_),
    .ZN(_09100_));
 AOI221_X1 _28031_ (.A(_09099_),
    .B1(_09100_),
    .B2(_08855_),
    .C1(_09049_),
    .C2(_05521_),
    .ZN(_09101_));
 NAND2_X1 _28032_ (.A1(_08862_),
    .A2(_09098_),
    .ZN(_09102_));
 OAI22_X1 _28033_ (.A1(_08646_),
    .A2(_08864_),
    .B1(_09102_),
    .B2(_05521_),
    .ZN(_09103_));
 NAND2_X1 _28034_ (.A1(_09054_),
    .A2(_09103_),
    .ZN(_09104_));
 NAND2_X1 _28035_ (.A1(_09101_),
    .A2(_09104_),
    .ZN(_02786_));
 NAND2_X1 _28036_ (.A1(_05521_),
    .A2(_09095_),
    .ZN(_09105_));
 AND3_X1 _28037_ (.A1(_05604_),
    .A2(_08895_),
    .A3(_09105_),
    .ZN(_09106_));
 AND2_X1 _28038_ (.A1(_05604_),
    .A2(_09052_),
    .ZN(_09107_));
 AOI221_X1 _28039_ (.A(_09106_),
    .B1(_09107_),
    .B2(_08855_),
    .C1(_09049_),
    .C2(_05604_),
    .ZN(_09108_));
 NOR3_X1 _28040_ (.A1(_05604_),
    .A2(_09055_),
    .A3(_09105_),
    .ZN(_09109_));
 NOR2_X1 _28041_ (.A1(_08655_),
    .A2(_08864_),
    .ZN(_09110_));
 OAI21_X1 _28042_ (.A(_09054_),
    .B1(_09109_),
    .B2(_09110_),
    .ZN(_09111_));
 NAND2_X1 _28043_ (.A1(_09108_),
    .A2(_09111_),
    .ZN(_02787_));
 AND2_X1 _28044_ (.A1(_05691_),
    .A2(_09048_),
    .ZN(_09112_));
 NAND2_X1 _28045_ (.A1(_05521_),
    .A2(_05604_),
    .ZN(_09113_));
 INV_X1 _28046_ (.A(_09113_),
    .ZN(_09114_));
 AOI21_X1 _28047_ (.A(_08856_),
    .B1(_09098_),
    .B2(_09114_),
    .ZN(_09115_));
 AND2_X1 _28048_ (.A1(_05691_),
    .A2(_09052_),
    .ZN(_09116_));
 AOI221_X1 _28049_ (.A(_09112_),
    .B1(_09115_),
    .B2(_05691_),
    .C1(_09116_),
    .C2(_08855_),
    .ZN(_09117_));
 NOR3_X1 _28050_ (.A1(_05691_),
    .A2(_09102_),
    .A3(_09113_),
    .ZN(_09118_));
 AOI21_X1 _28051_ (.A(_09118_),
    .B1(_09000_),
    .B2(_08666_),
    .ZN(_09119_));
 OAI21_X1 _28052_ (.A(_09117_),
    .B1(_09119_),
    .B2(_09078_),
    .ZN(_02788_));
 AND2_X1 _28053_ (.A1(_06596_),
    .A2(_08844_),
    .ZN(_09120_));
 NAND2_X1 _28054_ (.A1(_06560_),
    .A2(_08892_),
    .ZN(_09121_));
 OAI21_X1 _28055_ (.A(_09120_),
    .B1(_09121_),
    .B2(_08920_),
    .ZN(_09122_));
 NAND3_X1 _28056_ (.A1(_06560_),
    .A2(_08923_),
    .A3(_08892_),
    .ZN(_09123_));
 OAI221_X1 _28057_ (.A(_09122_),
    .B1(_08922_),
    .B2(_08629_),
    .C1(_06596_),
    .C2(_09123_),
    .ZN(_02789_));
 NAND3_X1 _28058_ (.A1(_05691_),
    .A2(_09095_),
    .A3(_09114_),
    .ZN(_09124_));
 AND3_X1 _28059_ (.A1(_04929_),
    .A2(_08895_),
    .A3(_09124_),
    .ZN(_09125_));
 AND2_X1 _28060_ (.A1(_04929_),
    .A2(_09052_),
    .ZN(_09126_));
 AOI221_X1 _28061_ (.A(_09125_),
    .B1(_09126_),
    .B2(_08855_),
    .C1(_09049_),
    .C2(_04929_),
    .ZN(_09127_));
 NOR3_X1 _28062_ (.A1(_04929_),
    .A2(_09055_),
    .A3(_09124_),
    .ZN(_09128_));
 NOR2_X1 _28063_ (.A1(_04942_),
    .A2(_08864_),
    .ZN(_09129_));
 OAI21_X1 _28064_ (.A(_09054_),
    .B1(_09128_),
    .B2(_09129_),
    .ZN(_09130_));
 NAND2_X1 _28065_ (.A1(_09127_),
    .A2(_09130_),
    .ZN(_02790_));
 NAND4_X2 _28066_ (.A1(_05691_),
    .A2(_04929_),
    .A3(_09098_),
    .A4(_09114_),
    .ZN(_09131_));
 AND3_X1 _28067_ (.A1(_04946_),
    .A2(_08895_),
    .A3(_09131_),
    .ZN(_09132_));
 AND2_X1 _28068_ (.A1(_04946_),
    .A2(_09052_),
    .ZN(_09133_));
 BUF_X4 _28069_ (.A(_08854_),
    .Z(_09134_));
 AOI221_X2 _28070_ (.A(_09132_),
    .B1(_09133_),
    .B2(_09134_),
    .C1(_09049_),
    .C2(_04946_),
    .ZN(_09135_));
 CLKBUF_X3 _28071_ (.A(_09053_),
    .Z(_09136_));
 NOR2_X1 _28072_ (.A1(_04960_),
    .A2(_08896_),
    .ZN(_09137_));
 NOR3_X1 _28073_ (.A1(_04946_),
    .A2(_08886_),
    .A3(_09131_),
    .ZN(_09138_));
 OAI21_X1 _28074_ (.A(_09136_),
    .B1(_09137_),
    .B2(_09138_),
    .ZN(_09139_));
 NAND2_X1 _28075_ (.A1(_09135_),
    .A2(_09139_),
    .ZN(_02791_));
 INV_X1 _28076_ (.A(_09124_),
    .ZN(_09140_));
 NAND3_X2 _28077_ (.A1(_04929_),
    .A2(_04946_),
    .A3(_09140_),
    .ZN(_09141_));
 AND3_X1 _28078_ (.A1(_05830_),
    .A2(_09066_),
    .A3(_09141_),
    .ZN(_09142_));
 INV_X1 _28079_ (.A(_05830_),
    .ZN(_09143_));
 AOI21_X1 _28080_ (.A(_09143_),
    .B1(_08835_),
    .B2(_09045_),
    .ZN(_09144_));
 AOI221_X2 _28081_ (.A(_09142_),
    .B1(_09144_),
    .B2(_09072_),
    .C1(_09073_),
    .C2(_05830_),
    .ZN(_09145_));
 NOR3_X1 _28082_ (.A1(_05830_),
    .A2(_08886_),
    .A3(_09141_),
    .ZN(_09146_));
 AOI21_X1 _28083_ (.A(_09146_),
    .B1(_09000_),
    .B2(_08867_),
    .ZN(_09147_));
 OAI21_X1 _28084_ (.A(_09145_),
    .B1(_09147_),
    .B2(_09078_),
    .ZN(_02792_));
 NAND2_X1 _28085_ (.A1(_04946_),
    .A2(_05830_),
    .ZN(_09148_));
 OR2_X2 _28086_ (.A1(_09131_),
    .A2(_09148_),
    .ZN(_09149_));
 AND3_X1 _28087_ (.A1(_04394_),
    .A2(_08895_),
    .A3(_09149_),
    .ZN(_09150_));
 INV_X2 _28088_ (.A(_04394_),
    .ZN(_09151_));
 AOI21_X1 _28089_ (.A(_09151_),
    .B1(_09044_),
    .B2(_09045_),
    .ZN(_09152_));
 AOI221_X2 _28090_ (.A(_09150_),
    .B1(_09152_),
    .B2(_09134_),
    .C1(_09049_),
    .C2(_04394_),
    .ZN(_09153_));
 NOR3_X1 _28091_ (.A1(_04394_),
    .A2(_09055_),
    .A3(_09149_),
    .ZN(_09154_));
 OAI21_X1 _28092_ (.A(_09136_),
    .B1(_09154_),
    .B2(_08897_),
    .ZN(_09155_));
 NAND2_X1 _28093_ (.A1(_09153_),
    .A2(_09155_),
    .ZN(_02793_));
 NOR3_X2 _28094_ (.A1(_09151_),
    .A2(_09143_),
    .A3(_09141_),
    .ZN(_09156_));
 AND2_X1 _28095_ (.A1(\cs_registers_i.mhpmcounter[2][44] ),
    .A2(_09156_),
    .ZN(_09157_));
 MUX2_X1 _28096_ (.A(_04527_),
    .B(_09157_),
    .S(_08895_),
    .Z(_09158_));
 AND2_X1 _28097_ (.A1(_09053_),
    .A2(_09158_),
    .ZN(_09159_));
 OR2_X1 _28098_ (.A1(_08871_),
    .A2(_09156_),
    .ZN(_09160_));
 NOR2_X2 _28099_ (.A1(\id_stage_i.branch_set_d ),
    .A2(_08873_),
    .ZN(_09161_));
 OAI221_X2 _28100_ (.A(_09160_),
    .B1(_08869_),
    .B2(_09161_),
    .C1(_08427_),
    .C2(_08923_),
    .ZN(_09162_));
 INV_X1 _28101_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .ZN(_09163_));
 AOI21_X1 _28102_ (.A(_09159_),
    .B1(_09162_),
    .B2(_09163_),
    .ZN(_02794_));
 INV_X1 _28103_ (.A(_04547_),
    .ZN(_09164_));
 NOR3_X4 _28104_ (.A1(_09163_),
    .A2(_09151_),
    .A3(_09149_),
    .ZN(_09165_));
 NOR3_X1 _28105_ (.A1(_09164_),
    .A2(_08856_),
    .A3(_09165_),
    .ZN(_09166_));
 AOI21_X1 _28106_ (.A(_09164_),
    .B1(_09044_),
    .B2(_09045_),
    .ZN(_09167_));
 AOI221_X1 _28107_ (.A(_09166_),
    .B1(_09167_),
    .B2(_09134_),
    .C1(_09049_),
    .C2(_04547_),
    .ZN(_09168_));
 NAND2_X1 _28108_ (.A1(_08862_),
    .A2(_09165_),
    .ZN(_09169_));
 OAI22_X1 _28109_ (.A1(_04562_),
    .A2(_08864_),
    .B1(_09169_),
    .B2(_04547_),
    .ZN(_09170_));
 NAND2_X1 _28110_ (.A1(_09054_),
    .A2(_09170_),
    .ZN(_09171_));
 NAND2_X1 _28111_ (.A1(_09168_),
    .A2(_09171_),
    .ZN(_02795_));
 NAND2_X1 _28112_ (.A1(_04547_),
    .A2(_09157_),
    .ZN(_09172_));
 AND3_X1 _28113_ (.A1(_04593_),
    .A2(_08895_),
    .A3(_09172_),
    .ZN(_09173_));
 AND2_X1 _28114_ (.A1(_04593_),
    .A2(_09052_),
    .ZN(_09174_));
 AOI221_X1 _28115_ (.A(_09173_),
    .B1(_09174_),
    .B2(_09134_),
    .C1(_09049_),
    .C2(_04593_),
    .ZN(_09175_));
 NOR3_X1 _28116_ (.A1(_04593_),
    .A2(_09055_),
    .A3(_09172_),
    .ZN(_09176_));
 NOR2_X1 _28117_ (.A1(_04597_),
    .A2(_08896_),
    .ZN(_09177_));
 OAI21_X1 _28118_ (.A(_09136_),
    .B1(_09176_),
    .B2(_09177_),
    .ZN(_09178_));
 NAND2_X1 _28119_ (.A1(_09175_),
    .A2(_09178_),
    .ZN(_02796_));
 AND2_X2 _28120_ (.A1(_04547_),
    .A2(_04593_),
    .ZN(_09179_));
 AOI21_X1 _28121_ (.A(_08856_),
    .B1(_09165_),
    .B2(_09179_),
    .ZN(_09180_));
 AND2_X1 _28122_ (.A1(_04603_),
    .A2(_09180_),
    .ZN(_09181_));
 AND2_X1 _28123_ (.A1(_04603_),
    .A2(_09058_),
    .ZN(_09182_));
 AOI221_X1 _28124_ (.A(_09181_),
    .B1(_09182_),
    .B2(_09072_),
    .C1(_09073_),
    .C2(_04603_),
    .ZN(_09183_));
 NAND2_X1 _28125_ (.A1(_04547_),
    .A2(_04593_),
    .ZN(_09184_));
 NOR3_X1 _28126_ (.A1(_04603_),
    .A2(_09169_),
    .A3(_09184_),
    .ZN(_09185_));
 AOI21_X1 _28127_ (.A(_09185_),
    .B1(_09000_),
    .B2(_08936_),
    .ZN(_09186_));
 OAI21_X1 _28128_ (.A(_09183_),
    .B1(_09186_),
    .B2(_09078_),
    .ZN(_02797_));
 NAND3_X2 _28129_ (.A1(_04603_),
    .A2(_09157_),
    .A3(_09179_),
    .ZN(_09187_));
 AND3_X1 _28130_ (.A1(_04624_),
    .A2(_08895_),
    .A3(_09187_),
    .ZN(_09188_));
 INV_X1 _28131_ (.A(_04624_),
    .ZN(_09189_));
 AOI21_X1 _28132_ (.A(_09189_),
    .B1(_09044_),
    .B2(_09045_),
    .ZN(_09190_));
 AOI221_X1 _28133_ (.A(_09188_),
    .B1(_09190_),
    .B2(_09134_),
    .C1(_09049_),
    .C2(_04624_),
    .ZN(_09191_));
 NOR3_X1 _28134_ (.A1(_04624_),
    .A2(_09055_),
    .A3(_09187_),
    .ZN(_09192_));
 NOR2_X1 _28135_ (.A1(_04645_),
    .A2(_08896_),
    .ZN(_09193_));
 OAI21_X1 _28136_ (.A(_09136_),
    .B1(_09192_),
    .B2(_09193_),
    .ZN(_09194_));
 NAND2_X1 _28137_ (.A1(_09191_),
    .A2(_09194_),
    .ZN(_02798_));
 NAND4_X4 _28138_ (.A1(_04603_),
    .A2(_04624_),
    .A3(_09165_),
    .A4(_09179_),
    .ZN(_09195_));
 AND3_X1 _28139_ (.A1(_04662_),
    .A2(_09066_),
    .A3(_09195_),
    .ZN(_09196_));
 AND2_X1 _28140_ (.A1(_04662_),
    .A2(_09058_),
    .ZN(_09197_));
 AOI221_X1 _28141_ (.A(_09196_),
    .B1(_09197_),
    .B2(_09072_),
    .C1(_09073_),
    .C2(_04662_),
    .ZN(_09198_));
 NOR3_X1 _28142_ (.A1(_04662_),
    .A2(_08886_),
    .A3(_09195_),
    .ZN(_09199_));
 INV_X2 _28143_ (.A(_04665_),
    .ZN(_09200_));
 AOI21_X1 _28144_ (.A(_09199_),
    .B1(_09000_),
    .B2(_09200_),
    .ZN(_09201_));
 OAI21_X1 _28145_ (.A(_09198_),
    .B1(_09201_),
    .B2(_09078_),
    .ZN(_02799_));
 NAND2_X1 _28146_ (.A1(_06560_),
    .A2(_06596_),
    .ZN(_09202_));
 OAI221_X1 _28147_ (.A(\cs_registers_i.mhpmcounter[2][4] ),
    .B1(_08427_),
    .B2(_09018_),
    .C1(_09202_),
    .C2(_09027_),
    .ZN(_09203_));
 OR2_X1 _28148_ (.A1(\cs_registers_i.mhpmcounter[2][4] ),
    .A2(_09202_),
    .ZN(_09204_));
 OAI221_X1 _28149_ (.A(_09203_),
    .B1(_09204_),
    .B2(_09027_),
    .C1(_08907_),
    .C2(_08639_),
    .ZN(_02800_));
 NOR2_X2 _28150_ (.A1(_09189_),
    .A2(_09187_),
    .ZN(_09205_));
 AOI21_X1 _28151_ (.A(_08842_),
    .B1(_09205_),
    .B2(_04662_),
    .ZN(_09206_));
 AND2_X1 _28152_ (.A1(_04671_),
    .A2(_09206_),
    .ZN(_09207_));
 INV_X1 _28153_ (.A(_04671_),
    .ZN(_09208_));
 AOI21_X1 _28154_ (.A(_09208_),
    .B1(_08835_),
    .B2(_09045_),
    .ZN(_09209_));
 AOI221_X2 _28155_ (.A(_09207_),
    .B1(_09209_),
    .B2(_09072_),
    .C1(_09073_),
    .C2(_04671_),
    .ZN(_09210_));
 AND4_X1 _28156_ (.A1(_04603_),
    .A2(_04624_),
    .A3(_09157_),
    .A4(_09179_),
    .ZN(_09211_));
 NAND3_X1 _28157_ (.A1(_04662_),
    .A2(_09208_),
    .A3(_09211_),
    .ZN(_09212_));
 MUX2_X1 _28158_ (.A(_09212_),
    .B(_04685_),
    .S(_08871_),
    .Z(_09213_));
 OAI22_X4 _28159_ (.A1(_09161_),
    .A2(_08869_),
    .B1(_08923_),
    .B2(_08427_),
    .ZN(_09214_));
 OAI21_X1 _28160_ (.A(_09210_),
    .B1(_09213_),
    .B2(_09214_),
    .ZN(_02801_));
 INV_X1 _28161_ (.A(_04697_),
    .ZN(_09215_));
 NAND2_X1 _28162_ (.A1(_04662_),
    .A2(_04671_),
    .ZN(_09216_));
 NOR2_X1 _28163_ (.A1(_09195_),
    .A2(_09216_),
    .ZN(_09217_));
 NOR3_X1 _28164_ (.A1(_09215_),
    .A2(_08856_),
    .A3(_09217_),
    .ZN(_09218_));
 AND2_X1 _28165_ (.A1(_04697_),
    .A2(_09058_),
    .ZN(_09219_));
 AOI221_X1 _28166_ (.A(_09218_),
    .B1(_09219_),
    .B2(_09072_),
    .C1(_09073_),
    .C2(_04697_),
    .ZN(_09220_));
 NOR4_X1 _28167_ (.A1(_04697_),
    .A2(_08857_),
    .A3(_09195_),
    .A4(_09216_),
    .ZN(_09221_));
 INV_X1 _28168_ (.A(_04700_),
    .ZN(_09222_));
 AOI21_X1 _28169_ (.A(_09221_),
    .B1(_09000_),
    .B2(_09222_),
    .ZN(_09223_));
 OAI21_X1 _28170_ (.A(_09220_),
    .B1(_09223_),
    .B2(_09078_),
    .ZN(_02802_));
 AND3_X1 _28171_ (.A1(_04662_),
    .A2(_04671_),
    .A3(_04697_),
    .ZN(_09224_));
 AOI21_X1 _28172_ (.A(_08842_),
    .B1(_09205_),
    .B2(_09224_),
    .ZN(_09225_));
 AND2_X1 _28173_ (.A1(_04703_),
    .A2(_09225_),
    .ZN(_09226_));
 INV_X1 _28174_ (.A(_04703_),
    .ZN(_09227_));
 AOI21_X1 _28175_ (.A(_09227_),
    .B1(_08835_),
    .B2(_08840_),
    .ZN(_09228_));
 AOI221_X2 _28176_ (.A(_09226_),
    .B1(_09228_),
    .B2(_09072_),
    .C1(_09073_),
    .C2(_04703_),
    .ZN(_09229_));
 NAND3_X1 _28177_ (.A1(_09227_),
    .A2(_09211_),
    .A3(_09224_),
    .ZN(_09230_));
 MUX2_X1 _28178_ (.A(_09230_),
    .B(_04720_),
    .S(_08871_),
    .Z(_09231_));
 OAI21_X1 _28179_ (.A(_09229_),
    .B1(_09231_),
    .B2(_09214_),
    .ZN(_02803_));
 INV_X1 _28180_ (.A(_09195_),
    .ZN(_09232_));
 NAND3_X1 _28181_ (.A1(_04703_),
    .A2(_09232_),
    .A3(_09224_),
    .ZN(_09233_));
 AND3_X1 _28182_ (.A1(_04739_),
    .A2(_09066_),
    .A3(_09233_),
    .ZN(_09234_));
 AND2_X1 _28183_ (.A1(_04739_),
    .A2(_09058_),
    .ZN(_09235_));
 AOI221_X1 _28184_ (.A(_09234_),
    .B1(_09235_),
    .B2(_08854_),
    .C1(_09073_),
    .C2(_04739_),
    .ZN(_09236_));
 NOR3_X1 _28185_ (.A1(_04739_),
    .A2(_08871_),
    .A3(_09233_),
    .ZN(_09237_));
 AOI21_X1 _28186_ (.A(_09237_),
    .B1(_09000_),
    .B2(_08971_),
    .ZN(_09238_));
 OAI21_X1 _28187_ (.A(_09236_),
    .B1(_09238_),
    .B2(_09078_),
    .ZN(_02804_));
 AND3_X1 _28188_ (.A1(_04703_),
    .A2(_04739_),
    .A3(_09224_),
    .ZN(_09239_));
 AOI21_X1 _28189_ (.A(_08856_),
    .B1(_09205_),
    .B2(_09239_),
    .ZN(_09240_));
 AND2_X1 _28190_ (.A1(_04758_),
    .A2(_09240_),
    .ZN(_09241_));
 INV_X1 _28191_ (.A(_04758_),
    .ZN(_09242_));
 AOI21_X1 _28192_ (.A(_09242_),
    .B1(_09044_),
    .B2(_09045_),
    .ZN(_09243_));
 AOI221_X1 _28193_ (.A(_09241_),
    .B1(_09243_),
    .B2(_09134_),
    .C1(_09062_),
    .C2(_04758_),
    .ZN(_09244_));
 NAND4_X1 _28194_ (.A1(_09242_),
    .A2(_08862_),
    .A3(_09205_),
    .A4(_09239_),
    .ZN(_09245_));
 OAI21_X1 _28195_ (.A(_09245_),
    .B1(_08864_),
    .B2(_04762_),
    .ZN(_09246_));
 NAND2_X1 _28196_ (.A1(_09054_),
    .A2(_09246_),
    .ZN(_09247_));
 NAND2_X1 _28197_ (.A1(_09244_),
    .A2(_09247_),
    .ZN(_02805_));
 NAND2_X1 _28198_ (.A1(_04758_),
    .A2(_09239_),
    .ZN(_09248_));
 OR2_X2 _28199_ (.A1(_09195_),
    .A2(_09248_),
    .ZN(_09249_));
 AND3_X1 _28200_ (.A1(_04777_),
    .A2(_09066_),
    .A3(_09249_),
    .ZN(_09250_));
 AND2_X1 _28201_ (.A1(_04777_),
    .A2(_09052_),
    .ZN(_09251_));
 AOI221_X1 _28202_ (.A(_09250_),
    .B1(_09251_),
    .B2(_09134_),
    .C1(_09062_),
    .C2(_04777_),
    .ZN(_09252_));
 NOR3_X1 _28203_ (.A1(_04777_),
    .A2(_09055_),
    .A3(_09249_),
    .ZN(_09253_));
 NOR2_X1 _28204_ (.A1(_04783_),
    .A2(_08896_),
    .ZN(_09254_));
 OAI21_X1 _28205_ (.A(_09136_),
    .B1(_09253_),
    .B2(_09254_),
    .ZN(_09255_));
 NAND2_X1 _28206_ (.A1(_09252_),
    .A2(_09255_),
    .ZN(_02806_));
 NOR3_X2 _28207_ (.A1(_09189_),
    .A2(_09187_),
    .A3(_09248_),
    .ZN(_09256_));
 NAND2_X1 _28208_ (.A1(_04777_),
    .A2(_09256_),
    .ZN(_09257_));
 AND3_X1 _28209_ (.A1(_04789_),
    .A2(_09066_),
    .A3(_09257_),
    .ZN(_09258_));
 AND2_X1 _28210_ (.A1(_04789_),
    .A2(_09052_),
    .ZN(_09259_));
 AOI221_X1 _28211_ (.A(_09258_),
    .B1(_09259_),
    .B2(_09134_),
    .C1(_09062_),
    .C2(_04789_),
    .ZN(_09260_));
 NOR3_X1 _28212_ (.A1(_04789_),
    .A2(_09055_),
    .A3(_09257_),
    .ZN(_09261_));
 NOR2_X1 _28213_ (.A1(_04805_),
    .A2(_08864_),
    .ZN(_09262_));
 OAI21_X1 _28214_ (.A(_09136_),
    .B1(_09261_),
    .B2(_09262_),
    .ZN(_09263_));
 NAND2_X1 _28215_ (.A1(_09260_),
    .A2(_09263_),
    .ZN(_02807_));
 INV_X1 _28216_ (.A(_04819_),
    .ZN(_09264_));
 NAND2_X1 _28217_ (.A1(_04777_),
    .A2(_04789_),
    .ZN(_09265_));
 NOR2_X1 _28218_ (.A1(_09249_),
    .A2(_09265_),
    .ZN(_09266_));
 NOR3_X1 _28219_ (.A1(_09264_),
    .A2(_08856_),
    .A3(_09266_),
    .ZN(_09267_));
 AND2_X1 _28220_ (.A1(_04819_),
    .A2(_09051_),
    .ZN(_09268_));
 AOI221_X2 _28221_ (.A(_09267_),
    .B1(_09268_),
    .B2(_08854_),
    .C1(_09073_),
    .C2(_04819_),
    .ZN(_09269_));
 NOR4_X1 _28222_ (.A1(_04819_),
    .A2(_08857_),
    .A3(_09249_),
    .A4(_09265_),
    .ZN(_09270_));
 INV_X1 _28223_ (.A(_04822_),
    .ZN(_09271_));
 AOI21_X1 _28224_ (.A(_09270_),
    .B1(_09000_),
    .B2(_09271_),
    .ZN(_09272_));
 OAI21_X1 _28225_ (.A(_09269_),
    .B1(_09272_),
    .B2(_09078_),
    .ZN(_02808_));
 NAND4_X1 _28226_ (.A1(_04777_),
    .A2(_04789_),
    .A3(_04819_),
    .A4(_09256_),
    .ZN(_09273_));
 AND3_X1 _28227_ (.A1(_04834_),
    .A2(_09066_),
    .A3(_09273_),
    .ZN(_09274_));
 AND2_X1 _28228_ (.A1(_04834_),
    .A2(_09058_),
    .ZN(_09275_));
 AOI221_X1 _28229_ (.A(_09274_),
    .B1(_09275_),
    .B2(_09134_),
    .C1(_09062_),
    .C2(_04834_),
    .ZN(_09276_));
 NOR3_X1 _28230_ (.A1(_04834_),
    .A2(_08886_),
    .A3(_09273_),
    .ZN(_09277_));
 NOR2_X1 _28231_ (.A1(_04838_),
    .A2(_08896_),
    .ZN(_09278_));
 OAI21_X1 _28232_ (.A(_09136_),
    .B1(_09277_),
    .B2(_09278_),
    .ZN(_09279_));
 NAND2_X1 _28233_ (.A1(_09276_),
    .A2(_09279_),
    .ZN(_02809_));
 INV_X1 _28234_ (.A(_04849_),
    .ZN(_09280_));
 NAND4_X1 _28235_ (.A1(_04777_),
    .A2(_04789_),
    .A3(_04819_),
    .A4(_04834_),
    .ZN(_09281_));
 NOR2_X2 _28236_ (.A1(_09249_),
    .A2(_09281_),
    .ZN(_09282_));
 NOR3_X1 _28237_ (.A1(_09280_),
    .A2(_08856_),
    .A3(_09282_),
    .ZN(_09283_));
 AOI21_X1 _28238_ (.A(_09280_),
    .B1(_09044_),
    .B2(_09045_),
    .ZN(_09284_));
 AOI221_X1 _28239_ (.A(_09283_),
    .B1(_09284_),
    .B2(_09134_),
    .C1(_09062_),
    .C2(_04849_),
    .ZN(_09285_));
 NAND2_X1 _28240_ (.A1(_08895_),
    .A2(_09282_),
    .ZN(_09286_));
 OAI22_X1 _28241_ (.A1(_04853_),
    .A2(_08864_),
    .B1(_09286_),
    .B2(_04849_),
    .ZN(_09287_));
 NAND2_X1 _28242_ (.A1(_09054_),
    .A2(_09287_),
    .ZN(_09288_));
 NAND2_X1 _28243_ (.A1(_09285_),
    .A2(_09288_),
    .ZN(_02810_));
 AND2_X1 _28244_ (.A1(_05519_),
    .A2(_08844_),
    .ZN(_09289_));
 AND3_X1 _28245_ (.A1(_06560_),
    .A2(_06596_),
    .A3(\cs_registers_i.mhpmcounter[2][4] ),
    .ZN(_09290_));
 NAND2_X1 _28246_ (.A1(_09290_),
    .A2(_08892_),
    .ZN(_09291_));
 OAI21_X1 _28247_ (.A(_09289_),
    .B1(_09291_),
    .B2(_08920_),
    .ZN(_09292_));
 NAND3_X1 _28248_ (.A1(_08923_),
    .A2(_09290_),
    .A3(_08892_),
    .ZN(_09293_));
 OAI221_X1 _28249_ (.A(_09292_),
    .B1(_08922_),
    .B2(_08646_),
    .C1(_05519_),
    .C2(_09293_),
    .ZN(_02811_));
 AND4_X1 _28250_ (.A1(_04777_),
    .A2(_04789_),
    .A3(_04819_),
    .A4(_09256_),
    .ZN(_09294_));
 NAND3_X1 _28251_ (.A1(_04834_),
    .A2(_04849_),
    .A3(_09294_),
    .ZN(_09295_));
 AND3_X1 _28252_ (.A1(_04864_),
    .A2(_09066_),
    .A3(_09295_),
    .ZN(_09296_));
 AND2_X1 _28253_ (.A1(_04864_),
    .A2(_09058_),
    .ZN(_09297_));
 AOI221_X1 _28254_ (.A(_09296_),
    .B1(_09297_),
    .B2(_09072_),
    .C1(_09062_),
    .C2(_04864_),
    .ZN(_09298_));
 NOR3_X1 _28255_ (.A1(_04864_),
    .A2(_08886_),
    .A3(_09295_),
    .ZN(_09299_));
 NOR2_X1 _28256_ (.A1(_04868_),
    .A2(_08896_),
    .ZN(_09300_));
 OAI21_X1 _28257_ (.A(_09136_),
    .B1(_09299_),
    .B2(_09300_),
    .ZN(_09301_));
 NAND2_X1 _28258_ (.A1(_09298_),
    .A2(_09301_),
    .ZN(_02812_));
 NAND3_X1 _28259_ (.A1(_04849_),
    .A2(_04864_),
    .A3(_09282_),
    .ZN(_09302_));
 AND3_X1 _28260_ (.A1(_04882_),
    .A2(_08861_),
    .A3(_09302_),
    .ZN(_09303_));
 AND2_X1 _28261_ (.A1(_04882_),
    .A2(_09051_),
    .ZN(_09304_));
 AOI221_X1 _28262_ (.A(_09303_),
    .B1(_09304_),
    .B2(_08854_),
    .C1(_09073_),
    .C2(_04882_),
    .ZN(_09305_));
 NAND2_X1 _28263_ (.A1(_04849_),
    .A2(_04864_),
    .ZN(_09306_));
 NOR3_X1 _28264_ (.A1(_04882_),
    .A2(_09286_),
    .A3(_09306_),
    .ZN(_09307_));
 INV_X1 _28265_ (.A(_04885_),
    .ZN(_09308_));
 AOI21_X1 _28266_ (.A(_09307_),
    .B1(_09000_),
    .B2(_09308_),
    .ZN(_09309_));
 OAI21_X1 _28267_ (.A(_09305_),
    .B1(_09309_),
    .B2(_09078_),
    .ZN(_02813_));
 AND3_X1 _28268_ (.A1(_04849_),
    .A2(_04864_),
    .A3(_04882_),
    .ZN(_09310_));
 NAND3_X1 _28269_ (.A1(_04834_),
    .A2(_09294_),
    .A3(_09310_),
    .ZN(_09311_));
 AND3_X1 _28270_ (.A1(_04888_),
    .A2(_09066_),
    .A3(_09311_),
    .ZN(_09312_));
 AND2_X1 _28271_ (.A1(_04888_),
    .A2(_09058_),
    .ZN(_09313_));
 AOI221_X1 _28272_ (.A(_09312_),
    .B1(_09313_),
    .B2(_09072_),
    .C1(_09062_),
    .C2(_04888_),
    .ZN(_09314_));
 NOR3_X1 _28273_ (.A1(_04888_),
    .A2(_08886_),
    .A3(_09311_),
    .ZN(_09315_));
 NOR2_X1 _28274_ (.A1(_04905_),
    .A2(_08896_),
    .ZN(_09316_));
 OAI21_X1 _28275_ (.A(_09136_),
    .B1(_09315_),
    .B2(_09316_),
    .ZN(_09317_));
 NAND2_X1 _28276_ (.A1(_09314_),
    .A2(_09317_),
    .ZN(_02814_));
 NAND3_X1 _28277_ (.A1(_04888_),
    .A2(_09282_),
    .A3(_09310_),
    .ZN(_09318_));
 AND3_X1 _28278_ (.A1(_04909_),
    .A2(_09066_),
    .A3(_09318_),
    .ZN(_09319_));
 AND2_X1 _28279_ (.A1(_04909_),
    .A2(_09058_),
    .ZN(_09320_));
 AOI221_X1 _28280_ (.A(_09319_),
    .B1(_09320_),
    .B2(_09072_),
    .C1(_09062_),
    .C2(_04909_),
    .ZN(_09321_));
 NOR3_X1 _28281_ (.A1(_04909_),
    .A2(_08886_),
    .A3(_09318_),
    .ZN(_09322_));
 NOR2_X1 _28282_ (.A1(_04924_),
    .A2(_08896_),
    .ZN(_09323_));
 OAI21_X1 _28283_ (.A(_09136_),
    .B1(_09322_),
    .B2(_09323_),
    .ZN(_09324_));
 NAND2_X1 _28284_ (.A1(_09321_),
    .A2(_09324_),
    .ZN(_02815_));
 NAND4_X1 _28285_ (.A1(_08876_),
    .A2(_07226_),
    .A3(_08914_),
    .A4(_08877_),
    .ZN(_09325_));
 NAND3_X1 _28286_ (.A1(\cs_registers_i.mhpmcounter[2][6] ),
    .A2(_08907_),
    .A3(_09325_),
    .ZN(_09326_));
 INV_X1 _28287_ (.A(\cs_registers_i.mhpmcounter[2][6] ),
    .ZN(_09327_));
 NAND3_X1 _28288_ (.A1(_05519_),
    .A2(_09327_),
    .A3(_09290_),
    .ZN(_09328_));
 OAI221_X1 _28289_ (.A(_09326_),
    .B1(_09328_),
    .B2(_09027_),
    .C1(_08907_),
    .C2(_08655_),
    .ZN(_02816_));
 NOR2_X1 _28290_ (.A1(_05694_),
    .A2(_08893_),
    .ZN(_09329_));
 AOI22_X1 _28291_ (.A1(_08666_),
    .A2(_08935_),
    .B1(_09329_),
    .B2(_08912_),
    .ZN(_09330_));
 NAND2_X1 _28292_ (.A1(_05694_),
    .A2(_08884_),
    .ZN(_09331_));
 NOR2_X1 _28293_ (.A1(_08920_),
    .A2(_08893_),
    .ZN(_09332_));
 OAI21_X1 _28294_ (.A(_09330_),
    .B1(_09331_),
    .B2(_09332_),
    .ZN(_02817_));
 OAI221_X1 _28295_ (.A(_04932_),
    .B1(_08427_),
    .B2(_09018_),
    .C1(_08915_),
    .C2(_08880_),
    .ZN(_09333_));
 OR2_X1 _28296_ (.A1(_04932_),
    .A2(_08880_),
    .ZN(_09334_));
 OAI221_X1 _28297_ (.A(_09333_),
    .B1(_09334_),
    .B2(_08899_),
    .C1(_08922_),
    .C2(_04942_),
    .ZN(_02818_));
 NOR4_X1 _28298_ (.A1(_04948_),
    .A2(_08886_),
    .A3(_08888_),
    .A4(_08893_),
    .ZN(_09335_));
 OAI21_X1 _28299_ (.A(_08858_),
    .B1(_09137_),
    .B2(_09335_),
    .ZN(_09336_));
 NOR3_X1 _28300_ (.A1(_08899_),
    .A2(_08888_),
    .A3(_08893_),
    .ZN(_09337_));
 NAND2_X1 _28301_ (.A1(_04948_),
    .A2(_08884_),
    .ZN(_09338_));
 OAI21_X1 _28302_ (.A(_09336_),
    .B1(_09337_),
    .B2(_09338_),
    .ZN(_02819_));
 AOI21_X2 _28303_ (.A(_07835_),
    .B1(_07249_),
    .B2(_04021_),
    .ZN(_09339_));
 NOR2_X2 _28304_ (.A1(_04009_),
    .A2(_07285_),
    .ZN(_09340_));
 OAI21_X2 _28305_ (.A(_09340_),
    .B1(_03998_),
    .B2(_03997_),
    .ZN(_09341_));
 AND2_X1 _28306_ (.A1(_04044_),
    .A2(_09341_),
    .ZN(_09342_));
 BUF_X2 _28307_ (.A(_09342_),
    .Z(_09343_));
 NAND4_X4 _28308_ (.A1(_04009_),
    .A2(_03975_),
    .A3(_04018_),
    .A4(_04035_),
    .ZN(_09344_));
 NAND2_X1 _28309_ (.A1(_09343_),
    .A2(_09344_),
    .ZN(_09345_));
 NOR2_X4 _28310_ (.A1(_09339_),
    .A2(_09345_),
    .ZN(_09346_));
 MUX2_X1 _28311_ (.A(_03660_),
    .B(\cs_registers_i.mstack_d[0] ),
    .S(_07289_),
    .Z(_09347_));
 NOR2_X1 _28312_ (.A1(_07751_),
    .A2(_09347_),
    .ZN(_09348_));
 NOR2_X1 _28313_ (.A1(\cs_registers_i.dcsr_q[0] ),
    .A2(_07284_),
    .ZN(_09349_));
 OAI21_X1 _28314_ (.A(_09346_),
    .B1(_09348_),
    .B2(_09349_),
    .ZN(_02820_));
 MUX2_X1 _28315_ (.A(_03661_),
    .B(\cs_registers_i.mstack_d[1] ),
    .S(_07289_),
    .Z(_09350_));
 NOR2_X1 _28316_ (.A1(_07751_),
    .A2(_09350_),
    .ZN(_09351_));
 NOR2_X1 _28317_ (.A1(\cs_registers_i.dcsr_q[1] ),
    .A2(_07284_),
    .ZN(_09352_));
 OAI21_X1 _28318_ (.A(_09346_),
    .B1(_09351_),
    .B2(_09352_),
    .ZN(_02821_));
 INV_X1 _28319_ (.A(_04472_),
    .ZN(_09353_));
 OR3_X1 _28320_ (.A1(_04383_),
    .A2(_03546_),
    .A3(_04404_),
    .ZN(_09354_));
 NOR3_X4 _28321_ (.A1(_03576_),
    .A2(_09354_),
    .A3(_04542_),
    .ZN(_09355_));
 MUX2_X1 _28322_ (.A(\cs_registers_i.dcsr_q[11] ),
    .B(_09353_),
    .S(_09355_),
    .Z(_02823_));
 INV_X1 _28323_ (.A(_04528_),
    .ZN(_09356_));
 MUX2_X1 _28324_ (.A(\cs_registers_i.dcsr_q[12] ),
    .B(_09356_),
    .S(_09355_),
    .Z(_02824_));
 MUX2_X1 _28325_ (.A(\cs_registers_i.dcsr_q[13] ),
    .B(_04563_),
    .S(_09355_),
    .Z(_02825_));
 MUX2_X1 _28326_ (.A(\cs_registers_i.dcsr_q[15] ),
    .B(_08936_),
    .S(_09355_),
    .Z(_02826_));
 MUX2_X1 _28327_ (.A(_03997_),
    .B(_08402_),
    .S(_09355_),
    .Z(_02828_));
 AND2_X1 _28328_ (.A1(_09341_),
    .A2(_09344_),
    .ZN(_09357_));
 BUF_X2 _28329_ (.A(_09357_),
    .Z(_09358_));
 INV_X1 _28330_ (.A(\cs_registers_i.dcsr_q[6] ),
    .ZN(_09359_));
 AOI22_X1 _28331_ (.A1(_03997_),
    .A2(_09340_),
    .B1(_09358_),
    .B2(_09359_),
    .ZN(_02829_));
 AOI22_X1 _28332_ (.A1(_03998_),
    .A2(_09340_),
    .B1(_09344_),
    .B2(\cs_registers_i.dcsr_q[7] ),
    .ZN(_09360_));
 AOI21_X1 _28333_ (.A(_09360_),
    .B1(_09340_),
    .B2(_03997_),
    .ZN(_02830_));
 NAND2_X4 _28334_ (.A1(_09341_),
    .A2(_09344_),
    .ZN(_09361_));
 CLKBUF_X3 _28335_ (.A(_09361_),
    .Z(_09362_));
 INV_X1 _28336_ (.A(\cs_registers_i.dcsr_q[8] ),
    .ZN(_09363_));
 OAI22_X1 _28337_ (.A1(_01164_),
    .A2(_09341_),
    .B1(_09362_),
    .B2(_09363_),
    .ZN(_02831_));
 CLKBUF_X3 _28338_ (.A(_09361_),
    .Z(_09364_));
 BUF_X4 _28339_ (.A(_09343_),
    .Z(_09365_));
 MUX2_X1 _28340_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(\cs_registers_i.pc_id_i[10] ),
    .S(_09365_),
    .Z(_09366_));
 NAND2_X1 _28341_ (.A1(_04518_),
    .A2(net12),
    .ZN(_09367_));
 INV_X1 _28342_ (.A(_09367_),
    .ZN(_09368_));
 AOI22_X1 _28343_ (.A1(_09364_),
    .A2(_09366_),
    .B1(_09368_),
    .B2(_08867_),
    .ZN(_09369_));
 NAND2_X1 _28344_ (.A1(_09358_),
    .A2(_09367_),
    .ZN(_09370_));
 CLKBUF_X3 _28345_ (.A(_09370_),
    .Z(_09371_));
 INV_X1 _28346_ (.A(\cs_registers_i.csr_depc_o[10] ),
    .ZN(_09372_));
 OAI21_X1 _28347_ (.A(_09369_),
    .B1(_09371_),
    .B2(_09372_),
    .ZN(_02832_));
 MUX2_X1 _28348_ (.A(_08083_),
    .B(\cs_registers_i.pc_id_i[11] ),
    .S(_09365_),
    .Z(_09373_));
 NAND2_X1 _28349_ (.A1(_09362_),
    .A2(_09373_),
    .ZN(_09374_));
 CLKBUF_X3 _28350_ (.A(_09367_),
    .Z(_09375_));
 CLKBUF_X3 _28351_ (.A(_09375_),
    .Z(_09376_));
 INV_X1 _28352_ (.A(\cs_registers_i.csr_depc_o[11] ),
    .ZN(_09377_));
 OAI221_X1 _28353_ (.A(_09374_),
    .B1(_09376_),
    .B2(_04472_),
    .C1(_09377_),
    .C2(_09371_),
    .ZN(_02833_));
 MUX2_X1 _28354_ (.A(\cs_registers_i.pc_if_i[12] ),
    .B(\cs_registers_i.pc_id_i[12] ),
    .S(_09365_),
    .Z(_09378_));
 NAND2_X1 _28355_ (.A1(_09362_),
    .A2(_09378_),
    .ZN(_09379_));
 INV_X1 _28356_ (.A(\cs_registers_i.csr_depc_o[12] ),
    .ZN(_09380_));
 OAI221_X1 _28357_ (.A(_09379_),
    .B1(_09376_),
    .B2(_04528_),
    .C1(_09380_),
    .C2(_09371_),
    .ZN(_02834_));
 MUX2_X1 _28358_ (.A(\cs_registers_i.pc_if_i[13] ),
    .B(_12512_),
    .S(_09365_),
    .Z(_09381_));
 OAI22_X1 _28359_ (.A1(_04563_),
    .A2(_09375_),
    .B1(_09381_),
    .B2(_09358_),
    .ZN(_09382_));
 CLKBUF_X3 _28360_ (.A(_09370_),
    .Z(_09383_));
 NOR2_X1 _28361_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_09383_),
    .ZN(_09384_));
 NOR2_X1 _28362_ (.A1(_09382_),
    .A2(_09384_),
    .ZN(_02835_));
 MUX2_X1 _28363_ (.A(\cs_registers_i.pc_if_i[14] ),
    .B(_12618_),
    .S(_09365_),
    .Z(_09385_));
 NAND2_X1 _28364_ (.A1(_09362_),
    .A2(_09385_),
    .ZN(_09386_));
 INV_X1 _28365_ (.A(\cs_registers_i.csr_depc_o[14] ),
    .ZN(_09387_));
 OAI221_X1 _28366_ (.A(_09386_),
    .B1(_09376_),
    .B2(_04597_),
    .C1(_09387_),
    .C2(_09371_),
    .ZN(_02836_));
 MUX2_X1 _28367_ (.A(_08123_),
    .B(\cs_registers_i.pc_id_i[15] ),
    .S(_09365_),
    .Z(_09388_));
 NAND2_X1 _28368_ (.A1(_09362_),
    .A2(_09388_),
    .ZN(_09389_));
 OAI221_X1 _28369_ (.A(_09389_),
    .B1(_09376_),
    .B2(_04620_),
    .C1(_07824_),
    .C2(_09371_),
    .ZN(_02837_));
 MUX2_X2 _28370_ (.A(\cs_registers_i.pc_if_i[16] ),
    .B(\cs_registers_i.pc_id_i[16] ),
    .S(_09365_),
    .Z(_09390_));
 NAND2_X1 _28371_ (.A1(_09362_),
    .A2(_09390_),
    .ZN(_09391_));
 INV_X1 _28372_ (.A(\cs_registers_i.csr_depc_o[16] ),
    .ZN(_09392_));
 OAI221_X1 _28373_ (.A(_09391_),
    .B1(_09376_),
    .B2(_04645_),
    .C1(_09392_),
    .C2(_09371_),
    .ZN(_02838_));
 MUX2_X2 _28374_ (.A(_08138_),
    .B(_12868_),
    .S(_09365_),
    .Z(_09393_));
 OAI22_X1 _28375_ (.A1(_09200_),
    .A2(_09375_),
    .B1(_09393_),
    .B2(_09358_),
    .ZN(_09394_));
 NOR2_X1 _28376_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(_09383_),
    .ZN(_09395_));
 NOR2_X1 _28377_ (.A1(_09394_),
    .A2(_09395_),
    .ZN(_02839_));
 MUX2_X1 _28378_ (.A(\cs_registers_i.pc_if_i[18] ),
    .B(_12973_),
    .S(_09365_),
    .Z(_09396_));
 NAND2_X1 _28379_ (.A1(_09362_),
    .A2(_09396_),
    .ZN(_09397_));
 INV_X1 _28380_ (.A(\cs_registers_i.csr_depc_o[18] ),
    .ZN(_09398_));
 OAI221_X1 _28381_ (.A(_09397_),
    .B1(_09376_),
    .B2(_04685_),
    .C1(_09398_),
    .C2(_09371_),
    .ZN(_02840_));
 BUF_X4 _28382_ (.A(_09343_),
    .Z(_09399_));
 MUX2_X2 _28383_ (.A(_08151_),
    .B(\cs_registers_i.pc_id_i[19] ),
    .S(_09399_),
    .Z(_09400_));
 NAND2_X1 _28384_ (.A1(_09362_),
    .A2(_09400_),
    .ZN(_09401_));
 INV_X1 _28385_ (.A(\cs_registers_i.csr_depc_o[19] ),
    .ZN(_09402_));
 OAI221_X1 _28386_ (.A(_09401_),
    .B1(_09376_),
    .B2(_04700_),
    .C1(_09402_),
    .C2(_09371_),
    .ZN(_02841_));
 CLKBUF_X3 _28387_ (.A(_09343_),
    .Z(_09403_));
 MUX2_X1 _28388_ (.A(_04123_),
    .B(_11116_),
    .S(_09403_),
    .Z(_09404_));
 NAND2_X1 _28389_ (.A1(_09362_),
    .A2(_09404_),
    .ZN(_09405_));
 INV_X1 _28390_ (.A(\cs_registers_i.csr_depc_o[1] ),
    .ZN(_09406_));
 OAI221_X1 _28391_ (.A(_09405_),
    .B1(_09376_),
    .B2(_08519_),
    .C1(_09406_),
    .C2(_09371_),
    .ZN(_02842_));
 MUX2_X2 _28392_ (.A(\cs_registers_i.pc_if_i[20] ),
    .B(\cs_registers_i.pc_id_i[20] ),
    .S(_09399_),
    .Z(_09407_));
 NAND2_X1 _28393_ (.A1(_09362_),
    .A2(_09407_),
    .ZN(_09408_));
 INV_X1 _28394_ (.A(\cs_registers_i.csr_depc_o[20] ),
    .ZN(_09409_));
 CLKBUF_X3 _28395_ (.A(_09370_),
    .Z(_09410_));
 OAI221_X1 _28396_ (.A(_09408_),
    .B1(_09376_),
    .B2(_04721_),
    .C1(_09409_),
    .C2(_09410_),
    .ZN(_02843_));
 CLKBUF_X3 _28397_ (.A(_09361_),
    .Z(_09411_));
 MUX2_X2 _28398_ (.A(_08168_),
    .B(_13237_),
    .S(_09399_),
    .Z(_09412_));
 NAND2_X1 _28399_ (.A1(_09411_),
    .A2(_09412_),
    .ZN(_09413_));
 INV_X1 _28400_ (.A(\cs_registers_i.csr_depc_o[21] ),
    .ZN(_09414_));
 OAI221_X1 _28401_ (.A(_09413_),
    .B1(_09376_),
    .B2(_04742_),
    .C1(_09414_),
    .C2(_09410_),
    .ZN(_02844_));
 MUX2_X2 _28402_ (.A(\cs_registers_i.pc_if_i[22] ),
    .B(_13347_),
    .S(_09399_),
    .Z(_09415_));
 NAND2_X1 _28403_ (.A1(_09411_),
    .A2(_09415_),
    .ZN(_09416_));
 CLKBUF_X3 _28404_ (.A(_09375_),
    .Z(_09417_));
 INV_X1 _28405_ (.A(\cs_registers_i.csr_depc_o[22] ),
    .ZN(_09418_));
 OAI221_X1 _28406_ (.A(_09416_),
    .B1(_09417_),
    .B2(_04762_),
    .C1(_09418_),
    .C2(_09410_),
    .ZN(_02845_));
 MUX2_X2 _28407_ (.A(\cs_registers_i.pc_if_i[23] ),
    .B(_13423_),
    .S(_09399_),
    .Z(_09419_));
 NAND2_X1 _28408_ (.A1(_09411_),
    .A2(_09419_),
    .ZN(_09420_));
 INV_X1 _28409_ (.A(\cs_registers_i.csr_depc_o[23] ),
    .ZN(_09421_));
 OAI221_X1 _28410_ (.A(_09420_),
    .B1(_09417_),
    .B2(_04783_),
    .C1(_09421_),
    .C2(_09410_),
    .ZN(_02846_));
 MUX2_X2 _28411_ (.A(\cs_registers_i.pc_if_i[24] ),
    .B(\cs_registers_i.pc_id_i[24] ),
    .S(_09399_),
    .Z(_09422_));
 NAND2_X1 _28412_ (.A1(_09411_),
    .A2(_09422_),
    .ZN(_09423_));
 INV_X1 _28413_ (.A(\cs_registers_i.csr_depc_o[24] ),
    .ZN(_09424_));
 OAI221_X1 _28414_ (.A(_09423_),
    .B1(_09417_),
    .B2(_04805_),
    .C1(_09424_),
    .C2(_09410_),
    .ZN(_02847_));
 MUX2_X2 _28415_ (.A(\cs_registers_i.pc_if_i[25] ),
    .B(\cs_registers_i.pc_id_i[25] ),
    .S(_09399_),
    .Z(_09425_));
 NAND2_X1 _28416_ (.A1(_09411_),
    .A2(_09425_),
    .ZN(_09426_));
 INV_X1 _28417_ (.A(\cs_registers_i.csr_depc_o[25] ),
    .ZN(_09427_));
 OAI221_X1 _28418_ (.A(_09426_),
    .B1(_09417_),
    .B2(_04822_),
    .C1(_09427_),
    .C2(_09410_),
    .ZN(_02848_));
 MUX2_X2 _28419_ (.A(_08194_),
    .B(_13688_),
    .S(_09399_),
    .Z(_09428_));
 NAND2_X1 _28420_ (.A1(_09411_),
    .A2(_09428_),
    .ZN(_09429_));
 INV_X1 _28421_ (.A(\cs_registers_i.csr_depc_o[26] ),
    .ZN(_09430_));
 OAI221_X1 _28422_ (.A(_09429_),
    .B1(_09417_),
    .B2(_04838_),
    .C1(_09430_),
    .C2(_09410_),
    .ZN(_02849_));
 MUX2_X1 _28423_ (.A(\cs_registers_i.pc_if_i[27] ),
    .B(_03142_),
    .S(_09399_),
    .Z(_09431_));
 NAND2_X1 _28424_ (.A1(_09411_),
    .A2(_09431_),
    .ZN(_09432_));
 INV_X1 _28425_ (.A(\cs_registers_i.csr_depc_o[27] ),
    .ZN(_09433_));
 OAI221_X1 _28426_ (.A(_09432_),
    .B1(_09417_),
    .B2(_04853_),
    .C1(_09433_),
    .C2(_09410_),
    .ZN(_02850_));
 MUX2_X2 _28427_ (.A(\cs_registers_i.pc_if_i[28] ),
    .B(_03238_),
    .S(_09399_),
    .Z(_09434_));
 NAND2_X1 _28428_ (.A1(_09411_),
    .A2(_09434_),
    .ZN(_09435_));
 INV_X1 _28429_ (.A(\cs_registers_i.csr_depc_o[28] ),
    .ZN(_09436_));
 OAI221_X1 _28430_ (.A(_09435_),
    .B1(_09417_),
    .B2(_04868_),
    .C1(_09436_),
    .C2(_09410_),
    .ZN(_02851_));
 MUX2_X1 _28431_ (.A(_08209_),
    .B(\cs_registers_i.pc_id_i[29] ),
    .S(_09403_),
    .Z(_09437_));
 NAND2_X1 _28432_ (.A1(_09411_),
    .A2(_09437_),
    .ZN(_09438_));
 INV_X1 _28433_ (.A(\cs_registers_i.csr_depc_o[29] ),
    .ZN(_09439_));
 OAI221_X1 _28434_ (.A(_09438_),
    .B1(_09417_),
    .B2(_04885_),
    .C1(_09439_),
    .C2(_09410_),
    .ZN(_02852_));
 MUX2_X1 _28435_ (.A(_15754_),
    .B(_00012_),
    .S(_09343_),
    .Z(_09440_));
 OR2_X1 _28436_ (.A1(_09358_),
    .A2(_09440_),
    .ZN(_09441_));
 INV_X1 _28437_ (.A(\cs_registers_i.csr_depc_o[2] ),
    .ZN(_09442_));
 OAI221_X1 _28438_ (.A(_09441_),
    .B1(_09417_),
    .B2(_09029_),
    .C1(_09442_),
    .C2(_09383_),
    .ZN(_02853_));
 MUX2_X2 _28439_ (.A(\cs_registers_i.pc_if_i[30] ),
    .B(\cs_registers_i.pc_id_i[30] ),
    .S(_09403_),
    .Z(_09443_));
 NAND2_X1 _28440_ (.A1(_09411_),
    .A2(_09443_),
    .ZN(_09444_));
 INV_X1 _28441_ (.A(\cs_registers_i.csr_depc_o[30] ),
    .ZN(_09445_));
 OAI221_X1 _28442_ (.A(_09444_),
    .B1(_09417_),
    .B2(_04905_),
    .C1(_09445_),
    .C2(_09383_),
    .ZN(_02854_));
 MUX2_X1 _28443_ (.A(\cs_registers_i.pc_if_i[31] ),
    .B(\cs_registers_i.pc_id_i[31] ),
    .S(_09403_),
    .Z(_09446_));
 NAND2_X1 _28444_ (.A1(_09364_),
    .A2(_09446_),
    .ZN(_09447_));
 INV_X1 _28445_ (.A(\cs_registers_i.csr_depc_o[31] ),
    .ZN(_09448_));
 OAI221_X1 _28446_ (.A(_09447_),
    .B1(_09375_),
    .B2(_04924_),
    .C1(_09448_),
    .C2(_09383_),
    .ZN(_02855_));
 MUX2_X1 _28447_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(_11969_),
    .S(_09403_),
    .Z(_09449_));
 NAND2_X1 _28448_ (.A1(_09364_),
    .A2(_09449_),
    .ZN(_09450_));
 INV_X1 _28449_ (.A(\cs_registers_i.csr_depc_o[3] ),
    .ZN(_09451_));
 OAI221_X1 _28450_ (.A(_09450_),
    .B1(_09375_),
    .B2(_08629_),
    .C1(_09451_),
    .C2(_09383_),
    .ZN(_02856_));
 MUX2_X1 _28451_ (.A(\cs_registers_i.pc_if_i[4] ),
    .B(_12011_),
    .S(_09403_),
    .Z(_09452_));
 NAND2_X1 _28452_ (.A1(_09364_),
    .A2(_09452_),
    .ZN(_09453_));
 INV_X1 _28453_ (.A(\cs_registers_i.csr_depc_o[4] ),
    .ZN(_09454_));
 OAI221_X1 _28454_ (.A(_09453_),
    .B1(_09375_),
    .B2(_08639_),
    .C1(_09454_),
    .C2(_09383_),
    .ZN(_02857_));
 NAND2_X1 _28455_ (.A1(_08646_),
    .A2(_09368_),
    .ZN(_09455_));
 MUX2_X1 _28456_ (.A(\cs_registers_i.pc_if_i[5] ),
    .B(\cs_registers_i.pc_id_i[5] ),
    .S(_09365_),
    .Z(_09456_));
 OAI21_X1 _28457_ (.A(_09455_),
    .B1(_09456_),
    .B2(_09358_),
    .ZN(_09457_));
 NOR2_X1 _28458_ (.A1(\cs_registers_i.csr_depc_o[5] ),
    .A2(_09370_),
    .ZN(_09458_));
 NOR2_X1 _28459_ (.A1(_09457_),
    .A2(_09458_),
    .ZN(_02858_));
 MUX2_X1 _28460_ (.A(\cs_registers_i.pc_if_i[6] ),
    .B(\cs_registers_i.pc_id_i[6] ),
    .S(_09403_),
    .Z(_09459_));
 NAND2_X1 _28461_ (.A1(_09364_),
    .A2(_09459_),
    .ZN(_09460_));
 INV_X1 _28462_ (.A(\cs_registers_i.csr_depc_o[6] ),
    .ZN(_09461_));
 OAI221_X1 _28463_ (.A(_09460_),
    .B1(_09375_),
    .B2(_08655_),
    .C1(_09461_),
    .C2(_09383_),
    .ZN(_02859_));
 MUX2_X1 _28464_ (.A(_08093_),
    .B(\cs_registers_i.pc_id_i[7] ),
    .S(_09403_),
    .Z(_09462_));
 AOI22_X1 _28465_ (.A1(_08666_),
    .A2(_09368_),
    .B1(_09462_),
    .B2(_09364_),
    .ZN(_09463_));
 INV_X1 _28466_ (.A(\cs_registers_i.csr_depc_o[7] ),
    .ZN(_09464_));
 OAI21_X1 _28467_ (.A(_09463_),
    .B1(_09371_),
    .B2(_09464_),
    .ZN(_02860_));
 MUX2_X1 _28468_ (.A(\cs_registers_i.pc_if_i[8] ),
    .B(_12218_),
    .S(_09403_),
    .Z(_09465_));
 NAND2_X1 _28469_ (.A1(_09364_),
    .A2(_09465_),
    .ZN(_09466_));
 INV_X1 _28470_ (.A(\cs_registers_i.csr_depc_o[8] ),
    .ZN(_09467_));
 OAI221_X1 _28471_ (.A(_09466_),
    .B1(_09375_),
    .B2(_04942_),
    .C1(_09467_),
    .C2(_09383_),
    .ZN(_02861_));
 MUX2_X1 _28472_ (.A(_08086_),
    .B(_12261_),
    .S(_09403_),
    .Z(_09468_));
 NAND2_X1 _28473_ (.A1(_09364_),
    .A2(_09468_),
    .ZN(_09469_));
 INV_X1 _28474_ (.A(\cs_registers_i.csr_depc_o[9] ),
    .ZN(_09470_));
 OAI221_X1 _28475_ (.A(_09469_),
    .B1(_09375_),
    .B2(_04960_),
    .C1(_09470_),
    .C2(_09383_),
    .ZN(_02862_));
 NAND2_X1 _28476_ (.A1(_04583_),
    .A2(_09044_),
    .ZN(_09471_));
 CLKBUF_X3 _28477_ (.A(_09471_),
    .Z(_09472_));
 MUX2_X1 _28478_ (.A(_08396_),
    .B(\cs_registers_i.dscratch0_q[0] ),
    .S(_09472_),
    .Z(_02863_));
 MUX2_X1 _28479_ (.A(_08867_),
    .B(\cs_registers_i.dscratch0_q[10] ),
    .S(_09472_),
    .Z(_02864_));
 CLKBUF_X3 _28480_ (.A(_09471_),
    .Z(_09473_));
 NAND2_X1 _28481_ (.A1(\cs_registers_i.dscratch0_q[11] ),
    .A2(_09473_),
    .ZN(_09474_));
 CLKBUF_X3 _28482_ (.A(_09472_),
    .Z(_09475_));
 OAI21_X1 _28483_ (.A(_09474_),
    .B1(_09475_),
    .B2(_04472_),
    .ZN(_02865_));
 NAND2_X1 _28484_ (.A1(\cs_registers_i.dscratch0_q[12] ),
    .A2(_09473_),
    .ZN(_09476_));
 OAI21_X1 _28485_ (.A(_09476_),
    .B1(_09475_),
    .B2(_04528_),
    .ZN(_02866_));
 NAND2_X1 _28486_ (.A1(\cs_registers_i.dscratch0_q[13] ),
    .A2(_09473_),
    .ZN(_09477_));
 OAI21_X1 _28487_ (.A(_09477_),
    .B1(_09475_),
    .B2(_04562_),
    .ZN(_02867_));
 CLKBUF_X3 _28488_ (.A(_09471_),
    .Z(_09478_));
 NAND2_X1 _28489_ (.A1(\cs_registers_i.dscratch0_q[14] ),
    .A2(_09478_),
    .ZN(_09479_));
 OAI21_X1 _28490_ (.A(_09479_),
    .B1(_09475_),
    .B2(_04597_),
    .ZN(_02868_));
 NAND2_X1 _28491_ (.A1(\cs_registers_i.dscratch0_q[15] ),
    .A2(_09478_),
    .ZN(_09480_));
 OAI21_X1 _28492_ (.A(_09480_),
    .B1(_09475_),
    .B2(_04620_),
    .ZN(_02869_));
 MUX2_X1 _28493_ (.A(_08493_),
    .B(\cs_registers_i.dscratch0_q[16] ),
    .S(_09472_),
    .Z(_02870_));
 NAND2_X1 _28494_ (.A1(\cs_registers_i.dscratch0_q[17] ),
    .A2(_09478_),
    .ZN(_09481_));
 OAI21_X1 _28495_ (.A(_09481_),
    .B1(_09475_),
    .B2(_04665_),
    .ZN(_02871_));
 NAND2_X1 _28496_ (.A1(\cs_registers_i.dscratch0_q[18] ),
    .A2(_09478_),
    .ZN(_09482_));
 OAI21_X1 _28497_ (.A(_09482_),
    .B1(_09475_),
    .B2(_04685_),
    .ZN(_02872_));
 NAND2_X1 _28498_ (.A1(\cs_registers_i.dscratch0_q[19] ),
    .A2(_09478_),
    .ZN(_09483_));
 OAI21_X1 _28499_ (.A(_09483_),
    .B1(_09475_),
    .B2(_04700_),
    .ZN(_02873_));
 NAND2_X1 _28500_ (.A1(\cs_registers_i.dscratch0_q[1] ),
    .A2(_09478_),
    .ZN(_09484_));
 OAI21_X1 _28501_ (.A(_09484_),
    .B1(_09475_),
    .B2(_08519_),
    .ZN(_02874_));
 NAND2_X1 _28502_ (.A1(\cs_registers_i.dscratch0_q[20] ),
    .A2(_09478_),
    .ZN(_09485_));
 OAI21_X1 _28503_ (.A(_09485_),
    .B1(_09475_),
    .B2(_04721_),
    .ZN(_02875_));
 NAND2_X1 _28504_ (.A1(\cs_registers_i.dscratch0_q[21] ),
    .A2(_09478_),
    .ZN(_09486_));
 CLKBUF_X3 _28505_ (.A(_09471_),
    .Z(_09487_));
 OAI21_X1 _28506_ (.A(_09486_),
    .B1(_09487_),
    .B2(_04742_),
    .ZN(_02876_));
 NAND2_X1 _28507_ (.A1(\cs_registers_i.dscratch0_q[22] ),
    .A2(_09478_),
    .ZN(_09488_));
 OAI21_X1 _28508_ (.A(_09488_),
    .B1(_09487_),
    .B2(_04762_),
    .ZN(_02877_));
 NAND2_X1 _28509_ (.A1(\cs_registers_i.dscratch0_q[23] ),
    .A2(_09478_),
    .ZN(_09489_));
 OAI21_X1 _28510_ (.A(_09489_),
    .B1(_09487_),
    .B2(_04783_),
    .ZN(_02878_));
 CLKBUF_X3 _28511_ (.A(_09471_),
    .Z(_09490_));
 NAND2_X1 _28512_ (.A1(\cs_registers_i.dscratch0_q[24] ),
    .A2(_09490_),
    .ZN(_09491_));
 OAI21_X1 _28513_ (.A(_09491_),
    .B1(_09487_),
    .B2(_04805_),
    .ZN(_02879_));
 NAND2_X1 _28514_ (.A1(\cs_registers_i.dscratch0_q[25] ),
    .A2(_09490_),
    .ZN(_09492_));
 OAI21_X1 _28515_ (.A(_09492_),
    .B1(_09487_),
    .B2(_04822_),
    .ZN(_02880_));
 NAND2_X1 _28516_ (.A1(\cs_registers_i.dscratch0_q[26] ),
    .A2(_09490_),
    .ZN(_09493_));
 OAI21_X1 _28517_ (.A(_09493_),
    .B1(_09487_),
    .B2(_04838_),
    .ZN(_02881_));
 NAND2_X1 _28518_ (.A1(\cs_registers_i.dscratch0_q[27] ),
    .A2(_09490_),
    .ZN(_09494_));
 OAI21_X1 _28519_ (.A(_09494_),
    .B1(_09487_),
    .B2(_04853_),
    .ZN(_02882_));
 NAND2_X1 _28520_ (.A1(\cs_registers_i.dscratch0_q[28] ),
    .A2(_09490_),
    .ZN(_09495_));
 OAI21_X1 _28521_ (.A(_09495_),
    .B1(_09487_),
    .B2(_04868_),
    .ZN(_02883_));
 NAND2_X1 _28522_ (.A1(\cs_registers_i.dscratch0_q[29] ),
    .A2(_09490_),
    .ZN(_09496_));
 OAI21_X1 _28523_ (.A(_09496_),
    .B1(_09487_),
    .B2(_04885_),
    .ZN(_02884_));
 MUX2_X1 _28524_ (.A(_08402_),
    .B(\cs_registers_i.dscratch0_q[2] ),
    .S(_09472_),
    .Z(_02885_));
 NAND2_X1 _28525_ (.A1(\cs_registers_i.dscratch0_q[30] ),
    .A2(_09490_),
    .ZN(_09497_));
 OAI21_X1 _28526_ (.A(_09497_),
    .B1(_09487_),
    .B2(_04905_),
    .ZN(_02886_));
 NAND2_X1 _28527_ (.A1(\cs_registers_i.dscratch0_q[31] ),
    .A2(_09490_),
    .ZN(_09498_));
 OAI21_X1 _28528_ (.A(_09498_),
    .B1(_09473_),
    .B2(_04924_),
    .ZN(_02887_));
 NAND2_X1 _28529_ (.A1(\cs_registers_i.dscratch0_q[3] ),
    .A2(_09490_),
    .ZN(_09499_));
 OAI21_X1 _28530_ (.A(_09499_),
    .B1(_09473_),
    .B2(_08629_),
    .ZN(_02888_));
 NAND2_X1 _28531_ (.A1(\cs_registers_i.dscratch0_q[4] ),
    .A2(_09490_),
    .ZN(_09500_));
 OAI21_X1 _28532_ (.A(_09500_),
    .B1(_09473_),
    .B2(_08639_),
    .ZN(_02889_));
 NAND2_X1 _28533_ (.A1(\cs_registers_i.dscratch0_q[5] ),
    .A2(_09472_),
    .ZN(_09501_));
 OAI21_X1 _28534_ (.A(_09501_),
    .B1(_09473_),
    .B2(_08646_),
    .ZN(_02890_));
 NAND2_X1 _28535_ (.A1(\cs_registers_i.dscratch0_q[6] ),
    .A2(_09472_),
    .ZN(_09502_));
 OAI21_X1 _28536_ (.A(_09502_),
    .B1(_09473_),
    .B2(_08655_),
    .ZN(_02891_));
 MUX2_X1 _28537_ (.A(_08666_),
    .B(\cs_registers_i.dscratch0_q[7] ),
    .S(_09472_),
    .Z(_02892_));
 NAND2_X1 _28538_ (.A1(\cs_registers_i.dscratch0_q[8] ),
    .A2(_09472_),
    .ZN(_09503_));
 OAI21_X1 _28539_ (.A(_09503_),
    .B1(_09473_),
    .B2(_04942_),
    .ZN(_02893_));
 NAND2_X1 _28540_ (.A1(\cs_registers_i.dscratch0_q[9] ),
    .A2(_09472_),
    .ZN(_09504_));
 OAI21_X1 _28541_ (.A(_09504_),
    .B1(_09473_),
    .B2(_04960_),
    .ZN(_02894_));
 NAND2_X2 _28542_ (.A1(_04584_),
    .A2(_09044_),
    .ZN(_09505_));
 BUF_X4 _28543_ (.A(_09505_),
    .Z(_09506_));
 MUX2_X1 _28544_ (.A(_08396_),
    .B(\cs_registers_i.dscratch1_q[0] ),
    .S(_09506_),
    .Z(_02895_));
 MUX2_X1 _28545_ (.A(_08867_),
    .B(\cs_registers_i.dscratch1_q[10] ),
    .S(_09506_),
    .Z(_02896_));
 CLKBUF_X3 _28546_ (.A(_09505_),
    .Z(_09507_));
 NAND2_X1 _28547_ (.A1(\cs_registers_i.dscratch1_q[11] ),
    .A2(_09507_),
    .ZN(_09508_));
 BUF_X4 _28548_ (.A(_09506_),
    .Z(_09509_));
 OAI21_X1 _28549_ (.A(_09508_),
    .B1(_09509_),
    .B2(_04472_),
    .ZN(_02897_));
 NAND2_X1 _28550_ (.A1(\cs_registers_i.dscratch1_q[12] ),
    .A2(_09507_),
    .ZN(_09510_));
 OAI21_X1 _28551_ (.A(_09510_),
    .B1(_09509_),
    .B2(_04528_),
    .ZN(_02898_));
 NAND2_X1 _28552_ (.A1(\cs_registers_i.dscratch1_q[13] ),
    .A2(_09507_),
    .ZN(_09511_));
 OAI21_X1 _28553_ (.A(_09511_),
    .B1(_09509_),
    .B2(_04562_),
    .ZN(_02899_));
 BUF_X4 _28554_ (.A(_09505_),
    .Z(_09512_));
 NAND2_X1 _28555_ (.A1(\cs_registers_i.dscratch1_q[14] ),
    .A2(_09512_),
    .ZN(_09513_));
 OAI21_X1 _28556_ (.A(_09513_),
    .B1(_09509_),
    .B2(_04597_),
    .ZN(_02900_));
 NAND2_X1 _28557_ (.A1(\cs_registers_i.dscratch1_q[15] ),
    .A2(_09512_),
    .ZN(_09514_));
 OAI21_X1 _28558_ (.A(_09514_),
    .B1(_09509_),
    .B2(_04620_),
    .ZN(_02901_));
 MUX2_X1 _28559_ (.A(_08493_),
    .B(\cs_registers_i.dscratch1_q[16] ),
    .S(_09506_),
    .Z(_02902_));
 NAND2_X1 _28560_ (.A1(\cs_registers_i.dscratch1_q[17] ),
    .A2(_09512_),
    .ZN(_09515_));
 OAI21_X1 _28561_ (.A(_09515_),
    .B1(_09509_),
    .B2(_04665_),
    .ZN(_02903_));
 NAND2_X1 _28562_ (.A1(\cs_registers_i.dscratch1_q[18] ),
    .A2(_09512_),
    .ZN(_09516_));
 OAI21_X1 _28563_ (.A(_09516_),
    .B1(_09509_),
    .B2(_04685_),
    .ZN(_02904_));
 NAND2_X1 _28564_ (.A1(\cs_registers_i.dscratch1_q[19] ),
    .A2(_09512_),
    .ZN(_09517_));
 OAI21_X1 _28565_ (.A(_09517_),
    .B1(_09509_),
    .B2(_04700_),
    .ZN(_02905_));
 NAND2_X1 _28566_ (.A1(\cs_registers_i.dscratch1_q[1] ),
    .A2(_09512_),
    .ZN(_09518_));
 OAI21_X1 _28567_ (.A(_09518_),
    .B1(_09509_),
    .B2(_08519_),
    .ZN(_02906_));
 NAND2_X1 _28568_ (.A1(\cs_registers_i.dscratch1_q[20] ),
    .A2(_09512_),
    .ZN(_09519_));
 OAI21_X1 _28569_ (.A(_09519_),
    .B1(_09509_),
    .B2(_04721_),
    .ZN(_02907_));
 NAND2_X1 _28570_ (.A1(\cs_registers_i.dscratch1_q[21] ),
    .A2(_09512_),
    .ZN(_09520_));
 CLKBUF_X3 _28571_ (.A(_09505_),
    .Z(_09521_));
 OAI21_X1 _28572_ (.A(_09520_),
    .B1(_09521_),
    .B2(_04742_),
    .ZN(_02908_));
 NAND2_X1 _28573_ (.A1(\cs_registers_i.dscratch1_q[22] ),
    .A2(_09512_),
    .ZN(_09522_));
 OAI21_X1 _28574_ (.A(_09522_),
    .B1(_09521_),
    .B2(_04762_),
    .ZN(_02909_));
 NAND2_X1 _28575_ (.A1(\cs_registers_i.dscratch1_q[23] ),
    .A2(_09512_),
    .ZN(_09523_));
 OAI21_X1 _28576_ (.A(_09523_),
    .B1(_09521_),
    .B2(_04783_),
    .ZN(_02910_));
 CLKBUF_X3 _28577_ (.A(_09505_),
    .Z(_09524_));
 NAND2_X1 _28578_ (.A1(\cs_registers_i.dscratch1_q[24] ),
    .A2(_09524_),
    .ZN(_09525_));
 OAI21_X1 _28579_ (.A(_09525_),
    .B1(_09521_),
    .B2(_04805_),
    .ZN(_02911_));
 NAND2_X1 _28580_ (.A1(\cs_registers_i.dscratch1_q[25] ),
    .A2(_09524_),
    .ZN(_09526_));
 OAI21_X1 _28581_ (.A(_09526_),
    .B1(_09521_),
    .B2(_04822_),
    .ZN(_02912_));
 NAND2_X1 _28582_ (.A1(\cs_registers_i.dscratch1_q[26] ),
    .A2(_09524_),
    .ZN(_09527_));
 OAI21_X1 _28583_ (.A(_09527_),
    .B1(_09521_),
    .B2(_04838_),
    .ZN(_02913_));
 NAND2_X1 _28584_ (.A1(\cs_registers_i.dscratch1_q[27] ),
    .A2(_09524_),
    .ZN(_09528_));
 OAI21_X1 _28585_ (.A(_09528_),
    .B1(_09521_),
    .B2(_04853_),
    .ZN(_02914_));
 NAND2_X1 _28586_ (.A1(\cs_registers_i.dscratch1_q[28] ),
    .A2(_09524_),
    .ZN(_09529_));
 OAI21_X1 _28587_ (.A(_09529_),
    .B1(_09521_),
    .B2(_04868_),
    .ZN(_02915_));
 NAND2_X1 _28588_ (.A1(\cs_registers_i.dscratch1_q[29] ),
    .A2(_09524_),
    .ZN(_09530_));
 OAI21_X1 _28589_ (.A(_09530_),
    .B1(_09521_),
    .B2(_04885_),
    .ZN(_02916_));
 MUX2_X1 _28590_ (.A(_08402_),
    .B(\cs_registers_i.dscratch1_q[2] ),
    .S(_09506_),
    .Z(_02917_));
 NAND2_X1 _28591_ (.A1(\cs_registers_i.dscratch1_q[30] ),
    .A2(_09524_),
    .ZN(_09531_));
 OAI21_X1 _28592_ (.A(_09531_),
    .B1(_09521_),
    .B2(_04905_),
    .ZN(_02918_));
 NAND2_X1 _28593_ (.A1(\cs_registers_i.dscratch1_q[31] ),
    .A2(_09524_),
    .ZN(_09532_));
 OAI21_X1 _28594_ (.A(_09532_),
    .B1(_09507_),
    .B2(_04924_),
    .ZN(_02919_));
 NAND2_X1 _28595_ (.A1(\cs_registers_i.dscratch1_q[3] ),
    .A2(_09524_),
    .ZN(_09533_));
 OAI21_X1 _28596_ (.A(_09533_),
    .B1(_09507_),
    .B2(_08629_),
    .ZN(_02920_));
 NAND2_X1 _28597_ (.A1(\cs_registers_i.dscratch1_q[4] ),
    .A2(_09524_),
    .ZN(_09534_));
 OAI21_X1 _28598_ (.A(_09534_),
    .B1(_09507_),
    .B2(_08639_),
    .ZN(_02921_));
 NAND2_X1 _28599_ (.A1(\cs_registers_i.dscratch1_q[5] ),
    .A2(_09506_),
    .ZN(_09535_));
 OAI21_X1 _28600_ (.A(_09535_),
    .B1(_09507_),
    .B2(_08646_),
    .ZN(_02922_));
 NAND2_X1 _28601_ (.A1(\cs_registers_i.dscratch1_q[6] ),
    .A2(_09506_),
    .ZN(_09536_));
 OAI21_X1 _28602_ (.A(_09536_),
    .B1(_09507_),
    .B2(_08655_),
    .ZN(_02923_));
 MUX2_X1 _28603_ (.A(_08666_),
    .B(\cs_registers_i.dscratch1_q[7] ),
    .S(_09506_),
    .Z(_02924_));
 NAND2_X1 _28604_ (.A1(\cs_registers_i.dscratch1_q[8] ),
    .A2(_09506_),
    .ZN(_09537_));
 OAI21_X1 _28605_ (.A(_09537_),
    .B1(_09507_),
    .B2(_04942_),
    .ZN(_02925_));
 NAND2_X1 _28606_ (.A1(\cs_registers_i.dscratch1_q[9] ),
    .A2(_09506_),
    .ZN(_09538_));
 OAI21_X1 _28607_ (.A(_09538_),
    .B1(_09507_),
    .B2(_04960_),
    .ZN(_02926_));
 NOR3_X2 _28608_ (.A1(_03564_),
    .A2(_09346_),
    .A3(_09361_),
    .ZN(_09539_));
 BUF_X4 _28609_ (.A(_09539_),
    .Z(_09540_));
 BUF_X4 _28610_ (.A(_09540_),
    .Z(_09541_));
 BUF_X4 _28611_ (.A(_04016_),
    .Z(_09542_));
 CLKBUF_X3 _28612_ (.A(_09542_),
    .Z(_09543_));
 NOR2_X1 _28613_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.load_err_q ),
    .ZN(_09544_));
 NOR3_X2 _28614_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_03681_),
    .A3(_09544_),
    .ZN(_09545_));
 NAND2_X1 _28615_ (.A1(_12368_),
    .A2(_04016_),
    .ZN(_09546_));
 NOR3_X1 _28616_ (.A1(_03647_),
    .A2(_03662_),
    .A3(_09546_),
    .ZN(_09547_));
 NAND2_X1 _28617_ (.A1(_04023_),
    .A2(_09547_),
    .ZN(_09548_));
 OAI21_X1 _28618_ (.A(_09548_),
    .B1(_04025_),
    .B2(_04019_),
    .ZN(_09549_));
 OAI21_X1 _28619_ (.A(_09543_),
    .B1(_09545_),
    .B2(_09549_),
    .ZN(_09550_));
 BUF_X4 _28620_ (.A(_04020_),
    .Z(_09551_));
 AOI21_X2 _28621_ (.A(_07835_),
    .B1(_09550_),
    .B2(_09551_),
    .ZN(_09552_));
 OAI21_X1 _28622_ (.A(_09541_),
    .B1(_09552_),
    .B2(_04063_),
    .ZN(_09553_));
 NAND2_X1 _28623_ (.A1(\cs_registers_i.nmi_mode_i ),
    .A2(_04070_),
    .ZN(_09554_));
 CLKBUF_X3 _28624_ (.A(_09554_),
    .Z(_09555_));
 OR3_X1 _28625_ (.A1(_03564_),
    .A2(_09346_),
    .A3(_09361_),
    .ZN(_09556_));
 BUF_X4 _28626_ (.A(_09556_),
    .Z(_09557_));
 NAND2_X4 _28627_ (.A1(_09555_),
    .A2(_09557_),
    .ZN(_09558_));
 INV_X1 _28628_ (.A(\cs_registers_i.mstack_cause_q[0] ),
    .ZN(_09559_));
 OAI221_X1 _28629_ (.A(_09553_),
    .B1(_09558_),
    .B2(_08860_),
    .C1(_09555_),
    .C2(_09559_),
    .ZN(_09560_));
 NOR3_X4 _28630_ (.A1(_04086_),
    .A2(_09346_),
    .A3(_09361_),
    .ZN(_09561_));
 INV_X1 _28631_ (.A(_04070_),
    .ZN(_09562_));
 NOR2_X4 _28632_ (.A1(_03977_),
    .A2(_09562_),
    .ZN(_09563_));
 OR2_X1 _28633_ (.A1(_09561_),
    .A2(_09563_),
    .ZN(_09564_));
 AOI21_X4 _28634_ (.A(_09564_),
    .B1(_04918_),
    .B2(net12),
    .ZN(_09565_));
 MUX2_X1 _28635_ (.A(_09560_),
    .B(\cs_registers_i.mcause_q[0] ),
    .S(_09565_),
    .Z(_02927_));
 NOR2_X1 _28636_ (.A1(_04011_),
    .A2(_07835_),
    .ZN(_09566_));
 NAND2_X1 _28637_ (.A1(_10794_),
    .A2(_03679_),
    .ZN(_09567_));
 NAND3_X1 _28638_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(_04024_),
    .A3(_09567_),
    .ZN(_09568_));
 NAND2_X1 _28639_ (.A1(_09543_),
    .A2(_09568_),
    .ZN(_09569_));
 OAI21_X1 _28640_ (.A(_09566_),
    .B1(_09569_),
    .B2(_09549_),
    .ZN(_09570_));
 NAND3_X1 _28641_ (.A1(_04096_),
    .A2(_09540_),
    .A3(_09570_),
    .ZN(_09571_));
 OAI21_X1 _28642_ (.A(_09571_),
    .B1(_09555_),
    .B2(\cs_registers_i.mstack_cause_q[1] ),
    .ZN(_09572_));
 NOR2_X4 _28643_ (.A1(_09563_),
    .A2(_09540_),
    .ZN(_09573_));
 AOI21_X1 _28644_ (.A(_09572_),
    .B1(_09573_),
    .B2(_08519_),
    .ZN(_09574_));
 MUX2_X1 _28645_ (.A(_09574_),
    .B(\cs_registers_i.mcause_q[1] ),
    .S(_09565_),
    .Z(_02928_));
 NAND2_X1 _28646_ (.A1(\cs_registers_i.mcause_q[2] ),
    .A2(_09565_),
    .ZN(_09575_));
 INV_X1 _28647_ (.A(_04016_),
    .ZN(_09576_));
 NAND2_X1 _28648_ (.A1(_09576_),
    .A2(_04020_),
    .ZN(_09577_));
 AND2_X1 _28649_ (.A1(_09545_),
    .A2(_09577_),
    .ZN(_09578_));
 CLKBUF_X3 _28650_ (.A(_09578_),
    .Z(_09579_));
 CLKBUF_X3 _28651_ (.A(_09579_),
    .Z(_09580_));
 AOI21_X2 _28652_ (.A(_09557_),
    .B1(_09566_),
    .B2(_09580_),
    .ZN(_09581_));
 NAND2_X1 _28653_ (.A1(_07739_),
    .A2(_09581_),
    .ZN(_09582_));
 CLKBUF_X3 _28654_ (.A(_09558_),
    .Z(_09583_));
 OAI221_X1 _28655_ (.A(_09582_),
    .B1(_09583_),
    .B2(_08402_),
    .C1(\cs_registers_i.mstack_cause_q[2] ),
    .C2(_09555_),
    .ZN(_09584_));
 OAI21_X1 _28656_ (.A(_09575_),
    .B1(_09584_),
    .B2(_09565_),
    .ZN(_02929_));
 NAND2_X1 _28657_ (.A1(\cs_registers_i.mcause_q[3] ),
    .A2(_09565_),
    .ZN(_09585_));
 BUF_X4 _28658_ (.A(_09540_),
    .Z(_09586_));
 CLKBUF_X3 _28659_ (.A(_04011_),
    .Z(_09587_));
 OR4_X1 _28660_ (.A1(_09587_),
    .A2(_07835_),
    .A3(_09546_),
    .A4(_09567_),
    .ZN(_09588_));
 NAND3_X1 _28661_ (.A1(_07728_),
    .A2(_09586_),
    .A3(_09588_),
    .ZN(_09589_));
 OAI221_X1 _28662_ (.A(_09589_),
    .B1(_09583_),
    .B2(_08630_),
    .C1(\cs_registers_i.mstack_cause_q[3] ),
    .C2(_09555_),
    .ZN(_09590_));
 OAI21_X1 _28663_ (.A(_09585_),
    .B1(_09590_),
    .B2(_09565_),
    .ZN(_02930_));
 NOR2_X1 _28664_ (.A1(\cs_registers_i.mstack_cause_q[4] ),
    .A2(_09554_),
    .ZN(_09591_));
 AOI221_X1 _28665_ (.A(_09591_),
    .B1(_09573_),
    .B2(_08639_),
    .C1(_07746_),
    .C2(_09540_),
    .ZN(_09592_));
 MUX2_X1 _28666_ (.A(_09592_),
    .B(\cs_registers_i.mcause_q[4] ),
    .S(_09565_),
    .Z(_02931_));
 INV_X1 _28667_ (.A(\cs_registers_i.mcause_q[5] ),
    .ZN(_09593_));
 BUF_X4 _28668_ (.A(_09563_),
    .Z(_09594_));
 NOR3_X1 _28669_ (.A1(_04923_),
    .A2(_09594_),
    .A3(_09586_),
    .ZN(_09595_));
 AOI21_X1 _28670_ (.A(_09595_),
    .B1(_09594_),
    .B2(\cs_registers_i.mstack_cause_q[5] ),
    .ZN(_09596_));
 NOR2_X1 _28671_ (.A1(_03995_),
    .A2(_09565_),
    .ZN(_09597_));
 AOI22_X1 _28672_ (.A1(_09593_),
    .A2(_09565_),
    .B1(_09596_),
    .B2(_09597_),
    .ZN(_02932_));
 NAND2_X1 _28673_ (.A1(\cs_registers_i.mstack_epc_q[0] ),
    .A2(_09594_),
    .ZN(_09598_));
 AND2_X1 _28674_ (.A1(_04571_),
    .A2(_08835_),
    .ZN(_09599_));
 OR2_X1 _28675_ (.A1(_09564_),
    .A2(_09599_),
    .ZN(_09600_));
 CLKBUF_X3 _28676_ (.A(_09600_),
    .Z(_09601_));
 BUF_X4 _28677_ (.A(_09601_),
    .Z(_09602_));
 INV_X1 _28678_ (.A(\cs_registers_i.csr_mepc_o[0] ),
    .ZN(_09603_));
 OAI21_X1 _28679_ (.A(_09598_),
    .B1(_09602_),
    .B2(_09603_),
    .ZN(_02933_));
 AOI22_X1 _28680_ (.A1(\cs_registers_i.mstack_epc_q[10] ),
    .A2(_09594_),
    .B1(_09541_),
    .B2(_09366_),
    .ZN(_09604_));
 OAI21_X1 _28681_ (.A(_09604_),
    .B1(_09583_),
    .B2(_08437_),
    .ZN(_09605_));
 MUX2_X1 _28682_ (.A(\cs_registers_i.csr_mepc_o[10] ),
    .B(_09605_),
    .S(_09602_),
    .Z(_02934_));
 AOI22_X1 _28683_ (.A1(\cs_registers_i.mstack_epc_q[11] ),
    .A2(_09594_),
    .B1(_09541_),
    .B2(_09373_),
    .ZN(_09606_));
 OAI21_X1 _28684_ (.A(_09606_),
    .B1(_09583_),
    .B2(_04472_),
    .ZN(_09607_));
 MUX2_X1 _28685_ (.A(\cs_registers_i.csr_mepc_o[11] ),
    .B(_09607_),
    .S(_09602_),
    .Z(_02935_));
 AOI22_X1 _28686_ (.A1(\cs_registers_i.mstack_epc_q[12] ),
    .A2(_09594_),
    .B1(_09541_),
    .B2(_09378_),
    .ZN(_09608_));
 OAI21_X1 _28687_ (.A(_09608_),
    .B1(_09583_),
    .B2(_04528_),
    .ZN(_09609_));
 MUX2_X1 _28688_ (.A(\cs_registers_i.csr_mepc_o[12] ),
    .B(_09609_),
    .S(_09602_),
    .Z(_02936_));
 CLKBUF_X3 _28689_ (.A(_09563_),
    .Z(_09610_));
 AOI22_X1 _28690_ (.A1(\cs_registers_i.mstack_epc_q[13] ),
    .A2(_09610_),
    .B1(_09541_),
    .B2(_09381_),
    .ZN(_09611_));
 OAI21_X1 _28691_ (.A(_09611_),
    .B1(_09583_),
    .B2(_04562_),
    .ZN(_09612_));
 MUX2_X1 _28692_ (.A(\cs_registers_i.csr_mepc_o[13] ),
    .B(_09612_),
    .S(_09602_),
    .Z(_02937_));
 AOI22_X1 _28693_ (.A1(\cs_registers_i.mstack_epc_q[14] ),
    .A2(_09610_),
    .B1(_09541_),
    .B2(_09385_),
    .ZN(_09613_));
 OAI21_X1 _28694_ (.A(_09613_),
    .B1(_09583_),
    .B2(_04596_),
    .ZN(_09614_));
 MUX2_X1 _28695_ (.A(\cs_registers_i.csr_mepc_o[14] ),
    .B(_09614_),
    .S(_09602_),
    .Z(_02938_));
 AOI22_X1 _28696_ (.A1(\cs_registers_i.mstack_epc_q[15] ),
    .A2(_09610_),
    .B1(_09541_),
    .B2(_09388_),
    .ZN(_09615_));
 OAI21_X1 _28697_ (.A(_09615_),
    .B1(_09583_),
    .B2(_04620_),
    .ZN(_09616_));
 MUX2_X1 _28698_ (.A(\cs_registers_i.csr_mepc_o[15] ),
    .B(_09616_),
    .S(_09602_),
    .Z(_02939_));
 AOI22_X1 _28699_ (.A1(\cs_registers_i.mstack_epc_q[16] ),
    .A2(_09610_),
    .B1(_09541_),
    .B2(_09390_),
    .ZN(_09617_));
 OAI21_X1 _28700_ (.A(_09617_),
    .B1(_09583_),
    .B2(_04645_),
    .ZN(_09618_));
 MUX2_X1 _28701_ (.A(\cs_registers_i.csr_mepc_o[16] ),
    .B(_09618_),
    .S(_09602_),
    .Z(_02940_));
 AOI22_X1 _28702_ (.A1(\cs_registers_i.mstack_epc_q[17] ),
    .A2(_09610_),
    .B1(_09541_),
    .B2(_09393_),
    .ZN(_09619_));
 OAI21_X1 _28703_ (.A(_09619_),
    .B1(_09583_),
    .B2(_04665_),
    .ZN(_09620_));
 BUF_X4 _28704_ (.A(_09601_),
    .Z(_09621_));
 MUX2_X1 _28705_ (.A(\cs_registers_i.csr_mepc_o[17] ),
    .B(_09620_),
    .S(_09621_),
    .Z(_02941_));
 AOI22_X1 _28706_ (.A1(\cs_registers_i.mstack_epc_q[18] ),
    .A2(_09610_),
    .B1(_09541_),
    .B2(_09396_),
    .ZN(_09622_));
 CLKBUF_X3 _28707_ (.A(_09558_),
    .Z(_09623_));
 OAI21_X1 _28708_ (.A(_09622_),
    .B1(_09623_),
    .B2(_04685_),
    .ZN(_09624_));
 MUX2_X1 _28709_ (.A(\cs_registers_i.csr_mepc_o[18] ),
    .B(_09624_),
    .S(_09621_),
    .Z(_02942_));
 BUF_X2 _28710_ (.A(_09540_),
    .Z(_09625_));
 AOI22_X1 _28711_ (.A1(\cs_registers_i.mstack_epc_q[19] ),
    .A2(_09610_),
    .B1(_09625_),
    .B2(_09400_),
    .ZN(_09626_));
 OAI21_X1 _28712_ (.A(_09626_),
    .B1(_09623_),
    .B2(_04700_),
    .ZN(_09627_));
 MUX2_X1 _28713_ (.A(\cs_registers_i.csr_mepc_o[19] ),
    .B(_09627_),
    .S(_09621_),
    .Z(_02943_));
 OAI22_X1 _28714_ (.A1(\cs_registers_i.mstack_epc_q[1] ),
    .A2(_09555_),
    .B1(_09557_),
    .B2(_09404_),
    .ZN(_09628_));
 AOI21_X1 _28715_ (.A(_09628_),
    .B1(_09573_),
    .B2(_08519_),
    .ZN(_09629_));
 MUX2_X1 _28716_ (.A(\cs_registers_i.csr_mepc_o[1] ),
    .B(_09629_),
    .S(_09621_),
    .Z(_02944_));
 AOI22_X1 _28717_ (.A1(\cs_registers_i.mstack_epc_q[20] ),
    .A2(_09610_),
    .B1(_09625_),
    .B2(_09407_),
    .ZN(_09630_));
 OAI21_X1 _28718_ (.A(_09630_),
    .B1(_09623_),
    .B2(_04721_),
    .ZN(_09631_));
 MUX2_X1 _28719_ (.A(\cs_registers_i.csr_mepc_o[20] ),
    .B(_09631_),
    .S(_09621_),
    .Z(_02945_));
 AOI22_X1 _28720_ (.A1(\cs_registers_i.mstack_epc_q[21] ),
    .A2(_09610_),
    .B1(_09625_),
    .B2(_09412_),
    .ZN(_09632_));
 OAI21_X1 _28721_ (.A(_09632_),
    .B1(_09623_),
    .B2(_04742_),
    .ZN(_09633_));
 MUX2_X1 _28722_ (.A(\cs_registers_i.csr_mepc_o[21] ),
    .B(_09633_),
    .S(_09621_),
    .Z(_02946_));
 AOI22_X1 _28723_ (.A1(\cs_registers_i.mstack_epc_q[22] ),
    .A2(_09610_),
    .B1(_09625_),
    .B2(_09415_),
    .ZN(_09634_));
 OAI21_X1 _28724_ (.A(_09634_),
    .B1(_09623_),
    .B2(_04762_),
    .ZN(_09635_));
 MUX2_X1 _28725_ (.A(\cs_registers_i.csr_mepc_o[22] ),
    .B(_09635_),
    .S(_09621_),
    .Z(_02947_));
 CLKBUF_X3 _28726_ (.A(_09563_),
    .Z(_09636_));
 AOI22_X1 _28727_ (.A1(\cs_registers_i.mstack_epc_q[23] ),
    .A2(_09636_),
    .B1(_09625_),
    .B2(_09419_),
    .ZN(_09637_));
 OAI21_X1 _28728_ (.A(_09637_),
    .B1(_09623_),
    .B2(_04783_),
    .ZN(_09638_));
 MUX2_X1 _28729_ (.A(\cs_registers_i.csr_mepc_o[23] ),
    .B(_09638_),
    .S(_09621_),
    .Z(_02948_));
 AOI22_X1 _28730_ (.A1(\cs_registers_i.mstack_epc_q[24] ),
    .A2(_09636_),
    .B1(_09625_),
    .B2(_09422_),
    .ZN(_09639_));
 OAI21_X1 _28731_ (.A(_09639_),
    .B1(_09623_),
    .B2(_04805_),
    .ZN(_09640_));
 MUX2_X1 _28732_ (.A(\cs_registers_i.csr_mepc_o[24] ),
    .B(_09640_),
    .S(_09621_),
    .Z(_02949_));
 AOI22_X1 _28733_ (.A1(\cs_registers_i.mstack_epc_q[25] ),
    .A2(_09636_),
    .B1(_09625_),
    .B2(_09425_),
    .ZN(_09641_));
 OAI21_X1 _28734_ (.A(_09641_),
    .B1(_09623_),
    .B2(_04822_),
    .ZN(_09642_));
 MUX2_X1 _28735_ (.A(\cs_registers_i.csr_mepc_o[25] ),
    .B(_09642_),
    .S(_09621_),
    .Z(_02950_));
 AOI22_X1 _28736_ (.A1(\cs_registers_i.mstack_epc_q[26] ),
    .A2(_09636_),
    .B1(_09625_),
    .B2(_09428_),
    .ZN(_09643_));
 OAI21_X1 _28737_ (.A(_09643_),
    .B1(_09623_),
    .B2(_04838_),
    .ZN(_09644_));
 BUF_X4 _28738_ (.A(_09601_),
    .Z(_09645_));
 MUX2_X1 _28739_ (.A(\cs_registers_i.csr_mepc_o[26] ),
    .B(_09644_),
    .S(_09645_),
    .Z(_02951_));
 AOI22_X1 _28740_ (.A1(\cs_registers_i.mstack_epc_q[27] ),
    .A2(_09636_),
    .B1(_09625_),
    .B2(_09431_),
    .ZN(_09646_));
 OAI21_X1 _28741_ (.A(_09646_),
    .B1(_09623_),
    .B2(_04852_),
    .ZN(_09647_));
 MUX2_X1 _28742_ (.A(\cs_registers_i.csr_mepc_o[27] ),
    .B(_09647_),
    .S(_09645_),
    .Z(_02952_));
 AOI22_X1 _28743_ (.A1(\cs_registers_i.mstack_epc_q[28] ),
    .A2(_09636_),
    .B1(_09625_),
    .B2(_09434_),
    .ZN(_09648_));
 OAI21_X1 _28744_ (.A(_09648_),
    .B1(_09558_),
    .B2(_04868_),
    .ZN(_09649_));
 MUX2_X1 _28745_ (.A(\cs_registers_i.csr_mepc_o[28] ),
    .B(_09649_),
    .S(_09645_),
    .Z(_02953_));
 BUF_X4 _28746_ (.A(_09540_),
    .Z(_09650_));
 AOI22_X1 _28747_ (.A1(\cs_registers_i.mstack_epc_q[29] ),
    .A2(_09636_),
    .B1(_09650_),
    .B2(_09437_),
    .ZN(_09651_));
 OAI21_X1 _28748_ (.A(_09651_),
    .B1(_09558_),
    .B2(_04885_),
    .ZN(_09652_));
 MUX2_X1 _28749_ (.A(\cs_registers_i.csr_mepc_o[29] ),
    .B(_09652_),
    .S(_09645_),
    .Z(_02954_));
 NOR2_X1 _28750_ (.A1(\cs_registers_i.mstack_epc_q[2] ),
    .A2(_09555_),
    .ZN(_09653_));
 AOI221_X1 _28751_ (.A(_09653_),
    .B1(_09540_),
    .B2(_09440_),
    .C1(_09029_),
    .C2(_09573_),
    .ZN(_09654_));
 MUX2_X1 _28752_ (.A(\cs_registers_i.csr_mepc_o[2] ),
    .B(_09654_),
    .S(_09645_),
    .Z(_02955_));
 AOI22_X1 _28753_ (.A1(\cs_registers_i.mstack_epc_q[30] ),
    .A2(_09636_),
    .B1(_09650_),
    .B2(_09443_),
    .ZN(_09655_));
 OAI21_X1 _28754_ (.A(_09655_),
    .B1(_09558_),
    .B2(_04904_),
    .ZN(_09656_));
 MUX2_X1 _28755_ (.A(\cs_registers_i.csr_mepc_o[30] ),
    .B(_09656_),
    .S(_09645_),
    .Z(_02956_));
 OAI22_X1 _28756_ (.A1(\cs_registers_i.mstack_epc_q[31] ),
    .A2(_09555_),
    .B1(_09557_),
    .B2(_09446_),
    .ZN(_09657_));
 AOI21_X1 _28757_ (.A(_09657_),
    .B1(_09573_),
    .B2(_04924_),
    .ZN(_09658_));
 MUX2_X1 _28758_ (.A(\cs_registers_i.csr_mepc_o[31] ),
    .B(_09658_),
    .S(_09645_),
    .Z(_02957_));
 OAI22_X1 _28759_ (.A1(\cs_registers_i.mstack_epc_q[3] ),
    .A2(_09555_),
    .B1(_09557_),
    .B2(_09449_),
    .ZN(_09659_));
 AOI21_X1 _28760_ (.A(_09659_),
    .B1(_09573_),
    .B2(_08629_),
    .ZN(_09660_));
 MUX2_X1 _28761_ (.A(\cs_registers_i.csr_mepc_o[3] ),
    .B(_09660_),
    .S(_09645_),
    .Z(_02958_));
 OAI22_X1 _28762_ (.A1(\cs_registers_i.mstack_epc_q[4] ),
    .A2(_09555_),
    .B1(_09557_),
    .B2(_09452_),
    .ZN(_09661_));
 AOI21_X1 _28763_ (.A(_09661_),
    .B1(_09573_),
    .B2(_08639_),
    .ZN(_09662_));
 MUX2_X1 _28764_ (.A(\cs_registers_i.csr_mepc_o[4] ),
    .B(_09662_),
    .S(_09645_),
    .Z(_02959_));
 AOI22_X1 _28765_ (.A1(\cs_registers_i.mstack_epc_q[5] ),
    .A2(_09636_),
    .B1(_09650_),
    .B2(_09456_),
    .ZN(_09663_));
 OAI21_X1 _28766_ (.A(_09663_),
    .B1(_09558_),
    .B2(_08646_),
    .ZN(_09664_));
 MUX2_X1 _28767_ (.A(\cs_registers_i.csr_mepc_o[5] ),
    .B(_09664_),
    .S(_09645_),
    .Z(_02960_));
 AOI22_X1 _28768_ (.A1(\cs_registers_i.mstack_epc_q[6] ),
    .A2(_09636_),
    .B1(_09650_),
    .B2(_09459_),
    .ZN(_09665_));
 OAI21_X1 _28769_ (.A(_09665_),
    .B1(_09558_),
    .B2(_08655_),
    .ZN(_09666_));
 MUX2_X1 _28770_ (.A(\cs_registers_i.csr_mepc_o[6] ),
    .B(_09666_),
    .S(_09601_),
    .Z(_02961_));
 NOR2_X1 _28771_ (.A1(\cs_registers_i.csr_mepc_o[7] ),
    .A2(_09602_),
    .ZN(_09667_));
 AND2_X1 _28772_ (.A1(_09462_),
    .A2(_09540_),
    .ZN(_09668_));
 AOI221_X2 _28773_ (.A(_09668_),
    .B1(_09573_),
    .B2(_08665_),
    .C1(\cs_registers_i.mstack_epc_q[7] ),
    .C2(_09594_),
    .ZN(_09669_));
 AOI21_X1 _28774_ (.A(_09667_),
    .B1(_09669_),
    .B2(_09602_),
    .ZN(_02962_));
 AOI22_X1 _28775_ (.A1(\cs_registers_i.mstack_epc_q[8] ),
    .A2(_09563_),
    .B1(_09650_),
    .B2(_09465_),
    .ZN(_09670_));
 OAI21_X1 _28776_ (.A(_09670_),
    .B1(_09558_),
    .B2(_04942_),
    .ZN(_09671_));
 MUX2_X1 _28777_ (.A(\cs_registers_i.csr_mepc_o[8] ),
    .B(_09671_),
    .S(_09601_),
    .Z(_02963_));
 AOI22_X1 _28778_ (.A1(\cs_registers_i.mstack_epc_q[9] ),
    .A2(_09563_),
    .B1(_09650_),
    .B2(_09468_),
    .ZN(_09672_));
 OAI21_X1 _28779_ (.A(_09672_),
    .B1(_09558_),
    .B2(_04960_),
    .ZN(_09673_));
 MUX2_X1 _28780_ (.A(\cs_registers_i.csr_mepc_o[9] ),
    .B(_09673_),
    .S(_09601_),
    .Z(_02964_));
 NOR3_X4 _28781_ (.A1(_04429_),
    .A2(_04656_),
    .A3(_04542_),
    .ZN(_09674_));
 BUF_X4 _28782_ (.A(_09674_),
    .Z(_09675_));
 MUX2_X1 _28783_ (.A(\cs_registers_i.mie_q[0] ),
    .B(_08493_),
    .S(_09675_),
    .Z(_02965_));
 INV_X1 _28784_ (.A(_04838_),
    .ZN(_09676_));
 MUX2_X1 _28785_ (.A(\cs_registers_i.mie_q[10] ),
    .B(_09676_),
    .S(_09675_),
    .Z(_02966_));
 INV_X1 _28786_ (.A(_04853_),
    .ZN(_09677_));
 MUX2_X1 _28787_ (.A(\cs_registers_i.mie_q[11] ),
    .B(_09677_),
    .S(_09675_),
    .Z(_02967_));
 INV_X1 _28788_ (.A(_04868_),
    .ZN(_09678_));
 MUX2_X1 _28789_ (.A(\cs_registers_i.mie_q[12] ),
    .B(_09678_),
    .S(_09675_),
    .Z(_02968_));
 MUX2_X1 _28790_ (.A(\cs_registers_i.mie_q[13] ),
    .B(_09308_),
    .S(_09675_),
    .Z(_02969_));
 INV_X1 _28791_ (.A(_04905_),
    .ZN(_09679_));
 MUX2_X1 _28792_ (.A(\cs_registers_i.mie_q[14] ),
    .B(_09679_),
    .S(_09675_),
    .Z(_02970_));
 MUX2_X1 _28793_ (.A(\cs_registers_i.mie_q[15] ),
    .B(_09353_),
    .S(_09675_),
    .Z(_02971_));
 MUX2_X1 _28794_ (.A(\cs_registers_i.mie_q[16] ),
    .B(_08666_),
    .S(_09675_),
    .Z(_02972_));
 MUX2_X1 _28795_ (.A(\cs_registers_i.mie_q[17] ),
    .B(_08630_),
    .S(_09675_),
    .Z(_02973_));
 MUX2_X1 _28796_ (.A(\cs_registers_i.mie_q[1] ),
    .B(_09200_),
    .S(_09675_),
    .Z(_02974_));
 MUX2_X1 _28797_ (.A(\cs_registers_i.mie_q[2] ),
    .B(_08743_),
    .S(_09674_),
    .Z(_02975_));
 MUX2_X1 _28798_ (.A(\cs_registers_i.mie_q[3] ),
    .B(_09222_),
    .S(_09674_),
    .Z(_02976_));
 INV_X1 _28799_ (.A(\cs_registers_i.mie_q[4] ),
    .ZN(_09680_));
 MUX2_X1 _28800_ (.A(_09680_),
    .B(_04721_),
    .S(_09674_),
    .Z(_09681_));
 INV_X1 _28801_ (.A(_09681_),
    .ZN(_02977_));
 MUX2_X1 _28802_ (.A(\cs_registers_i.mie_q[5] ),
    .B(_08971_),
    .S(_09674_),
    .Z(_02978_));
 MUX2_X1 _28803_ (.A(\cs_registers_i.mie_q[6] ),
    .B(_08765_),
    .S(_09674_),
    .Z(_02979_));
 MUX2_X1 _28804_ (.A(\cs_registers_i.mie_q[7] ),
    .B(_08982_),
    .S(_09674_),
    .Z(_02980_));
 INV_X1 _28805_ (.A(_04805_),
    .ZN(_09682_));
 MUX2_X1 _28806_ (.A(\cs_registers_i.mie_q[8] ),
    .B(_09682_),
    .S(_09674_),
    .Z(_02981_));
 MUX2_X1 _28807_ (.A(\cs_registers_i.mie_q[9] ),
    .B(_09271_),
    .S(_09674_),
    .Z(_02982_));
 NAND2_X2 _28808_ (.A1(_04575_),
    .A2(_09044_),
    .ZN(_09683_));
 BUF_X4 _28809_ (.A(_09683_),
    .Z(_09684_));
 MUX2_X1 _28810_ (.A(_08396_),
    .B(\cs_registers_i.mscratch_q[0] ),
    .S(_09684_),
    .Z(_02983_));
 MUX2_X1 _28811_ (.A(_08867_),
    .B(\cs_registers_i.mscratch_q[10] ),
    .S(_09684_),
    .Z(_02984_));
 BUF_X4 _28812_ (.A(_09683_),
    .Z(_09685_));
 NAND2_X1 _28813_ (.A1(\cs_registers_i.mscratch_q[11] ),
    .A2(_09685_),
    .ZN(_09686_));
 BUF_X4 _28814_ (.A(_09684_),
    .Z(_09687_));
 OAI21_X1 _28815_ (.A(_09686_),
    .B1(_09687_),
    .B2(_04472_),
    .ZN(_02985_));
 NAND2_X1 _28816_ (.A1(\cs_registers_i.mscratch_q[12] ),
    .A2(_09685_),
    .ZN(_09688_));
 OAI21_X1 _28817_ (.A(_09688_),
    .B1(_09687_),
    .B2(_04528_),
    .ZN(_02986_));
 NAND2_X1 _28818_ (.A1(\cs_registers_i.mscratch_q[13] ),
    .A2(_09685_),
    .ZN(_09689_));
 OAI21_X1 _28819_ (.A(_09689_),
    .B1(_09687_),
    .B2(_04562_),
    .ZN(_02987_));
 CLKBUF_X3 _28820_ (.A(_09683_),
    .Z(_09690_));
 NAND2_X1 _28821_ (.A1(\cs_registers_i.mscratch_q[14] ),
    .A2(_09690_),
    .ZN(_09691_));
 OAI21_X1 _28822_ (.A(_09691_),
    .B1(_09687_),
    .B2(_04597_),
    .ZN(_02988_));
 NAND2_X1 _28823_ (.A1(\cs_registers_i.mscratch_q[15] ),
    .A2(_09690_),
    .ZN(_09692_));
 OAI21_X1 _28824_ (.A(_09692_),
    .B1(_09687_),
    .B2(_04620_),
    .ZN(_02989_));
 MUX2_X1 _28825_ (.A(_08493_),
    .B(\cs_registers_i.mscratch_q[16] ),
    .S(_09684_),
    .Z(_02990_));
 NAND2_X1 _28826_ (.A1(\cs_registers_i.mscratch_q[17] ),
    .A2(_09690_),
    .ZN(_09693_));
 OAI21_X1 _28827_ (.A(_09693_),
    .B1(_09687_),
    .B2(_04665_),
    .ZN(_02991_));
 NAND2_X1 _28828_ (.A1(\cs_registers_i.mscratch_q[18] ),
    .A2(_09690_),
    .ZN(_09694_));
 OAI21_X1 _28829_ (.A(_09694_),
    .B1(_09687_),
    .B2(_04685_),
    .ZN(_02992_));
 NAND2_X1 _28830_ (.A1(\cs_registers_i.mscratch_q[19] ),
    .A2(_09690_),
    .ZN(_09695_));
 OAI21_X1 _28831_ (.A(_09695_),
    .B1(_09687_),
    .B2(_04700_),
    .ZN(_02993_));
 NAND2_X1 _28832_ (.A1(\cs_registers_i.mscratch_q[1] ),
    .A2(_09690_),
    .ZN(_09696_));
 OAI21_X1 _28833_ (.A(_09696_),
    .B1(_09687_),
    .B2(_08519_),
    .ZN(_02994_));
 NAND2_X1 _28834_ (.A1(\cs_registers_i.mscratch_q[20] ),
    .A2(_09690_),
    .ZN(_09697_));
 OAI21_X1 _28835_ (.A(_09697_),
    .B1(_09687_),
    .B2(_04721_),
    .ZN(_02995_));
 NAND2_X1 _28836_ (.A1(\cs_registers_i.mscratch_q[21] ),
    .A2(_09690_),
    .ZN(_09698_));
 CLKBUF_X3 _28837_ (.A(_09683_),
    .Z(_09699_));
 OAI21_X1 _28838_ (.A(_09698_),
    .B1(_09699_),
    .B2(_04742_),
    .ZN(_02996_));
 NAND2_X1 _28839_ (.A1(\cs_registers_i.mscratch_q[22] ),
    .A2(_09690_),
    .ZN(_09700_));
 OAI21_X1 _28840_ (.A(_09700_),
    .B1(_09699_),
    .B2(_04762_),
    .ZN(_02997_));
 NAND2_X1 _28841_ (.A1(\cs_registers_i.mscratch_q[23] ),
    .A2(_09690_),
    .ZN(_09701_));
 OAI21_X1 _28842_ (.A(_09701_),
    .B1(_09699_),
    .B2(_04783_),
    .ZN(_02998_));
 CLKBUF_X3 _28843_ (.A(_09683_),
    .Z(_09702_));
 NAND2_X1 _28844_ (.A1(\cs_registers_i.mscratch_q[24] ),
    .A2(_09702_),
    .ZN(_09703_));
 OAI21_X1 _28845_ (.A(_09703_),
    .B1(_09699_),
    .B2(_04805_),
    .ZN(_02999_));
 NAND2_X1 _28846_ (.A1(\cs_registers_i.mscratch_q[25] ),
    .A2(_09702_),
    .ZN(_09704_));
 OAI21_X1 _28847_ (.A(_09704_),
    .B1(_09699_),
    .B2(_04822_),
    .ZN(_03000_));
 NAND2_X1 _28848_ (.A1(\cs_registers_i.mscratch_q[26] ),
    .A2(_09702_),
    .ZN(_09705_));
 OAI21_X1 _28849_ (.A(_09705_),
    .B1(_09699_),
    .B2(_04838_),
    .ZN(_03001_));
 NAND2_X1 _28850_ (.A1(\cs_registers_i.mscratch_q[27] ),
    .A2(_09702_),
    .ZN(_09706_));
 OAI21_X1 _28851_ (.A(_09706_),
    .B1(_09699_),
    .B2(_04853_),
    .ZN(_03002_));
 NAND2_X1 _28852_ (.A1(\cs_registers_i.mscratch_q[28] ),
    .A2(_09702_),
    .ZN(_09707_));
 OAI21_X1 _28853_ (.A(_09707_),
    .B1(_09699_),
    .B2(_04868_),
    .ZN(_03003_));
 NAND2_X1 _28854_ (.A1(\cs_registers_i.mscratch_q[29] ),
    .A2(_09702_),
    .ZN(_09708_));
 OAI21_X1 _28855_ (.A(_09708_),
    .B1(_09699_),
    .B2(_04885_),
    .ZN(_03004_));
 MUX2_X1 _28856_ (.A(_08402_),
    .B(\cs_registers_i.mscratch_q[2] ),
    .S(_09684_),
    .Z(_03005_));
 NAND2_X1 _28857_ (.A1(\cs_registers_i.mscratch_q[30] ),
    .A2(_09702_),
    .ZN(_09709_));
 OAI21_X1 _28858_ (.A(_09709_),
    .B1(_09699_),
    .B2(_04905_),
    .ZN(_03006_));
 NAND2_X1 _28859_ (.A1(\cs_registers_i.mscratch_q[31] ),
    .A2(_09702_),
    .ZN(_09710_));
 OAI21_X1 _28860_ (.A(_09710_),
    .B1(_09685_),
    .B2(_04924_),
    .ZN(_03007_));
 NAND2_X1 _28861_ (.A1(\cs_registers_i.mscratch_q[3] ),
    .A2(_09702_),
    .ZN(_09711_));
 OAI21_X1 _28862_ (.A(_09711_),
    .B1(_09685_),
    .B2(_08629_),
    .ZN(_03008_));
 NAND2_X1 _28863_ (.A1(\cs_registers_i.mscratch_q[4] ),
    .A2(_09702_),
    .ZN(_09712_));
 OAI21_X1 _28864_ (.A(_09712_),
    .B1(_09685_),
    .B2(_08639_),
    .ZN(_03009_));
 NAND2_X1 _28865_ (.A1(\cs_registers_i.mscratch_q[5] ),
    .A2(_09684_),
    .ZN(_09713_));
 OAI21_X1 _28866_ (.A(_09713_),
    .B1(_09685_),
    .B2(_08646_),
    .ZN(_03010_));
 NAND2_X1 _28867_ (.A1(\cs_registers_i.mscratch_q[6] ),
    .A2(_09684_),
    .ZN(_09714_));
 OAI21_X1 _28868_ (.A(_09714_),
    .B1(_09685_),
    .B2(_08655_),
    .ZN(_03011_));
 MUX2_X1 _28869_ (.A(_08666_),
    .B(\cs_registers_i.mscratch_q[7] ),
    .S(_09684_),
    .Z(_03012_));
 NAND2_X1 _28870_ (.A1(\cs_registers_i.mscratch_q[8] ),
    .A2(_09684_),
    .ZN(_09715_));
 OAI21_X1 _28871_ (.A(_09715_),
    .B1(_09685_),
    .B2(_04942_),
    .ZN(_03013_));
 NAND2_X1 _28872_ (.A1(\cs_registers_i.mscratch_q[9] ),
    .A2(_09684_),
    .ZN(_09716_));
 OAI21_X1 _28873_ (.A(_09716_),
    .B1(_09685_),
    .B2(_04960_),
    .ZN(_03014_));
 CLKBUF_X3 _28874_ (.A(_09586_),
    .Z(_09717_));
 MUX2_X1 _28875_ (.A(\cs_registers_i.mstack_cause_q[0] ),
    .B(\cs_registers_i.mcause_q[0] ),
    .S(_09717_),
    .Z(_03015_));
 MUX2_X1 _28876_ (.A(\cs_registers_i.mstack_cause_q[1] ),
    .B(\cs_registers_i.mcause_q[1] ),
    .S(_09717_),
    .Z(_03016_));
 MUX2_X1 _28877_ (.A(\cs_registers_i.mstack_cause_q[2] ),
    .B(\cs_registers_i.mcause_q[2] ),
    .S(_09717_),
    .Z(_03017_));
 MUX2_X1 _28878_ (.A(\cs_registers_i.mstack_cause_q[3] ),
    .B(\cs_registers_i.mcause_q[3] ),
    .S(_09717_),
    .Z(_03018_));
 MUX2_X1 _28879_ (.A(\cs_registers_i.mstack_cause_q[4] ),
    .B(\cs_registers_i.mcause_q[4] ),
    .S(_09717_),
    .Z(_03019_));
 MUX2_X1 _28880_ (.A(\cs_registers_i.mstack_cause_q[5] ),
    .B(\cs_registers_i.mcause_q[5] ),
    .S(_09717_),
    .Z(_03020_));
 MUX2_X1 _28881_ (.A(\cs_registers_i.mstack_q[0] ),
    .B(\cs_registers_i.mstack_d[0] ),
    .S(_09717_),
    .Z(_03021_));
 MUX2_X1 _28882_ (.A(\cs_registers_i.mstack_q[1] ),
    .B(\cs_registers_i.mstack_d[1] ),
    .S(_09717_),
    .Z(_03022_));
 MUX2_X1 _28883_ (.A(\cs_registers_i.mstack_q[2] ),
    .B(\cs_registers_i.mstack_d[2] ),
    .S(_09717_),
    .Z(_03023_));
 MUX2_X1 _28884_ (.A(\cs_registers_i.mstack_epc_q[0] ),
    .B(\cs_registers_i.csr_mepc_o[0] ),
    .S(_09717_),
    .Z(_03024_));
 BUF_X4 _28885_ (.A(_09586_),
    .Z(_09718_));
 MUX2_X1 _28886_ (.A(\cs_registers_i.mstack_epc_q[10] ),
    .B(\cs_registers_i.csr_mepc_o[10] ),
    .S(_09718_),
    .Z(_03025_));
 MUX2_X1 _28887_ (.A(\cs_registers_i.mstack_epc_q[11] ),
    .B(\cs_registers_i.csr_mepc_o[11] ),
    .S(_09718_),
    .Z(_03026_));
 MUX2_X1 _28888_ (.A(\cs_registers_i.mstack_epc_q[12] ),
    .B(\cs_registers_i.csr_mepc_o[12] ),
    .S(_09718_),
    .Z(_03027_));
 MUX2_X1 _28889_ (.A(\cs_registers_i.mstack_epc_q[13] ),
    .B(\cs_registers_i.csr_mepc_o[13] ),
    .S(_09718_),
    .Z(_03028_));
 MUX2_X1 _28890_ (.A(\cs_registers_i.mstack_epc_q[14] ),
    .B(\cs_registers_i.csr_mepc_o[14] ),
    .S(_09718_),
    .Z(_03029_));
 MUX2_X1 _28891_ (.A(\cs_registers_i.mstack_epc_q[15] ),
    .B(\cs_registers_i.csr_mepc_o[15] ),
    .S(_09718_),
    .Z(_03030_));
 MUX2_X1 _28892_ (.A(\cs_registers_i.mstack_epc_q[16] ),
    .B(\cs_registers_i.csr_mepc_o[16] ),
    .S(_09718_),
    .Z(_03031_));
 MUX2_X1 _28893_ (.A(\cs_registers_i.mstack_epc_q[17] ),
    .B(\cs_registers_i.csr_mepc_o[17] ),
    .S(_09718_),
    .Z(_03032_));
 MUX2_X1 _28894_ (.A(\cs_registers_i.mstack_epc_q[18] ),
    .B(\cs_registers_i.csr_mepc_o[18] ),
    .S(_09718_),
    .Z(_03033_));
 MUX2_X1 _28895_ (.A(\cs_registers_i.mstack_epc_q[19] ),
    .B(\cs_registers_i.csr_mepc_o[19] ),
    .S(_09718_),
    .Z(_03034_));
 BUF_X4 _28896_ (.A(_09586_),
    .Z(_09719_));
 MUX2_X1 _28897_ (.A(\cs_registers_i.mstack_epc_q[1] ),
    .B(\cs_registers_i.csr_mepc_o[1] ),
    .S(_09719_),
    .Z(_03035_));
 MUX2_X1 _28898_ (.A(\cs_registers_i.mstack_epc_q[20] ),
    .B(\cs_registers_i.csr_mepc_o[20] ),
    .S(_09719_),
    .Z(_03036_));
 MUX2_X1 _28899_ (.A(\cs_registers_i.mstack_epc_q[21] ),
    .B(\cs_registers_i.csr_mepc_o[21] ),
    .S(_09719_),
    .Z(_03037_));
 MUX2_X1 _28900_ (.A(\cs_registers_i.mstack_epc_q[22] ),
    .B(\cs_registers_i.csr_mepc_o[22] ),
    .S(_09719_),
    .Z(_03038_));
 MUX2_X1 _28901_ (.A(\cs_registers_i.mstack_epc_q[23] ),
    .B(\cs_registers_i.csr_mepc_o[23] ),
    .S(_09719_),
    .Z(_03039_));
 MUX2_X1 _28902_ (.A(\cs_registers_i.mstack_epc_q[24] ),
    .B(\cs_registers_i.csr_mepc_o[24] ),
    .S(_09719_),
    .Z(_03040_));
 MUX2_X1 _28903_ (.A(\cs_registers_i.mstack_epc_q[25] ),
    .B(\cs_registers_i.csr_mepc_o[25] ),
    .S(_09719_),
    .Z(_03041_));
 MUX2_X1 _28904_ (.A(\cs_registers_i.mstack_epc_q[26] ),
    .B(\cs_registers_i.csr_mepc_o[26] ),
    .S(_09719_),
    .Z(_03042_));
 MUX2_X1 _28905_ (.A(\cs_registers_i.mstack_epc_q[27] ),
    .B(\cs_registers_i.csr_mepc_o[27] ),
    .S(_09719_),
    .Z(_03043_));
 MUX2_X1 _28906_ (.A(\cs_registers_i.mstack_epc_q[28] ),
    .B(\cs_registers_i.csr_mepc_o[28] ),
    .S(_09719_),
    .Z(_03044_));
 BUF_X4 _28907_ (.A(_09586_),
    .Z(_09720_));
 MUX2_X1 _28908_ (.A(\cs_registers_i.mstack_epc_q[29] ),
    .B(\cs_registers_i.csr_mepc_o[29] ),
    .S(_09720_),
    .Z(_03045_));
 MUX2_X1 _28909_ (.A(\cs_registers_i.mstack_epc_q[2] ),
    .B(\cs_registers_i.csr_mepc_o[2] ),
    .S(_09720_),
    .Z(_03046_));
 MUX2_X1 _28910_ (.A(\cs_registers_i.mstack_epc_q[30] ),
    .B(\cs_registers_i.csr_mepc_o[30] ),
    .S(_09720_),
    .Z(_03047_));
 MUX2_X1 _28911_ (.A(\cs_registers_i.mstack_epc_q[31] ),
    .B(\cs_registers_i.csr_mepc_o[31] ),
    .S(_09720_),
    .Z(_03048_));
 MUX2_X1 _28912_ (.A(\cs_registers_i.mstack_epc_q[3] ),
    .B(\cs_registers_i.csr_mepc_o[3] ),
    .S(_09720_),
    .Z(_03049_));
 MUX2_X1 _28913_ (.A(\cs_registers_i.mstack_epc_q[4] ),
    .B(\cs_registers_i.csr_mepc_o[4] ),
    .S(_09720_),
    .Z(_03050_));
 MUX2_X1 _28914_ (.A(\cs_registers_i.mstack_epc_q[5] ),
    .B(\cs_registers_i.csr_mepc_o[5] ),
    .S(_09720_),
    .Z(_03051_));
 MUX2_X1 _28915_ (.A(\cs_registers_i.mstack_epc_q[6] ),
    .B(\cs_registers_i.csr_mepc_o[6] ),
    .S(_09720_),
    .Z(_03052_));
 MUX2_X1 _28916_ (.A(\cs_registers_i.mstack_epc_q[7] ),
    .B(\cs_registers_i.csr_mepc_o[7] ),
    .S(_09720_),
    .Z(_03053_));
 MUX2_X1 _28917_ (.A(\cs_registers_i.mstack_epc_q[8] ),
    .B(\cs_registers_i.csr_mepc_o[8] ),
    .S(_09720_),
    .Z(_03054_));
 CLKBUF_X3 _28918_ (.A(_09650_),
    .Z(_09721_));
 MUX2_X1 _28919_ (.A(\cs_registers_i.mstack_epc_q[9] ),
    .B(\cs_registers_i.csr_mepc_o[9] ),
    .S(_09721_),
    .Z(_03055_));
 NAND2_X1 _28920_ (.A1(_15908_),
    .A2(_04451_),
    .ZN(_09722_));
 NOR2_X1 _28921_ (.A1(_04542_),
    .A2(_09722_),
    .ZN(_09723_));
 MUX2_X1 _28922_ (.A(\cs_registers_i.csr_mstatus_tw_o ),
    .B(_08971_),
    .S(_09723_),
    .Z(_03056_));
 MUX2_X1 _28923_ (.A(\cs_registers_i.mstatus_q[1] ),
    .B(_09200_),
    .S(_09723_),
    .Z(_03057_));
 NOR2_X1 _28924_ (.A1(_07289_),
    .A2(_09561_),
    .ZN(_09724_));
 INV_X1 _28925_ (.A(_04404_),
    .ZN(_09725_));
 CLKBUF_X3 _28926_ (.A(_03618_),
    .Z(_09726_));
 NAND3_X1 _28927_ (.A1(_03555_),
    .A2(_11379_),
    .A3(_03596_),
    .ZN(_09727_));
 AOI21_X1 _28928_ (.A(_03552_),
    .B1(_09726_),
    .B2(_09727_),
    .ZN(_09728_));
 NOR2_X1 _28929_ (.A1(_11490_),
    .A2(_11379_),
    .ZN(_09729_));
 OAI21_X1 _28930_ (.A(_08404_),
    .B1(_03552_),
    .B2(_03636_),
    .ZN(_09730_));
 AND3_X1 _28931_ (.A1(_09726_),
    .A2(_09729_),
    .A3(_09730_),
    .ZN(_09731_));
 NOR3_X1 _28932_ (.A1(_04410_),
    .A2(_09728_),
    .A3(_09731_),
    .ZN(_09732_));
 AND4_X1 _28933_ (.A1(_03564_),
    .A2(_11492_),
    .A3(_03606_),
    .A4(_04437_),
    .ZN(_09733_));
 OAI21_X1 _28934_ (.A(_09725_),
    .B1(_09732_),
    .B2(_09733_),
    .ZN(_09734_));
 AOI21_X1 _28935_ (.A(_03632_),
    .B1(_03634_),
    .B2(_03596_),
    .ZN(_09735_));
 NOR2_X1 _28936_ (.A1(_03631_),
    .A2(_09735_),
    .ZN(_09736_));
 NAND2_X1 _28937_ (.A1(_04409_),
    .A2(_16262_),
    .ZN(_09737_));
 AOI21_X1 _28938_ (.A(_03554_),
    .B1(_04577_),
    .B2(_09737_),
    .ZN(_09738_));
 OR4_X2 _28939_ (.A1(_03631_),
    .A2(_16330_),
    .A3(_03560_),
    .A4(_04411_),
    .ZN(_09739_));
 NOR3_X1 _28940_ (.A1(_09736_),
    .A2(_09738_),
    .A3(_09739_),
    .ZN(_09740_));
 NAND2_X1 _28941_ (.A1(_11379_),
    .A2(_03618_),
    .ZN(_09741_));
 NAND3_X1 _28942_ (.A1(_03584_),
    .A2(_04439_),
    .A3(_09741_),
    .ZN(_09742_));
 NAND2_X1 _28943_ (.A1(_03556_),
    .A2(_03640_),
    .ZN(_09743_));
 AOI221_X1 _28944_ (.A(_09742_),
    .B1(_09726_),
    .B2(_04409_),
    .C1(_03589_),
    .C2(_09743_),
    .ZN(_09744_));
 NAND3_X1 _28945_ (.A1(_04437_),
    .A2(_04439_),
    .A3(_04444_),
    .ZN(_09745_));
 AOI21_X1 _28946_ (.A(_04429_),
    .B1(_04420_),
    .B2(_09745_),
    .ZN(_09746_));
 NOR3_X1 _28947_ (.A1(_09740_),
    .A2(_09744_),
    .A3(_09746_),
    .ZN(_09747_));
 OR2_X2 _28948_ (.A1(_16270_),
    .A2(_04410_),
    .ZN(_09748_));
 NOR4_X4 _28949_ (.A1(_03560_),
    .A2(_03561_),
    .A3(_04373_),
    .A4(_09748_),
    .ZN(_09749_));
 INV_X1 _28950_ (.A(_03618_),
    .ZN(_09750_));
 NOR2_X1 _28951_ (.A1(_04409_),
    .A2(_09750_),
    .ZN(_09751_));
 NOR4_X4 _28952_ (.A1(_03561_),
    .A2(_04373_),
    .A3(_03566_),
    .A4(_09748_),
    .ZN(_09752_));
 AOI22_X1 _28953_ (.A1(_15908_),
    .A2(_09749_),
    .B1(_09751_),
    .B2(_09752_),
    .ZN(_09753_));
 NAND2_X1 _28954_ (.A1(_16270_),
    .A2(_04455_),
    .ZN(_09754_));
 OAI21_X1 _28955_ (.A(_03555_),
    .B1(_04577_),
    .B2(_04409_),
    .ZN(_09755_));
 NOR2_X1 _28956_ (.A1(_03552_),
    .A2(_03551_),
    .ZN(_09756_));
 OAI21_X1 _28957_ (.A(_16266_),
    .B1(_09756_),
    .B2(_11379_),
    .ZN(_09757_));
 AOI22_X1 _28958_ (.A1(_09750_),
    .A2(_09755_),
    .B1(_09757_),
    .B2(_03581_),
    .ZN(_09758_));
 OAI21_X1 _28959_ (.A(_09753_),
    .B1(_09754_),
    .B2(_09758_),
    .ZN(_09759_));
 NOR2_X1 _28960_ (.A1(_04410_),
    .A2(_04404_),
    .ZN(_09760_));
 NAND3_X1 _28961_ (.A1(_16266_),
    .A2(_08404_),
    .A3(_09760_),
    .ZN(_09761_));
 AOI221_X2 _28962_ (.A(_04410_),
    .B1(_04440_),
    .B2(_04404_),
    .C1(_09761_),
    .C2(_04383_),
    .ZN(_09762_));
 AOI21_X1 _28963_ (.A(_09759_),
    .B1(_09762_),
    .B2(_03633_),
    .ZN(_09763_));
 AOI22_X2 _28964_ (.A1(_11490_),
    .A2(_03632_),
    .B1(_03634_),
    .B2(_03554_),
    .ZN(_09764_));
 OAI22_X2 _28965_ (.A1(_04409_),
    .A2(_09726_),
    .B1(_09764_),
    .B2(_03631_),
    .ZN(_09765_));
 NAND3_X1 _28966_ (.A1(_03554_),
    .A2(_11379_),
    .A3(_09726_),
    .ZN(_09766_));
 AOI22_X1 _28967_ (.A1(_03640_),
    .A2(_09741_),
    .B1(_09766_),
    .B2(_03589_),
    .ZN(_09767_));
 OAI21_X1 _28968_ (.A(_09752_),
    .B1(_09765_),
    .B2(_09767_),
    .ZN(_09768_));
 NAND4_X1 _28969_ (.A1(_09734_),
    .A2(_09747_),
    .A3(_09763_),
    .A4(_09768_),
    .ZN(_09769_));
 NAND2_X1 _28970_ (.A1(_09726_),
    .A2(_08404_),
    .ZN(_09770_));
 NOR2_X1 _28971_ (.A1(_16270_),
    .A2(_06499_),
    .ZN(_09771_));
 OR3_X1 _28972_ (.A1(_09752_),
    .A2(_09760_),
    .A3(_09771_),
    .ZN(_09772_));
 AOI222_X2 _28973_ (.A1(_03636_),
    .A2(_04399_),
    .B1(_09752_),
    .B2(_03551_),
    .C1(_09772_),
    .C2(_03554_),
    .ZN(_09773_));
 INV_X1 _28974_ (.A(_04385_),
    .ZN(_09774_));
 AOI21_X1 _28975_ (.A(_11490_),
    .B1(_04452_),
    .B2(_09774_),
    .ZN(_09775_));
 AOI21_X1 _28976_ (.A(_09775_),
    .B1(_09739_),
    .B2(_04420_),
    .ZN(_09776_));
 OAI21_X1 _28977_ (.A(_09754_),
    .B1(_04537_),
    .B2(_04373_),
    .ZN(_09777_));
 AOI221_X2 _28978_ (.A(_09776_),
    .B1(_09777_),
    .B2(_03551_),
    .C1(_03556_),
    .C2(_09749_),
    .ZN(_09778_));
 OAI22_X1 _28979_ (.A1(_09770_),
    .A2(_09773_),
    .B1(_09778_),
    .B2(_04383_),
    .ZN(_09779_));
 NAND3_X1 _28980_ (.A1(_04383_),
    .A2(_03584_),
    .A3(_04439_),
    .ZN(_09780_));
 AOI22_X1 _28981_ (.A1(_03576_),
    .A2(_04409_),
    .B1(_03618_),
    .B2(_08404_),
    .ZN(_09781_));
 OAI22_X1 _28982_ (.A1(_03552_),
    .A2(_09726_),
    .B1(_09781_),
    .B2(_03636_),
    .ZN(_09782_));
 AOI21_X1 _28983_ (.A(_09780_),
    .B1(_09782_),
    .B2(_03555_),
    .ZN(_09783_));
 NOR3_X1 _28984_ (.A1(_11490_),
    .A2(_03554_),
    .A3(_09726_),
    .ZN(_09784_));
 AOI21_X1 _28985_ (.A(_09729_),
    .B1(_03637_),
    .B2(_03632_),
    .ZN(_09785_));
 NOR2_X1 _28986_ (.A1(_03631_),
    .A2(_09785_),
    .ZN(_09786_));
 OAI221_X1 _28987_ (.A(_04409_),
    .B1(_03631_),
    .B2(_03635_),
    .C1(_09784_),
    .C2(_09786_),
    .ZN(_09787_));
 AOI21_X1 _28988_ (.A(_09783_),
    .B1(_09787_),
    .B2(_09771_),
    .ZN(_09788_));
 MUX2_X1 _28989_ (.A(_03556_),
    .B(_03551_),
    .S(_04577_),
    .Z(_09789_));
 AOI21_X1 _28990_ (.A(_09765_),
    .B1(_09789_),
    .B2(_09726_),
    .ZN(_09790_));
 OAI21_X1 _28991_ (.A(_09788_),
    .B1(_09790_),
    .B2(_09739_),
    .ZN(_09791_));
 NOR2_X1 _28992_ (.A1(_04410_),
    .A2(_04440_),
    .ZN(_09792_));
 NOR2_X1 _28993_ (.A1(_11379_),
    .A2(_03577_),
    .ZN(_09793_));
 AOI21_X1 _28994_ (.A(_04385_),
    .B1(_16262_),
    .B2(_16253_),
    .ZN(_09794_));
 OAI221_X1 _28995_ (.A(_11329_),
    .B1(_16262_),
    .B2(_09793_),
    .C1(_09794_),
    .C2(_11490_),
    .ZN(_09795_));
 NAND2_X1 _28996_ (.A1(_03555_),
    .A2(_16262_),
    .ZN(_09796_));
 AOI21_X1 _28997_ (.A(_03552_),
    .B1(_04577_),
    .B2(_09796_),
    .ZN(_09797_));
 OAI21_X1 _28998_ (.A(_09795_),
    .B1(_09797_),
    .B2(_09736_),
    .ZN(_09798_));
 OAI21_X1 _28999_ (.A(_11492_),
    .B1(_04451_),
    .B2(_09749_),
    .ZN(_09799_));
 OAI21_X1 _29000_ (.A(_09799_),
    .B1(_09741_),
    .B2(_09739_),
    .ZN(_09800_));
 AOI22_X1 _29001_ (.A1(_09792_),
    .A2(_09798_),
    .B1(_09800_),
    .B2(_03636_),
    .ZN(_09801_));
 NOR3_X1 _29002_ (.A1(_03589_),
    .A2(_03631_),
    .A3(_03603_),
    .ZN(_09802_));
 AOI22_X1 _29003_ (.A1(_11490_),
    .A2(_04511_),
    .B1(_09802_),
    .B2(_04451_),
    .ZN(_09803_));
 AND3_X1 _29004_ (.A1(_03584_),
    .A2(_04439_),
    .A3(_09741_),
    .ZN(_09804_));
 NOR2_X1 _29005_ (.A1(_09762_),
    .A2(_09804_),
    .ZN(_09805_));
 OAI221_X1 _29006_ (.A(_09801_),
    .B1(_09803_),
    .B2(_09726_),
    .C1(_09805_),
    .C2(_03576_),
    .ZN(_09806_));
 OR4_X1 _29007_ (.A1(_09769_),
    .A2(_09779_),
    .A3(_09791_),
    .A4(_09806_),
    .ZN(_09807_));
 NAND4_X2 _29008_ (.A1(_15908_),
    .A2(_03541_),
    .A3(_04531_),
    .A4(_09807_),
    .ZN(_09808_));
 OAI21_X1 _29009_ (.A(_09724_),
    .B1(_09808_),
    .B2(_04656_),
    .ZN(_09809_));
 AOI22_X1 _29010_ (.A1(\cs_registers_i.mstack_q[0] ),
    .A2(_09594_),
    .B1(_09586_),
    .B2(_03660_),
    .ZN(_09810_));
 INV_X1 _29011_ (.A(_09810_),
    .ZN(_09811_));
 OR2_X2 _29012_ (.A1(_04542_),
    .A2(_09722_),
    .ZN(_09812_));
 AOI21_X1 _29013_ (.A(_09812_),
    .B1(_04527_),
    .B2(_04471_),
    .ZN(_09813_));
 OAI21_X1 _29014_ (.A(_09809_),
    .B1(_09811_),
    .B2(_09813_),
    .ZN(_09814_));
 AOI21_X1 _29015_ (.A(_07289_),
    .B1(_09561_),
    .B2(_09721_),
    .ZN(_09815_));
 NAND2_X1 _29016_ (.A1(_09812_),
    .A2(_09815_),
    .ZN(_09816_));
 INV_X1 _29017_ (.A(\cs_registers_i.mstack_d[0] ),
    .ZN(_09817_));
 OAI21_X1 _29018_ (.A(_09814_),
    .B1(_09816_),
    .B2(_09817_),
    .ZN(_03058_));
 AOI22_X1 _29019_ (.A1(\cs_registers_i.mstack_q[1] ),
    .A2(_09594_),
    .B1(_09586_),
    .B2(_03661_),
    .ZN(_09818_));
 INV_X1 _29020_ (.A(_09818_),
    .ZN(_09819_));
 OAI21_X1 _29021_ (.A(_09809_),
    .B1(_09813_),
    .B2(_09819_),
    .ZN(_09820_));
 OAI21_X1 _29022_ (.A(_09820_),
    .B1(_09816_),
    .B2(_04515_),
    .ZN(_03059_));
 OR2_X1 _29023_ (.A1(_07289_),
    .A2(_09561_),
    .ZN(_09821_));
 AND2_X1 _29024_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_09540_),
    .ZN(_09822_));
 INV_X1 _29025_ (.A(\cs_registers_i.mstack_q[2] ),
    .ZN(_09823_));
 NAND2_X1 _29026_ (.A1(\cs_registers_i.nmi_mode_i ),
    .A2(_09823_),
    .ZN(_09824_));
 AOI221_X2 _29027_ (.A(\cs_registers_i.mstack_d[2] ),
    .B1(_09821_),
    .B2(_09822_),
    .C1(_09824_),
    .C2(_04070_),
    .ZN(_09825_));
 AOI21_X1 _29028_ (.A(_09586_),
    .B1(_09594_),
    .B2(_09823_),
    .ZN(_09826_));
 OR2_X1 _29029_ (.A1(_08666_),
    .A2(_09812_),
    .ZN(_09827_));
 AOI21_X1 _29030_ (.A(_09822_),
    .B1(_09826_),
    .B2(_09827_),
    .ZN(_09828_));
 AOI22_X1 _29031_ (.A1(_09812_),
    .A2(_09825_),
    .B1(_09828_),
    .B2(_09809_),
    .ZN(_03060_));
 AOI21_X1 _29032_ (.A(_09724_),
    .B1(_09346_),
    .B2(\cs_registers_i.mstack_d[2] ),
    .ZN(_09829_));
 NOR2_X1 _29033_ (.A1(_08629_),
    .A2(_09812_),
    .ZN(_09830_));
 AOI21_X1 _29034_ (.A(_09830_),
    .B1(_09812_),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .ZN(_09831_));
 AOI21_X1 _29035_ (.A(_09829_),
    .B1(_09831_),
    .B2(_09562_),
    .ZN(_03061_));
 AOI21_X1 _29036_ (.A(_09576_),
    .B1(_09545_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .ZN(_09832_));
 BUF_X4 _29037_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_09833_));
 BUF_X4 _29038_ (.A(_09833_),
    .Z(_09834_));
 MUX2_X1 _29039_ (.A(_10787_),
    .B(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .S(_09834_),
    .Z(_09835_));
 NOR2_X1 _29040_ (.A1(_09543_),
    .A2(_09835_),
    .ZN(_09836_));
 NOR4_X1 _29041_ (.A1(_09587_),
    .A2(_07835_),
    .A3(_09832_),
    .A4(_09836_),
    .ZN(_09837_));
 MUX2_X1 _29042_ (.A(_08396_),
    .B(_09837_),
    .S(_09650_),
    .Z(_09838_));
 AOI21_X4 _29043_ (.A(_09561_),
    .B1(_08835_),
    .B2(_04570_),
    .ZN(_09839_));
 CLKBUF_X3 _29044_ (.A(_09839_),
    .Z(_09840_));
 MUX2_X1 _29045_ (.A(_09838_),
    .B(\cs_registers_i.mtval_q[0] ),
    .S(_09840_),
    .Z(_03062_));
 CLKBUF_X3 _29046_ (.A(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_09841_));
 NAND3_X1 _29047_ (.A1(_11116_),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(_09841_),
    .ZN(_09842_));
 INV_X1 _29048_ (.A(\cs_registers_i.pc_id_i[6] ),
    .ZN(_09843_));
 NAND3_X1 _29049_ (.A1(_11969_),
    .A2(_12011_),
    .A3(\cs_registers_i.pc_id_i[5] ),
    .ZN(_09844_));
 NOR2_X1 _29050_ (.A1(_09843_),
    .A2(_09844_),
    .ZN(_09845_));
 NAND2_X1 _29051_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_09845_),
    .ZN(_09846_));
 NOR2_X2 _29052_ (.A1(_09842_),
    .A2(_09846_),
    .ZN(_09847_));
 NAND3_X1 _29053_ (.A1(_12218_),
    .A2(_12261_),
    .A3(_09847_),
    .ZN(_09848_));
 XNOR2_X1 _29054_ (.A(_00038_),
    .B(_09848_),
    .ZN(_09849_));
 MUX2_X1 _29055_ (.A(_00036_),
    .B(_00037_),
    .S(_09834_),
    .Z(_09850_));
 NOR2_X1 _29056_ (.A1(_09543_),
    .A2(_09850_),
    .ZN(_09851_));
 AOI21_X1 _29057_ (.A(_09851_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .ZN(_09852_));
 MUX2_X1 _29058_ (.A(_09849_),
    .B(_09852_),
    .S(_09551_),
    .Z(_09853_));
 NAND2_X1 _29059_ (.A1(_04084_),
    .A2(_09539_),
    .ZN(_09854_));
 CLKBUF_X3 _29060_ (.A(_09854_),
    .Z(_09855_));
 OAI22_X1 _29061_ (.A1(_08437_),
    .A2(_09721_),
    .B1(_09853_),
    .B2(_09855_),
    .ZN(_09856_));
 MUX2_X1 _29062_ (.A(_09856_),
    .B(\cs_registers_i.mtval_q[10] ),
    .S(_09840_),
    .Z(_03063_));
 CLKBUF_X3 _29063_ (.A(_09855_),
    .Z(_09857_));
 NAND2_X1 _29064_ (.A1(_09841_),
    .A2(_15938_),
    .ZN(_09858_));
 NOR2_X1 _29065_ (.A1(_09846_),
    .A2(_09858_),
    .ZN(_09859_));
 NAND4_X1 _29066_ (.A1(_12218_),
    .A2(_12261_),
    .A3(\cs_registers_i.pc_id_i[10] ),
    .A4(_09859_),
    .ZN(_09860_));
 XNOR2_X1 _29067_ (.A(_00041_),
    .B(_09860_),
    .ZN(_09861_));
 MUX2_X1 _29068_ (.A(_06878_),
    .B(_00040_),
    .S(_09834_),
    .Z(_09862_));
 NOR2_X1 _29069_ (.A1(_09543_),
    .A2(_09862_),
    .ZN(_09863_));
 AOI21_X1 _29070_ (.A(_09863_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .ZN(_09864_));
 MUX2_X1 _29071_ (.A(_09861_),
    .B(_09864_),
    .S(_09551_),
    .Z(_09865_));
 OAI22_X1 _29072_ (.A1(_04472_),
    .A2(_09721_),
    .B1(_09857_),
    .B2(_09865_),
    .ZN(_09866_));
 MUX2_X1 _29073_ (.A(_09866_),
    .B(\cs_registers_i.mtval_q[11] ),
    .S(_09840_),
    .Z(_03064_));
 AND4_X1 _29074_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_12218_),
    .A3(_12261_),
    .A4(\cs_registers_i.pc_id_i[10] ),
    .ZN(_09867_));
 NAND2_X1 _29075_ (.A1(_09847_),
    .A2(_09867_),
    .ZN(_09868_));
 XNOR2_X1 _29076_ (.A(_00043_),
    .B(_09868_),
    .ZN(_09869_));
 NOR2_X1 _29077_ (.A1(_09551_),
    .A2(_09869_),
    .ZN(_09870_));
 NAND3_X1 _29078_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(_09543_),
    .A3(_09545_),
    .ZN(_09871_));
 MUX2_X1 _29079_ (.A(_00176_),
    .B(_00042_),
    .S(_09834_),
    .Z(_09872_));
 OAI21_X1 _29080_ (.A(_09871_),
    .B1(_09872_),
    .B2(_09543_),
    .ZN(_09873_));
 AOI21_X1 _29081_ (.A(_09870_),
    .B1(_09873_),
    .B2(_09551_),
    .ZN(_09874_));
 OAI22_X1 _29082_ (.A1(_04528_),
    .A2(_09721_),
    .B1(_09857_),
    .B2(_09874_),
    .ZN(_09875_));
 MUX2_X1 _29083_ (.A(_09875_),
    .B(\cs_registers_i.mtval_q[12] ),
    .S(_09840_),
    .Z(_03065_));
 AND3_X1 _29084_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_09859_),
    .A3(_09867_),
    .ZN(_09876_));
 XOR2_X1 _29085_ (.A(_00045_),
    .B(_09876_),
    .Z(_09877_));
 MUX2_X1 _29086_ (.A(_00175_),
    .B(_00044_),
    .S(_09834_),
    .Z(_09878_));
 NOR2_X1 _29087_ (.A1(_09543_),
    .A2(_09878_),
    .ZN(_09879_));
 AOI21_X1 _29088_ (.A(_09879_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .ZN(_09880_));
 MUX2_X1 _29089_ (.A(_09877_),
    .B(_09880_),
    .S(_09551_),
    .Z(_09881_));
 OAI22_X1 _29090_ (.A1(_04562_),
    .A2(_09721_),
    .B1(_09857_),
    .B2(_09881_),
    .ZN(_09882_));
 MUX2_X1 _29091_ (.A(_09882_),
    .B(\cs_registers_i.mtval_q[13] ),
    .S(_09840_),
    .Z(_03066_));
 MUX2_X1 _29092_ (.A(_10917_),
    .B(_00046_),
    .S(_09833_),
    .Z(_09883_));
 NOR2_X1 _29093_ (.A1(_09542_),
    .A2(_09883_),
    .ZN(_09884_));
 AOI21_X1 _29094_ (.A(_09884_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .ZN(_09885_));
 AND4_X1 _29095_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_12512_),
    .A3(_09847_),
    .A4(_09867_),
    .ZN(_09886_));
 XOR2_X1 _29096_ (.A(_00047_),
    .B(_09886_),
    .Z(_09887_));
 MUX2_X1 _29097_ (.A(_09885_),
    .B(_09887_),
    .S(_09587_),
    .Z(_09888_));
 OAI22_X1 _29098_ (.A1(_04597_),
    .A2(_09721_),
    .B1(_09857_),
    .B2(_09888_),
    .ZN(_09889_));
 MUX2_X1 _29099_ (.A(_09889_),
    .B(\cs_registers_i.mtval_q[14] ),
    .S(_09840_),
    .Z(_03067_));
 NAND3_X1 _29100_ (.A1(_12512_),
    .A2(_12618_),
    .A3(_09876_),
    .ZN(_09890_));
 XNOR2_X1 _29101_ (.A(_00049_),
    .B(_09890_),
    .ZN(_09891_));
 MUX2_X1 _29102_ (.A(_00184_),
    .B(_00048_),
    .S(_09834_),
    .Z(_09892_));
 NOR2_X1 _29103_ (.A1(_09543_),
    .A2(_09892_),
    .ZN(_09893_));
 AOI21_X1 _29104_ (.A(_09893_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .ZN(_09894_));
 MUX2_X1 _29105_ (.A(_09891_),
    .B(_09894_),
    .S(_09551_),
    .Z(_09895_));
 OAI22_X1 _29106_ (.A1(_04620_),
    .A2(_09721_),
    .B1(_09857_),
    .B2(_09895_),
    .ZN(_09896_));
 MUX2_X1 _29107_ (.A(_09896_),
    .B(\cs_registers_i.mtval_q[15] ),
    .S(_09840_),
    .Z(_03068_));
 NAND3_X1 _29108_ (.A1(_12618_),
    .A2(\cs_registers_i.pc_id_i[15] ),
    .A3(_09886_),
    .ZN(_09897_));
 XNOR2_X1 _29109_ (.A(_00050_),
    .B(_09897_),
    .ZN(_09898_));
 CLKBUF_X3 _29110_ (.A(_09578_),
    .Z(_09899_));
 NOR2_X4 _29111_ (.A1(_09834_),
    .A2(_09542_),
    .ZN(_09900_));
 CLKBUF_X3 _29112_ (.A(_09900_),
    .Z(_09901_));
 AOI22_X1 _29113_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(_09899_),
    .B1(_09901_),
    .B2(_11081_),
    .ZN(_09902_));
 MUX2_X1 _29114_ (.A(_09898_),
    .B(_09902_),
    .S(_09551_),
    .Z(_09903_));
 OAI22_X1 _29115_ (.A1(_04645_),
    .A2(_09721_),
    .B1(_09857_),
    .B2(_09903_),
    .ZN(_09904_));
 MUX2_X1 _29116_ (.A(_09904_),
    .B(\cs_registers_i.mtval_q[16] ),
    .S(_09840_),
    .Z(_03069_));
 AOI22_X1 _29117_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(_09579_),
    .B1(_09900_),
    .B2(_10989_),
    .ZN(_09905_));
 AND3_X1 _29118_ (.A1(_12618_),
    .A2(\cs_registers_i.pc_id_i[15] ),
    .A3(\cs_registers_i.pc_id_i[16] ),
    .ZN(_09906_));
 NAND3_X2 _29119_ (.A1(_12512_),
    .A2(_09876_),
    .A3(_09906_),
    .ZN(_09907_));
 XNOR2_X1 _29120_ (.A(_00051_),
    .B(_09907_),
    .ZN(_09908_));
 MUX2_X1 _29121_ (.A(_09905_),
    .B(_09908_),
    .S(_09587_),
    .Z(_09909_));
 OAI22_X1 _29122_ (.A1(_04665_),
    .A2(_09721_),
    .B1(_09857_),
    .B2(_09909_),
    .ZN(_09910_));
 CLKBUF_X3 _29123_ (.A(_09839_),
    .Z(_09911_));
 MUX2_X1 _29124_ (.A(_09910_),
    .B(\cs_registers_i.mtval_q[17] ),
    .S(_09911_),
    .Z(_03070_));
 CLKBUF_X3 _29125_ (.A(_09650_),
    .Z(_09912_));
 AND2_X1 _29126_ (.A1(_09886_),
    .A2(_09906_),
    .ZN(_09913_));
 NAND2_X1 _29127_ (.A1(_12868_),
    .A2(_09913_),
    .ZN(_09914_));
 XNOR2_X1 _29128_ (.A(_00052_),
    .B(_09914_),
    .ZN(_09915_));
 AOI22_X1 _29129_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(_09899_),
    .B1(_09901_),
    .B2(_11056_),
    .ZN(_09916_));
 MUX2_X1 _29130_ (.A(_09915_),
    .B(_09916_),
    .S(_09551_),
    .Z(_09917_));
 OAI22_X1 _29131_ (.A1(_04685_),
    .A2(_09912_),
    .B1(_09857_),
    .B2(_09917_),
    .ZN(_09918_));
 MUX2_X1 _29132_ (.A(_09918_),
    .B(\cs_registers_i.mtval_q[18] ),
    .S(_09911_),
    .Z(_03071_));
 NAND2_X1 _29133_ (.A1(_12868_),
    .A2(_12973_),
    .ZN(_09919_));
 NOR2_X1 _29134_ (.A1(_09907_),
    .A2(_09919_),
    .ZN(_09920_));
 XOR2_X1 _29135_ (.A(_00053_),
    .B(_09920_),
    .Z(_09921_));
 AOI22_X1 _29136_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(_09899_),
    .B1(_09901_),
    .B2(_11054_),
    .ZN(_09922_));
 MUX2_X1 _29137_ (.A(_09921_),
    .B(_09922_),
    .S(_09551_),
    .Z(_09923_));
 OAI22_X1 _29138_ (.A1(_04700_),
    .A2(_09912_),
    .B1(_09857_),
    .B2(_09923_),
    .ZN(_09924_));
 MUX2_X1 _29139_ (.A(_09924_),
    .B(\cs_registers_i.mtval_q[19] ),
    .S(_09911_),
    .Z(_03072_));
 MUX2_X1 _29140_ (.A(_00013_),
    .B(_00014_),
    .S(_09833_),
    .Z(_09925_));
 NOR2_X1 _29141_ (.A1(_09542_),
    .A2(_09925_),
    .ZN(_09926_));
 AOI21_X1 _29142_ (.A(_09926_),
    .B1(_09899_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .ZN(_09927_));
 XNOR2_X1 _29143_ (.A(_11116_),
    .B(_09841_),
    .ZN(_09928_));
 MUX2_X1 _29144_ (.A(_09927_),
    .B(_09928_),
    .S(_09587_),
    .Z(_09929_));
 OAI22_X1 _29145_ (.A1(_08519_),
    .A2(_09912_),
    .B1(_09857_),
    .B2(_09929_),
    .ZN(_09930_));
 MUX2_X1 _29146_ (.A(_09930_),
    .B(\cs_registers_i.mtval_q[1] ),
    .S(_09911_),
    .Z(_03073_));
 BUF_X4 _29147_ (.A(_09854_),
    .Z(_09931_));
 NAND4_X1 _29148_ (.A1(_12868_),
    .A2(_12973_),
    .A3(\cs_registers_i.pc_id_i[19] ),
    .A4(_09913_),
    .ZN(_09932_));
 XNOR2_X1 _29149_ (.A(_00054_),
    .B(_09932_),
    .ZN(_09933_));
 AOI22_X1 _29150_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(_09899_),
    .B1(_09901_),
    .B2(_12426_),
    .ZN(_09934_));
 CLKBUF_X3 _29151_ (.A(_04020_),
    .Z(_09935_));
 MUX2_X1 _29152_ (.A(_09933_),
    .B(_09934_),
    .S(_09935_),
    .Z(_09936_));
 OAI22_X1 _29153_ (.A1(_04721_),
    .A2(_09912_),
    .B1(_09931_),
    .B2(_09936_),
    .ZN(_09937_));
 MUX2_X1 _29154_ (.A(_09937_),
    .B(\cs_registers_i.mtval_q[20] ),
    .S(_09911_),
    .Z(_03074_));
 AND4_X1 _29155_ (.A1(_12868_),
    .A2(_12973_),
    .A3(\cs_registers_i.pc_id_i[19] ),
    .A4(\cs_registers_i.pc_id_i[20] ),
    .ZN(_09938_));
 NAND4_X1 _29156_ (.A1(_12512_),
    .A2(_09876_),
    .A3(_09906_),
    .A4(_09938_),
    .ZN(_09939_));
 XNOR2_X1 _29157_ (.A(_00055_),
    .B(_09939_),
    .ZN(_09940_));
 AOI22_X1 _29158_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(_09899_),
    .B1(_09901_),
    .B2(_12438_),
    .ZN(_09941_));
 MUX2_X1 _29159_ (.A(_09940_),
    .B(_09941_),
    .S(_09935_),
    .Z(_09942_));
 OAI22_X1 _29160_ (.A1(_04742_),
    .A2(_09912_),
    .B1(_09931_),
    .B2(_09942_),
    .ZN(_09943_));
 MUX2_X1 _29161_ (.A(_09943_),
    .B(\cs_registers_i.mtval_q[21] ),
    .S(_09911_),
    .Z(_03075_));
 AOI22_X1 _29162_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(_09579_),
    .B1(_09900_),
    .B2(_12424_),
    .ZN(_09944_));
 AND3_X1 _29163_ (.A1(_13237_),
    .A2(_09913_),
    .A3(_09938_),
    .ZN(_09945_));
 XOR2_X1 _29164_ (.A(_00056_),
    .B(_09945_),
    .Z(_09946_));
 MUX2_X1 _29165_ (.A(_09944_),
    .B(_09946_),
    .S(_09587_),
    .Z(_09947_));
 OAI22_X1 _29166_ (.A1(_04762_),
    .A2(_09912_),
    .B1(_09931_),
    .B2(_09947_),
    .ZN(_09948_));
 MUX2_X1 _29167_ (.A(_09948_),
    .B(\cs_registers_i.mtval_q[22] ),
    .S(_09911_),
    .Z(_03076_));
 NAND2_X1 _29168_ (.A1(_13237_),
    .A2(_09938_),
    .ZN(_09949_));
 NOR2_X1 _29169_ (.A1(_09907_),
    .A2(_09949_),
    .ZN(_09950_));
 NAND2_X1 _29170_ (.A1(_13347_),
    .A2(_09950_),
    .ZN(_09951_));
 XNOR2_X1 _29171_ (.A(_00057_),
    .B(_09951_),
    .ZN(_09952_));
 AOI22_X1 _29172_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(_09899_),
    .B1(_09901_),
    .B2(_12432_),
    .ZN(_09953_));
 MUX2_X1 _29173_ (.A(_09952_),
    .B(_09953_),
    .S(_09935_),
    .Z(_09954_));
 OAI22_X1 _29174_ (.A1(_04783_),
    .A2(_09912_),
    .B1(_09931_),
    .B2(_09954_),
    .ZN(_09955_));
 MUX2_X1 _29175_ (.A(_09955_),
    .B(\cs_registers_i.mtval_q[23] ),
    .S(_09911_),
    .Z(_03077_));
 NAND3_X1 _29176_ (.A1(_13347_),
    .A2(_13423_),
    .A3(_09945_),
    .ZN(_09956_));
 XNOR2_X1 _29177_ (.A(_00058_),
    .B(_09956_),
    .ZN(_09957_));
 AOI22_X1 _29178_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(_09899_),
    .B1(_09901_),
    .B2(_12419_),
    .ZN(_09958_));
 MUX2_X1 _29179_ (.A(_09957_),
    .B(_09958_),
    .S(_09935_),
    .Z(_09959_));
 OAI22_X1 _29180_ (.A1(_04805_),
    .A2(_09912_),
    .B1(_09931_),
    .B2(_09959_),
    .ZN(_09960_));
 MUX2_X1 _29181_ (.A(_09960_),
    .B(\cs_registers_i.mtval_q[24] ),
    .S(_09911_),
    .Z(_03078_));
 NAND4_X1 _29182_ (.A1(_13347_),
    .A2(_13423_),
    .A3(\cs_registers_i.pc_id_i[24] ),
    .A4(_09950_),
    .ZN(_09961_));
 XNOR2_X1 _29183_ (.A(_00059_),
    .B(_09961_),
    .ZN(_09962_));
 AOI22_X1 _29184_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(_09579_),
    .B1(_09901_),
    .B2(_10945_),
    .ZN(_09963_));
 MUX2_X1 _29185_ (.A(_09962_),
    .B(_09963_),
    .S(_09935_),
    .Z(_09964_));
 OAI22_X1 _29186_ (.A1(_04822_),
    .A2(_09912_),
    .B1(_09931_),
    .B2(_09964_),
    .ZN(_09965_));
 MUX2_X1 _29187_ (.A(_09965_),
    .B(\cs_registers_i.mtval_q[25] ),
    .S(_09911_),
    .Z(_03079_));
 AOI22_X1 _29188_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(_09579_),
    .B1(_09900_),
    .B2(_10869_),
    .ZN(_09966_));
 AND4_X1 _29189_ (.A1(_13347_),
    .A2(_13423_),
    .A3(\cs_registers_i.pc_id_i[24] ),
    .A4(\cs_registers_i.pc_id_i[25] ),
    .ZN(_09967_));
 NAND2_X1 _29190_ (.A1(_09945_),
    .A2(_09967_),
    .ZN(_09968_));
 XNOR2_X1 _29191_ (.A(_00060_),
    .B(_09968_),
    .ZN(_09969_));
 MUX2_X1 _29192_ (.A(_09966_),
    .B(_09969_),
    .S(_09587_),
    .Z(_09970_));
 OAI22_X2 _29193_ (.A1(_04838_),
    .A2(_09912_),
    .B1(_09931_),
    .B2(_09970_),
    .ZN(_09971_));
 BUF_X4 _29194_ (.A(_09839_),
    .Z(_09972_));
 MUX2_X1 _29195_ (.A(_09971_),
    .B(\cs_registers_i.mtval_q[26] ),
    .S(_09972_),
    .Z(_03080_));
 BUF_X4 _29196_ (.A(_09650_),
    .Z(_09973_));
 NAND2_X1 _29197_ (.A1(_09950_),
    .A2(_09967_),
    .ZN(_09974_));
 INV_X1 _29198_ (.A(_09974_),
    .ZN(_09975_));
 NAND2_X1 _29199_ (.A1(_13688_),
    .A2(_09975_),
    .ZN(_09976_));
 XNOR2_X1 _29200_ (.A(_00061_),
    .B(_09976_),
    .ZN(_09977_));
 AOI22_X1 _29201_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(_09579_),
    .B1(_09901_),
    .B2(_10873_),
    .ZN(_09978_));
 MUX2_X1 _29202_ (.A(_09977_),
    .B(_09978_),
    .S(_09935_),
    .Z(_09979_));
 OAI22_X2 _29203_ (.A1(_04853_),
    .A2(_09973_),
    .B1(_09931_),
    .B2(_09979_),
    .ZN(_09980_));
 MUX2_X1 _29204_ (.A(_09980_),
    .B(\cs_registers_i.mtval_q[27] ),
    .S(_09972_),
    .Z(_03081_));
 NAND4_X1 _29205_ (.A1(_13688_),
    .A2(_03142_),
    .A3(_09945_),
    .A4(_09967_),
    .ZN(_09981_));
 XNOR2_X1 _29206_ (.A(_00062_),
    .B(_09981_),
    .ZN(_09982_));
 AOI22_X1 _29207_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(_09579_),
    .B1(_09901_),
    .B2(_10876_),
    .ZN(_09983_));
 MUX2_X1 _29208_ (.A(_09982_),
    .B(_09983_),
    .S(_09935_),
    .Z(_09984_));
 OAI22_X2 _29209_ (.A1(_04868_),
    .A2(_09973_),
    .B1(_09931_),
    .B2(_09984_),
    .ZN(_09985_));
 MUX2_X1 _29210_ (.A(_09985_),
    .B(\cs_registers_i.mtval_q[28] ),
    .S(_09972_),
    .Z(_03082_));
 NAND4_X1 _29211_ (.A1(_13688_),
    .A2(_03142_),
    .A3(_03238_),
    .A4(_09975_),
    .ZN(_09986_));
 XNOR2_X1 _29212_ (.A(_00063_),
    .B(_09986_),
    .ZN(_09987_));
 AOI22_X1 _29213_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(_09579_),
    .B1(_09900_),
    .B2(_10875_),
    .ZN(_09988_));
 MUX2_X1 _29214_ (.A(_09987_),
    .B(_09988_),
    .S(_09935_),
    .Z(_09989_));
 OAI22_X1 _29215_ (.A1(_04885_),
    .A2(_09973_),
    .B1(_09931_),
    .B2(_09989_),
    .ZN(_09990_));
 MUX2_X1 _29216_ (.A(_09990_),
    .B(\cs_registers_i.mtval_q[29] ),
    .S(_09972_),
    .Z(_03083_));
 INV_X1 _29217_ (.A(_09854_),
    .ZN(_09991_));
 MUX2_X1 _29218_ (.A(_00015_),
    .B(_00016_),
    .S(_09833_),
    .Z(_09992_));
 NOR2_X1 _29219_ (.A1(_09542_),
    .A2(_09992_),
    .ZN(_09993_));
 AOI221_X2 _29220_ (.A(_09993_),
    .B1(_09578_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .C1(_10794_),
    .C2(_03647_),
    .ZN(_09994_));
 NOR2_X1 _29221_ (.A1(_00012_),
    .A2(_09841_),
    .ZN(_09995_));
 AOI21_X1 _29222_ (.A(_09995_),
    .B1(_15939_),
    .B2(_09841_),
    .ZN(_09996_));
 AOI21_X1 _29223_ (.A(_09994_),
    .B1(_09996_),
    .B2(_09587_),
    .ZN(_09997_));
 AOI221_X1 _29224_ (.A(_09839_),
    .B1(_09991_),
    .B2(_09997_),
    .C1(_09557_),
    .C2(_08402_),
    .ZN(_09998_));
 INV_X1 _29225_ (.A(\cs_registers_i.mtval_q[2] ),
    .ZN(_09999_));
 AOI21_X1 _29226_ (.A(_09998_),
    .B1(_09840_),
    .B2(_09999_),
    .ZN(_03084_));
 NAND4_X1 _29227_ (.A1(_13688_),
    .A2(_03142_),
    .A3(_03238_),
    .A4(\cs_registers_i.pc_id_i[29] ),
    .ZN(_10000_));
 NOR2_X1 _29228_ (.A1(_09968_),
    .A2(_10000_),
    .ZN(_10001_));
 XOR2_X1 _29229_ (.A(_00064_),
    .B(_10001_),
    .Z(_10002_));
 AOI22_X2 _29230_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(_09579_),
    .B1(_09900_),
    .B2(_10884_),
    .ZN(_10003_));
 MUX2_X1 _29231_ (.A(_10002_),
    .B(_10003_),
    .S(_09935_),
    .Z(_10004_));
 OAI22_X2 _29232_ (.A1(_04905_),
    .A2(_09973_),
    .B1(_09855_),
    .B2(_10004_),
    .ZN(_10005_));
 MUX2_X1 _29233_ (.A(_10005_),
    .B(\cs_registers_i.mtval_q[30] ),
    .S(_09972_),
    .Z(_03085_));
 INV_X1 _29234_ (.A(\cs_registers_i.pc_id_i[30] ),
    .ZN(_10006_));
 NOR3_X1 _29235_ (.A1(_10006_),
    .A2(_09974_),
    .A3(_10000_),
    .ZN(_10007_));
 XOR2_X1 _29236_ (.A(_00065_),
    .B(_10007_),
    .Z(_10008_));
 AOI22_X1 _29237_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(_09579_),
    .B1(_09900_),
    .B2(_10878_),
    .ZN(_10009_));
 MUX2_X1 _29238_ (.A(_10008_),
    .B(_10009_),
    .S(_09935_),
    .Z(_10010_));
 OAI22_X1 _29239_ (.A1(_04924_),
    .A2(_09973_),
    .B1(_09855_),
    .B2(_10010_),
    .ZN(_10011_));
 MUX2_X1 _29240_ (.A(_10011_),
    .B(\cs_registers_i.mtval_q[31] ),
    .S(_09972_),
    .Z(_03086_));
 MUX2_X1 _29241_ (.A(_00017_),
    .B(_00018_),
    .S(_09833_),
    .Z(_10012_));
 NOR2_X1 _29242_ (.A1(_09542_),
    .A2(_10012_),
    .ZN(_10013_));
 AOI21_X1 _29243_ (.A(_10013_),
    .B1(_09899_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .ZN(_10014_));
 XNOR2_X1 _29244_ (.A(_00019_),
    .B(_09858_),
    .ZN(_10015_));
 MUX2_X1 _29245_ (.A(_10014_),
    .B(_10015_),
    .S(_09587_),
    .Z(_10016_));
 OAI22_X1 _29246_ (.A1(_08629_),
    .A2(_09973_),
    .B1(_09855_),
    .B2(_10016_),
    .ZN(_10017_));
 MUX2_X1 _29247_ (.A(_10017_),
    .B(\cs_registers_i.mtval_q[3] ),
    .S(_09972_),
    .Z(_03087_));
 NAND4_X1 _29248_ (.A1(_11116_),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(_11969_),
    .A4(_09841_),
    .ZN(_10018_));
 XNOR2_X1 _29249_ (.A(_00022_),
    .B(_10018_),
    .ZN(_10019_));
 MUX2_X1 _29250_ (.A(_00020_),
    .B(_00021_),
    .S(_09834_),
    .Z(_10020_));
 NOR2_X1 _29251_ (.A1(_09543_),
    .A2(_10020_),
    .ZN(_10021_));
 AOI21_X1 _29252_ (.A(_10021_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .ZN(_10022_));
 MUX2_X1 _29253_ (.A(_10019_),
    .B(_10022_),
    .S(_04020_),
    .Z(_10023_));
 OAI22_X2 _29254_ (.A1(_08639_),
    .A2(_09973_),
    .B1(_09855_),
    .B2(_10023_),
    .ZN(_10024_));
 MUX2_X1 _29255_ (.A(_10024_),
    .B(\cs_registers_i.mtval_q[4] ),
    .S(_09972_),
    .Z(_03088_));
 NAND4_X1 _29256_ (.A1(_11969_),
    .A2(_12011_),
    .A3(_09841_),
    .A4(_15938_),
    .ZN(_10025_));
 XNOR2_X1 _29257_ (.A(_00025_),
    .B(_10025_),
    .ZN(_10026_));
 MUX2_X1 _29258_ (.A(_00023_),
    .B(_00024_),
    .S(_09834_),
    .Z(_10027_));
 NOR2_X1 _29259_ (.A1(_09542_),
    .A2(_10027_),
    .ZN(_10028_));
 AOI21_X1 _29260_ (.A(_10028_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .ZN(_10029_));
 MUX2_X1 _29261_ (.A(_10026_),
    .B(_10029_),
    .S(_04020_),
    .Z(_10030_));
 OAI22_X2 _29262_ (.A1(_08646_),
    .A2(_09973_),
    .B1(_09855_),
    .B2(_10030_),
    .ZN(_10031_));
 MUX2_X1 _29263_ (.A(_10031_),
    .B(\cs_registers_i.mtval_q[5] ),
    .S(_09972_),
    .Z(_03089_));
 NOR2_X1 _29264_ (.A1(_09842_),
    .A2(_09844_),
    .ZN(_10032_));
 XOR2_X1 _29265_ (.A(_00027_),
    .B(_10032_),
    .Z(_10033_));
 MUX2_X1 _29266_ (.A(_00172_),
    .B(_00026_),
    .S(_09833_),
    .Z(_10034_));
 NOR2_X1 _29267_ (.A1(_09542_),
    .A2(_10034_),
    .ZN(_10035_));
 AOI21_X1 _29268_ (.A(_10035_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .ZN(_10036_));
 MUX2_X1 _29269_ (.A(_10033_),
    .B(_10036_),
    .S(_04020_),
    .Z(_10037_));
 OAI22_X1 _29270_ (.A1(_08655_),
    .A2(_09973_),
    .B1(_09855_),
    .B2(_10037_),
    .ZN(_10038_));
 MUX2_X1 _29271_ (.A(_10038_),
    .B(\cs_registers_i.mtval_q[6] ),
    .S(_09972_),
    .Z(_03090_));
 INV_X1 _29272_ (.A(_00028_),
    .ZN(_10039_));
 NAND2_X1 _29273_ (.A1(_09833_),
    .A2(_10039_),
    .ZN(_10040_));
 OAI21_X2 _29274_ (.A(_10040_),
    .B1(_00216_),
    .B2(_09833_),
    .ZN(_10041_));
 AOI221_X2 _29275_ (.A(_04011_),
    .B1(_09578_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .C1(_10041_),
    .C2(_09576_),
    .ZN(_10042_));
 NAND3_X1 _29276_ (.A1(_09841_),
    .A2(_15938_),
    .A3(_09845_),
    .ZN(_10043_));
 XNOR2_X1 _29277_ (.A(_00029_),
    .B(_10043_),
    .ZN(_10044_));
 AOI21_X1 _29278_ (.A(_10042_),
    .B1(_10044_),
    .B2(_04011_),
    .ZN(_10045_));
 AOI221_X1 _29279_ (.A(_09839_),
    .B1(_09991_),
    .B2(_10045_),
    .C1(_09557_),
    .C2(_08665_),
    .ZN(_10046_));
 INV_X1 _29280_ (.A(\cs_registers_i.mtval_q[7] ),
    .ZN(_10047_));
 AOI21_X1 _29281_ (.A(_10046_),
    .B1(_09840_),
    .B2(_10047_),
    .ZN(_03091_));
 MUX2_X1 _29282_ (.A(_00030_),
    .B(_00031_),
    .S(_09833_),
    .Z(_10048_));
 NOR2_X1 _29283_ (.A1(_09542_),
    .A2(_10048_),
    .ZN(_10049_));
 AOI21_X1 _29284_ (.A(_10049_),
    .B1(_09899_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .ZN(_10050_));
 XOR2_X1 _29285_ (.A(_00032_),
    .B(_09847_),
    .Z(_10051_));
 MUX2_X1 _29286_ (.A(_10050_),
    .B(_10051_),
    .S(_09587_),
    .Z(_10052_));
 OAI22_X1 _29287_ (.A1(_04942_),
    .A2(_09973_),
    .B1(_09855_),
    .B2(_10052_),
    .ZN(_10053_));
 MUX2_X1 _29288_ (.A(_10053_),
    .B(\cs_registers_i.mtval_q[8] ),
    .S(_09839_),
    .Z(_03092_));
 NAND2_X1 _29289_ (.A1(_12218_),
    .A2(_09859_),
    .ZN(_10054_));
 XNOR2_X1 _29290_ (.A(_00035_),
    .B(_10054_),
    .ZN(_10055_));
 MUX2_X1 _29291_ (.A(_00033_),
    .B(_00034_),
    .S(_09833_),
    .Z(_10056_));
 NOR2_X1 _29292_ (.A1(_09542_),
    .A2(_10056_),
    .ZN(_10057_));
 AOI21_X1 _29293_ (.A(_10057_),
    .B1(_09580_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .ZN(_10058_));
 MUX2_X1 _29294_ (.A(_10055_),
    .B(_10058_),
    .S(_04020_),
    .Z(_10059_));
 OAI22_X1 _29295_ (.A1(_04960_),
    .A2(_09586_),
    .B1(_09855_),
    .B2(_10059_),
    .ZN(_10060_));
 MUX2_X1 _29296_ (.A(_10060_),
    .B(\cs_registers_i.mtval_q[9] ),
    .S(_09839_),
    .Z(_03093_));
 NAND2_X1 _29297_ (.A1(net1),
    .A2(_04370_),
    .ZN(_10061_));
 INV_X1 _29298_ (.A(\cs_registers_i.csr_mtvec_o[10] ),
    .ZN(_10062_));
 OAI221_X1 _29299_ (.A(_10061_),
    .B1(_08437_),
    .B2(_04491_),
    .C1(_10062_),
    .C2(_04493_),
    .ZN(_03094_));
 CLKBUF_X3 _29300_ (.A(_08076_),
    .Z(_10063_));
 NAND2_X1 _29301_ (.A1(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .A2(_10063_),
    .ZN(_10064_));
 MUX2_X1 _29302_ (.A(net94),
    .B(_04110_),
    .S(_04105_),
    .Z(_10065_));
 MUX2_X1 _29303_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .S(_04105_),
    .Z(_10066_));
 MUX2_X1 _29304_ (.A(_10065_),
    .B(_10066_),
    .S(_04120_),
    .Z(_10067_));
 BUF_X4 _29305_ (.A(_10067_),
    .Z(_10068_));
 MUX2_X1 _29306_ (.A(net103),
    .B(_04109_),
    .S(_04105_),
    .Z(_10069_));
 MUX2_X1 _29307_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(_04105_),
    .Z(_10070_));
 MUX2_X1 _29308_ (.A(_10069_),
    .B(_10070_),
    .S(_04120_),
    .Z(_10071_));
 BUF_X4 _29309_ (.A(_10071_),
    .Z(_10072_));
 NOR2_X4 _29310_ (.A1(_10068_),
    .A2(_10072_),
    .ZN(_10073_));
 MUX2_X1 _29311_ (.A(net99),
    .B(net115),
    .S(_04103_),
    .Z(_10074_));
 MUX2_X1 _29312_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .S(_04103_),
    .Z(_10075_));
 MUX2_X2 _29313_ (.A(_10074_),
    .B(_10075_),
    .S(_04106_),
    .Z(_10076_));
 BUF_X4 _29314_ (.A(_10076_),
    .Z(_10077_));
 BUF_X4 _29315_ (.A(_04103_),
    .Z(_10078_));
 MUX2_X1 _29316_ (.A(net98),
    .B(net113),
    .S(_10078_),
    .Z(_10079_));
 OR2_X1 _29317_ (.A1(_04119_),
    .A2(_10079_),
    .ZN(_10080_));
 MUX2_X1 _29318_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(_10078_),
    .Z(_10081_));
 OAI21_X2 _29319_ (.A(_10080_),
    .B1(_10081_),
    .B2(_04107_),
    .ZN(_10082_));
 BUF_X4 _29320_ (.A(_10082_),
    .Z(_10083_));
 NAND2_X4 _29321_ (.A1(_10077_),
    .A2(_10083_),
    .ZN(_10084_));
 NAND2_X2 _29322_ (.A1(_10073_),
    .A2(_10084_),
    .ZN(_10085_));
 MUX2_X1 _29323_ (.A(net95),
    .B(net110),
    .S(_10078_),
    .Z(_10086_));
 MUX2_X2 _29324_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(_04103_),
    .Z(_10087_));
 MUX2_X2 _29325_ (.A(_10086_),
    .B(_10087_),
    .S(_04106_),
    .Z(_10088_));
 MUX2_X1 _29326_ (.A(net96),
    .B(net111),
    .S(_04103_),
    .Z(_10089_));
 MUX2_X1 _29327_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(_04103_),
    .Z(_10090_));
 MUX2_X2 _29328_ (.A(_10089_),
    .B(_10090_),
    .S(_04106_),
    .Z(_10091_));
 MUX2_X1 _29329_ (.A(net123),
    .B(net109),
    .S(_04103_),
    .Z(_10092_));
 MUX2_X1 _29330_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(_04103_),
    .Z(_10093_));
 MUX2_X2 _29331_ (.A(_10092_),
    .B(_10093_),
    .S(_04106_),
    .Z(_10094_));
 MUX2_X1 _29332_ (.A(net121),
    .B(net107),
    .S(\cs_registers_i.pc_if_i[1] ),
    .Z(_10095_));
 MUX2_X1 _29333_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(\cs_registers_i.pc_if_i[1] ),
    .Z(_10096_));
 MUX2_X1 _29334_ (.A(_10095_),
    .B(_10096_),
    .S(_04106_),
    .Z(_10097_));
 BUF_X4 _29335_ (.A(_10097_),
    .Z(_10098_));
 NOR4_X4 _29336_ (.A1(_10088_),
    .A2(_10091_),
    .A3(_10094_),
    .A4(_10098_),
    .ZN(_10099_));
 MUX2_X1 _29337_ (.A(net122),
    .B(net108),
    .S(_04104_),
    .Z(_10100_));
 MUX2_X1 _29338_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(_04104_),
    .Z(_10101_));
 MUX2_X1 _29339_ (.A(_10100_),
    .B(_10101_),
    .S(_04119_),
    .Z(_10102_));
 BUF_X4 _29340_ (.A(_10102_),
    .Z(_10103_));
 INV_X1 _29341_ (.A(_10103_),
    .ZN(_10104_));
 MUX2_X1 _29342_ (.A(net97),
    .B(net112),
    .S(_04104_),
    .Z(_10105_));
 OR2_X1 _29343_ (.A1(_04119_),
    .A2(_10105_),
    .ZN(_10106_));
 MUX2_X2 _29344_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(_04104_),
    .Z(_10107_));
 OAI21_X4 _29345_ (.A(_10106_),
    .B1(_10107_),
    .B2(_04107_),
    .ZN(_10108_));
 BUF_X4 _29346_ (.A(_10108_),
    .Z(_10109_));
 BUF_X4 _29347_ (.A(_10109_),
    .Z(_10110_));
 MUX2_X1 _29348_ (.A(net119),
    .B(net105),
    .S(_10078_),
    .Z(_10111_));
 MUX2_X1 _29349_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(_10078_),
    .Z(_10112_));
 MUX2_X1 _29350_ (.A(_10111_),
    .B(_10112_),
    .S(_04119_),
    .Z(_10113_));
 BUF_X4 _29351_ (.A(_10113_),
    .Z(_10114_));
 NAND2_X1 _29352_ (.A1(_04104_),
    .A2(net106),
    .ZN(_10115_));
 NAND2_X1 _29353_ (.A1(_08073_),
    .A2(net120),
    .ZN(_10116_));
 NAND3_X1 _29354_ (.A1(_04107_),
    .A2(_10115_),
    .A3(_10116_),
    .ZN(_10117_));
 MUX2_X1 _29355_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(_04104_),
    .Z(_10118_));
 OAI21_X2 _29356_ (.A(_10117_),
    .B1(_10118_),
    .B2(_04107_),
    .ZN(_10119_));
 INV_X1 _29357_ (.A(_10119_),
    .ZN(_10120_));
 NOR2_X4 _29358_ (.A1(_10114_),
    .A2(_10120_),
    .ZN(_10121_));
 NAND4_X1 _29359_ (.A1(_10099_),
    .A2(_10104_),
    .A3(_10110_),
    .A4(_10121_),
    .ZN(_10122_));
 MUX2_X1 _29360_ (.A(net100),
    .B(net116),
    .S(_04103_),
    .Z(_10123_));
 MUX2_X1 _29361_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(_10078_),
    .Z(_10124_));
 MUX2_X2 _29362_ (.A(_10123_),
    .B(_10124_),
    .S(_04106_),
    .Z(_10125_));
 MUX2_X1 _29363_ (.A(_10079_),
    .B(_10081_),
    .S(_04119_),
    .Z(_10126_));
 BUF_X4 _29364_ (.A(_10126_),
    .Z(_10127_));
 NOR2_X2 _29365_ (.A1(_10125_),
    .A2(_10127_),
    .ZN(_10128_));
 CLKBUF_X3 _29366_ (.A(_10128_),
    .Z(_10129_));
 AOI21_X1 _29367_ (.A(_10085_),
    .B1(_10122_),
    .B2(_10129_),
    .ZN(_10130_));
 MUX2_X1 _29368_ (.A(net114),
    .B(net101),
    .S(_04104_),
    .Z(_10131_));
 MUX2_X1 _29369_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(_04104_),
    .Z(_10132_));
 MUX2_X2 _29370_ (.A(_10131_),
    .B(_10132_),
    .S(_04119_),
    .Z(_10133_));
 MUX2_X1 _29371_ (.A(net118),
    .B(net104),
    .S(_10078_),
    .Z(_10134_));
 MUX2_X2 _29372_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(_10078_),
    .Z(_10135_));
 MUX2_X2 _29373_ (.A(_10134_),
    .B(_10135_),
    .S(_04119_),
    .Z(_10136_));
 MUX2_X1 _29374_ (.A(net117),
    .B(net102),
    .S(_10078_),
    .Z(_10137_));
 MUX2_X1 _29375_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S(_10078_),
    .Z(_10138_));
 MUX2_X2 _29376_ (.A(_10137_),
    .B(_10138_),
    .S(_04119_),
    .Z(_10139_));
 NOR3_X4 _29377_ (.A1(_10133_),
    .A2(_10136_),
    .A3(_10139_),
    .ZN(_10140_));
 NAND3_X1 _29378_ (.A1(_10109_),
    .A2(_10121_),
    .A3(_10140_),
    .ZN(_10141_));
 BUF_X4 _29379_ (.A(_10083_),
    .Z(_10142_));
 CLKBUF_X3 _29380_ (.A(_10142_),
    .Z(_10143_));
 OR2_X1 _29381_ (.A1(_04119_),
    .A2(_10123_),
    .ZN(_10144_));
 OAI21_X4 _29382_ (.A(_10144_),
    .B1(_10124_),
    .B2(_04107_),
    .ZN(_10145_));
 NAND2_X4 _29383_ (.A1(_10145_),
    .A2(_10077_),
    .ZN(_10146_));
 NOR2_X4 _29384_ (.A1(_10145_),
    .A2(_10076_),
    .ZN(_10147_));
 NAND2_X4 _29385_ (.A1(_10083_),
    .A2(_10147_),
    .ZN(_10148_));
 CLKBUF_X3 _29386_ (.A(_10088_),
    .Z(_10149_));
 OR2_X1 _29387_ (.A1(_04120_),
    .A2(_10089_),
    .ZN(_10150_));
 OAI21_X4 _29388_ (.A(_10150_),
    .B1(_10090_),
    .B2(_04107_),
    .ZN(_10151_));
 NOR2_X1 _29389_ (.A1(_10149_),
    .A2(_10151_),
    .ZN(_10152_));
 OAI33_X1 _29390_ (.A1(_10141_),
    .A2(_10143_),
    .A3(_10146_),
    .B1(_10148_),
    .B2(_10152_),
    .B3(_10110_),
    .ZN(_10153_));
 OR2_X1 _29391_ (.A1(_04120_),
    .A2(_10065_),
    .ZN(_10154_));
 OAI21_X4 _29392_ (.A(_10154_),
    .B1(_10066_),
    .B2(_08033_),
    .ZN(_10155_));
 NOR2_X4 _29393_ (.A1(_10155_),
    .A2(_10072_),
    .ZN(_10156_));
 CLKBUF_X3 _29394_ (.A(_10077_),
    .Z(_10157_));
 CLKBUF_X3 _29395_ (.A(_10157_),
    .Z(_10158_));
 BUF_X4 _29396_ (.A(_10125_),
    .Z(_10159_));
 NAND2_X1 _29397_ (.A1(_10099_),
    .A2(_10104_),
    .ZN(_10160_));
 CLKBUF_X3 _29398_ (.A(_10145_),
    .Z(_10161_));
 BUF_X4 _29399_ (.A(_10161_),
    .Z(_10162_));
 NOR2_X1 _29400_ (.A1(_10141_),
    .A2(_10158_),
    .ZN(_10163_));
 NOR2_X1 _29401_ (.A1(_10162_),
    .A2(_10163_),
    .ZN(_10164_));
 OAI221_X2 _29402_ (.A(_10143_),
    .B1(_10158_),
    .B2(_10159_),
    .C1(_10160_),
    .C2(_10164_),
    .ZN(_10165_));
 NAND2_X1 _29403_ (.A1(_10155_),
    .A2(_10071_),
    .ZN(_10166_));
 CLKBUF_X3 _29404_ (.A(_10166_),
    .Z(_10167_));
 NAND2_X1 _29405_ (.A1(_10161_),
    .A2(_10083_),
    .ZN(_10168_));
 NOR2_X2 _29406_ (.A1(_10077_),
    .A2(_10168_),
    .ZN(_10169_));
 BUF_X4 _29407_ (.A(_10169_),
    .Z(_10170_));
 BUF_X4 _29408_ (.A(_10110_),
    .Z(_10171_));
 AOI21_X1 _29409_ (.A(_10167_),
    .B1(_10170_),
    .B2(_10171_),
    .ZN(_10172_));
 AOI221_X2 _29410_ (.A(_10130_),
    .B1(_10153_),
    .B2(_10156_),
    .C1(_10165_),
    .C2(_10172_),
    .ZN(_10173_));
 BUF_X4 _29411_ (.A(_08076_),
    .Z(_10174_));
 OAI21_X1 _29412_ (.A(_10064_),
    .B1(_10173_),
    .B2(_10174_),
    .ZN(_02535_));
 NAND2_X1 _29413_ (.A1(_03647_),
    .A2(_10063_),
    .ZN(_10175_));
 INV_X1 _29414_ (.A(_04108_),
    .ZN(_10176_));
 NOR3_X1 _29415_ (.A1(_08040_),
    .A2(_04123_),
    .A3(_10176_),
    .ZN(_10177_));
 OAI21_X1 _29416_ (.A(_04108_),
    .B1(_00136_),
    .B2(_04115_),
    .ZN(_10178_));
 OR2_X1 _29417_ (.A1(_04308_),
    .A2(_10178_),
    .ZN(_10179_));
 AOI21_X1 _29418_ (.A(_04113_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B2(_04115_),
    .ZN(_10180_));
 OAI21_X1 _29419_ (.A(_10179_),
    .B1(_10180_),
    .B2(_08061_),
    .ZN(_10181_));
 AOI221_X2 _29420_ (.A(_10177_),
    .B1(_10181_),
    .B2(_04123_),
    .C1(_08040_),
    .C2(_04113_),
    .ZN(_10182_));
 OAI21_X1 _29421_ (.A(_10175_),
    .B1(_10182_),
    .B2(_10174_),
    .ZN(_02536_));
 NOR3_X1 _29422_ (.A1(_08033_),
    .A2(_08029_),
    .A3(_10176_),
    .ZN(_10183_));
 AOI21_X1 _29423_ (.A(_10183_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B2(_08029_),
    .ZN(_10184_));
 NOR3_X1 _29424_ (.A1(_08074_),
    .A2(_04113_),
    .A3(_10184_),
    .ZN(_10185_));
 BUF_X4 _29425_ (.A(_08153_),
    .Z(_10186_));
 MUX2_X1 _29426_ (.A(_09841_),
    .B(_10185_),
    .S(_10186_),
    .Z(_02537_));
 NAND2_X4 _29427_ (.A1(_10068_),
    .A2(_10072_),
    .ZN(_10187_));
 MUX2_X1 _29428_ (.A(_09834_),
    .B(_10187_),
    .S(_10186_),
    .Z(_02538_));
 BUF_X4 _29429_ (.A(_10155_),
    .Z(_10188_));
 OR2_X1 _29430_ (.A1(_04106_),
    .A2(_10074_),
    .ZN(_10189_));
 OAI21_X4 _29431_ (.A(_10189_),
    .B1(_10075_),
    .B2(_04107_),
    .ZN(_10190_));
 NAND2_X2 _29432_ (.A1(_10125_),
    .A2(_10190_),
    .ZN(_10191_));
 OAI21_X1 _29433_ (.A(_10142_),
    .B1(_10072_),
    .B2(_10191_),
    .ZN(_10192_));
 NAND2_X2 _29434_ (.A1(_10188_),
    .A2(_10192_),
    .ZN(_10193_));
 MUX2_X1 _29435_ (.A(_10787_),
    .B(_10193_),
    .S(_10186_),
    .Z(_02539_));
 NAND2_X1 _29436_ (.A1(_11308_),
    .A2(_10063_),
    .ZN(_10194_));
 CLKBUF_X3 _29437_ (.A(_10127_),
    .Z(_10195_));
 CLKBUF_X3 _29438_ (.A(_10195_),
    .Z(_10196_));
 AOI21_X1 _29439_ (.A(_10149_),
    .B1(_10156_),
    .B2(_10147_),
    .ZN(_10197_));
 OR2_X1 _29440_ (.A1(_04120_),
    .A2(_10069_),
    .ZN(_10198_));
 OAI21_X4 _29441_ (.A(_10198_),
    .B1(_10070_),
    .B2(_08033_),
    .ZN(_10199_));
 BUF_X4 _29442_ (.A(_10199_),
    .Z(_10200_));
 AOI21_X1 _29443_ (.A(_10149_),
    .B1(_10200_),
    .B2(_10129_),
    .ZN(_10201_));
 BUF_X4 _29444_ (.A(_10068_),
    .Z(_10202_));
 NOR2_X2 _29445_ (.A1(_10157_),
    .A2(_10072_),
    .ZN(_10203_));
 OR2_X1 _29446_ (.A1(_04120_),
    .A2(_10086_),
    .ZN(_10204_));
 OAI21_X4 _29447_ (.A(_10204_),
    .B1(_10087_),
    .B2(_04107_),
    .ZN(_10205_));
 OAI222_X2 _29448_ (.A1(_10196_),
    .A2(_10197_),
    .B1(_10201_),
    .B2(_10202_),
    .C1(_10203_),
    .C2(_10205_),
    .ZN(_10206_));
 NOR2_X2 _29449_ (.A1(_10127_),
    .A2(_10191_),
    .ZN(_10207_));
 BUF_X4 _29450_ (.A(_10207_),
    .Z(_10208_));
 NAND3_X1 _29451_ (.A1(_10121_),
    .A2(_10140_),
    .A3(_10208_),
    .ZN(_10209_));
 OAI21_X1 _29452_ (.A(_10206_),
    .B1(_10209_),
    .B2(_10167_),
    .ZN(_10210_));
 OAI21_X1 _29453_ (.A(_10194_),
    .B1(_10210_),
    .B2(_10174_),
    .ZN(_02540_));
 NAND2_X2 _29454_ (.A1(_10088_),
    .A2(_10091_),
    .ZN(_10211_));
 NOR2_X4 _29455_ (.A1(_10108_),
    .A2(_10211_),
    .ZN(_10212_));
 NAND2_X2 _29456_ (.A1(_10208_),
    .A2(_10212_),
    .ZN(_10213_));
 NAND2_X4 _29457_ (.A1(_10068_),
    .A2(_10199_),
    .ZN(_10214_));
 NOR3_X1 _29458_ (.A1(_10158_),
    .A2(_10128_),
    .A3(_10214_),
    .ZN(_10215_));
 NAND2_X1 _29459_ (.A1(_10199_),
    .A2(_10129_),
    .ZN(_10216_));
 OAI21_X1 _29460_ (.A(_10216_),
    .B1(_10209_),
    .B2(_10199_),
    .ZN(_10217_));
 AOI221_X2 _29461_ (.A(_10151_),
    .B1(_10213_),
    .B2(_10215_),
    .C1(_10217_),
    .C2(_10188_),
    .ZN(_10218_));
 MUX2_X1 _29462_ (.A(_11310_),
    .B(_10218_),
    .S(_10186_),
    .Z(_02541_));
 CLKBUF_X3 _29463_ (.A(_10190_),
    .Z(_10219_));
 NAND2_X4 _29464_ (.A1(_10099_),
    .A2(_10103_),
    .ZN(_10220_));
 CLKBUF_X3 _29465_ (.A(_10133_),
    .Z(_10221_));
 AOI21_X1 _29466_ (.A(_10219_),
    .B1(_10220_),
    .B2(_10221_),
    .ZN(_10222_));
 OAI21_X1 _29467_ (.A(_10162_),
    .B1(_10143_),
    .B2(_10222_),
    .ZN(_10223_));
 INV_X1 _29468_ (.A(_10114_),
    .ZN(_10224_));
 NOR2_X1 _29469_ (.A1(_10224_),
    .A2(_10119_),
    .ZN(_10225_));
 OAI21_X1 _29470_ (.A(_10143_),
    .B1(_10211_),
    .B2(_10225_),
    .ZN(_10226_));
 NAND3_X1 _29471_ (.A1(_10171_),
    .A2(_10219_),
    .A3(_10226_),
    .ZN(_10227_));
 NOR2_X2 _29472_ (.A1(_10170_),
    .A2(_10214_),
    .ZN(_10228_));
 NAND4_X2 _29473_ (.A1(_10084_),
    .A2(_10223_),
    .A3(_10227_),
    .A4(_10228_),
    .ZN(_10229_));
 MUX2_X1 _29474_ (.A(_10105_),
    .B(_10107_),
    .S(_04120_),
    .Z(_10230_));
 BUF_X4 _29475_ (.A(_10230_),
    .Z(_10231_));
 NAND2_X4 _29476_ (.A1(_10142_),
    .A2(_10188_),
    .ZN(_10232_));
 NOR2_X1 _29477_ (.A1(_10158_),
    .A2(_10232_),
    .ZN(_10233_));
 AOI22_X2 _29478_ (.A1(_10231_),
    .A2(_10202_),
    .B1(_10233_),
    .B2(_10162_),
    .ZN(_10234_));
 OAI221_X2 _29479_ (.A(_10229_),
    .B1(_10234_),
    .B2(_10200_),
    .C1(_10193_),
    .C2(_10171_),
    .ZN(_10235_));
 MUX2_X1 _29480_ (.A(_10914_),
    .B(_10235_),
    .S(_10186_),
    .Z(_02542_));
 CLKBUF_X3 _29481_ (.A(_10072_),
    .Z(_10236_));
 NAND2_X1 _29482_ (.A1(_10190_),
    .A2(_10142_),
    .ZN(_10237_));
 AOI22_X1 _29483_ (.A1(_10196_),
    .A2(_10236_),
    .B1(_10237_),
    .B2(_10188_),
    .ZN(_10238_));
 NAND2_X4 _29484_ (.A1(_10190_),
    .A2(_10127_),
    .ZN(_10239_));
 NOR2_X1 _29485_ (.A1(_10110_),
    .A2(_10239_),
    .ZN(_10240_));
 NAND2_X2 _29486_ (.A1(_10091_),
    .A2(_10207_),
    .ZN(_10241_));
 INV_X1 _29487_ (.A(_10241_),
    .ZN(_10242_));
 CLKBUF_X3 _29488_ (.A(_10119_),
    .Z(_10243_));
 OAI21_X1 _29489_ (.A(_10149_),
    .B1(_10231_),
    .B2(_10243_),
    .ZN(_10244_));
 NOR2_X4 _29490_ (.A1(_10082_),
    .A2(_10146_),
    .ZN(_10245_));
 AND2_X2 _29491_ (.A1(_10245_),
    .A2(_10220_),
    .ZN(_10246_));
 AOI221_X2 _29492_ (.A(_10240_),
    .B1(_10242_),
    .B2(_10244_),
    .C1(_10246_),
    .C2(_10139_),
    .ZN(_10247_));
 NAND2_X1 _29493_ (.A1(_10190_),
    .A2(_10128_),
    .ZN(_10248_));
 CLKBUF_X3 _29494_ (.A(_10248_),
    .Z(_10249_));
 NAND2_X2 _29495_ (.A1(_10249_),
    .A2(_10156_),
    .ZN(_10250_));
 OAI21_X1 _29496_ (.A(_10238_),
    .B1(_10247_),
    .B2(_10250_),
    .ZN(_10251_));
 MUX2_X1 _29497_ (.A(_10882_),
    .B(_10251_),
    .S(_10186_),
    .Z(_02543_));
 OAI21_X2 _29498_ (.A(_10187_),
    .B1(_10068_),
    .B2(_10142_),
    .ZN(_10252_));
 NAND2_X1 _29499_ (.A1(_10158_),
    .A2(_10252_),
    .ZN(_10253_));
 NOR2_X2 _29500_ (.A1(_10205_),
    .A2(_10151_),
    .ZN(_10254_));
 OAI21_X1 _29501_ (.A(_10254_),
    .B1(_10121_),
    .B2(_10231_),
    .ZN(_10255_));
 AOI221_X1 _29502_ (.A(_10240_),
    .B1(_10246_),
    .B2(_10136_),
    .C1(_10255_),
    .C2(_10208_),
    .ZN(_10256_));
 OAI21_X1 _29503_ (.A(_10253_),
    .B1(_10256_),
    .B2(_10250_),
    .ZN(_10257_));
 MUX2_X1 _29504_ (.A(_10924_),
    .B(_10257_),
    .S(_10186_),
    .Z(_02544_));
 NAND2_X1 _29505_ (.A1(_11002_),
    .A2(_10063_),
    .ZN(_10258_));
 NAND2_X2 _29506_ (.A1(_10121_),
    .A2(_10140_),
    .ZN(_10259_));
 AOI21_X2 _29507_ (.A(_10148_),
    .B1(_10259_),
    .B2(_10109_),
    .ZN(_10260_));
 AOI221_X2 _29508_ (.A(_10169_),
    .B1(_10260_),
    .B2(_10098_),
    .C1(_10159_),
    .C2(_10195_),
    .ZN(_10261_));
 OR2_X1 _29509_ (.A1(_10167_),
    .A2(_10261_),
    .ZN(_10262_));
 NOR2_X2 _29510_ (.A1(_10077_),
    .A2(_10083_),
    .ZN(_10263_));
 NOR2_X1 _29511_ (.A1(_10148_),
    .A2(_10211_),
    .ZN(_10264_));
 OAI21_X1 _29512_ (.A(_10231_),
    .B1(_10263_),
    .B2(_10264_),
    .ZN(_10265_));
 NAND2_X2 _29513_ (.A1(_10245_),
    .A2(_10220_),
    .ZN(_10266_));
 OAI21_X1 _29514_ (.A(_10265_),
    .B1(_10266_),
    .B2(_10224_),
    .ZN(_10267_));
 AOI21_X1 _29515_ (.A(_10127_),
    .B1(_10212_),
    .B2(_10125_),
    .ZN(_10268_));
 MUX2_X1 _29516_ (.A(_10159_),
    .B(_10268_),
    .S(_10219_),
    .Z(_10269_));
 OAI21_X1 _29517_ (.A(_10156_),
    .B1(_10267_),
    .B2(_10269_),
    .ZN(_10270_));
 NOR2_X1 _29518_ (.A1(_10167_),
    .A2(_10261_),
    .ZN(_10271_));
 OAI21_X1 _29519_ (.A(_10249_),
    .B1(_10271_),
    .B2(_10267_),
    .ZN(_10272_));
 INV_X1 _29520_ (.A(_10098_),
    .ZN(_10273_));
 AOI22_X1 _29521_ (.A1(_10262_),
    .A2(_10270_),
    .B1(_10272_),
    .B2(_10273_),
    .ZN(_10274_));
 NAND2_X4 _29522_ (.A1(_10155_),
    .A2(_10199_),
    .ZN(_10275_));
 NOR3_X1 _29523_ (.A1(_10273_),
    .A2(_10275_),
    .A3(_10084_),
    .ZN(_10276_));
 AOI21_X1 _29524_ (.A(_10162_),
    .B1(_10085_),
    .B2(_10187_),
    .ZN(_10277_));
 NOR3_X1 _29525_ (.A1(_10274_),
    .A2(_10276_),
    .A3(_10277_),
    .ZN(_10278_));
 OAI21_X1 _29526_ (.A(_10258_),
    .B1(_10278_),
    .B2(_10174_),
    .ZN(_02545_));
 NAND2_X1 _29527_ (.A1(_11081_),
    .A2(_10063_),
    .ZN(_10279_));
 NAND2_X4 _29528_ (.A1(_10083_),
    .A2(_10191_),
    .ZN(_10280_));
 NAND2_X1 _29529_ (.A1(_04120_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .ZN(_10281_));
 NAND2_X1 _29530_ (.A1(_08033_),
    .A2(_04110_),
    .ZN(_10282_));
 NAND3_X1 _29531_ (.A1(_08073_),
    .A2(_10281_),
    .A3(_10282_),
    .ZN(_10283_));
 OAI21_X2 _29532_ (.A(_10283_),
    .B1(_08251_),
    .B2(_08073_),
    .ZN(_10284_));
 OAI21_X1 _29533_ (.A(_10280_),
    .B1(_10284_),
    .B2(_10083_),
    .ZN(_10285_));
 AOI21_X1 _29534_ (.A(_10285_),
    .B1(_10260_),
    .B2(_10103_),
    .ZN(_10286_));
 NOR2_X1 _29535_ (.A1(_10166_),
    .A2(_10286_),
    .ZN(_10287_));
 OAI21_X1 _29536_ (.A(_10146_),
    .B1(_10268_),
    .B2(_10157_),
    .ZN(_10288_));
 INV_X1 _29537_ (.A(_10264_),
    .ZN(_10289_));
 OAI21_X1 _29538_ (.A(_10239_),
    .B1(_10289_),
    .B2(_10284_),
    .ZN(_10290_));
 NAND2_X1 _29539_ (.A1(_10119_),
    .A2(_10220_),
    .ZN(_10291_));
 AOI22_X2 _29540_ (.A1(_10231_),
    .A2(_10290_),
    .B1(_10291_),
    .B2(_10245_),
    .ZN(_10292_));
 AOI21_X1 _29541_ (.A(_10214_),
    .B1(_10288_),
    .B2(_10292_),
    .ZN(_10293_));
 OAI21_X1 _29542_ (.A(_10292_),
    .B1(_10286_),
    .B2(_10166_),
    .ZN(_10294_));
 AND2_X1 _29543_ (.A1(_10249_),
    .A2(_10294_),
    .ZN(_10295_));
 OAI22_X2 _29544_ (.A1(_10287_),
    .A2(_10293_),
    .B1(_10295_),
    .B2(_10103_),
    .ZN(_10296_));
 NOR2_X1 _29545_ (.A1(_10200_),
    .A2(_10296_),
    .ZN(_10297_));
 NOR2_X4 _29546_ (.A1(_10127_),
    .A2(_10147_),
    .ZN(_10298_));
 OAI221_X2 _29547_ (.A(_10249_),
    .B1(_10298_),
    .B2(_10284_),
    .C1(_10084_),
    .C2(_10104_),
    .ZN(_10299_));
 OAI21_X1 _29548_ (.A(_10296_),
    .B1(_10284_),
    .B2(_10200_),
    .ZN(_10300_));
 AOI221_X2 _29549_ (.A(_10297_),
    .B1(_10299_),
    .B2(_10073_),
    .C1(_10202_),
    .C2(_10300_),
    .ZN(_10301_));
 OAI21_X1 _29550_ (.A(_10279_),
    .B1(_10301_),
    .B2(_10174_),
    .ZN(_02546_));
 MUX2_X1 _29551_ (.A(_04109_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(_04121_),
    .Z(_10302_));
 MUX2_X2 _29552_ (.A(_08263_),
    .B(_10302_),
    .S(_08073_),
    .Z(_10303_));
 OAI21_X2 _29553_ (.A(_10187_),
    .B1(_10085_),
    .B2(_10129_),
    .ZN(_10304_));
 INV_X2 _29554_ (.A(_10094_),
    .ZN(_10305_));
 NOR2_X2 _29555_ (.A1(_10305_),
    .A2(_10275_),
    .ZN(_10306_));
 NOR2_X1 _29556_ (.A1(_10190_),
    .A2(_10195_),
    .ZN(_10307_));
 AOI22_X2 _29557_ (.A1(_10303_),
    .A2(_10304_),
    .B1(_10306_),
    .B2(_10307_),
    .ZN(_10308_));
 NOR2_X2 _29558_ (.A1(_10263_),
    .A2(_10246_),
    .ZN(_10309_));
 NOR2_X1 _29559_ (.A1(_10109_),
    .A2(_10309_),
    .ZN(_10310_));
 OAI21_X1 _29560_ (.A(_10254_),
    .B1(_10225_),
    .B2(_10230_),
    .ZN(_10311_));
 AOI21_X1 _29561_ (.A(_10157_),
    .B1(_10208_),
    .B2(_10311_),
    .ZN(_10312_));
 NAND2_X1 _29562_ (.A1(_10109_),
    .A2(_10225_),
    .ZN(_10313_));
 NOR3_X1 _29563_ (.A1(_10305_),
    .A2(_10121_),
    .A3(_10313_),
    .ZN(_10314_));
 AOI21_X1 _29564_ (.A(_10314_),
    .B1(_10303_),
    .B2(_10212_),
    .ZN(_10315_));
 OAI22_X2 _29565_ (.A1(_10305_),
    .A2(_10312_),
    .B1(_10315_),
    .B2(_10148_),
    .ZN(_10316_));
 AOI221_X2 _29566_ (.A(_10310_),
    .B1(_10316_),
    .B2(_10159_),
    .C1(_10094_),
    .C2(_10170_),
    .ZN(_10317_));
 BUF_X4 _29567_ (.A(_10214_),
    .Z(_10318_));
 OR2_X1 _29568_ (.A1(_10170_),
    .A2(_10260_),
    .ZN(_10319_));
 AOI22_X1 _29569_ (.A1(_10094_),
    .A2(_10319_),
    .B1(_10303_),
    .B2(_10196_),
    .ZN(_10320_));
 OAI221_X2 _29570_ (.A(_10308_),
    .B1(_10317_),
    .B2(_10318_),
    .C1(_10320_),
    .C2(_10167_),
    .ZN(_10321_));
 MUX2_X1 _29571_ (.A(_10989_),
    .B(_10321_),
    .S(_10186_),
    .Z(_02547_));
 MUX2_X1 _29572_ (.A(net101),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(_04121_),
    .Z(_10322_));
 MUX2_X2 _29573_ (.A(_08275_),
    .B(_10322_),
    .S(_08073_),
    .Z(_10323_));
 AOI22_X1 _29574_ (.A1(_10149_),
    .A2(_10319_),
    .B1(_10323_),
    .B2(_10195_),
    .ZN(_10324_));
 NAND2_X1 _29575_ (.A1(_10230_),
    .A2(_10254_),
    .ZN(_10325_));
 NOR3_X1 _29576_ (.A1(_10161_),
    .A2(_10325_),
    .A3(_10323_),
    .ZN(_10326_));
 OAI21_X1 _29577_ (.A(_10190_),
    .B1(_10195_),
    .B2(_10326_),
    .ZN(_10327_));
 AOI21_X1 _29578_ (.A(_10310_),
    .B1(_10327_),
    .B2(_10146_),
    .ZN(_10328_));
 OAI22_X1 _29579_ (.A1(_10167_),
    .A2(_10324_),
    .B1(_10328_),
    .B2(_10318_),
    .ZN(_10329_));
 OAI21_X1 _29580_ (.A(_10329_),
    .B1(_10249_),
    .B2(_10149_),
    .ZN(_10330_));
 NOR2_X1 _29581_ (.A1(_10236_),
    .A2(_10170_),
    .ZN(_10331_));
 OAI21_X1 _29582_ (.A(_10331_),
    .B1(_10323_),
    .B2(_10307_),
    .ZN(_10332_));
 INV_X1 _29583_ (.A(_10323_),
    .ZN(_10333_));
 OAI221_X2 _29584_ (.A(_10330_),
    .B1(_10332_),
    .B2(_10202_),
    .C1(_10187_),
    .C2(_10333_),
    .ZN(_10334_));
 BUF_X8 _29585_ (.A(_08153_),
    .Z(_10335_));
 MUX2_X1 _29586_ (.A(_11056_),
    .B(_10334_),
    .S(_10335_),
    .Z(_02548_));
 NOR2_X1 _29587_ (.A1(_10202_),
    .A2(_10199_),
    .ZN(_10336_));
 AOI21_X1 _29588_ (.A(_10241_),
    .B1(_10259_),
    .B2(_10110_),
    .ZN(_10337_));
 NAND2_X1 _29589_ (.A1(_08040_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .ZN(_10338_));
 NAND2_X1 _29590_ (.A1(_08033_),
    .A2(net102),
    .ZN(_10339_));
 AOI21_X1 _29591_ (.A(_04105_),
    .B1(_10338_),
    .B2(_10339_),
    .ZN(_10340_));
 AOI21_X2 _29592_ (.A(_10340_),
    .B1(_08286_),
    .B2(_04123_),
    .ZN(_10341_));
 OAI21_X1 _29593_ (.A(_10249_),
    .B1(_10341_),
    .B2(_10142_),
    .ZN(_10342_));
 OAI21_X1 _29594_ (.A(_10336_),
    .B1(_10337_),
    .B2(_10342_),
    .ZN(_10343_));
 OAI21_X1 _29595_ (.A(_10248_),
    .B1(_10309_),
    .B2(_10109_),
    .ZN(_10344_));
 NOR2_X1 _29596_ (.A1(_10213_),
    .A2(_10341_),
    .ZN(_10345_));
 NOR2_X1 _29597_ (.A1(_10344_),
    .A2(_10345_),
    .ZN(_10346_));
 OAI21_X1 _29598_ (.A(_10343_),
    .B1(_10346_),
    .B2(_10318_),
    .ZN(_10347_));
 OAI21_X1 _29599_ (.A(_10347_),
    .B1(_10249_),
    .B2(_10091_),
    .ZN(_10348_));
 INV_X1 _29600_ (.A(_10304_),
    .ZN(_10349_));
 OAI21_X1 _29601_ (.A(_10348_),
    .B1(_10341_),
    .B2(_10349_),
    .ZN(_10350_));
 MUX2_X1 _29602_ (.A(_11054_),
    .B(_10350_),
    .S(_10335_),
    .Z(_02549_));
 OAI221_X1 _29603_ (.A(_10186_),
    .B1(_10129_),
    .B2(_10085_),
    .C1(_10213_),
    .C2(_10318_),
    .ZN(_10351_));
 INV_X1 _29604_ (.A(_10786_),
    .ZN(_10352_));
 OAI21_X1 _29605_ (.A(_10351_),
    .B1(_10186_),
    .B2(_10352_),
    .ZN(_02550_));
 MUX2_X1 _29606_ (.A(net104),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(_04121_),
    .Z(_10353_));
 MUX2_X2 _29607_ (.A(_08299_),
    .B(_10353_),
    .S(_08074_),
    .Z(_10354_));
 NOR2_X1 _29608_ (.A1(_10148_),
    .A2(_10325_),
    .ZN(_10355_));
 OAI22_X1 _29609_ (.A1(_10125_),
    .A2(_10084_),
    .B1(_10212_),
    .B2(_10148_),
    .ZN(_10356_));
 AOI221_X1 _29610_ (.A(_10344_),
    .B1(_10354_),
    .B2(_10355_),
    .C1(_10356_),
    .C2(_10221_),
    .ZN(_10357_));
 INV_X1 _29611_ (.A(_10354_),
    .ZN(_10358_));
 NOR4_X1 _29612_ (.A1(_10160_),
    .A2(_10109_),
    .A3(_10077_),
    .A4(_10259_),
    .ZN(_10359_));
 AOI21_X1 _29613_ (.A(_10359_),
    .B1(_10146_),
    .B2(_10221_),
    .ZN(_10360_));
 MUX2_X1 _29614_ (.A(_10358_),
    .B(_10360_),
    .S(_10142_),
    .Z(_10361_));
 OAI22_X1 _29615_ (.A1(_10318_),
    .A2(_10357_),
    .B1(_10361_),
    .B2(_10167_),
    .ZN(_10362_));
 OAI21_X1 _29616_ (.A(_10362_),
    .B1(_10249_),
    .B2(_10221_),
    .ZN(_10363_));
 NAND2_X1 _29617_ (.A1(_10188_),
    .A2(_10331_),
    .ZN(_10364_));
 NOR2_X1 _29618_ (.A1(_10161_),
    .A2(_10084_),
    .ZN(_10365_));
 AOI22_X2 _29619_ (.A1(_10280_),
    .A2(_10354_),
    .B1(_10365_),
    .B2(_10221_),
    .ZN(_10366_));
 OAI221_X2 _29620_ (.A(_10363_),
    .B1(_10364_),
    .B2(_10366_),
    .C1(_10187_),
    .C2(_10358_),
    .ZN(_10367_));
 MUX2_X1 _29621_ (.A(_12426_),
    .B(_10367_),
    .S(_10335_),
    .Z(_02551_));
 INV_X2 _29622_ (.A(_10139_),
    .ZN(_10368_));
 NAND2_X1 _29623_ (.A1(_10208_),
    .A2(_10311_),
    .ZN(_10369_));
 OAI21_X1 _29624_ (.A(_10190_),
    .B1(_10195_),
    .B2(_10161_),
    .ZN(_10370_));
 AOI21_X1 _29625_ (.A(_10214_),
    .B1(_10369_),
    .B2(_10370_),
    .ZN(_10371_));
 OAI21_X1 _29626_ (.A(_10146_),
    .B1(_10191_),
    .B2(_10313_),
    .ZN(_10372_));
 NAND2_X1 _29627_ (.A1(_10156_),
    .A2(_10372_),
    .ZN(_10373_));
 NAND2_X2 _29628_ (.A1(_10125_),
    .A2(_10077_),
    .ZN(_10374_));
 OAI21_X1 _29629_ (.A(_10373_),
    .B1(_10374_),
    .B2(_10166_),
    .ZN(_10375_));
 AOI21_X1 _29630_ (.A(_10371_),
    .B1(_10375_),
    .B2(_10143_),
    .ZN(_10376_));
 NOR2_X1 _29631_ (.A1(_10368_),
    .A2(_10376_),
    .ZN(_10377_));
 NOR3_X1 _29632_ (.A1(_10368_),
    .A2(_10157_),
    .A3(_10232_),
    .ZN(_10378_));
 MUX2_X1 _29633_ (.A(net105),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(_04121_),
    .Z(_10379_));
 MUX2_X2 _29634_ (.A(_08312_),
    .B(_10379_),
    .S(_08074_),
    .Z(_10380_));
 AOI21_X1 _29635_ (.A(_10378_),
    .B1(_10380_),
    .B2(_10232_),
    .ZN(_10381_));
 NAND2_X1 _29636_ (.A1(_10190_),
    .A2(_10380_),
    .ZN(_10382_));
 OAI21_X1 _29637_ (.A(_10382_),
    .B1(_10084_),
    .B2(_10368_),
    .ZN(_10383_));
 AOI22_X1 _29638_ (.A1(_10195_),
    .A2(_10380_),
    .B1(_10383_),
    .B2(_10159_),
    .ZN(_10384_));
 OAI22_X1 _29639_ (.A1(_10200_),
    .A2(_10381_),
    .B1(_10384_),
    .B2(_10275_),
    .ZN(_10385_));
 AOI21_X1 _29640_ (.A(_10246_),
    .B1(_10264_),
    .B2(_10380_),
    .ZN(_10386_));
 NOR3_X1 _29641_ (.A1(_10171_),
    .A2(_10250_),
    .A3(_10386_),
    .ZN(_10387_));
 OR3_X1 _29642_ (.A1(_10377_),
    .A2(_10385_),
    .A3(_10387_),
    .ZN(_10388_));
 MUX2_X1 _29643_ (.A(_12438_),
    .B(_10388_),
    .S(_10335_),
    .Z(_02552_));
 NAND2_X1 _29644_ (.A1(_12424_),
    .A2(_10063_),
    .ZN(_10389_));
 MUX2_X1 _29645_ (.A(net106),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(_08040_),
    .Z(_10390_));
 MUX2_X1 _29646_ (.A(_08317_),
    .B(_10390_),
    .S(_08074_),
    .Z(_10391_));
 OR2_X1 _29647_ (.A1(_04121_),
    .A2(_10134_),
    .ZN(_10392_));
 OAI21_X4 _29648_ (.A(_10392_),
    .B1(_10135_),
    .B2(_08033_),
    .ZN(_10393_));
 NOR2_X2 _29649_ (.A1(_10161_),
    .A2(_10190_),
    .ZN(_10394_));
 AOI22_X1 _29650_ (.A1(_10161_),
    .A2(_10243_),
    .B1(_10393_),
    .B2(_10394_),
    .ZN(_10395_));
 OAI221_X1 _29651_ (.A(_10188_),
    .B1(_10298_),
    .B2(_10391_),
    .C1(_10395_),
    .C2(_10195_),
    .ZN(_10396_));
 OR2_X1 _29652_ (.A1(_10236_),
    .A2(_10396_),
    .ZN(_10397_));
 NOR3_X1 _29653_ (.A1(_10393_),
    .A2(_10232_),
    .A3(_10365_),
    .ZN(_10398_));
 AOI21_X1 _29654_ (.A(_10398_),
    .B1(_10391_),
    .B2(_10232_),
    .ZN(_10399_));
 AOI21_X1 _29655_ (.A(_10214_),
    .B1(_10239_),
    .B2(_10369_),
    .ZN(_10400_));
 OAI22_X1 _29656_ (.A1(_10159_),
    .A2(_10214_),
    .B1(_10374_),
    .B2(_10167_),
    .ZN(_10401_));
 AOI21_X1 _29657_ (.A(_10400_),
    .B1(_10401_),
    .B2(_10143_),
    .ZN(_10402_));
 OAI221_X2 _29658_ (.A(_10397_),
    .B1(_10399_),
    .B2(_10200_),
    .C1(_10402_),
    .C2(_10393_),
    .ZN(_10403_));
 NAND2_X1 _29659_ (.A1(_10212_),
    .A2(_10391_),
    .ZN(_10404_));
 OAI21_X1 _29660_ (.A(_10404_),
    .B1(_10313_),
    .B2(_10393_),
    .ZN(_10405_));
 NAND2_X1 _29661_ (.A1(_10208_),
    .A2(_10405_),
    .ZN(_10406_));
 AOI21_X1 _29662_ (.A(_10246_),
    .B1(_10405_),
    .B2(_10208_),
    .ZN(_10407_));
 OAI22_X2 _29663_ (.A1(_10121_),
    .A2(_10406_),
    .B1(_10407_),
    .B2(_10171_),
    .ZN(_10408_));
 AOI21_X2 _29664_ (.A(_10403_),
    .B1(_10408_),
    .B2(_10228_),
    .ZN(_10409_));
 OAI21_X1 _29665_ (.A(_10389_),
    .B1(_10409_),
    .B2(_10174_),
    .ZN(_02553_));
 NAND2_X1 _29666_ (.A1(_12432_),
    .A2(_10063_),
    .ZN(_10410_));
 MUX2_X1 _29667_ (.A(net107),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(_08040_),
    .Z(_10411_));
 MUX2_X1 _29668_ (.A(_08319_),
    .B(_10411_),
    .S(_08074_),
    .Z(_10412_));
 NAND3_X1 _29669_ (.A1(_10236_),
    .A2(_10232_),
    .A3(_10412_),
    .ZN(_10413_));
 MUX2_X1 _29670_ (.A(_10114_),
    .B(_10088_),
    .S(_10157_),
    .Z(_10414_));
 OAI22_X1 _29671_ (.A1(_10298_),
    .A2(_10412_),
    .B1(_10414_),
    .B2(_10168_),
    .ZN(_10415_));
 OAI21_X1 _29672_ (.A(_10413_),
    .B1(_10415_),
    .B2(_10275_),
    .ZN(_10416_));
 OAI21_X1 _29673_ (.A(_10146_),
    .B1(_10191_),
    .B2(_10254_),
    .ZN(_10417_));
 NAND3_X1 _29674_ (.A1(_10114_),
    .A2(_10143_),
    .A3(_10417_),
    .ZN(_10418_));
 NOR2_X1 _29675_ (.A1(_10110_),
    .A2(_10412_),
    .ZN(_10419_));
 OAI221_X2 _29676_ (.A(_10418_),
    .B1(_10419_),
    .B2(_10289_),
    .C1(_10266_),
    .C2(_10110_),
    .ZN(_10420_));
 OAI21_X1 _29677_ (.A(_10203_),
    .B1(_10196_),
    .B2(_10162_),
    .ZN(_10421_));
 OAI22_X2 _29678_ (.A1(_10200_),
    .A2(_10232_),
    .B1(_10421_),
    .B2(_10188_),
    .ZN(_10422_));
 AOI221_X2 _29679_ (.A(_10416_),
    .B1(_10420_),
    .B2(_10228_),
    .C1(_10114_),
    .C2(_10422_),
    .ZN(_10423_));
 OAI21_X1 _29680_ (.A(_10410_),
    .B1(_10423_),
    .B2(_10174_),
    .ZN(_02554_));
 MUX2_X1 _29681_ (.A(net108),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(_04121_),
    .Z(_10424_));
 MUX2_X2 _29682_ (.A(_08321_),
    .B(_10424_),
    .S(_08074_),
    .Z(_10425_));
 AOI221_X1 _29683_ (.A(_10072_),
    .B1(_10280_),
    .B2(_10425_),
    .C1(_10128_),
    .C2(_10091_),
    .ZN(_10426_));
 NAND2_X1 _29684_ (.A1(_10243_),
    .A2(_10143_),
    .ZN(_10427_));
 OAI21_X1 _29685_ (.A(_10427_),
    .B1(_10425_),
    .B2(_10143_),
    .ZN(_10428_));
 AOI21_X1 _29686_ (.A(_10426_),
    .B1(_10428_),
    .B2(_10236_),
    .ZN(_10429_));
 NAND2_X1 _29687_ (.A1(_10188_),
    .A2(_10429_),
    .ZN(_10430_));
 NOR3_X1 _29688_ (.A1(_10151_),
    .A2(_10077_),
    .A3(_10083_),
    .ZN(_10431_));
 NAND2_X1 _29689_ (.A1(_10243_),
    .A2(_10157_),
    .ZN(_10432_));
 AOI221_X2 _29690_ (.A(_10431_),
    .B1(_10432_),
    .B2(_10128_),
    .C1(_10355_),
    .C2(_10425_),
    .ZN(_10433_));
 INV_X1 _29691_ (.A(_10220_),
    .ZN(_10434_));
 AOI22_X2 _29692_ (.A1(_10208_),
    .A2(_10211_),
    .B1(_10434_),
    .B2(_10245_),
    .ZN(_10435_));
 OAI221_X2 _29693_ (.A(_10433_),
    .B1(_10435_),
    .B2(_10243_),
    .C1(_10266_),
    .C2(_10171_),
    .ZN(_10436_));
 AOI21_X1 _29694_ (.A(_10318_),
    .B1(_10170_),
    .B2(_10243_),
    .ZN(_10437_));
 AOI22_X2 _29695_ (.A1(_10236_),
    .A2(_10425_),
    .B1(_10436_),
    .B2(_10437_),
    .ZN(_10438_));
 OAI21_X2 _29696_ (.A(_10430_),
    .B1(_10438_),
    .B2(_10188_),
    .ZN(_10439_));
 MUX2_X1 _29697_ (.A(_12419_),
    .B(_10439_),
    .S(_10335_),
    .Z(_02555_));
 NAND3_X1 _29698_ (.A1(_10231_),
    .A2(_10157_),
    .A3(_10142_),
    .ZN(_10440_));
 AOI21_X1 _29699_ (.A(_10068_),
    .B1(_10072_),
    .B2(_10440_),
    .ZN(_10441_));
 NOR2_X2 _29700_ (.A1(_10108_),
    .A2(_10241_),
    .ZN(_10442_));
 MUX2_X1 _29701_ (.A(net109),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(_04121_),
    .Z(_10443_));
 MUX2_X2 _29702_ (.A(_08322_),
    .B(_10443_),
    .S(_08074_),
    .Z(_10444_));
 OAI21_X1 _29703_ (.A(_10442_),
    .B1(_10444_),
    .B2(_10205_),
    .ZN(_10445_));
 AOI21_X1 _29704_ (.A(_10083_),
    .B1(_10220_),
    .B2(_10157_),
    .ZN(_10446_));
 OAI21_X1 _29705_ (.A(_10133_),
    .B1(_10394_),
    .B2(_10446_),
    .ZN(_10447_));
 AOI21_X1 _29706_ (.A(_10109_),
    .B1(_10168_),
    .B2(_10266_),
    .ZN(_10448_));
 NOR2_X1 _29707_ (.A1(_10169_),
    .A2(_10448_),
    .ZN(_10449_));
 NAND3_X1 _29708_ (.A1(_10445_),
    .A2(_10447_),
    .A3(_10449_),
    .ZN(_10450_));
 AOI21_X4 _29709_ (.A(_10214_),
    .B1(_10170_),
    .B2(_10109_),
    .ZN(_10451_));
 AOI221_X2 _29710_ (.A(_10441_),
    .B1(_10450_),
    .B2(_10451_),
    .C1(_10252_),
    .C2(_10444_),
    .ZN(_10452_));
 NAND2_X1 _29711_ (.A1(_10171_),
    .A2(_10298_),
    .ZN(_10453_));
 OAI21_X1 _29712_ (.A(_10453_),
    .B1(_10444_),
    .B2(_10298_),
    .ZN(_10454_));
 AOI21_X2 _29713_ (.A(_10452_),
    .B1(_10454_),
    .B2(_10073_),
    .ZN(_10455_));
 MUX2_X1 _29714_ (.A(_10945_),
    .B(_10455_),
    .S(_10335_),
    .Z(_02556_));
 NAND2_X1 _29715_ (.A1(_10869_),
    .A2(_10063_),
    .ZN(_10456_));
 MUX2_X1 _29716_ (.A(_10221_),
    .B(_10098_),
    .S(_10159_),
    .Z(_10457_));
 AND3_X1 _29717_ (.A1(_10336_),
    .A2(_10307_),
    .A3(_10457_),
    .ZN(_10458_));
 NOR2_X1 _29718_ (.A1(_10195_),
    .A2(_10068_),
    .ZN(_10459_));
 NAND2_X1 _29719_ (.A1(_08040_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .ZN(_10460_));
 NAND2_X1 _29720_ (.A1(_08033_),
    .A2(net110),
    .ZN(_10461_));
 AOI21_X2 _29721_ (.A(_04105_),
    .B1(_10460_),
    .B2(_10461_),
    .ZN(_10462_));
 AOI21_X4 _29722_ (.A(_10462_),
    .B1(_08252_),
    .B2(_04123_),
    .ZN(_10463_));
 NOR2_X1 _29723_ (.A1(_10098_),
    .A2(_10249_),
    .ZN(_10464_));
 NOR2_X1 _29724_ (.A1(_10114_),
    .A2(_10084_),
    .ZN(_10465_));
 OAI33_X1 _29725_ (.A1(_10200_),
    .A2(_10459_),
    .A3(_10463_),
    .B1(_10464_),
    .B2(_10465_),
    .B3(_10275_),
    .ZN(_10466_));
 NAND2_X1 _29726_ (.A1(_10280_),
    .A2(_10463_),
    .ZN(_10467_));
 OAI21_X1 _29727_ (.A(_10161_),
    .B1(_10142_),
    .B2(_10220_),
    .ZN(_10468_));
 NAND3_X1 _29728_ (.A1(_10114_),
    .A2(_10158_),
    .A3(_10468_),
    .ZN(_10469_));
 AOI21_X1 _29729_ (.A(_10241_),
    .B1(_10463_),
    .B2(_10149_),
    .ZN(_10470_));
 NOR3_X1 _29730_ (.A1(_10129_),
    .A2(_10246_),
    .A3(_10470_),
    .ZN(_10471_));
 OAI221_X2 _29731_ (.A(_10469_),
    .B1(_10471_),
    .B2(_10171_),
    .C1(_10273_),
    .C2(_10239_),
    .ZN(_10472_));
 AOI221_X2 _29732_ (.A(_10458_),
    .B1(_10466_),
    .B2(_10467_),
    .C1(_10472_),
    .C2(_10156_),
    .ZN(_10473_));
 OAI21_X1 _29733_ (.A(_10456_),
    .B1(_10473_),
    .B2(_10063_),
    .ZN(_02557_));
 OAI21_X1 _29734_ (.A(_10156_),
    .B1(_10248_),
    .B2(_10231_),
    .ZN(_10474_));
 MUX2_X1 _29735_ (.A(net111),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(_04120_),
    .Z(_10475_));
 MUX2_X1 _29736_ (.A(_08253_),
    .B(_10475_),
    .S(_08073_),
    .Z(_10476_));
 OAI21_X1 _29737_ (.A(_10442_),
    .B1(_10476_),
    .B2(_10205_),
    .ZN(_10477_));
 OAI21_X1 _29738_ (.A(_10477_),
    .B1(_10374_),
    .B2(_10243_),
    .ZN(_10478_));
 NAND3_X1 _29739_ (.A1(_10161_),
    .A2(_10139_),
    .A3(_10077_),
    .ZN(_10479_));
 OAI22_X1 _29740_ (.A1(_10243_),
    .A2(_10157_),
    .B1(_10220_),
    .B2(_10479_),
    .ZN(_10480_));
 AOI21_X1 _29741_ (.A(_10478_),
    .B1(_10480_),
    .B2(_10127_),
    .ZN(_10481_));
 AOI21_X1 _29742_ (.A(_10474_),
    .B1(_10449_),
    .B2(_10481_),
    .ZN(_10482_));
 MUX2_X1 _29743_ (.A(_10104_),
    .B(_10368_),
    .S(_10161_),
    .Z(_10483_));
 OAI21_X1 _29744_ (.A(_10072_),
    .B1(_10084_),
    .B2(_10483_),
    .ZN(_10484_));
 AOI221_X1 _29745_ (.A(_10482_),
    .B1(_10476_),
    .B2(_10252_),
    .C1(_10188_),
    .C2(_10484_),
    .ZN(_10485_));
 AOI22_X1 _29746_ (.A1(_10103_),
    .A2(_10170_),
    .B1(_10280_),
    .B2(_10476_),
    .ZN(_10486_));
 AOI21_X1 _29747_ (.A(_10485_),
    .B1(_10486_),
    .B2(_10073_),
    .ZN(_10487_));
 MUX2_X1 _29748_ (.A(_10873_),
    .B(_10487_),
    .S(_10335_),
    .Z(_02558_));
 NAND2_X1 _29749_ (.A1(_10876_),
    .A2(_08077_),
    .ZN(_10488_));
 MUX2_X1 _29750_ (.A(net112),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(_08040_),
    .Z(_10489_));
 MUX2_X2 _29751_ (.A(_08254_),
    .B(_10489_),
    .S(_08074_),
    .Z(_10490_));
 OAI21_X1 _29752_ (.A(_10442_),
    .B1(_10490_),
    .B2(_10205_),
    .ZN(_10491_));
 AOI22_X1 _29753_ (.A1(_10094_),
    .A2(_10263_),
    .B1(_10394_),
    .B2(_10231_),
    .ZN(_10492_));
 NAND3_X1 _29754_ (.A1(_10136_),
    .A2(_10245_),
    .A3(_10434_),
    .ZN(_10493_));
 NAND4_X1 _29755_ (.A1(_10449_),
    .A2(_10491_),
    .A3(_10492_),
    .A4(_10493_),
    .ZN(_10494_));
 NAND2_X2 _29756_ (.A1(_10187_),
    .A2(_10193_),
    .ZN(_10495_));
 AOI222_X2 _29757_ (.A1(_10170_),
    .A2(_10306_),
    .B1(_10451_),
    .B2(_10494_),
    .C1(_10495_),
    .C2(_10490_),
    .ZN(_10496_));
 OAI21_X1 _29758_ (.A(_10488_),
    .B1(_10496_),
    .B2(_10063_),
    .ZN(_02559_));
 NAND3_X1 _29759_ (.A1(_10149_),
    .A2(_10170_),
    .A3(_10073_),
    .ZN(_10497_));
 NAND2_X1 _29760_ (.A1(_08040_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .ZN(_10498_));
 NAND2_X1 _29761_ (.A1(_08033_),
    .A2(net113),
    .ZN(_10499_));
 AOI21_X1 _29762_ (.A(_04123_),
    .B1(_10498_),
    .B2(_10499_),
    .ZN(_10500_));
 AOI21_X2 _29763_ (.A(_10500_),
    .B1(_08255_),
    .B2(_04123_),
    .ZN(_10501_));
 AND2_X1 _29764_ (.A1(_10187_),
    .A2(_10193_),
    .ZN(_10502_));
 OAI221_X1 _29765_ (.A(_10249_),
    .B1(_10239_),
    .B2(_10205_),
    .C1(_10110_),
    .C2(_10219_),
    .ZN(_10503_));
 NAND2_X1 _29766_ (.A1(_10149_),
    .A2(_10501_),
    .ZN(_10504_));
 AOI21_X1 _29767_ (.A(_10503_),
    .B1(_10504_),
    .B2(_10442_),
    .ZN(_10505_));
 OAI221_X2 _29768_ (.A(_10497_),
    .B1(_10501_),
    .B2(_10502_),
    .C1(_10474_),
    .C2(_10505_),
    .ZN(_10506_));
 MUX2_X1 _29769_ (.A(_10875_),
    .B(_10506_),
    .S(_10335_),
    .Z(_02560_));
 NOR2_X1 _29770_ (.A1(_10213_),
    .A2(_10250_),
    .ZN(_10507_));
 OAI21_X1 _29771_ (.A(_10221_),
    .B1(_10304_),
    .B2(_10507_),
    .ZN(_10508_));
 NAND4_X1 _29772_ (.A1(_10160_),
    .A2(_10231_),
    .A3(_10121_),
    .A4(_10140_),
    .ZN(_10509_));
 AND2_X1 _29773_ (.A1(_10141_),
    .A2(_10509_),
    .ZN(_10510_));
 NOR2_X1 _29774_ (.A1(_10148_),
    .A2(_10510_),
    .ZN(_10511_));
 AOI21_X1 _29775_ (.A(_10511_),
    .B1(_10196_),
    .B2(_10221_),
    .ZN(_10512_));
 OAI221_X1 _29776_ (.A(_10508_),
    .B1(_10512_),
    .B2(_10167_),
    .C1(_10250_),
    .C2(_10309_),
    .ZN(_10513_));
 MUX2_X1 _29777_ (.A(_10790_),
    .B(_10513_),
    .S(_10335_),
    .Z(_02561_));
 NAND2_X1 _29778_ (.A1(_04121_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .ZN(_10514_));
 NAND2_X1 _29779_ (.A1(_08033_),
    .A2(net115),
    .ZN(_10515_));
 AOI21_X1 _29780_ (.A(_04105_),
    .B1(_10514_),
    .B2(_10515_),
    .ZN(_10516_));
 AOI21_X2 _29781_ (.A(_10516_),
    .B1(_08256_),
    .B2(_04105_),
    .ZN(_10517_));
 INV_X1 _29782_ (.A(_10517_),
    .ZN(_10518_));
 NOR2_X1 _29783_ (.A1(_10088_),
    .A2(_10091_),
    .ZN(_10519_));
 OAI21_X1 _29784_ (.A(_10088_),
    .B1(_10151_),
    .B2(_10121_),
    .ZN(_10520_));
 AOI221_X1 _29785_ (.A(_10519_),
    .B1(_10109_),
    .B2(_10520_),
    .C1(_10517_),
    .C2(_10212_),
    .ZN(_10521_));
 NOR3_X1 _29786_ (.A1(_10162_),
    .A2(_10195_),
    .A3(_10521_),
    .ZN(_10522_));
 OAI21_X1 _29787_ (.A(_10219_),
    .B1(_10143_),
    .B2(_10103_),
    .ZN(_10523_));
 OAI22_X1 _29788_ (.A1(_10171_),
    .A2(_10219_),
    .B1(_10522_),
    .B2(_10523_),
    .ZN(_10524_));
 AOI221_X2 _29789_ (.A(_08076_),
    .B1(_10495_),
    .B2(_10518_),
    .C1(_10524_),
    .C2(_10451_),
    .ZN(_10525_));
 AOI21_X1 _29790_ (.A(_10525_),
    .B1(_10174_),
    .B2(_10888_),
    .ZN(_02562_));
 MUX2_X1 _29791_ (.A(net116),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(_08040_),
    .Z(_10526_));
 MUX2_X1 _29792_ (.A(_08257_),
    .B(_10526_),
    .S(_08074_),
    .Z(_10527_));
 OAI21_X1 _29793_ (.A(_10091_),
    .B1(_10527_),
    .B2(_10205_),
    .ZN(_10528_));
 NAND2_X1 _29794_ (.A1(_10208_),
    .A2(_10528_),
    .ZN(_10529_));
 NOR2_X1 _29795_ (.A1(_10171_),
    .A2(_10318_),
    .ZN(_10530_));
 AOI221_X2 _29796_ (.A(_08076_),
    .B1(_10495_),
    .B2(_10527_),
    .C1(_10529_),
    .C2(_10530_),
    .ZN(_10531_));
 AOI21_X1 _29797_ (.A(_10531_),
    .B1(_10174_),
    .B2(_11727_),
    .ZN(_02563_));
 NOR2_X1 _29798_ (.A1(_10495_),
    .A2(_10507_),
    .ZN(_10532_));
 OAI22_X1 _29799_ (.A1(_10318_),
    .A2(_10239_),
    .B1(_10532_),
    .B2(_10368_),
    .ZN(_10533_));
 MUX2_X1 _29800_ (.A(_10798_),
    .B(_10533_),
    .S(_10335_),
    .Z(_02564_));
 OAI221_X1 _29801_ (.A(_10073_),
    .B1(_10196_),
    .B2(_10219_),
    .C1(_10136_),
    .C2(_10129_),
    .ZN(_10534_));
 NOR3_X1 _29802_ (.A1(_10393_),
    .A2(_10083_),
    .A3(_10068_),
    .ZN(_10535_));
 NOR2_X1 _29803_ (.A1(_10263_),
    .A2(_10394_),
    .ZN(_10536_));
 MUX2_X1 _29804_ (.A(_10136_),
    .B(_10536_),
    .S(_10199_),
    .Z(_10537_));
 AOI21_X1 _29805_ (.A(_10535_),
    .B1(_10537_),
    .B2(_10068_),
    .ZN(_10538_));
 AOI21_X1 _29806_ (.A(_10538_),
    .B1(_10212_),
    .B2(_10393_),
    .ZN(_10539_));
 OAI21_X1 _29807_ (.A(_10538_),
    .B1(_10232_),
    .B2(_10158_),
    .ZN(_10540_));
 AOI221_X1 _29808_ (.A(_10539_),
    .B1(_10540_),
    .B2(_10162_),
    .C1(_10233_),
    .C2(_10510_),
    .ZN(_10541_));
 OAI21_X1 _29809_ (.A(_10534_),
    .B1(_10541_),
    .B2(_10073_),
    .ZN(_10542_));
 BUF_X8 _29810_ (.A(_08153_),
    .Z(_10543_));
 MUX2_X1 _29811_ (.A(_10778_),
    .B(_10542_),
    .S(_10543_),
    .Z(_02565_));
 NAND3_X1 _29812_ (.A1(_10114_),
    .A2(_10202_),
    .A3(_10236_),
    .ZN(_10544_));
 OAI21_X1 _29813_ (.A(_10544_),
    .B1(_10129_),
    .B2(_10202_),
    .ZN(_10545_));
 OAI21_X1 _29814_ (.A(_10224_),
    .B1(_10196_),
    .B2(_10203_),
    .ZN(_10546_));
 NAND2_X1 _29815_ (.A1(_10545_),
    .A2(_10546_),
    .ZN(_10547_));
 OAI21_X1 _29816_ (.A(_10254_),
    .B1(_10114_),
    .B2(_10110_),
    .ZN(_10548_));
 AOI21_X1 _29817_ (.A(_10162_),
    .B1(_10219_),
    .B2(_10548_),
    .ZN(_10549_));
 OAI221_X1 _29818_ (.A(_10156_),
    .B1(_10146_),
    .B2(_10220_),
    .C1(_10549_),
    .C2(_10196_),
    .ZN(_10550_));
 NAND2_X1 _29819_ (.A1(_10547_),
    .A2(_10550_),
    .ZN(_10551_));
 MUX2_X1 _29820_ (.A(_10785_),
    .B(_10551_),
    .S(_10543_),
    .Z(_02566_));
 NAND4_X1 _29821_ (.A1(_10121_),
    .A2(_10140_),
    .A3(_10336_),
    .A4(_10208_),
    .ZN(_10552_));
 OAI221_X2 _29822_ (.A(_10552_),
    .B1(_10536_),
    .B2(_10318_),
    .C1(_10243_),
    .C2(_10532_),
    .ZN(_10553_));
 MUX2_X1 _29823_ (.A(_10779_),
    .B(_10553_),
    .S(_10543_),
    .Z(_02567_));
 NAND2_X1 _29824_ (.A1(_10147_),
    .A2(_10259_),
    .ZN(_10554_));
 NAND3_X1 _29825_ (.A1(_10146_),
    .A2(_10459_),
    .A3(_10554_),
    .ZN(_10555_));
 NAND3_X1 _29826_ (.A1(_10098_),
    .A2(_10236_),
    .A3(_10555_),
    .ZN(_10556_));
 AOI22_X2 _29827_ (.A1(_10221_),
    .A2(_10129_),
    .B1(_10280_),
    .B2(_10098_),
    .ZN(_10557_));
 OAI21_X1 _29828_ (.A(_10162_),
    .B1(_10219_),
    .B2(_10098_),
    .ZN(_10558_));
 OAI221_X2 _29829_ (.A(_10558_),
    .B1(_10374_),
    .B2(_10110_),
    .C1(_10273_),
    .C2(_10237_),
    .ZN(_10559_));
 NAND2_X1 _29830_ (.A1(_10159_),
    .A2(_10509_),
    .ZN(_10560_));
 NOR2_X1 _29831_ (.A1(_10167_),
    .A2(_10237_),
    .ZN(_10561_));
 AOI22_X2 _29832_ (.A1(_10156_),
    .A2(_10559_),
    .B1(_10560_),
    .B2(_10561_),
    .ZN(_10562_));
 OAI221_X2 _29833_ (.A(_10556_),
    .B1(_10557_),
    .B2(_10275_),
    .C1(_10464_),
    .C2(_10562_),
    .ZN(_10563_));
 MUX2_X1 _29834_ (.A(_11306_),
    .B(_10563_),
    .S(_10543_),
    .Z(_02568_));
 AOI221_X1 _29835_ (.A(_10275_),
    .B1(_10280_),
    .B2(_10103_),
    .C1(_10139_),
    .C2(_10129_),
    .ZN(_10564_));
 AOI21_X1 _29836_ (.A(_10232_),
    .B1(_10259_),
    .B2(_10219_),
    .ZN(_10565_));
 AOI21_X1 _29837_ (.A(_10565_),
    .B1(_10200_),
    .B2(_10158_),
    .ZN(_10566_));
 OAI221_X1 _29838_ (.A(_10103_),
    .B1(_10236_),
    .B2(_10239_),
    .C1(_10566_),
    .C2(_10162_),
    .ZN(_10567_));
 OAI21_X1 _29839_ (.A(_10202_),
    .B1(_10374_),
    .B2(_10368_),
    .ZN(_10568_));
 NAND2_X1 _29840_ (.A1(_10200_),
    .A2(_10568_),
    .ZN(_10569_));
 AOI21_X1 _29841_ (.A(_10564_),
    .B1(_10567_),
    .B2(_10569_),
    .ZN(_10570_));
 MUX2_X1 _29842_ (.A(_10862_),
    .B(_10570_),
    .S(_10543_),
    .Z(_02569_));
 NOR3_X1 _29843_ (.A1(_10305_),
    .A2(_10158_),
    .A3(_10196_),
    .ZN(_10571_));
 AOI21_X1 _29844_ (.A(_10571_),
    .B1(_10394_),
    .B2(_10136_),
    .ZN(_10572_));
 NAND3_X1 _29845_ (.A1(_10125_),
    .A2(_10243_),
    .A3(_10077_),
    .ZN(_10573_));
 OAI21_X1 _29846_ (.A(_10573_),
    .B1(_10136_),
    .B2(_10159_),
    .ZN(_10574_));
 AOI21_X1 _29847_ (.A(_10275_),
    .B1(_10574_),
    .B2(_10142_),
    .ZN(_10575_));
 AOI21_X1 _29848_ (.A(_10094_),
    .B1(_10298_),
    .B2(_10575_),
    .ZN(_10576_));
 NAND2_X1 _29849_ (.A1(_10199_),
    .A2(_10146_),
    .ZN(_10577_));
 AOI221_X1 _29850_ (.A(_10575_),
    .B1(_10577_),
    .B2(_10202_),
    .C1(_10072_),
    .C2(_10209_),
    .ZN(_10578_));
 OAI22_X1 _29851_ (.A1(_10318_),
    .A2(_10572_),
    .B1(_10576_),
    .B2(_10578_),
    .ZN(_10579_));
 MUX2_X1 _29852_ (.A(_11309_),
    .B(_10579_),
    .S(_10543_),
    .Z(_02570_));
 MUX2_X1 _29853_ (.A(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .B(_10202_),
    .S(_10543_),
    .Z(_02571_));
 MUX2_X1 _29854_ (.A(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .B(_10149_),
    .S(_10543_),
    .Z(_02572_));
 MUX2_X1 _29855_ (.A(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .B(_10091_),
    .S(_10543_),
    .Z(_02573_));
 MUX2_X1 _29856_ (.A(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .B(_10231_),
    .S(_10543_),
    .Z(_02574_));
 BUF_X8 _29857_ (.A(_08153_),
    .Z(_10580_));
 MUX2_X1 _29858_ (.A(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .B(_10196_),
    .S(_10580_),
    .Z(_02575_));
 MUX2_X1 _29859_ (.A(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .B(_10158_),
    .S(_10580_),
    .Z(_02576_));
 MUX2_X1 _29860_ (.A(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .B(_10159_),
    .S(_10580_),
    .Z(_02577_));
 MUX2_X1 _29861_ (.A(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .B(_10236_),
    .S(_10580_),
    .Z(_02578_));
 MUX2_X1 _29862_ (.A(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .B(_10221_),
    .S(_10580_),
    .Z(_02579_));
 MUX2_X1 _29863_ (.A(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .B(_10139_),
    .S(_10580_),
    .Z(_02580_));
 MUX2_X1 _29864_ (.A(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .B(_10136_),
    .S(_10580_),
    .Z(_02581_));
 MUX2_X1 _29865_ (.A(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .B(_10114_),
    .S(_10580_),
    .Z(_02582_));
 MUX2_X1 _29866_ (.A(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .B(_10120_),
    .S(_10580_),
    .Z(_02583_));
 MUX2_X1 _29867_ (.A(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .B(_10098_),
    .S(_10580_),
    .Z(_02584_));
 BUF_X8 _29868_ (.A(_08153_),
    .Z(_10581_));
 MUX2_X1 _29869_ (.A(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .B(_10103_),
    .S(_10581_),
    .Z(_02585_));
 MUX2_X1 _29870_ (.A(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .B(_10094_),
    .S(_10581_),
    .Z(_02586_));
 MUX2_X1 _29871_ (.A(\cs_registers_i.pc_id_i[10] ),
    .B(\cs_registers_i.pc_if_i[10] ),
    .S(_10581_),
    .Z(_02587_));
 MUX2_X1 _29872_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_08083_),
    .S(_10581_),
    .Z(_02588_));
 MUX2_X1 _29873_ (.A(\cs_registers_i.pc_id_i[12] ),
    .B(\cs_registers_i.pc_if_i[12] ),
    .S(_10581_),
    .Z(_02589_));
 MUX2_X1 _29874_ (.A(_12512_),
    .B(\cs_registers_i.pc_if_i[13] ),
    .S(_10581_),
    .Z(_02590_));
 MUX2_X1 _29875_ (.A(_12618_),
    .B(\cs_registers_i.pc_if_i[14] ),
    .S(_10581_),
    .Z(_02591_));
 MUX2_X1 _29876_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(_08123_),
    .S(_10581_),
    .Z(_02592_));
 MUX2_X1 _29877_ (.A(\cs_registers_i.pc_id_i[16] ),
    .B(\cs_registers_i.pc_if_i[16] ),
    .S(_10581_),
    .Z(_02593_));
 MUX2_X1 _29878_ (.A(_12868_),
    .B(_08138_),
    .S(_10581_),
    .Z(_02594_));
 BUF_X8 _29879_ (.A(_08153_),
    .Z(_10582_));
 MUX2_X1 _29880_ (.A(_12973_),
    .B(\cs_registers_i.pc_if_i[18] ),
    .S(_10582_),
    .Z(_02595_));
 MUX2_X1 _29881_ (.A(\cs_registers_i.pc_id_i[19] ),
    .B(_08151_),
    .S(_10582_),
    .Z(_02596_));
 MUX2_X1 _29882_ (.A(_04123_),
    .B(_11116_),
    .S(_08077_),
    .Z(_02597_));
 MUX2_X1 _29883_ (.A(\cs_registers_i.pc_id_i[20] ),
    .B(\cs_registers_i.pc_if_i[20] ),
    .S(_10582_),
    .Z(_02598_));
 MUX2_X1 _29884_ (.A(_13237_),
    .B(_08168_),
    .S(_10582_),
    .Z(_02599_));
 MUX2_X1 _29885_ (.A(_13347_),
    .B(\cs_registers_i.pc_if_i[22] ),
    .S(_10582_),
    .Z(_02600_));
 MUX2_X1 _29886_ (.A(_13423_),
    .B(\cs_registers_i.pc_if_i[23] ),
    .S(_10582_),
    .Z(_02601_));
 MUX2_X1 _29887_ (.A(\cs_registers_i.pc_id_i[24] ),
    .B(\cs_registers_i.pc_if_i[24] ),
    .S(_10582_),
    .Z(_02602_));
 MUX2_X1 _29888_ (.A(\cs_registers_i.pc_id_i[25] ),
    .B(\cs_registers_i.pc_if_i[25] ),
    .S(_10582_),
    .Z(_02603_));
 MUX2_X1 _29889_ (.A(_13688_),
    .B(_08194_),
    .S(_10582_),
    .Z(_02604_));
 MUX2_X1 _29890_ (.A(_03142_),
    .B(\cs_registers_i.pc_if_i[27] ),
    .S(_10582_),
    .Z(_02605_));
 CLKBUF_X3 _29891_ (.A(_08152_),
    .Z(_10583_));
 MUX2_X1 _29892_ (.A(_03238_),
    .B(\cs_registers_i.pc_if_i[28] ),
    .S(_10583_),
    .Z(_02606_));
 MUX2_X1 _29893_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(_08209_),
    .S(_10583_),
    .Z(_02607_));
 MUX2_X1 _29894_ (.A(\cs_registers_i.pc_id_i[2] ),
    .B(\cs_registers_i.pc_if_i[2] ),
    .S(_10583_),
    .Z(_02608_));
 MUX2_X1 _29895_ (.A(\cs_registers_i.pc_id_i[30] ),
    .B(\cs_registers_i.pc_if_i[30] ),
    .S(_10583_),
    .Z(_02609_));
 MUX2_X1 _29896_ (.A(\cs_registers_i.pc_id_i[31] ),
    .B(\cs_registers_i.pc_if_i[31] ),
    .S(_10583_),
    .Z(_02610_));
 MUX2_X1 _29897_ (.A(_11969_),
    .B(\cs_registers_i.pc_if_i[3] ),
    .S(_10583_),
    .Z(_02611_));
 MUX2_X1 _29898_ (.A(_12011_),
    .B(\cs_registers_i.pc_if_i[4] ),
    .S(_10583_),
    .Z(_02612_));
 MUX2_X1 _29899_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(\cs_registers_i.pc_if_i[5] ),
    .S(_10583_),
    .Z(_02613_));
 MUX2_X1 _29900_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(\cs_registers_i.pc_if_i[6] ),
    .S(_10583_),
    .Z(_02614_));
 MUX2_X1 _29901_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(_08093_),
    .S(_10583_),
    .Z(_02615_));
 MUX2_X1 _29902_ (.A(_12218_),
    .B(\cs_registers_i.pc_if_i[8] ),
    .S(_08153_),
    .Z(_02616_));
 MUX2_X1 _29903_ (.A(_12261_),
    .B(_08086_),
    .S(_08153_),
    .Z(_02617_));
 AND3_X1 _29904_ (.A1(_08860_),
    .A2(_08518_),
    .A3(_09358_),
    .ZN(_10584_));
 INV_X1 _29905_ (.A(_03660_),
    .ZN(_10585_));
 AOI21_X1 _29906_ (.A(_10584_),
    .B1(_09364_),
    .B2(_10585_),
    .ZN(_10586_));
 NAND2_X1 _29907_ (.A1(_04437_),
    .A2(_09725_),
    .ZN(_10587_));
 OAI21_X1 _29908_ (.A(_09358_),
    .B1(_09808_),
    .B2(_10587_),
    .ZN(_10588_));
 MUX2_X1 _29909_ (.A(\cs_registers_i.dcsr_q[0] ),
    .B(_10586_),
    .S(_10588_),
    .Z(_02822_));
 INV_X1 _29910_ (.A(_03661_),
    .ZN(_10589_));
 AOI21_X1 _29911_ (.A(_10584_),
    .B1(_09364_),
    .B2(_10589_),
    .ZN(_10590_));
 MUX2_X1 _29912_ (.A(\cs_registers_i.dcsr_q[1] ),
    .B(_10590_),
    .S(_10588_),
    .Z(_02827_));
 INV_X1 _29913_ (.A(_04312_),
    .ZN(_10591_));
 NAND2_X1 _29914_ (.A1(_03527_),
    .A2(_08045_),
    .ZN(_10592_));
 NOR3_X1 _29915_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(_04305_),
    .A3(_10592_),
    .ZN(_10593_));
 OAI21_X1 _29916_ (.A(_04009_),
    .B1(_03564_),
    .B2(_07255_),
    .ZN(_10594_));
 NAND4_X1 _29917_ (.A1(_00133_),
    .A2(_10591_),
    .A3(_10593_),
    .A4(_10594_),
    .ZN(core_busy_d));
 NAND2_X1 _29918_ (.A1(fetch_enable_q),
    .A2(_04125_),
    .ZN(net146));
 AND2_X1 _29919_ (.A1(clknet_1_0__leaf_clk_i),
    .A2(\core_clock_gate_i.en_latch ),
    .ZN(clk));
 NOR2_X1 _29920_ (.A1(_10914_),
    .A2(_03704_),
    .ZN(_10595_));
 AOI21_X1 _29921_ (.A(_10595_),
    .B1(_16487_),
    .B2(_10914_),
    .ZN(_10596_));
 MUX2_X2 _29922_ (.A(_16488_),
    .B(_10596_),
    .S(_08359_),
    .Z(net177));
 MUX2_X1 _29923_ (.A(_16498_),
    .B(_16492_),
    .S(_10914_),
    .Z(_10597_));
 MUX2_X2 _29924_ (.A(_16490_),
    .B(_10597_),
    .S(_08359_),
    .Z(net178));
 NAND3_X1 _29925_ (.A1(_10849_),
    .A2(_16503_),
    .A3(_08359_),
    .ZN(_10598_));
 BUF_X4 _29926_ (.A(_08358_),
    .Z(_10599_));
 BUF_X4 _29927_ (.A(_10599_),
    .Z(_10600_));
 NAND2_X1 _29928_ (.A1(_10600_),
    .A2(\load_store_unit_i.handle_misaligned_q ),
    .ZN(_10601_));
 NAND2_X1 _29929_ (.A1(_10914_),
    .A2(_16495_),
    .ZN(_10602_));
 MUX2_X1 _29930_ (.A(_16494_),
    .B(_10602_),
    .S(_08359_),
    .Z(_10603_));
 OAI221_X2 _29931_ (.A(_10598_),
    .B1(_10601_),
    .B2(_08359_),
    .C1(_10603_),
    .C2(\load_store_unit_i.handle_misaligned_q ),
    .ZN(net179));
 MUX2_X1 _29932_ (.A(_10599_),
    .B(_16489_),
    .S(_10914_),
    .Z(_10604_));
 MUX2_X2 _29933_ (.A(_16486_),
    .B(_10604_),
    .S(_08359_),
    .Z(net180));
 AOI21_X4 _29934_ (.A(_03523_),
    .B1(_03525_),
    .B2(_08343_),
    .ZN(net181));
 BUF_X4 _29935_ (.A(_04302_),
    .Z(_10605_));
 NOR2_X1 _29936_ (.A1(_10605_),
    .A2(net277),
    .ZN(_10606_));
 BUF_X4 _29937_ (.A(_16505_),
    .Z(_10607_));
 BUF_X4 _29938_ (.A(_10607_),
    .Z(_10608_));
 BUF_X1 _29939_ (.A(_16500_),
    .Z(_10609_));
 BUF_X4 _29940_ (.A(_10609_),
    .Z(_10610_));
 AOI222_X2 _29941_ (.A1(_10600_),
    .A2(_11648_),
    .B1(_12752_),
    .B2(_10608_),
    .C1(_13480_),
    .C2(_10610_),
    .ZN(_10611_));
 AOI21_X4 _29942_ (.A(_10606_),
    .B1(_10611_),
    .B2(_16485_),
    .ZN(net182));
 NOR2_X1 _29943_ (.A1(_10605_),
    .A2(_11724_),
    .ZN(_10612_));
 BUF_X4 _29944_ (.A(_10609_),
    .Z(_10613_));
 BUF_X4 _29945_ (.A(_10613_),
    .Z(_10614_));
 AOI222_X2 _29946_ (.A1(_10600_),
    .A2(net287),
    .B1(_13648_),
    .B2(_10608_),
    .C1(_10614_),
    .C2(net365),
    .ZN(_10615_));
 AOI21_X2 _29947_ (.A(_10612_),
    .B1(_10615_),
    .B2(_16485_),
    .ZN(net183));
 AOI22_X1 _29948_ (.A1(_10599_),
    .A2(net283),
    .B1(_03104_),
    .B2(_10607_),
    .ZN(_10616_));
 INV_X1 _29949_ (.A(_10609_),
    .ZN(_10617_));
 OAI21_X1 _29950_ (.A(_10616_),
    .B1(_03815_),
    .B2(_10617_),
    .ZN(_10618_));
 MUX2_X1 _29951_ (.A(_11769_),
    .B(_10618_),
    .S(_04302_),
    .Z(net184));
 NOR2_X1 _29952_ (.A1(_10605_),
    .A2(_12420_),
    .ZN(_10619_));
 AOI222_X2 _29953_ (.A1(_10600_),
    .A2(_13118_),
    .B1(_03198_),
    .B2(_10608_),
    .C1(_10614_),
    .C2(net331),
    .ZN(_10620_));
 AOI21_X2 _29954_ (.A(_10619_),
    .B1(_10620_),
    .B2(_16485_),
    .ZN(net185));
 NOR2_X1 _29955_ (.A1(_10605_),
    .A2(net325),
    .ZN(_10621_));
 AOI222_X2 _29956_ (.A1(_10600_),
    .A2(_13198_),
    .B1(_03276_),
    .B2(_10608_),
    .C1(_10614_),
    .C2(_03831_),
    .ZN(_10622_));
 AOI21_X2 _29957_ (.A(_10621_),
    .B1(_10622_),
    .B2(_16485_),
    .ZN(net186));
 CLKBUF_X3 _29958_ (.A(_04302_),
    .Z(_10623_));
 NOR2_X1 _29959_ (.A1(_10623_),
    .A2(_12580_),
    .ZN(_10624_));
 BUF_X4 _29960_ (.A(_10607_),
    .Z(_10625_));
 AOI222_X2 _29961_ (.A1(_10600_),
    .A2(net323),
    .B1(_03372_),
    .B2(_10625_),
    .C1(_10614_),
    .C2(net362),
    .ZN(_10626_));
 AOI21_X2 _29962_ (.A(_10624_),
    .B1(_10626_),
    .B2(_16485_),
    .ZN(net187));
 NOR2_X1 _29963_ (.A1(_10623_),
    .A2(net318),
    .ZN(_10627_));
 AOI222_X2 _29964_ (.A1(_10600_),
    .A2(net319),
    .B1(_03452_),
    .B2(_10625_),
    .C1(_10610_),
    .C2(_03849_),
    .ZN(_10628_));
 AOI21_X2 _29965_ (.A(_10627_),
    .B1(_10628_),
    .B2(_16485_),
    .ZN(net188));
 NOR2_X1 _29966_ (.A1(_10623_),
    .A2(_12752_),
    .ZN(_10629_));
 AOI222_X2 _29967_ (.A1(_10608_),
    .A2(net277),
    .B1(_11648_),
    .B2(_10614_),
    .C1(_13480_),
    .C2(_10599_),
    .ZN(_10630_));
 AOI21_X2 _29968_ (.A(_10629_),
    .B1(_10630_),
    .B2(_16485_),
    .ZN(net189));
 AOI22_X1 _29969_ (.A1(_10613_),
    .A2(_03867_),
    .B1(_13555_),
    .B2(_08358_),
    .ZN(_10631_));
 INV_X1 _29970_ (.A(_16505_),
    .ZN(_10632_));
 OAI21_X1 _29971_ (.A(_10631_),
    .B1(net301),
    .B2(_10632_),
    .ZN(_10633_));
 NOR2_X1 _29972_ (.A1(_03704_),
    .A2(_10633_),
    .ZN(_10634_));
 AOI21_X2 _29973_ (.A(_10634_),
    .B1(_12825_),
    .B2(_03704_),
    .ZN(net190));
 NOR2_X1 _29974_ (.A1(_10623_),
    .A2(net286),
    .ZN(_10635_));
 AOI222_X2 _29975_ (.A1(_10608_),
    .A2(net365),
    .B1(_11724_),
    .B2(_10614_),
    .C1(_13648_),
    .C2(_10599_),
    .ZN(_10636_));
 AOI21_X2 _29976_ (.A(_10635_),
    .B1(_10636_),
    .B2(_16485_),
    .ZN(net191));
 AOI22_X1 _29977_ (.A1(_10613_),
    .A2(_11769_),
    .B1(_03104_),
    .B2(_08358_),
    .ZN(_10637_));
 OAI21_X1 _29978_ (.A(_10637_),
    .B1(_03815_),
    .B2(_10632_),
    .ZN(_10638_));
 MUX2_X2 _29979_ (.A(net283),
    .B(_10638_),
    .S(_04302_),
    .Z(net192));
 AOI22_X1 _29980_ (.A1(_08358_),
    .A2(_03867_),
    .B1(_13555_),
    .B2(_10613_),
    .ZN(_10639_));
 OAI21_X1 _29981_ (.A(_10639_),
    .B1(_12825_),
    .B2(_10632_),
    .ZN(_10640_));
 NOR2_X1 _29982_ (.A1(_03704_),
    .A2(_10640_),
    .ZN(_10641_));
 AOI21_X2 _29983_ (.A(_10641_),
    .B1(net301),
    .B2(_03704_),
    .ZN(net193));
 NOR2_X1 _29984_ (.A1(_10623_),
    .A2(_13118_),
    .ZN(_10642_));
 AOI222_X2 _29985_ (.A1(_10608_),
    .A2(net331),
    .B1(_12420_),
    .B2(_10614_),
    .C1(_03198_),
    .C2(_10599_),
    .ZN(_10643_));
 AOI21_X2 _29986_ (.A(_10642_),
    .B1(_10643_),
    .B2(_16485_),
    .ZN(net194));
 NOR2_X1 _29987_ (.A1(_10623_),
    .A2(_13198_),
    .ZN(_10644_));
 AOI222_X2 _29988_ (.A1(_10608_),
    .A2(_03831_),
    .B1(net325),
    .B2(_10614_),
    .C1(_03276_),
    .C2(_10599_),
    .ZN(_10645_));
 BUF_X4 _29989_ (.A(_04302_),
    .Z(_10646_));
 AOI21_X2 _29990_ (.A(_10644_),
    .B1(_10645_),
    .B2(_10646_),
    .ZN(net195));
 NOR2_X1 _29991_ (.A1(_10623_),
    .A2(net323),
    .ZN(_10647_));
 AOI222_X2 _29992_ (.A1(_10608_),
    .A2(net362),
    .B1(_12580_),
    .B2(_10614_),
    .C1(_03372_),
    .C2(_10599_),
    .ZN(_10648_));
 AOI21_X2 _29993_ (.A(_10647_),
    .B1(_10648_),
    .B2(_10646_),
    .ZN(net196));
 NOR2_X1 _29994_ (.A1(_10623_),
    .A2(net319),
    .ZN(_10649_));
 AOI222_X2 _29995_ (.A1(_10608_),
    .A2(_03849_),
    .B1(net318),
    .B2(_10614_),
    .C1(_03452_),
    .C2(_10599_),
    .ZN(_10650_));
 AOI21_X2 _29996_ (.A(_10649_),
    .B1(_10650_),
    .B2(_10646_),
    .ZN(net197));
 NOR2_X1 _29997_ (.A1(_10623_),
    .A2(_13480_),
    .ZN(_10651_));
 AOI222_X2 _29998_ (.A1(_10600_),
    .A2(net277),
    .B1(_11648_),
    .B2(_10625_),
    .C1(_12752_),
    .C2(_10610_),
    .ZN(_10652_));
 AOI21_X2 _29999_ (.A(_10651_),
    .B1(_10652_),
    .B2(_10646_),
    .ZN(net198));
 INV_X1 _30000_ (.A(_08358_),
    .ZN(_10653_));
 OAI222_X2 _30001_ (.A1(_10653_),
    .A2(net302),
    .B1(_11686_),
    .B2(_10632_),
    .C1(_12825_),
    .C2(_10617_),
    .ZN(_10654_));
 MUX2_X2 _30002_ (.A(_13555_),
    .B(_10654_),
    .S(_04302_),
    .Z(net199));
 NOR2_X1 _30003_ (.A1(_10623_),
    .A2(_13648_),
    .ZN(_10655_));
 AOI222_X2 _30004_ (.A1(_10600_),
    .A2(net364),
    .B1(_11724_),
    .B2(_10625_),
    .C1(net286),
    .C2(_10610_),
    .ZN(_10656_));
 AOI21_X2 _30005_ (.A(_10655_),
    .B1(_10656_),
    .B2(_10646_),
    .ZN(net200));
 AOI22_X1 _30006_ (.A1(_10607_),
    .A2(_11769_),
    .B1(net284),
    .B2(_10613_),
    .ZN(_10657_));
 OAI21_X1 _30007_ (.A(_10657_),
    .B1(_03815_),
    .B2(_10653_),
    .ZN(_10658_));
 MUX2_X2 _30008_ (.A(_03104_),
    .B(_10658_),
    .S(_04302_),
    .Z(net201));
 CLKBUF_X3 _30009_ (.A(_03705_),
    .Z(_10659_));
 NOR2_X1 _30010_ (.A1(_10659_),
    .A2(_03198_),
    .ZN(_10660_));
 AOI222_X2 _30011_ (.A1(_10600_),
    .A2(net331),
    .B1(_12420_),
    .B2(_10625_),
    .C1(_13118_),
    .C2(_10610_),
    .ZN(_10661_));
 AOI21_X2 _30012_ (.A(_10660_),
    .B1(_10661_),
    .B2(_10646_),
    .ZN(net202));
 NOR2_X1 _30013_ (.A1(_10659_),
    .A2(_03276_),
    .ZN(_10662_));
 BUF_X4 _30014_ (.A(_10599_),
    .Z(_10663_));
 AOI222_X2 _30015_ (.A1(_10663_),
    .A2(_03831_),
    .B1(net325),
    .B2(_10625_),
    .C1(_13198_),
    .C2(_10610_),
    .ZN(_10664_));
 AOI21_X2 _30016_ (.A(_10662_),
    .B1(_10664_),
    .B2(_10646_),
    .ZN(net203));
 NOR2_X1 _30017_ (.A1(_10659_),
    .A2(net364),
    .ZN(_10665_));
 AOI222_X2 _30018_ (.A1(_10663_),
    .A2(_11724_),
    .B1(net286),
    .B2(_10625_),
    .C1(_13648_),
    .C2(_10610_),
    .ZN(_10666_));
 AOI21_X2 _30019_ (.A(_10665_),
    .B1(_10666_),
    .B2(_10646_),
    .ZN(net204));
 NOR2_X1 _30020_ (.A1(_10659_),
    .A2(_03372_),
    .ZN(_10667_));
 AOI222_X2 _30021_ (.A1(_10663_),
    .A2(net362),
    .B1(_12580_),
    .B2(_10625_),
    .C1(_13307_),
    .C2(_10610_),
    .ZN(_10668_));
 AOI21_X2 _30022_ (.A(_10667_),
    .B1(_10668_),
    .B2(_10646_),
    .ZN(net205));
 NOR2_X1 _30023_ (.A1(_10659_),
    .A2(_03452_),
    .ZN(_10669_));
 AOI222_X2 _30024_ (.A1(_10663_),
    .A2(_03849_),
    .B1(net318),
    .B2(_10625_),
    .C1(_13384_),
    .C2(_10610_),
    .ZN(_10670_));
 AOI21_X2 _30025_ (.A(_10669_),
    .B1(_10670_),
    .B2(_10646_),
    .ZN(net206));
 NOR2_X1 _30026_ (.A1(_10659_),
    .A2(_11427_),
    .ZN(_10671_));
 AOI222_X2 _30027_ (.A1(_10663_),
    .A2(_11769_),
    .B1(net283),
    .B2(_10625_),
    .C1(_03104_),
    .C2(_10613_),
    .ZN(_10672_));
 AOI21_X2 _30028_ (.A(_10671_),
    .B1(_10672_),
    .B2(_10605_),
    .ZN(net207));
 NOR2_X1 _30029_ (.A1(_10659_),
    .A2(net331),
    .ZN(_10673_));
 AOI222_X2 _30030_ (.A1(_10663_),
    .A2(_12420_),
    .B1(net368),
    .B2(_10607_),
    .C1(_03198_),
    .C2(_10613_),
    .ZN(_10674_));
 AOI21_X2 _30031_ (.A(_10673_),
    .B1(_10674_),
    .B2(_10605_),
    .ZN(net208));
 NOR2_X1 _30032_ (.A1(_10659_),
    .A2(_03831_),
    .ZN(_10675_));
 AOI222_X2 _30033_ (.A1(_10663_),
    .A2(net325),
    .B1(_13198_),
    .B2(_10607_),
    .C1(_03276_),
    .C2(_10613_),
    .ZN(_10676_));
 AOI21_X2 _30034_ (.A(_10675_),
    .B1(_10676_),
    .B2(_10605_),
    .ZN(net209));
 NOR2_X1 _30035_ (.A1(_10659_),
    .A2(net362),
    .ZN(_10677_));
 AOI222_X2 _30036_ (.A1(_10663_),
    .A2(_12580_),
    .B1(net323),
    .B2(_10607_),
    .C1(_03372_),
    .C2(_10613_),
    .ZN(_10678_));
 AOI21_X2 _30037_ (.A(_10677_),
    .B1(_10678_),
    .B2(_10605_),
    .ZN(net210));
 NOR2_X1 _30038_ (.A1(_10659_),
    .A2(_03849_),
    .ZN(_10679_));
 AOI222_X2 _30039_ (.A1(_10663_),
    .A2(net318),
    .B1(net319),
    .B2(_10607_),
    .C1(_03452_),
    .C2(_10613_),
    .ZN(_10680_));
 AOI21_X4 _30040_ (.A(_10679_),
    .B1(_10680_),
    .B2(_10605_),
    .ZN(net211));
 NOR2_X1 _30041_ (.A1(_04302_),
    .A2(_11648_),
    .ZN(_10681_));
 AOI222_X2 _30042_ (.A1(_10663_),
    .A2(_12752_),
    .B1(_13480_),
    .B2(_10607_),
    .C1(_10610_),
    .C2(net277),
    .ZN(_10682_));
 AOI21_X2 _30043_ (.A(_10681_),
    .B1(_10682_),
    .B2(_10605_),
    .ZN(net212));
 NAND2_X1 _30044_ (.A1(_10607_),
    .A2(_13555_),
    .ZN(_10683_));
 OAI221_X1 _30045_ (.A(_10683_),
    .B1(net302),
    .B2(_10617_),
    .C1(_10653_),
    .C2(_12825_),
    .ZN(_10684_));
 MUX2_X2 _30046_ (.A(_03867_),
    .B(_10684_),
    .S(_04302_),
    .Z(net213));
 NAND2_X2 _30047_ (.A1(_00133_),
    .A2(_10591_),
    .ZN(net245));
 NAND2_X1 _30048_ (.A1(net93),
    .A2(net245),
    .ZN(_10685_));
 NOR2_X1 _30049_ (.A1(_04102_),
    .A2(_10685_),
    .ZN(_10686_));
 OAI21_X1 _30050_ (.A(_04305_),
    .B1(net124),
    .B2(_04081_),
    .ZN(_10687_));
 AOI21_X1 _30051_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .B1(_04081_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_10688_));
 AOI22_X1 _30052_ (.A1(_08034_),
    .A2(_10687_),
    .B1(_10688_),
    .B2(_08036_),
    .ZN(_10689_));
 OR2_X1 _30053_ (.A1(_10686_),
    .A2(_10689_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 NAND2_X1 _30054_ (.A1(_04305_),
    .A2(_10686_),
    .ZN(_10690_));
 AOI21_X1 _30055_ (.A(_08036_),
    .B1(_10688_),
    .B2(_10690_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 MUX2_X1 _30056_ (.A(_08039_),
    .B(_08050_),
    .S(_08054_),
    .Z(_10691_));
 AND2_X1 _30057_ (.A1(_07858_),
    .A2(_10691_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 MUX2_X1 _30058_ (.A(_08062_),
    .B(_08039_),
    .S(_08054_),
    .Z(_10692_));
 AND2_X1 _30059_ (.A1(_07858_),
    .A2(_10692_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 AND3_X1 _30060_ (.A1(_07858_),
    .A2(_08054_),
    .A3(_08062_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 NAND2_X1 _30061_ (.A1(_00134_),
    .A2(net124),
    .ZN(_10693_));
 NAND2_X1 _30062_ (.A1(_04305_),
    .A2(_10693_),
    .ZN(_10694_));
 NAND2_X1 _30063_ (.A1(_10685_),
    .A2(_10694_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 NAND3_X1 _30064_ (.A1(_04305_),
    .A2(net93),
    .A3(net245),
    .ZN(_10695_));
 AOI21_X1 _30065_ (.A(_08036_),
    .B1(_10695_),
    .B2(_00134_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 AOI21_X1 _30066_ (.A(net93),
    .B1(_10591_),
    .B2(_00133_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 NOR2_X1 _30067_ (.A1(_03999_),
    .A2(_07285_),
    .ZN(_10696_));
 NOR4_X2 _30068_ (.A1(_10810_),
    .A2(_04027_),
    .A3(_08045_),
    .A4(_10696_),
    .ZN(_10697_));
 NAND2_X1 _30069_ (.A1(_08079_),
    .A2(_10697_),
    .ZN(_10698_));
 OAI21_X1 _30070_ (.A(_10698_),
    .B1(_10174_),
    .B2(_08068_),
    .ZN(\if_stage_i.instr_valid_id_d ));
 FA_X1 _30071_ (.A(_14466_),
    .B(_14464_),
    .CI(_14465_),
    .CO(_14467_),
    .S(\alu_adder_result_ex[0] ));
 FA_X1 _30072_ (.A(_14468_),
    .B(_14469_),
    .CI(_14470_),
    .CO(_14471_),
    .S(_14472_));
 FA_X1 _30073_ (.A(_14473_),
    .B(_14474_),
    .CI(_14475_),
    .CO(_14476_),
    .S(_14477_));
 FA_X1 _30074_ (.A(_14478_),
    .B(_14479_),
    .CI(_14480_),
    .CO(_14481_),
    .S(_14482_));
 FA_X1 _30075_ (.A(_14483_),
    .B(_14484_),
    .CI(_14485_),
    .CO(_14486_),
    .S(_14487_));
 FA_X1 _30076_ (.A(_14488_),
    .B(_14489_),
    .CI(_14490_),
    .CO(_14491_),
    .S(_14492_));
 FA_X1 _30077_ (.A(_14493_),
    .B(_14494_),
    .CI(_14495_),
    .CO(_14496_),
    .S(_14497_));
 FA_X1 _30078_ (.A(_14498_),
    .B(_14499_),
    .CI(_14500_),
    .CO(_14501_),
    .S(_14502_));
 FA_X1 _30079_ (.A(_14503_),
    .B(_14504_),
    .CI(_14505_),
    .CO(_14506_),
    .S(_14507_));
 FA_X1 _30080_ (.A(_14508_),
    .B(_14509_),
    .CI(_14510_),
    .CO(_14511_),
    .S(_14512_));
 FA_X1 _30081_ (.A(_14491_),
    .B(_14513_),
    .CI(_14512_),
    .CO(_14514_),
    .S(_14515_));
 FA_X1 _30082_ (.A(_14516_),
    .B(_14517_),
    .CI(_14518_),
    .CO(_14519_),
    .S(_14520_));
 FA_X1 _30083_ (.A(_14521_),
    .B(_14522_),
    .CI(_14523_),
    .CO(_14524_),
    .S(_14525_));
 FA_X1 _30084_ (.A(_14526_),
    .B(_14527_),
    .CI(_14528_),
    .CO(_14529_),
    .S(_14530_));
 FA_X1 _30085_ (.A(_14531_),
    .B(_14532_),
    .CI(_14533_),
    .CO(_14534_),
    .S(_14535_));
 FA_X1 _30086_ (.A(_14536_),
    .B(_14535_),
    .CI(_14511_),
    .CO(_14537_),
    .S(_14538_));
 FA_X1 _30087_ (.A(_14539_),
    .B(_14540_),
    .CI(_14541_),
    .CO(_14542_),
    .S(_14543_));
 FA_X1 _30088_ (.A(_14544_),
    .B(_14545_),
    .CI(_14546_),
    .CO(_14547_),
    .S(_14548_));
 FA_X1 _30089_ (.A(_14549_),
    .B(_14550_),
    .CI(_14551_),
    .CO(_14552_),
    .S(_14553_));
 FA_X1 _30090_ (.A(_14554_),
    .B(_14553_),
    .CI(_14555_),
    .CO(_14556_),
    .S(_14557_));
 FA_X1 _30091_ (.A(_14558_),
    .B(_14559_),
    .CI(_14560_),
    .CO(_14561_),
    .S(_14562_));
 FA_X1 _30092_ (.A(_14534_),
    .B(_14563_),
    .CI(_14562_),
    .CO(_14564_),
    .S(_14565_));
 FA_X1 _30093_ (.A(_14566_),
    .B(_14567_),
    .CI(_14568_),
    .CO(_14569_),
    .S(_14570_));
 FA_X1 _30094_ (.A(_14571_),
    .B(_14572_),
    .CI(_14573_),
    .CO(_14574_),
    .S(_14575_));
 FA_X1 _30095_ (.A(_14576_),
    .B(_14577_),
    .CI(_14578_),
    .CO(_14579_),
    .S(_14580_));
 FA_X1 _30096_ (.A(_14581_),
    .B(_14582_),
    .CI(_14583_),
    .CO(_14584_),
    .S(_14585_));
 FA_X1 _30097_ (.A(_14586_),
    .B(_14580_),
    .CI(_14547_),
    .CO(_14587_),
    .S(_14588_));
 FA_X1 _30098_ (.A(_14589_),
    .B(_14590_),
    .CI(_14591_),
    .CO(_14592_),
    .S(_14593_));
 FA_X1 _30099_ (.A(_14594_),
    .B(_14593_),
    .CI(_14561_),
    .CO(_14595_),
    .S(_14596_));
 FA_X1 _30100_ (.A(_14597_),
    .B(_14598_),
    .CI(_14599_),
    .CO(_14600_),
    .S(_14601_));
 FA_X1 _30101_ (.A(_14602_),
    .B(_14603_),
    .CI(_14604_),
    .CO(_14605_),
    .S(_14606_));
 FA_X1 _30102_ (.A(_14607_),
    .B(_14608_),
    .CI(_14609_),
    .CO(_14610_),
    .S(_14611_));
 FA_X1 _30103_ (.A(_14612_),
    .B(_14613_),
    .CI(_14614_),
    .CO(_14615_),
    .S(_14616_));
 FA_X1 _30104_ (.A(_14579_),
    .B(_14617_),
    .CI(_14611_),
    .CO(_14618_),
    .S(_14619_));
 FA_X1 _30105_ (.A(_14620_),
    .B(_14621_),
    .CI(_14622_),
    .CO(_14623_),
    .S(_14624_));
 FA_X1 _30106_ (.A(_14625_),
    .B(_14624_),
    .CI(_14592_),
    .CO(_14626_),
    .S(_14627_));
 FA_X1 _30107_ (.A(_14628_),
    .B(_14629_),
    .CI(_14630_),
    .CO(_14631_),
    .S(_14632_));
 FA_X1 _30108_ (.A(_14633_),
    .B(_14634_),
    .CI(_14635_),
    .CO(_14636_),
    .S(_14637_));
 FA_X1 _30109_ (.A(_14638_),
    .B(_14639_),
    .CI(_14637_),
    .CO(_14640_),
    .S(_14641_));
 FA_X1 _30110_ (.A(_14642_),
    .B(_14643_),
    .CI(_14644_),
    .CO(_14645_),
    .S(_14646_));
 FA_X1 _30111_ (.A(_14647_),
    .B(_14648_),
    .CI(_14649_),
    .CO(_14650_),
    .S(_14651_));
 FA_X1 _30112_ (.A(_14652_),
    .B(_14653_),
    .CI(_14654_),
    .CO(_14655_),
    .S(_14656_));
 FA_X1 _30113_ (.A(_14610_),
    .B(_14657_),
    .CI(_14651_),
    .CO(_14658_),
    .S(_14659_));
 FA_X1 _30114_ (.A(_14660_),
    .B(_14661_),
    .CI(_14662_),
    .CO(_14663_),
    .S(_14664_));
 FA_X1 _30115_ (.A(_14665_),
    .B(_14664_),
    .CI(_14623_),
    .CO(_14666_),
    .S(_14667_));
 FA_X1 _30116_ (.A(_14668_),
    .B(_14669_),
    .CI(_14670_),
    .CO(_14671_),
    .S(_14672_));
 FA_X1 _30117_ (.A(_14673_),
    .B(_14674_),
    .CI(_14675_),
    .CO(_14676_),
    .S(_14677_));
 FA_X1 _30118_ (.A(_14678_),
    .B(_14679_),
    .CI(_14631_),
    .CO(_14680_),
    .S(_14681_));
 FA_X1 _30119_ (.A(_14682_),
    .B(_14683_),
    .CI(_14684_),
    .CO(_14685_),
    .S(_14686_));
 FA_X1 _30120_ (.A(_14687_),
    .B(_14688_),
    .CI(_14689_),
    .CO(_14690_),
    .S(_14691_));
 FA_X1 _30121_ (.A(_14692_),
    .B(_14693_),
    .CI(_14694_),
    .CO(_14695_),
    .S(_14696_));
 FA_X1 _30122_ (.A(_14650_),
    .B(_14697_),
    .CI(_14691_),
    .CO(_14698_),
    .S(_14699_));
 FA_X1 _30123_ (.A(_14700_),
    .B(_14699_),
    .CI(_14658_),
    .CO(_14701_),
    .S(_14702_));
 FA_X1 _30124_ (.A(_14703_),
    .B(_14704_),
    .CI(_14705_),
    .CO(_14706_),
    .S(_14707_));
 FA_X1 _30125_ (.A(_14708_),
    .B(_14707_),
    .CI(_14663_),
    .CO(_14709_),
    .S(_14710_));
 FA_X1 _30126_ (.A(_14711_),
    .B(_14712_),
    .CI(_14713_),
    .CO(_14714_),
    .S(_14715_));
 FA_X1 _30127_ (.A(_14716_),
    .B(_14717_),
    .CI(_14718_),
    .CO(_14719_),
    .S(_14720_));
 FA_X1 _30128_ (.A(_14721_),
    .B(_14722_),
    .CI(_14671_),
    .CO(_14723_),
    .S(_14724_));
 FA_X1 _30129_ (.A(_14725_),
    .B(_14726_),
    .CI(_14727_),
    .CO(_14728_),
    .S(_14729_));
 FA_X1 _30130_ (.A(_14730_),
    .B(_14732_),
    .CI(_14731_),
    .CO(_14733_),
    .S(_14734_));
 FA_X1 _30131_ (.A(_14735_),
    .B(_14736_),
    .CI(_14737_),
    .CO(_14738_),
    .S(_14739_));
 FA_X1 _30132_ (.A(_14690_),
    .B(_14734_),
    .CI(_14740_),
    .CO(_14741_),
    .S(_14742_));
 FA_X1 _30133_ (.A(_14743_),
    .B(_14742_),
    .CI(_14698_),
    .CO(_14744_),
    .S(_14745_));
 FA_X1 _30134_ (.A(_14746_),
    .B(_14747_),
    .CI(_14748_),
    .CO(_14749_),
    .S(_14750_));
 FA_X1 _30135_ (.A(_14751_),
    .B(_14752_),
    .CI(_14753_),
    .CO(_14754_),
    .S(_14755_));
 FA_X1 _30136_ (.A(_14756_),
    .B(_14755_),
    .CI(_14706_),
    .CO(_14757_),
    .S(_14758_));
 FA_X1 _30137_ (.A(_14759_),
    .B(_14760_),
    .CI(_14761_),
    .CO(_14762_),
    .S(_14763_));
 FA_X1 _30138_ (.A(_14763_),
    .B(_14764_),
    .CI(_14750_),
    .CO(_14765_),
    .S(_14766_));
 FA_X1 _30139_ (.A(_14767_),
    .B(_14768_),
    .CI(_14714_),
    .CO(_14769_),
    .S(_14770_));
 FA_X1 _30140_ (.A(_14771_),
    .B(_14772_),
    .CI(_14773_),
    .CO(_14774_),
    .S(_14775_));
 FA_X1 _30141_ (.A(_14776_),
    .B(_14777_),
    .CI(_14778_),
    .CO(_14779_),
    .S(_14780_));
 FA_X1 _30142_ (.A(_14781_),
    .B(_14780_),
    .CI(_14728_),
    .CO(_14782_),
    .S(_14783_));
 FA_X1 _30143_ (.A(_14784_),
    .B(_14785_),
    .CI(_14786_),
    .CO(_14787_),
    .S(_14788_));
 FA_X1 _30144_ (.A(_14789_),
    .B(_14790_),
    .CI(_14791_),
    .CO(_14792_),
    .S(_14793_));
 FA_X1 _30145_ (.A(_14794_),
    .B(_14733_),
    .CI(_14788_),
    .CO(_14795_),
    .S(_14796_));
 FA_X1 _30146_ (.A(_14797_),
    .B(_14741_),
    .CI(_14796_),
    .CO(_14798_),
    .S(_14799_));
 FA_X1 _30147_ (.A(_14800_),
    .B(_14801_),
    .CI(_14802_),
    .CO(_14803_),
    .S(_14804_));
 FA_X1 _30148_ (.A(_14805_),
    .B(_14806_),
    .CI(_14807_),
    .CO(_14808_),
    .S(_14809_));
 FA_X1 _30149_ (.A(_14810_),
    .B(_14809_),
    .CI(_14754_),
    .CO(_14811_),
    .S(_14812_));
 FA_X1 _30150_ (.A(_14813_),
    .B(_14814_),
    .CI(_14815_),
    .CO(_14816_),
    .S(_14817_));
 FA_X1 _30151_ (.A(_14818_),
    .B(_14819_),
    .CI(_14820_),
    .CO(_14821_),
    .S(_14822_));
 FA_X1 _30152_ (.A(_14823_),
    .B(_14824_),
    .CI(_14822_),
    .CO(_14825_),
    .S(_14826_));
 FA_X1 _30153_ (.A(_14827_),
    .B(_14828_),
    .CI(_14829_),
    .CO(_14830_),
    .S(_14831_));
 FA_X1 _30154_ (.A(_14832_),
    .B(_14833_),
    .CI(_14834_),
    .CO(_14835_),
    .S(_14836_));
 FA_X1 _30155_ (.A(_14836_),
    .B(_14779_),
    .CI(_14837_),
    .CO(_14838_),
    .S(_14839_));
 FA_X1 _30156_ (.A(_14840_),
    .B(_14841_),
    .CI(_14842_),
    .CO(_14843_),
    .S(_14844_));
 FA_X1 _30157_ (.A(_14845_),
    .B(_14846_),
    .CI(_14847_),
    .CO(_14848_),
    .S(_14849_));
 FA_X1 _30158_ (.A(_14844_),
    .B(_14787_),
    .CI(_14850_),
    .CO(_14851_),
    .S(_14852_));
 FA_X1 _30159_ (.A(_14782_),
    .B(_14852_),
    .CI(_14795_),
    .CO(_14853_),
    .S(_14854_));
 FA_X1 _30160_ (.A(_14855_),
    .B(_14856_),
    .CI(_14857_),
    .CO(_14858_),
    .S(_14859_));
 FA_X1 _30161_ (.A(_14860_),
    .B(_14861_),
    .CI(_14862_),
    .CO(_14863_),
    .S(_14864_));
 FA_X1 _30162_ (.A(_14865_),
    .B(_14864_),
    .CI(_14808_),
    .CO(_14866_),
    .S(_14867_));
 FA_X1 _30163_ (.A(_14868_),
    .B(_14869_),
    .CI(_14870_),
    .CO(_14871_),
    .S(_14872_));
 FA_X1 _30164_ (.A(_14873_),
    .B(_14874_),
    .CI(_14875_),
    .CO(_14876_),
    .S(_14877_));
 FA_X1 _30165_ (.A(_14821_),
    .B(_14878_),
    .CI(_14877_),
    .CO(_14879_),
    .S(_14880_));
 FA_X1 _30166_ (.A(_14881_),
    .B(_14882_),
    .CI(_14883_),
    .CO(_14884_),
    .S(_14885_));
 FA_X1 _30167_ (.A(_14886_),
    .B(_14887_),
    .CI(_14888_),
    .CO(_14889_),
    .S(_14890_));
 FA_X1 _30168_ (.A(_14890_),
    .B(_14835_),
    .CI(_14830_),
    .CO(_14891_),
    .S(_14892_));
 FA_X1 _30169_ (.A(_14893_),
    .B(_14894_),
    .CI(_14895_),
    .CO(_14896_),
    .S(_14897_));
 FA_X1 _30170_ (.A(_14898_),
    .B(_14899_),
    .CI(_14900_),
    .CO(_14901_),
    .S(_14902_));
 FA_X1 _30171_ (.A(_14903_),
    .B(_14904_),
    .CI(_14905_),
    .CO(_14906_),
    .S(_14907_));
 FA_X1 _30172_ (.A(_14908_),
    .B(_14902_),
    .CI(_14843_),
    .CO(_14909_),
    .S(_14910_));
 FA_X1 _30173_ (.A(_14838_),
    .B(_14910_),
    .CI(_14851_),
    .CO(_14911_),
    .S(_14912_));
 FA_X1 _30174_ (.A(_14897_),
    .B(_14913_),
    .CI(_14914_),
    .CO(_14915_),
    .S(_14916_));
 FA_X1 _30175_ (.A(_14917_),
    .B(_14918_),
    .CI(_14919_),
    .CO(_14920_),
    .S(_14921_));
 FA_X1 _30176_ (.A(_14922_),
    .B(_14921_),
    .CI(_14863_),
    .CO(_14923_),
    .S(_14924_));
 FA_X1 _30177_ (.A(_14925_),
    .B(_14926_),
    .CI(_14927_),
    .CO(_14928_),
    .S(_14929_));
 FA_X1 _30178_ (.A(_14930_),
    .B(_14931_),
    .CI(_14932_),
    .CO(_14933_),
    .S(_14934_));
 FA_X1 _30179_ (.A(_14934_),
    .B(_14876_),
    .CI(_14935_),
    .CO(_14936_),
    .S(_14937_));
 FA_X1 _30180_ (.A(_14938_),
    .B(_14939_),
    .CI(_14940_),
    .CO(_14941_),
    .S(_14942_));
 FA_X1 _30181_ (.A(_14943_),
    .B(_14944_),
    .CI(_14945_),
    .CO(_14946_),
    .S(_14947_));
 FA_X1 _30182_ (.A(_14947_),
    .B(_14948_),
    .CI(_14949_),
    .CO(_14950_),
    .S(_14951_));
 FA_X1 _30183_ (.A(_14952_),
    .B(_14953_),
    .CI(_14954_),
    .CO(_14955_),
    .S(_14956_));
 FA_X1 _30184_ (.A(_14956_),
    .B(_14889_),
    .CI(_14957_),
    .CO(_14958_),
    .S(_14959_));
 FA_X1 _30185_ (.A(_14960_),
    .B(_14961_),
    .CI(_14951_),
    .CO(_14962_),
    .S(_14963_));
 FA_X1 _30186_ (.A(_14964_),
    .B(_14965_),
    .CI(_14966_),
    .CO(_14967_),
    .S(_14968_));
 FA_X1 _30187_ (.A(_14969_),
    .B(_14970_),
    .CI(_14971_),
    .CO(_14972_),
    .S(_14973_));
 FA_X1 _30188_ (.A(_14901_),
    .B(_14974_),
    .CI(_14968_),
    .CO(_14975_),
    .S(_14976_));
 FA_X1 _30189_ (.A(_14891_),
    .B(_14976_),
    .CI(_14909_),
    .CO(_14977_),
    .S(_14978_));
 FA_X1 _30190_ (.A(_14979_),
    .B(_14978_),
    .CI(_14980_),
    .CO(_14981_),
    .S(_14982_));
 FA_X1 _30191_ (.A(_14983_),
    .B(_14984_),
    .CI(_14985_),
    .CO(_14986_),
    .S(_14987_));
 FA_X1 _30192_ (.A(_14988_),
    .B(_14920_),
    .CI(_14989_),
    .CO(_14990_),
    .S(_14991_));
 FA_X1 _30193_ (.A(_14992_),
    .B(_14993_),
    .CI(_14994_),
    .CO(_14995_),
    .S(_14996_));
 FA_X1 _30194_ (.A(_14997_),
    .B(_14998_),
    .CI(_14996_),
    .CO(_14999_),
    .S(_15000_));
 FA_X1 _30195_ (.A(_15001_),
    .B(_15002_),
    .CI(_14982_),
    .CO(_15003_),
    .S(_15004_));
 FA_X1 _30196_ (.A(_14933_),
    .B(_15005_),
    .CI(_15004_),
    .CO(_15006_),
    .S(_15007_));
 FA_X1 _30197_ (.A(_15008_),
    .B(_15009_),
    .CI(_15010_),
    .CO(_15011_),
    .S(_15012_));
 FA_X1 _30198_ (.A(_15013_),
    .B(_15014_),
    .CI(_15015_),
    .CO(_15016_),
    .S(_15017_));
 FA_X1 _30199_ (.A(_15012_),
    .B(_14941_),
    .CI(_15018_),
    .CO(_15019_),
    .S(_15020_));
 FA_X1 _30200_ (.A(_15021_),
    .B(_15022_),
    .CI(_15023_),
    .CO(_15024_),
    .S(_15025_));
 FA_X1 _30201_ (.A(_15025_),
    .B(_14955_),
    .CI(_15026_),
    .CO(_15027_),
    .S(_15028_));
 FA_X1 _30202_ (.A(_15028_),
    .B(_15020_),
    .CI(_15029_),
    .CO(_15030_),
    .S(_15031_));
 FA_X1 _30203_ (.A(_15032_),
    .B(_15033_),
    .CI(_15034_),
    .CO(_15035_),
    .S(_15036_));
 FA_X1 _30204_ (.A(_15037_),
    .B(_15038_),
    .CI(_15039_),
    .CO(_15040_),
    .S(_15041_));
 FA_X1 _30205_ (.A(_15036_),
    .B(_14967_),
    .CI(_15042_),
    .CO(_15043_),
    .S(_15044_));
 FA_X1 _30206_ (.A(_14958_),
    .B(_15044_),
    .CI(_14975_),
    .CO(_15045_),
    .S(_15046_));
 FA_X1 _30207_ (.A(_15031_),
    .B(_15047_),
    .CI(_15046_),
    .CO(_15048_),
    .S(_15049_));
 FA_X1 _30208_ (.A(_15050_),
    .B(_14983_),
    .CI(_15051_),
    .CO(_15052_),
    .S(_15053_));
 FA_X1 _30209_ (.A(_15054_),
    .B(_15055_),
    .CI(_15056_),
    .CO(_15057_),
    .S(_15058_));
 FA_X1 _30210_ (.A(_14977_),
    .B(_15059_),
    .CI(_15060_),
    .CO(_15061_),
    .S(_15062_));
 FA_X1 _30211_ (.A(_15049_),
    .B(_14981_),
    .CI(_15062_),
    .CO(_15063_),
    .S(_15064_));
 FA_X1 _30212_ (.A(_15064_),
    .B(_15003_),
    .CI(_15065_),
    .CO(_15066_),
    .S(_15067_));
 FA_X1 _30213_ (.A(_15068_),
    .B(_15069_),
    .CI(_15070_),
    .CO(_15071_),
    .S(_15072_));
 FA_X1 _30214_ (.A(_15073_),
    .B(_15074_),
    .CI(_15075_),
    .CO(_15076_),
    .S(_15077_));
 FA_X1 _30215_ (.A(_15078_),
    .B(_15072_),
    .CI(_15011_),
    .CO(_15079_),
    .S(_15080_));
 FA_X1 _30216_ (.A(_15081_),
    .B(_15082_),
    .CI(_15083_),
    .CO(_15084_),
    .S(_15085_));
 FA_X1 _30217_ (.A(_15085_),
    .B(_15024_),
    .CI(_15086_),
    .CO(_15087_),
    .S(_15088_));
 FA_X1 _30218_ (.A(_15080_),
    .B(_15019_),
    .CI(_15088_),
    .CO(_15089_),
    .S(_15090_));
 FA_X1 _30219_ (.A(_15091_),
    .B(_15092_),
    .CI(_15093_),
    .CO(_15094_),
    .S(_15095_));
 FA_X1 _30220_ (.A(_15096_),
    .B(_15097_),
    .CI(_15098_),
    .CO(_15099_),
    .S(_15100_));
 FA_X1 _30221_ (.A(_15101_),
    .B(_15095_),
    .CI(_15035_),
    .CO(_15102_),
    .S(_15103_));
 FA_X1 _30222_ (.A(_15103_),
    .B(_15043_),
    .CI(_15027_),
    .CO(_15104_),
    .S(_15105_));
 FA_X1 _30223_ (.A(_15090_),
    .B(_15030_),
    .CI(_15105_),
    .CO(_15106_),
    .S(_15107_));
 FA_X1 _30224_ (.A(_15050_),
    .B(_15108_),
    .CI(_14983_),
    .CO(_15109_),
    .S(_15110_));
 FA_X1 _30225_ (.A(_15111_),
    .B(_15112_),
    .CI(_15113_),
    .CO(_15114_),
    .S(_15115_));
 FA_X1 _30226_ (.A(_15116_),
    .B(_15117_),
    .CI(_15118_),
    .CO(_15119_),
    .S(_15120_));
 FA_X1 _30227_ (.A(_15107_),
    .B(_15121_),
    .CI(_15048_),
    .CO(_15122_),
    .S(_15123_));
 FA_X1 _30228_ (.A(_15123_),
    .B(_15063_),
    .CI(_15061_),
    .CO(_15124_),
    .S(_15125_));
 FA_X1 _30229_ (.A(_15126_),
    .B(_15127_),
    .CI(_15128_),
    .CO(_15129_),
    .S(_15130_));
 FA_X1 _30230_ (.A(_15131_),
    .B(_15132_),
    .CI(_15133_),
    .CO(_15134_),
    .S(_15135_));
 FA_X1 _30231_ (.A(_15136_),
    .B(_15130_),
    .CI(_15071_),
    .CO(_15137_),
    .S(_15138_));
 FA_X1 _30232_ (.A(_15139_),
    .B(_15140_),
    .CI(_15141_),
    .CO(_15142_),
    .S(_15143_));
 FA_X1 _30233_ (.A(_15143_),
    .B(_15084_),
    .CI(_15144_),
    .CO(_15145_),
    .S(_15146_));
 FA_X1 _30234_ (.A(_15138_),
    .B(_15079_),
    .CI(_15146_),
    .CO(_15147_),
    .S(_15148_));
 FA_X1 _30235_ (.A(_15149_),
    .B(_15150_),
    .CI(_15151_),
    .CO(_15152_),
    .S(_15153_));
 FA_X1 _30236_ (.A(_15154_),
    .B(_15155_),
    .CI(_15156_),
    .CO(_15157_),
    .S(_15158_));
 FA_X1 _30237_ (.A(_15153_),
    .B(_15158_),
    .CI(_15094_),
    .CO(_15159_),
    .S(_15160_));
 FA_X1 _30238_ (.A(_15160_),
    .B(_15102_),
    .CI(_15087_),
    .CO(_15161_),
    .S(_15162_));
 FA_X1 _30239_ (.A(_15162_),
    .B(_15148_),
    .CI(_15089_),
    .CO(_15163_),
    .S(_15164_));
 FA_X1 _30240_ (.A(_15050_),
    .B(_14983_),
    .CI(_15165_),
    .CO(_15166_),
    .S(_15167_));
 FA_X1 _30241_ (.A(_15168_),
    .B(_15169_),
    .CI(_15170_),
    .CO(_15171_),
    .S(_15172_));
 FA_X1 _30242_ (.A(_15173_),
    .B(_15174_),
    .CI(_15175_),
    .CO(_15176_),
    .S(_15177_));
 FA_X1 _30243_ (.A(_15106_),
    .B(_15178_),
    .CI(_15164_),
    .CO(_15179_),
    .S(_15180_));
 FA_X1 _30244_ (.A(_15122_),
    .B(_15181_),
    .CI(_15180_),
    .CO(_15182_),
    .S(_15183_));
 FA_X1 _30245_ (.A(_15184_),
    .B(_15185_),
    .CI(_15186_),
    .CO(_15187_),
    .S(_15188_));
 FA_X1 _30246_ (.A(_15189_),
    .B(_15190_),
    .CI(_15191_),
    .CO(_15192_),
    .S(_15193_));
 FA_X1 _30247_ (.A(_15188_),
    .B(_15129_),
    .CI(_15194_),
    .CO(_15195_),
    .S(_15196_));
 FA_X1 _30248_ (.A(_15197_),
    .B(_15198_),
    .CI(_15199_),
    .CO(_15200_),
    .S(_15201_));
 FA_X1 _30249_ (.A(_15201_),
    .B(_15142_),
    .CI(_15202_),
    .CO(_15203_),
    .S(_15204_));
 FA_X1 _30250_ (.A(_15204_),
    .B(_15196_),
    .CI(_15137_),
    .CO(_15205_),
    .S(_15206_));
 FA_X1 _30251_ (.A(_15207_),
    .B(_15208_),
    .CI(_15209_),
    .CO(_15210_),
    .S(_15211_));
 FA_X1 _30252_ (.A(_15212_),
    .B(_15098_),
    .CI(_15213_),
    .CO(_15214_),
    .S(_15215_));
 FA_X1 _30253_ (.A(_15211_),
    .B(_15152_),
    .CI(_15216_),
    .CO(_15217_),
    .S(_15218_));
 FA_X1 _30254_ (.A(_15218_),
    .B(_15159_),
    .CI(_15145_),
    .CO(_15219_),
    .S(_15220_));
 FA_X1 _30255_ (.A(_15206_),
    .B(_15147_),
    .CI(_15220_),
    .CO(_15221_),
    .S(_15222_));
 FA_X1 _30256_ (.A(_15050_),
    .B(_15223_),
    .CI(net326),
    .CO(_15224_),
    .S(_15225_));
 FA_X1 _30257_ (.A(_15157_),
    .B(_15226_),
    .CI(_15227_),
    .CO(_15228_),
    .S(_15229_));
 FA_X1 _30258_ (.A(_15230_),
    .B(_15231_),
    .CI(_15232_),
    .CO(_15233_),
    .S(_15234_));
 FA_X1 _30259_ (.A(_15222_),
    .B(_15163_),
    .CI(_15235_),
    .CO(_15236_),
    .S(_15237_));
 FA_X1 _30260_ (.A(_15237_),
    .B(_15179_),
    .CI(_15238_),
    .CO(_15239_),
    .S(_15240_));
 FA_X1 _30261_ (.A(_15241_),
    .B(_15242_),
    .CI(_15243_),
    .CO(_15244_),
    .S(_15245_));
 FA_X1 _30262_ (.A(_15246_),
    .B(_15247_),
    .CI(_15248_),
    .CO(_15249_),
    .S(_15250_));
 FA_X1 _30263_ (.A(_15187_),
    .B(_15251_),
    .CI(_15245_),
    .CO(_15252_),
    .S(_15253_));
 FA_X1 _30264_ (.A(_15254_),
    .B(_15255_),
    .CI(_15256_),
    .CO(_15257_),
    .S(_15258_));
 FA_X1 _30265_ (.A(_15258_),
    .B(_15200_),
    .CI(_15259_),
    .CO(_15260_),
    .S(_15261_));
 FA_X1 _30266_ (.A(_15261_),
    .B(_15253_),
    .CI(_15195_),
    .CO(_15262_),
    .S(_15263_));
 FA_X1 _30267_ (.A(_15264_),
    .B(_15265_),
    .CI(_15266_),
    .CO(_15267_),
    .S(_15268_));
 FA_X1 _30268_ (.A(_15210_),
    .B(_15216_),
    .CI(_15268_),
    .CO(_15269_),
    .S(_15270_));
 FA_X1 _30269_ (.A(_15203_),
    .B(_15270_),
    .CI(_15217_),
    .CO(_15271_),
    .S(_15272_));
 FA_X1 _30270_ (.A(_15205_),
    .B(_15272_),
    .CI(_15263_),
    .CO(_15273_),
    .S(_15274_));
 FA_X1 _30271_ (.A(_15050_),
    .B(net326),
    .CI(_15275_),
    .CO(_15276_),
    .S(_15277_));
 FA_X1 _30272_ (.A(_15278_),
    .B(_15279_),
    .CI(_15280_),
    .CO(_15281_),
    .S(_15282_));
 FA_X1 _30273_ (.A(_15283_),
    .B(_15284_),
    .CI(_15285_),
    .CO(_15286_),
    .S(_15287_));
 FA_X1 _30274_ (.A(_15274_),
    .B(_15221_),
    .CI(_15288_),
    .CO(_15289_),
    .S(_15290_));
 FA_X1 _30275_ (.A(_15290_),
    .B(_15236_),
    .CI(_15291_),
    .CO(_15292_),
    .S(_15293_));
 FA_X1 _30276_ (.A(_15294_),
    .B(_15295_),
    .CI(_15296_),
    .CO(_15297_),
    .S(_15298_));
 FA_X1 _30277_ (.A(_15299_),
    .B(_15300_),
    .CI(_15301_),
    .CO(_15302_),
    .S(_15303_));
 FA_X1 _30278_ (.A(_15304_),
    .B(_15298_),
    .CI(_15244_),
    .CO(_15305_),
    .S(_15306_));
 FA_X1 _30279_ (.A(_15307_),
    .B(_15308_),
    .CI(_15309_),
    .CO(_15310_),
    .S(_15311_));
 FA_X1 _30280_ (.A(_15311_),
    .B(_15257_),
    .CI(_15312_),
    .CO(_15313_),
    .S(_15314_));
 FA_X1 _30281_ (.A(_15306_),
    .B(_15252_),
    .CI(_15314_),
    .CO(_15315_),
    .S(_15316_));
 FA_X1 _30282_ (.A(_15264_),
    .B(_15317_),
    .CI(_15318_),
    .CO(_15319_),
    .S(_15320_));
 FA_X1 _30283_ (.A(_15215_),
    .B(_15321_),
    .CI(_15322_),
    .CO(_15323_),
    .S(_15324_));
 FA_X1 _30284_ (.A(_15325_),
    .B(_15269_),
    .CI(_15260_),
    .CO(_15326_),
    .S(_15327_));
 FA_X1 _30285_ (.A(_15327_),
    .B(_15262_),
    .CI(_15316_),
    .CO(_15328_),
    .S(_15329_));
 FA_X1 _30286_ (.A(_15050_),
    .B(_15330_),
    .CI(net326),
    .CO(_15331_),
    .S(_15332_));
 FA_X1 _30287_ (.A(_15333_),
    .B(_15279_),
    .CI(_15334_),
    .CO(_15335_),
    .S(_15336_));
 FA_X1 _30288_ (.A(_15337_),
    .B(_15338_),
    .CI(_15339_),
    .CO(_15340_),
    .S(_15341_));
 FA_X1 _30289_ (.A(_15273_),
    .B(_15329_),
    .CI(_15342_),
    .CO(_15343_),
    .S(_15344_));
 FA_X1 _30290_ (.A(_15344_),
    .B(_15289_),
    .CI(_15345_),
    .CO(_15346_),
    .S(_15347_));
 FA_X1 _30291_ (.A(_15348_),
    .B(_15349_),
    .CI(_15350_),
    .CO(_15351_),
    .S(_15352_));
 FA_X1 _30292_ (.A(_15353_),
    .B(_15354_),
    .CI(_15355_),
    .CO(_15356_),
    .S(_15357_));
 FA_X1 _30293_ (.A(_15352_),
    .B(_15297_),
    .CI(_15357_),
    .CO(_15358_),
    .S(_15359_));
 FA_X1 _30294_ (.A(_15360_),
    .B(_15361_),
    .CI(_15362_),
    .CO(_15363_),
    .S(_15364_));
 FA_X1 _30295_ (.A(_15364_),
    .B(_15310_),
    .CI(_15365_),
    .CO(_15366_),
    .S(_15367_));
 FA_X1 _30296_ (.A(_15367_),
    .B(_15359_),
    .CI(_15305_),
    .CO(_15368_),
    .S(_15369_));
 FA_X1 _30297_ (.A(_15370_),
    .B(_15371_),
    .CI(_15372_),
    .CO(_15373_),
    .S(_15374_));
 FA_X1 _30298_ (.A(_15216_),
    .B(_15375_),
    .CI(_15319_),
    .CO(_15376_),
    .S(_15377_));
 FA_X1 _30299_ (.A(_15377_),
    .B(_15378_),
    .CI(_15313_),
    .CO(_15379_),
    .S(_15380_));
 FA_X1 _30300_ (.A(_15369_),
    .B(_15315_),
    .CI(_15380_),
    .CO(_15381_),
    .S(_15382_));
 FA_X1 _30301_ (.A(_15050_),
    .B(net326),
    .CI(_15383_),
    .CO(_15384_),
    .S(_15385_));
 FA_X1 _30302_ (.A(_15279_),
    .B(_15386_),
    .CI(_15387_),
    .CO(_15388_),
    .S(_15389_));
 FA_X1 _30303_ (.A(_15390_),
    .B(_15391_),
    .CI(_15392_),
    .CO(_15393_),
    .S(_15394_));
 FA_X1 _30304_ (.A(_15382_),
    .B(_15395_),
    .CI(_15328_),
    .CO(_15396_),
    .S(_15397_));
 FA_X1 _30305_ (.A(_15397_),
    .B(_15343_),
    .CI(_15398_),
    .CO(_15399_),
    .S(_15400_));
 FA_X1 _30306_ (.A(_15401_),
    .B(_15402_),
    .CI(_15403_),
    .CO(_15404_),
    .S(_15405_));
 FA_X1 _30307_ (.A(_15406_),
    .B(_15407_),
    .CI(_15408_),
    .CO(_15409_),
    .S(_15410_));
 FA_X1 _30308_ (.A(_15351_),
    .B(_15410_),
    .CI(_15405_),
    .CO(_15411_),
    .S(_15412_));
 FA_X1 _30309_ (.A(_15413_),
    .B(_15414_),
    .CI(_15415_),
    .CO(_15416_),
    .S(_15417_));
 FA_X1 _30310_ (.A(_15417_),
    .B(_15363_),
    .CI(_15356_),
    .CO(_15418_),
    .S(_15419_));
 FA_X1 _30311_ (.A(_15419_),
    .B(_15412_),
    .CI(_15358_),
    .CO(_15420_),
    .S(_15421_));
 FA_X1 _30312_ (.A(_15215_),
    .B(_15374_),
    .CI(_15373_),
    .CO(_15422_),
    .S(_15423_));
 FA_X1 _30313_ (.A(_15366_),
    .B(_15424_),
    .CI(_15376_),
    .CO(_15425_),
    .S(_15426_));
 FA_X1 _30314_ (.A(_15368_),
    .B(_15426_),
    .CI(_15421_),
    .CO(_15427_),
    .S(_15428_));
 FA_X1 _30315_ (.A(_15050_),
    .B(net327),
    .CI(_15429_),
    .CO(_15430_),
    .S(_15431_));
 FA_X1 _30316_ (.A(_15432_),
    .B(_15279_),
    .CI(_15433_),
    .CO(_15434_),
    .S(_15435_));
 FA_X1 _30317_ (.A(_15436_),
    .B(_15437_),
    .CI(_15438_),
    .CO(_15439_),
    .S(_15440_));
 FA_X1 _30318_ (.A(_15428_),
    .B(_15441_),
    .CI(_15381_),
    .CO(_15442_),
    .S(_15443_));
 FA_X1 _30319_ (.A(_15443_),
    .B(_15396_),
    .CI(_15444_),
    .CO(_15445_),
    .S(_15446_));
 FA_X1 _30320_ (.A(_15447_),
    .B(_15448_),
    .CI(_15449_),
    .CO(_15450_),
    .S(_15451_));
 FA_X1 _30321_ (.A(_15452_),
    .B(_15453_),
    .CI(_15454_),
    .CO(_15455_),
    .S(_15456_));
 FA_X1 _30322_ (.A(_15456_),
    .B(_15451_),
    .CI(_15404_),
    .CO(_15457_),
    .S(_15458_));
 FA_X1 _30323_ (.A(_15459_),
    .B(_15415_),
    .CI(_15460_),
    .CO(_15461_),
    .S(_15462_));
 FA_X1 _30324_ (.A(_15409_),
    .B(_15462_),
    .CI(_15416_),
    .CO(_15463_),
    .S(_15464_));
 FA_X1 _30325_ (.A(_15458_),
    .B(_15464_),
    .CI(_15411_),
    .CO(_15465_),
    .S(_15466_));
 FA_X1 _30326_ (.A(_15418_),
    .B(_15467_),
    .CI(_15424_),
    .CO(_15468_),
    .S(_15469_));
 FA_X1 _30327_ (.A(_15420_),
    .B(_15469_),
    .CI(_15466_),
    .CO(_15470_),
    .S(_15471_));
 FA_X1 _30328_ (.A(_15050_),
    .B(net315),
    .CI(_15472_),
    .CO(_15473_),
    .S(_15474_));
 FA_X1 _30329_ (.A(_15475_),
    .B(_15279_),
    .CI(_15476_),
    .CO(_15477_),
    .S(_15478_));
 FA_X1 _30330_ (.A(_15479_),
    .B(_15480_),
    .CI(_15481_),
    .CO(_15482_),
    .S(_15483_));
 FA_X1 _30331_ (.A(_15471_),
    .B(_15484_),
    .CI(_15427_),
    .CO(_15485_),
    .S(_15486_));
 FA_X1 _30332_ (.A(_15486_),
    .B(_15442_),
    .CI(_15487_),
    .CO(_15488_),
    .S(_15489_));
 FA_X1 _30333_ (.A(_15490_),
    .B(_15491_),
    .CI(_15492_),
    .CO(_15493_),
    .S(_15494_));
 FA_X1 _30334_ (.A(_15495_),
    .B(_15496_),
    .CI(_15497_),
    .CO(_15498_),
    .S(_15499_));
 FA_X1 _30335_ (.A(_15499_),
    .B(_15450_),
    .CI(_15494_),
    .CO(_15500_),
    .S(_15501_));
 FA_X1 _30336_ (.A(_15502_),
    .B(_15503_),
    .CI(_15504_),
    .CO(_15505_),
    .S(_15506_));
 FA_X1 _30337_ (.A(_15461_),
    .B(_15455_),
    .CI(_15507_),
    .CO(_15508_),
    .S(_15509_));
 FA_X1 _30338_ (.A(_15457_),
    .B(_15501_),
    .CI(_15509_),
    .CO(_15510_),
    .S(_15511_));
 FA_X1 _30339_ (.A(_15463_),
    .B(_15467_),
    .CI(_15424_),
    .CO(_15512_),
    .S(_15513_));
 FA_X1 _30340_ (.A(_15465_),
    .B(_15511_),
    .CI(_15513_),
    .CO(_15514_),
    .S(_15515_));
 FA_X1 _30341_ (.A(_15050_),
    .B(net315),
    .CI(_15516_),
    .CO(_15517_),
    .S(_15518_));
 FA_X1 _30342_ (.A(_15519_),
    .B(_15279_),
    .CI(_15520_),
    .CO(_15521_),
    .S(_15522_));
 FA_X1 _30343_ (.A(_15523_),
    .B(_15524_),
    .CI(_15525_),
    .CO(_15526_),
    .S(_15527_));
 FA_X1 _30344_ (.A(_15470_),
    .B(_15515_),
    .CI(_15528_),
    .CO(_15529_),
    .S(_15530_));
 FA_X1 _30345_ (.A(_15485_),
    .B(_15531_),
    .CI(_15530_),
    .CO(_15532_),
    .S(_15533_));
 FA_X1 _30346_ (.A(_15534_),
    .B(_15535_),
    .CI(_15536_),
    .CO(_15537_),
    .S(_15538_));
 FA_X1 _30347_ (.A(_15539_),
    .B(_15540_),
    .CI(_15541_),
    .CO(_15542_),
    .S(_15543_));
 FA_X1 _30348_ (.A(_15538_),
    .B(_15543_),
    .CI(_15493_),
    .CO(_15544_),
    .S(_15545_));
 FA_X1 _30349_ (.A(_15498_),
    .B(_15546_),
    .CI(_15507_),
    .CO(_15547_),
    .S(_15548_));
 FA_X1 _30350_ (.A(_15548_),
    .B(_15545_),
    .CI(_15500_),
    .CO(_15549_),
    .S(_15550_));
 FA_X1 _30351_ (.A(_15467_),
    .B(_15508_),
    .CI(_15424_),
    .CO(_15551_),
    .S(_15552_));
 FA_X1 _30352_ (.A(_15552_),
    .B(_15510_),
    .CI(_15550_),
    .CO(_15553_),
    .S(_15554_));
 FA_X1 _30353_ (.A(_15050_),
    .B(net315),
    .CI(_15555_),
    .CO(_15556_),
    .S(_15557_));
 FA_X1 _30354_ (.A(_15558_),
    .B(_15279_),
    .CI(_15559_),
    .CO(_15560_),
    .S(_15561_));
 FA_X1 _30355_ (.A(_15562_),
    .B(_15563_),
    .CI(_15564_),
    .CO(_15565_),
    .S(_15566_));
 FA_X1 _30356_ (.A(_15567_),
    .B(_15514_),
    .CI(_15554_),
    .CO(_15568_),
    .S(_15569_));
 FA_X1 _30357_ (.A(_15529_),
    .B(_15570_),
    .CI(_15569_),
    .CO(_15571_),
    .S(_15572_));
 FA_X1 _30358_ (.A(_15573_),
    .B(_15574_),
    .CI(_15575_),
    .CO(_15576_),
    .S(_15577_));
 FA_X1 _30359_ (.A(_15578_),
    .B(_15579_),
    .CI(_15541_),
    .CO(_15580_),
    .S(_15581_));
 FA_X1 _30360_ (.A(_15537_),
    .B(_15581_),
    .CI(_15577_),
    .CO(_15582_),
    .S(_15583_));
 FA_X1 _30361_ (.A(_15546_),
    .B(_15542_),
    .CI(_15507_),
    .CO(_15584_),
    .S(_15585_));
 FA_X1 _30362_ (.A(_15585_),
    .B(_15544_),
    .CI(_15583_),
    .CO(_15586_),
    .S(_15587_));
 FA_X1 _30363_ (.A(_15467_),
    .B(_15547_),
    .CI(_15424_),
    .CO(_15588_),
    .S(_15589_));
 FA_X1 _30364_ (.A(_15589_),
    .B(_15549_),
    .CI(_15587_),
    .CO(_15590_),
    .S(_15591_));
 FA_X1 _30365_ (.A(_15592_),
    .B(_15050_),
    .CI(net315),
    .CO(_15593_),
    .S(_15594_));
 FA_X1 _30366_ (.A(_15595_),
    .B(_15279_),
    .CI(_15596_),
    .CO(_15597_),
    .S(_15598_));
 FA_X1 _30367_ (.A(_15599_),
    .B(_15600_),
    .CI(_15601_),
    .CO(_15602_),
    .S(_15603_));
 FA_X1 _30368_ (.A(_15553_),
    .B(_15591_),
    .CI(_15604_),
    .CO(_15605_),
    .S(_15606_));
 FA_X1 _30369_ (.A(_15606_),
    .B(_15568_),
    .CI(_15607_),
    .CO(_15608_),
    .S(_15609_));
 FA_X1 _30370_ (.A(_15610_),
    .B(_15611_),
    .CI(_15612_),
    .CO(_15613_),
    .S(_15614_));
 FA_X1 _30371_ (.A(_15615_),
    .B(_15616_),
    .CI(_15617_),
    .CO(_15618_),
    .S(_15619_));
 FA_X1 _30372_ (.A(_15614_),
    .B(_15576_),
    .CI(_15620_),
    .CO(_15621_),
    .S(_15622_));
 FA_X1 _30373_ (.A(_15546_),
    .B(_15580_),
    .CI(_15507_),
    .CO(_15623_),
    .S(_15624_));
 FA_X1 _30374_ (.A(_15582_),
    .B(_15624_),
    .CI(_15622_),
    .CO(_15625_),
    .S(_15626_));
 FA_X1 _30375_ (.A(_15584_),
    .B(_15467_),
    .CI(_15424_),
    .CO(_15627_),
    .S(_15628_));
 FA_X1 _30376_ (.A(_15586_),
    .B(_15628_),
    .CI(_15626_),
    .CO(_15629_),
    .S(_15630_));
 FA_X1 _30377_ (.A(_15050_),
    .B(net315),
    .CI(_15631_),
    .CO(_15632_),
    .S(_15633_));
 FA_X1 _30378_ (.A(_15634_),
    .B(_15635_),
    .CI(_15279_),
    .CO(_15636_),
    .S(_15637_));
 FA_X1 _30379_ (.A(_15638_),
    .B(_15639_),
    .CI(_15640_),
    .CO(_15641_),
    .S(_15642_));
 FA_X1 _30380_ (.A(_15630_),
    .B(_15643_),
    .CI(_15590_),
    .CO(_15644_),
    .S(_15645_));
 FA_X1 _30381_ (.A(_15645_),
    .B(_15605_),
    .CI(_15646_),
    .CO(_15647_),
    .S(_15648_));
 FA_X1 _30382_ (.A(_15649_),
    .B(_15650_),
    .CI(_15651_),
    .CO(_15652_),
    .S(_15653_));
 FA_X1 _30383_ (.A(_15619_),
    .B(_15654_),
    .CI(_15655_),
    .CO(_15656_),
    .S(_15657_));
 FA_X1 _30384_ (.A(_15546_),
    .B(_15658_),
    .CI(_15507_),
    .CO(_15659_),
    .S(_15660_));
 FA_X1 _30385_ (.A(_15660_),
    .B(_15661_),
    .CI(_15621_),
    .CO(_15662_),
    .S(_15663_));
 FA_X1 _30386_ (.A(_15423_),
    .B(_15664_),
    .CI(_15422_),
    .CO(_15665_),
    .S(_15666_));
 FA_X1 _30387_ (.A(_15663_),
    .B(_15625_),
    .CI(_15667_),
    .CO(_15668_),
    .S(_15669_));
 FA_X1 _30388_ (.A(_15050_),
    .B(net315),
    .CI(_15670_),
    .CO(_15671_),
    .S(_15672_));
 FA_X1 _30389_ (.A(_15673_),
    .B(_15279_),
    .CI(_15674_),
    .CO(_15675_),
    .S(_15676_));
 FA_X1 _30390_ (.A(_15677_),
    .B(_15678_),
    .CI(_15679_),
    .CO(_15680_),
    .S(_15681_));
 FA_X1 _30391_ (.A(_15669_),
    .B(_15682_),
    .CI(_15629_),
    .CO(_15683_),
    .S(_15684_));
 FA_X1 _30392_ (.A(_15684_),
    .B(_15644_),
    .CI(_15685_),
    .CO(_15686_),
    .S(_15687_));
 FA_X1 _30393_ (.A(_15688_),
    .B(_15689_),
    .CI(_15651_),
    .CO(_15690_),
    .S(_15691_));
 FA_X1 _30394_ (.A(_15619_),
    .B(_15692_),
    .CI(_15693_),
    .CO(_15694_),
    .S(_15695_));
 FA_X1 _30395_ (.A(_15660_),
    .B(_15696_),
    .CI(_15697_),
    .CO(_15698_),
    .S(_15699_));
 FA_X1 _30396_ (.A(_15700_),
    .B(_15422_),
    .CI(_15423_),
    .CO(_15701_),
    .S(_15702_));
 FA_X1 _30397_ (.A(_15699_),
    .B(_15662_),
    .CI(_15703_),
    .CO(_15704_),
    .S(_15705_));
 FA_X1 _30398_ (.A(_15706_),
    .B(_15050_),
    .CI(net315),
    .CO(_15707_),
    .S(_15708_));
 FA_X1 _30399_ (.A(_15709_),
    .B(_15710_),
    .CI(_15279_),
    .CO(_15711_),
    .S(_15712_));
 FA_X1 _30400_ (.A(_15713_),
    .B(_15665_),
    .CI(_15714_),
    .CO(_15715_),
    .S(_15716_));
 FA_X1 _30401_ (.A(_15705_),
    .B(_15668_),
    .CI(_15717_),
    .CO(_15718_),
    .S(_15719_));
 FA_X1 _30402_ (.A(_15720_),
    .B(_15719_),
    .CI(_15683_),
    .CO(_15721_),
    .S(_15722_));
 FA_X1 _30403_ (.A(_15688_),
    .B(_15723_),
    .CI(_15651_),
    .CO(_15724_),
    .S(_15725_));
 FA_X1 _30404_ (.A(_15619_),
    .B(_15726_),
    .CI(_15727_),
    .CO(_15728_),
    .S(_15729_));
 FA_X1 _30405_ (.A(_15660_),
    .B(_15730_),
    .CI(_15731_),
    .CO(_15732_),
    .S(_15733_));
 FA_X1 _30406_ (.A(_15702_),
    .B(_15734_),
    .CI(_15735_),
    .CO(_15736_),
    .S(_15737_));
 FA_X1 _30407_ (.A(_15050_),
    .B(net315),
    .CI(_15738_),
    .CO(_15739_),
    .S(_15740_));
 FA_X1 _30408_ (.A(_15740_),
    .B(_15707_),
    .CI(_15214_),
    .CO(_15741_),
    .S(_15742_));
 FA_X1 _30409_ (.A(_15701_),
    .B(_15743_),
    .CI(_15744_),
    .CO(_15745_),
    .S(_15746_));
 FA_X1 _30410_ (.A(_15747_),
    .B(_15704_),
    .CI(_15748_),
    .CO(_15749_),
    .S(_15750_));
 FA_X1 _30411_ (.A(_15751_),
    .B(_15750_),
    .CI(_15718_),
    .CO(_15752_),
    .S(_15753_));
 FA_X1 _30412_ (.A(_15754_),
    .B(_15755_),
    .CI(_15756_),
    .CO(_15757_),
    .S(_15758_));
 HA_X1 _30413_ (.A(_15760_),
    .B(_15759_),
    .CO(_15761_),
    .S(_15762_));
 HA_X1 _30414_ (.A(_15759_),
    .B(_15763_),
    .CO(_15764_),
    .S(_15765_));
 HA_X1 _30415_ (.A(_15766_),
    .B(_15760_),
    .CO(_15767_),
    .S(_15768_));
 HA_X1 _30416_ (.A(_15766_),
    .B(_15763_),
    .CO(_15769_),
    .S(_15770_));
 HA_X1 _30417_ (.A(_15772_),
    .B(_15771_),
    .CO(_15773_),
    .S(_15774_));
 HA_X1 _30418_ (.A(_14465_),
    .B(_14466_),
    .CO(_15775_),
    .S(_15776_));
 HA_X1 _30419_ (.A(_15777_),
    .B(_15778_),
    .CO(_15779_),
    .S(_15780_));
 HA_X1 _30420_ (.A(_15781_),
    .B(_15782_),
    .CO(_15783_),
    .S(_15784_));
 HA_X1 _30421_ (.A(_15785_),
    .B(_15786_),
    .CO(_15787_),
    .S(_15788_));
 HA_X1 _30422_ (.A(_15789_),
    .B(_15790_),
    .CO(_15791_),
    .S(_15792_));
 HA_X1 _30423_ (.A(_15793_),
    .B(_15794_),
    .CO(_15795_),
    .S(_15796_));
 HA_X1 _30424_ (.A(_15797_),
    .B(_15798_),
    .CO(_15799_),
    .S(_15800_));
 HA_X1 _30425_ (.A(_15801_),
    .B(_15802_),
    .CO(_15803_),
    .S(_15804_));
 HA_X1 _30426_ (.A(_15805_),
    .B(_15806_),
    .CO(_15807_),
    .S(_15808_));
 HA_X1 _30427_ (.A(_15809_),
    .B(_15810_),
    .CO(_15811_),
    .S(_15812_));
 HA_X1 _30428_ (.A(_15813_),
    .B(_15814_),
    .CO(_15815_),
    .S(_15816_));
 HA_X1 _30429_ (.A(_15817_),
    .B(_15818_),
    .CO(_15819_),
    .S(_15820_));
 HA_X1 _30430_ (.A(_15821_),
    .B(_15822_),
    .CO(_15823_),
    .S(_15824_));
 HA_X1 _30431_ (.A(_15825_),
    .B(_15826_),
    .CO(_15827_),
    .S(_15828_));
 HA_X1 _30432_ (.A(_15829_),
    .B(_15830_),
    .CO(_15831_),
    .S(_15832_));
 HA_X1 _30433_ (.A(_15833_),
    .B(_15834_),
    .CO(_15835_),
    .S(_15836_));
 HA_X1 _30434_ (.A(_15837_),
    .B(_15838_),
    .CO(_15839_),
    .S(_15840_));
 HA_X1 _30435_ (.A(_15841_),
    .B(_15842_),
    .CO(_15843_),
    .S(_15844_));
 HA_X1 _30436_ (.A(_15845_),
    .B(_15846_),
    .CO(_15847_),
    .S(_15848_));
 HA_X1 _30437_ (.A(_15849_),
    .B(_15850_),
    .CO(_15851_),
    .S(_15852_));
 HA_X1 _30438_ (.A(_15853_),
    .B(_15854_),
    .CO(_15855_),
    .S(_15856_));
 HA_X1 _30439_ (.A(_15857_),
    .B(_15858_),
    .CO(_15859_),
    .S(_15860_));
 HA_X1 _30440_ (.A(_15861_),
    .B(_15862_),
    .CO(_15863_),
    .S(_15864_));
 HA_X1 _30441_ (.A(_15865_),
    .B(_15866_),
    .CO(_15867_),
    .S(_15868_));
 HA_X1 _30442_ (.A(_15869_),
    .B(_15870_),
    .CO(_15871_),
    .S(_15872_));
 HA_X1 _30443_ (.A(_15873_),
    .B(_15874_),
    .CO(_15875_),
    .S(_15876_));
 HA_X1 _30444_ (.A(_15877_),
    .B(_15878_),
    .CO(_15879_),
    .S(_15880_));
 HA_X1 _30445_ (.A(_15881_),
    .B(_15882_),
    .CO(_15883_),
    .S(_15884_));
 HA_X1 _30446_ (.A(_15885_),
    .B(_15886_),
    .CO(_15887_),
    .S(_15888_));
 HA_X1 _30447_ (.A(_15889_),
    .B(_15890_),
    .CO(_15891_),
    .S(_15892_));
 HA_X1 _30448_ (.A(_15893_),
    .B(_15894_),
    .CO(_15895_),
    .S(_15896_));
 HA_X1 _30449_ (.A(_15897_),
    .B(_15898_),
    .CO(_15899_),
    .S(_15900_));
 HA_X1 _30450_ (.A(_15901_),
    .B(_15902_),
    .CO(_15903_),
    .S(_15904_));
 HA_X1 _30451_ (.A(_15905_),
    .B(\cs_registers_i.priv_lvl_q[0] ),
    .CO(_15906_),
    .S(_15907_));
 HA_X1 _30452_ (.A(_15908_),
    .B(_15909_),
    .CO(_15910_),
    .S(_15911_));
 HA_X1 _30453_ (.A(_15912_),
    .B(_15913_),
    .CO(_15914_),
    .S(_15915_));
 HA_X1 _30454_ (.A(_15912_),
    .B(_15916_),
    .CO(_15917_),
    .S(_15918_));
 HA_X1 _30455_ (.A(_15919_),
    .B(_15913_),
    .CO(_15920_),
    .S(_15921_));
 HA_X1 _30456_ (.A(_15919_),
    .B(_15916_),
    .CO(_15922_),
    .S(_15923_));
 HA_X1 _30457_ (.A(_15924_),
    .B(_15925_),
    .CO(_15926_),
    .S(_15927_));
 HA_X1 _30458_ (.A(_15924_),
    .B(_15928_),
    .CO(_15929_),
    .S(_15930_));
 HA_X1 _30459_ (.A(_15931_),
    .B(_15925_),
    .CO(_15932_),
    .S(_15933_));
 HA_X1 _30460_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(\cs_registers_i.mhpmcounter[2][1] ),
    .CO(_15934_),
    .S(_15935_));
 HA_X1 _30461_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .CO(_15936_),
    .S(_15937_));
 HA_X1 _30462_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CO(_15938_),
    .S(_15939_));
 HA_X1 _30463_ (.A(_15940_),
    .B(_15941_),
    .CO(_15942_),
    .S(_15943_));
 HA_X1 _30464_ (.A(_15940_),
    .B(_15941_),
    .CO(_15944_),
    .S(_15945_));
 HA_X1 _30465_ (.A(_15940_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_15946_),
    .S(_15947_));
 HA_X1 _30466_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_15941_),
    .CO(_15948_),
    .S(_15949_));
 HA_X1 _30467_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_15950_),
    .S(_15951_));
 HA_X1 _30468_ (.A(_15952_),
    .B(_15953_),
    .CO(_15954_),
    .S(_15955_));
 HA_X1 _30469_ (.A(_15956_),
    .B(_15954_),
    .CO(_15957_),
    .S(_15958_));
 HA_X1 _30470_ (.A(_15959_),
    .B(_15960_),
    .CO(_15961_),
    .S(_15962_));
 HA_X1 _30471_ (.A(_15962_),
    .B(_15957_),
    .CO(_15963_),
    .S(_15964_));
 HA_X1 _30472_ (.A(_15964_),
    .B(_15965_),
    .CO(_15966_),
    .S(_15967_));
 HA_X1 _30473_ (.A(_15968_),
    .B(_15969_),
    .CO(_14494_),
    .S(_15970_));
 HA_X1 _30474_ (.A(_15971_),
    .B(_15972_),
    .CO(_15973_),
    .S(_15974_));
 HA_X1 _30475_ (.A(_15961_),
    .B(_15974_),
    .CO(_15975_),
    .S(_15976_));
 HA_X1 _30476_ (.A(_15976_),
    .B(_15963_),
    .CO(_15977_),
    .S(_15978_));
 HA_X1 _30477_ (.A(_15978_),
    .B(_15970_),
    .CO(_15979_),
    .S(_15980_));
 HA_X1 _30478_ (.A(_15980_),
    .B(_15966_),
    .CO(_15981_),
    .S(_15982_));
 HA_X1 _30479_ (.A(_14497_),
    .B(_15973_),
    .CO(_15983_),
    .S(_15984_));
 HA_X1 _30480_ (.A(_15975_),
    .B(_15984_),
    .CO(_15985_),
    .S(_15986_));
 HA_X1 _30481_ (.A(_14487_),
    .B(_15986_),
    .CO(_15987_),
    .S(_15988_));
 HA_X1 _30482_ (.A(_15989_),
    .B(_15981_),
    .CO(_14521_),
    .S(_15990_));
 HA_X1 _30483_ (.A(_14507_),
    .B(_15991_),
    .CO(_15992_),
    .S(_15993_));
 HA_X1 _30484_ (.A(_14496_),
    .B(_15994_),
    .CO(_15995_),
    .S(_15996_));
 HA_X1 _30485_ (.A(_15996_),
    .B(_15983_),
    .CO(_15997_),
    .S(_15998_));
 HA_X1 _30486_ (.A(_15998_),
    .B(_15993_),
    .CO(_15999_),
    .S(_16000_));
 HA_X1 _30487_ (.A(_14522_),
    .B(_14523_),
    .CO(_16001_),
    .S(_16002_));
 HA_X1 _30488_ (.A(_16003_),
    .B(_16004_),
    .CO(_14554_),
    .S(_16005_));
 HA_X1 _30489_ (.A(_16005_),
    .B(_14530_),
    .CO(_16006_),
    .S(_16007_));
 HA_X1 _30490_ (.A(_16007_),
    .B(_15992_),
    .CO(_16008_),
    .S(_16009_));
 HA_X1 _30491_ (.A(_16010_),
    .B(_16011_),
    .CO(_16012_),
    .S(_16013_));
 HA_X1 _30492_ (.A(_15995_),
    .B(_16013_),
    .CO(_16014_),
    .S(_16015_));
 HA_X1 _30493_ (.A(_16015_),
    .B(_16009_),
    .CO(_16016_),
    .S(_16017_));
 HA_X1 _30494_ (.A(_16018_),
    .B(_16019_),
    .CO(_16020_),
    .S(_16021_));
 HA_X1 _30495_ (.A(_14557_),
    .B(_16006_),
    .CO(_16022_),
    .S(_16023_));
 HA_X1 _30496_ (.A(_16024_),
    .B(_16025_),
    .CO(_16026_),
    .S(_16027_));
 HA_X1 _30497_ (.A(_16023_),
    .B(_16028_),
    .CO(_14602_),
    .S(_16029_));
 HA_X1 _30498_ (.A(_16030_),
    .B(_16031_),
    .CO(_16032_),
    .S(_16033_));
 HA_X1 _30499_ (.A(_14556_),
    .B(_16034_),
    .CO(_16035_),
    .S(_16036_));
 HA_X1 _30500_ (.A(_16037_),
    .B(_16036_),
    .CO(_14633_),
    .S(_16038_));
 HA_X1 _30501_ (.A(_16039_),
    .B(_16040_),
    .CO(_16041_),
    .S(_16042_));
 HA_X1 _30502_ (.A(_16043_),
    .B(_16038_),
    .CO(_14638_),
    .S(_14604_));
 HA_X1 _30503_ (.A(_14606_),
    .B(_16044_),
    .CO(_16045_),
    .S(_16046_));
 HA_X1 _30504_ (.A(_16047_),
    .B(_16048_),
    .CO(_16049_),
    .S(_16050_));
 HA_X1 _30505_ (.A(_16051_),
    .B(_16052_),
    .CO(_16053_),
    .S(_16054_));
 HA_X1 _30506_ (.A(_16054_),
    .B(_16050_),
    .CO(_14673_),
    .S(_14634_));
 HA_X1 _30507_ (.A(_16055_),
    .B(_16056_),
    .CO(_16057_),
    .S(_16058_));
 HA_X1 _30508_ (.A(_14641_),
    .B(_14605_),
    .CO(_16059_),
    .S(_16060_));
 HA_X1 _30509_ (.A(_16049_),
    .B(_16061_),
    .CO(_16062_),
    .S(_16063_));
 HA_X1 _30510_ (.A(_16064_),
    .B(_16065_),
    .CO(_16066_),
    .S(_16067_));
 HA_X1 _30511_ (.A(_16067_),
    .B(_16063_),
    .CO(_14716_),
    .S(_14674_));
 HA_X1 _30512_ (.A(_16068_),
    .B(_16069_),
    .CO(_16070_),
    .S(_16071_));
 HA_X1 _30513_ (.A(_16072_),
    .B(_14640_),
    .CO(_16073_),
    .S(_16074_));
 HA_X1 _30514_ (.A(_16075_),
    .B(_16076_),
    .CO(_16077_),
    .S(_16078_));
 HA_X1 _30515_ (.A(_16079_),
    .B(_16078_),
    .CO(_14748_),
    .S(_16080_));
 HA_X1 _30516_ (.A(_16081_),
    .B(_16080_),
    .CO(_14764_),
    .S(_14717_));
 HA_X1 _30517_ (.A(_16082_),
    .B(_16083_),
    .CO(_14761_),
    .S(_16084_));
 HA_X1 _30518_ (.A(_16086_),
    .B(_16085_),
    .CO(_16087_),
    .S(_16088_));
 HA_X1 _30519_ (.A(_16089_),
    .B(_16090_),
    .CO(_16091_),
    .S(_16092_));
 HA_X1 _30520_ (.A(_16093_),
    .B(_16094_),
    .CO(_16095_),
    .S(_16096_));
 HA_X1 _30521_ (.A(_16096_),
    .B(_16092_),
    .CO(_14800_),
    .S(_14746_));
 HA_X1 _30522_ (.A(_16097_),
    .B(_16098_),
    .CO(_14814_),
    .S(_14759_));
 HA_X1 _30523_ (.A(_16100_),
    .B(_16099_),
    .CO(_16101_),
    .S(_16102_));
 HA_X1 _30524_ (.A(_14775_),
    .B(_16103_),
    .CO(_14855_),
    .S(_14801_));
 HA_X1 _30525_ (.A(_16104_),
    .B(_16105_),
    .CO(_14869_),
    .S(_14815_));
 HA_X1 _30526_ (.A(_16106_),
    .B(_16107_),
    .CO(_16108_),
    .S(_16109_));
 HA_X1 _30527_ (.A(_16110_),
    .B(_16111_),
    .CO(_14893_),
    .S(_16112_));
 HA_X1 _30528_ (.A(_16112_),
    .B(_16113_),
    .CO(_14914_),
    .S(_14857_));
 HA_X1 _30529_ (.A(_16114_),
    .B(_16115_),
    .CO(_14927_),
    .S(_14870_));
 HA_X1 _30530_ (.A(_16116_),
    .B(_16117_),
    .CO(_16118_),
    .S(_16119_));
 HA_X1 _30531_ (.A(_16120_),
    .B(_16121_),
    .CO(_14948_),
    .S(_16122_));
 HA_X1 _30532_ (.A(_16122_),
    .B(_14885_),
    .CO(_14961_),
    .S(_14894_));
 HA_X1 _30533_ (.A(_16123_),
    .B(_16124_),
    .CO(_14997_),
    .S(_14925_));
 HA_X1 _30534_ (.A(_16125_),
    .B(_16126_),
    .CO(_16127_),
    .S(_16128_));
 HA_X1 _30535_ (.A(_16129_),
    .B(_16130_),
    .CO(_16131_),
    .S(_16132_));
 HA_X1 _30536_ (.A(_15050_),
    .B(net315),
    .CO(_16133_),
    .S(_16134_));
 HA_X1 _30537_ (.A(_16135_),
    .B(_16136_),
    .CO(_15118_),
    .S(_16137_));
 HA_X1 _30538_ (.A(_16138_),
    .B(_16139_),
    .CO(_16140_),
    .S(_16141_));
 HA_X1 _30539_ (.A(_16142_),
    .B(_16143_),
    .CO(_15174_),
    .S(_15116_));
 HA_X1 _30540_ (.A(_16144_),
    .B(_16145_),
    .CO(_16146_),
    .S(_16147_));
 HA_X1 _30541_ (.A(_16148_),
    .B(_16149_),
    .CO(_15230_),
    .S(_15175_));
 HA_X1 _30542_ (.A(_16150_),
    .B(_16151_),
    .CO(_16152_),
    .S(_16153_));
 HA_X1 _30543_ (.A(_16154_),
    .B(_16155_),
    .CO(_15285_),
    .S(_15231_));
 HA_X1 _30544_ (.A(_16156_),
    .B(_16157_),
    .CO(_16158_),
    .S(_16159_));
 HA_X1 _30545_ (.A(_16160_),
    .B(_16161_),
    .CO(_15338_),
    .S(_15283_));
 HA_X1 _30546_ (.A(_16162_),
    .B(_16163_),
    .CO(_16164_),
    .S(_16165_));
 HA_X1 _30547_ (.A(_16166_),
    .B(_16167_),
    .CO(_15392_),
    .S(_15339_));
 HA_X1 _30548_ (.A(_16169_),
    .B(_16168_),
    .CO(_16170_),
    .S(_16171_));
 HA_X1 _30549_ (.A(_16172_),
    .B(_16173_),
    .CO(_15438_),
    .S(_15390_));
 HA_X1 _30550_ (.A(_16174_),
    .B(_16175_),
    .CO(_16176_),
    .S(_16177_));
 HA_X1 _30551_ (.A(_16178_),
    .B(_16179_),
    .CO(_15479_),
    .S(_15436_));
 HA_X1 _30552_ (.A(_16180_),
    .B(_16181_),
    .CO(_16182_),
    .S(_16183_));
 HA_X1 _30553_ (.A(_16184_),
    .B(_16185_),
    .CO(_15523_),
    .S(_15481_));
 HA_X1 _30554_ (.A(_16186_),
    .B(_16187_),
    .CO(_16188_),
    .S(_16189_));
 HA_X1 _30555_ (.A(_16190_),
    .B(_16191_),
    .CO(_15562_),
    .S(_15525_));
 HA_X1 _30556_ (.A(_16192_),
    .B(_16193_),
    .CO(_16194_),
    .S(_16195_));
 HA_X1 _30557_ (.A(_16196_),
    .B(_16197_),
    .CO(_15600_),
    .S(_15564_));
 HA_X1 _30558_ (.A(_16198_),
    .B(_16199_),
    .CO(_16200_),
    .S(_16201_));
 HA_X1 _30559_ (.A(_16202_),
    .B(_16203_),
    .CO(_15640_),
    .S(_15601_));
 HA_X1 _30560_ (.A(_16204_),
    .B(_16205_),
    .CO(_16206_),
    .S(_16207_));
 HA_X1 _30561_ (.A(_16208_),
    .B(_16209_),
    .CO(_15679_),
    .S(_15638_));
 HA_X1 _30562_ (.A(_16210_),
    .B(_16211_),
    .CO(_16212_),
    .S(_16213_));
 HA_X1 _30563_ (.A(_16214_),
    .B(_16215_),
    .CO(_15713_),
    .S(_15677_));
 HA_X1 _30564_ (.A(_16216_),
    .B(_16217_),
    .CO(_16218_),
    .S(_16219_));
 HA_X1 _30565_ (.A(_16220_),
    .B(_16221_),
    .CO(_15743_),
    .S(_15714_));
 HA_X1 _30566_ (.A(_16222_),
    .B(_16223_),
    .CO(_16224_),
    .S(_16225_));
 HA_X1 _30567_ (.A(_15742_),
    .B(_16226_),
    .CO(_16227_),
    .S(_15744_));
 HA_X1 _30568_ (.A(_16228_),
    .B(_16229_),
    .CO(_16230_),
    .S(_16231_));
 HA_X1 _30569_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_16232_),
    .CO(_16233_),
    .S(_16234_));
 HA_X1 _30570_ (.A(_11173_),
    .B(_16236_),
    .CO(_16237_),
    .S(_16238_));
 HA_X1 _30571_ (.A(_11173_),
    .B(_16239_),
    .CO(_16240_),
    .S(_16241_));
 HA_X1 _30572_ (.A(_16242_),
    .B(_16243_),
    .CO(_16244_),
    .S(_16245_));
 HA_X1 _30573_ (.A(_16246_),
    .B(_16247_),
    .CO(_16248_),
    .S(_16249_));
 HA_X1 _30574_ (.A(_16250_),
    .B(_16236_),
    .CO(_16251_),
    .S(_16252_));
 HA_X1 _30575_ (.A(_16253_),
    .B(_16254_),
    .CO(_16255_),
    .S(_16256_));
 HA_X1 _30576_ (.A(_11379_),
    .B(_16258_),
    .CO(_16259_),
    .S(_16260_));
 HA_X1 _30577_ (.A(_16261_),
    .B(_16262_),
    .CO(_16263_),
    .S(_16264_));
 HA_X1 _30578_ (.A(_16265_),
    .B(_16266_),
    .CO(_16267_),
    .S(_16268_));
 HA_X1 _30579_ (.A(_16269_),
    .B(_16270_),
    .CO(_16271_),
    .S(_16272_));
 HA_X1 _30580_ (.A(_16273_),
    .B(_16274_),
    .CO(_16275_),
    .S(_16276_));
 HA_X1 _30581_ (.A(_16277_),
    .B(_16278_),
    .CO(_16279_),
    .S(_16280_));
 HA_X1 _30582_ (.A(_16281_),
    .B(_16282_),
    .CO(_16283_),
    .S(_16284_));
 HA_X1 _30583_ (.A(_16285_),
    .B(_16286_),
    .CO(_16287_),
    .S(_16288_));
 HA_X1 _30584_ (.A(_16289_),
    .B(_16290_),
    .CO(_16291_),
    .S(_16292_));
 HA_X1 _30585_ (.A(_16293_),
    .B(_16294_),
    .CO(_16295_),
    .S(_16296_));
 HA_X1 _30586_ (.A(_16297_),
    .B(_16298_),
    .CO(_16299_),
    .S(_16300_));
 HA_X1 _30587_ (.A(_16301_),
    .B(_16302_),
    .CO(_16303_),
    .S(_16304_));
 HA_X1 _30588_ (.A(_16305_),
    .B(_16306_),
    .CO(_16307_),
    .S(_16308_));
 HA_X1 _30589_ (.A(_16309_),
    .B(_16310_),
    .CO(_16311_),
    .S(_16312_));
 HA_X1 _30590_ (.A(_16313_),
    .B(_16314_),
    .CO(_16315_),
    .S(_16316_));
 HA_X1 _30591_ (.A(_16317_),
    .B(_16318_),
    .CO(_16319_),
    .S(_16320_));
 HA_X1 _30592_ (.A(_16321_),
    .B(_16322_),
    .CO(_16323_),
    .S(_16324_));
 HA_X1 _30593_ (.A(_16325_),
    .B(_16326_),
    .CO(_16327_),
    .S(_16328_));
 HA_X1 _30594_ (.A(_16329_),
    .B(_16330_),
    .CO(_16331_),
    .S(_16332_));
 HA_X1 _30595_ (.A(_16333_),
    .B(_16334_),
    .CO(_16335_),
    .S(_16336_));
 HA_X1 _30596_ (.A(_16337_),
    .B(_16338_),
    .CO(_16339_),
    .S(_16340_));
 HA_X1 _30597_ (.A(_16341_),
    .B(_16342_),
    .CO(_16343_),
    .S(_16344_));
 HA_X1 _30598_ (.A(_16345_),
    .B(_16346_),
    .CO(_16347_),
    .S(_16348_));
 HA_X1 _30599_ (.A(_16349_),
    .B(_16350_),
    .CO(_16351_),
    .S(_16352_));
 HA_X1 _30600_ (.A(_16353_),
    .B(_16354_),
    .CO(_16355_),
    .S(_16356_));
 HA_X1 _30601_ (.A(_16357_),
    .B(_16358_),
    .CO(_16359_),
    .S(_16360_));
 HA_X1 _30602_ (.A(_16361_),
    .B(_16362_),
    .CO(_16363_),
    .S(_16364_));
 HA_X1 _30603_ (.A(_16365_),
    .B(_16366_),
    .CO(_16367_),
    .S(_16368_));
 HA_X1 _30604_ (.A(_16369_),
    .B(_16370_),
    .CO(_16371_),
    .S(_16372_));
 HA_X1 _30605_ (.A(_16373_),
    .B(_16374_),
    .CO(_16375_),
    .S(_16376_));
 HA_X1 _30606_ (.A(_16377_),
    .B(_16378_),
    .CO(_16379_),
    .S(_16380_));
 HA_X1 _30607_ (.A(_16381_),
    .B(_16382_),
    .CO(_16383_),
    .S(_16384_));
 HA_X1 _30608_ (.A(_16385_),
    .B(_16386_),
    .CO(_16387_),
    .S(_16388_));
 HA_X1 _30609_ (.A(_16389_),
    .B(_16390_),
    .CO(_16391_),
    .S(_16392_));
 HA_X1 _30610_ (.A(_16393_),
    .B(_16394_),
    .CO(_16395_),
    .S(_16396_));
 HA_X1 _30611_ (.A(_16397_),
    .B(_16398_),
    .CO(_16399_),
    .S(_16400_));
 HA_X1 _30612_ (.A(_16401_),
    .B(_16402_),
    .CO(_16403_),
    .S(_16404_));
 HA_X1 _30613_ (.A(_16405_),
    .B(_16406_),
    .CO(_16407_),
    .S(_16408_));
 HA_X1 _30614_ (.A(_16409_),
    .B(_16410_),
    .CO(_16411_),
    .S(_16412_));
 HA_X1 _30615_ (.A(_16413_),
    .B(_16414_),
    .CO(_16415_),
    .S(_16416_));
 HA_X1 _30616_ (.A(_16417_),
    .B(_16418_),
    .CO(_16419_),
    .S(_16420_));
 HA_X1 _30617_ (.A(_16421_),
    .B(_16422_),
    .CO(_16423_),
    .S(_16424_));
 HA_X1 _30618_ (.A(_16425_),
    .B(_16426_),
    .CO(_16427_),
    .S(_16428_));
 HA_X1 _30619_ (.A(_16429_),
    .B(_16430_),
    .CO(_16431_),
    .S(_16432_));
 HA_X1 _30620_ (.A(_16433_),
    .B(_16434_),
    .CO(_16435_),
    .S(_16436_));
 HA_X1 _30621_ (.A(_16437_),
    .B(_16438_),
    .CO(_16439_),
    .S(_16440_));
 HA_X1 _30622_ (.A(_16441_),
    .B(_16442_),
    .CO(_16443_),
    .S(_16444_));
 HA_X1 _30623_ (.A(_16445_),
    .B(_16446_),
    .CO(_16447_),
    .S(_16448_));
 HA_X1 _30624_ (.A(_16449_),
    .B(_16450_),
    .CO(_16451_),
    .S(_16452_));
 HA_X1 _30625_ (.A(_16453_),
    .B(_16454_),
    .CO(_16455_),
    .S(_16456_));
 HA_X1 _30626_ (.A(_16457_),
    .B(_16458_),
    .CO(_16459_),
    .S(_16460_));
 HA_X1 _30627_ (.A(_16461_),
    .B(_16462_),
    .CO(_16463_),
    .S(_16464_));
 HA_X1 _30628_ (.A(_16465_),
    .B(_16466_),
    .CO(_16467_),
    .S(_16468_));
 HA_X1 _30629_ (.A(_16469_),
    .B(_16470_),
    .CO(_16471_),
    .S(_16472_));
 HA_X1 _30630_ (.A(_16473_),
    .B(_16474_),
    .CO(_16475_),
    .S(_16476_));
 HA_X1 _30631_ (.A(_16477_),
    .B(_16478_),
    .CO(_16479_),
    .S(_16480_));
 HA_X1 _30632_ (.A(_16481_),
    .B(_16482_),
    .CO(_16483_),
    .S(_16484_));
 HA_X1 _30633_ (.A(_16485_),
    .B(_16486_),
    .CO(_16487_),
    .S(_16488_));
 HA_X1 _30634_ (.A(\alu_adder_result_ex[1] ),
    .B(_16486_),
    .CO(_16489_),
    .S(_16490_));
 HA_X1 _30635_ (.A(_16491_),
    .B(_16486_),
    .CO(_16492_),
    .S(_16493_));
 HA_X1 _30636_ (.A(\alu_adder_result_ex[0] ),
    .B(\alu_adder_result_ex[1] ),
    .CO(_16494_),
    .S(_16495_));
 HA_X1 _30637_ (.A(\alu_adder_result_ex[0] ),
    .B(\alu_adder_result_ex[1] ),
    .CO(_16496_),
    .S(_16497_));
 HA_X1 _30638_ (.A(\alu_adder_result_ex[0] ),
    .B(_16491_),
    .CO(_16498_),
    .S(_16499_));
 HA_X1 _30639_ (.A(\alu_adder_result_ex[0] ),
    .B(_16491_),
    .CO(_16500_),
    .S(_16501_));
 HA_X1 _30640_ (.A(_16502_),
    .B(\alu_adder_result_ex[1] ),
    .CO(_16503_),
    .S(_16504_));
 HA_X1 _30641_ (.A(_16502_),
    .B(\alu_adder_result_ex[1] ),
    .CO(_16505_),
    .S(_16506_));
 HA_X1 _30642_ (.A(_16502_),
    .B(_16491_),
    .CO(_16507_),
    .S(_16508_));
 HA_X1 _30643_ (.A(_16509_),
    .B(_16510_),
    .CO(_16511_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ));
 HA_X1 _30644_ (.A(_16511_),
    .B(_16512_),
    .CO(_16513_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ));
 DFFR_X2 _30645_ (.D(_02683_),
    .RN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .QN(_14449_));
 DFFR_X1 _30646_ (.D(_02684_),
    .RN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .QN(_14448_));
 DFFR_X2 _30647_ (.D(_02685_),
    .RN(net246),
    .CK(clknet_leaf_39_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .QN(_00179_));
 DFFR_X1 _30648_ (.D(_02686_),
    .RN(net246),
    .CK(clknet_leaf_39_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .QN(_14447_));
 DFFS_X1 _30649_ (.D(_02687_),
    .SN(net246),
    .CK(clknet_leaf_41_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .QN(_14446_));
 DFFR_X1 _30650_ (.D(_02688_),
    .RN(net265),
    .CK(clknet_leaf_19_clk),
    .Q(\load_store_unit_i.data_type_q[2] ),
    .QN(_14445_));
 DFFR_X1 _30651_ (.D(_02689_),
    .RN(net265),
    .CK(clknet_leaf_18_clk),
    .Q(\load_store_unit_i.data_type_q[1] ),
    .QN(_14450_));
 CLKBUF_X3 clkbuf_regs_0_core_clock (.A(clk_i),
    .Z(delaynet_0_core_clock));
 BUF_X1 _30653_ (.A(net269),
    .Z(alert_major_o));
 BUF_X1 _30654_ (.A(net270),
    .Z(alert_minor_o));
 BUF_X1 _30655_ (.A(net271),
    .Z(data_addr_o[0]));
 BUF_X1 _30656_ (.A(net272),
    .Z(data_addr_o[1]));
 BUF_X1 _30657_ (.A(\alu_adder_result_ex[2] ),
    .Z(net167));
 BUF_X1 _30658_ (.A(\alu_adder_result_ex[3] ),
    .Z(net170));
 BUF_X1 _30659_ (.A(\alu_adder_result_ex[4] ),
    .Z(net171));
 BUF_X1 _30660_ (.A(\alu_adder_result_ex[5] ),
    .Z(net172));
 CLKBUF_X2 _30661_ (.A(net8),
    .Z(net173));
 BUF_X1 _30662_ (.A(\alu_adder_result_ex[7] ),
    .Z(net174));
 BUF_X1 _30663_ (.A(\alu_adder_result_ex[8] ),
    .Z(net175));
 BUF_X2 _30664_ (.A(\alu_adder_result_ex[9] ),
    .Z(net176));
 BUF_X1 _30665_ (.A(\alu_adder_result_ex[10] ),
    .Z(net147));
 BUF_X2 _30666_ (.A(\alu_adder_result_ex[11] ),
    .Z(net148));
 BUF_X2 _30667_ (.A(\alu_adder_result_ex[12] ),
    .Z(net149));
 BUF_X1 _30668_ (.A(\alu_adder_result_ex[13] ),
    .Z(net150));
 BUF_X1 _30669_ (.A(net7),
    .Z(net151));
 BUF_X1 _30670_ (.A(net437),
    .Z(net152));
 BUF_X1 _30671_ (.A(\alu_adder_result_ex[16] ),
    .Z(net153));
 BUF_X1 _30672_ (.A(\alu_adder_result_ex[17] ),
    .Z(net154));
 BUF_X1 _30673_ (.A(\alu_adder_result_ex[18] ),
    .Z(net155));
 BUF_X1 _30674_ (.A(\alu_adder_result_ex[19] ),
    .Z(net156));
 BUF_X1 _30675_ (.A(\alu_adder_result_ex[20] ),
    .Z(net157));
 CLKBUF_X2 _30676_ (.A(\alu_adder_result_ex[21] ),
    .Z(net158));
 BUF_X1 _30677_ (.A(\alu_adder_result_ex[22] ),
    .Z(net159));
 BUF_X1 _30678_ (.A(net356),
    .Z(net160));
 CLKBUF_X2 _30679_ (.A(\alu_adder_result_ex[24] ),
    .Z(net161));
 BUF_X2 _30680_ (.A(net390),
    .Z(net162));
 BUF_X2 _30681_ (.A(\alu_adder_result_ex[26] ),
    .Z(net163));
 BUF_X1 _30682_ (.A(\alu_adder_result_ex[27] ),
    .Z(net164));
 BUF_X1 _30683_ (.A(\alu_adder_result_ex[28] ),
    .Z(net165));
 CLKBUF_X2 _30684_ (.A(\alu_adder_result_ex[29] ),
    .Z(net166));
 BUF_X1 _30685_ (.A(\alu_adder_result_ex[30] ),
    .Z(net168));
 BUF_X1 _30686_ (.A(_03517_),
    .Z(net169));
 BUF_X1 _30687_ (.A(net273),
    .Z(instr_addr_o[0]));
 BUF_X1 _30688_ (.A(net274),
    .Z(instr_addr_o[1]));
 DFFR_X1 \core_busy_q$_DFF_PN0_  (.D(core_busy_d),
    .RN(net254),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(core_busy_q),
    .QN(_14444_));
 DLL_X1 \core_clock_gate_i.en_latch$_DLATCH_N_  (.D(_00006_),
    .GN(clknet_leaf_118_clk_i_regs),
    .Q(\core_clock_gate_i.en_latch ));
 DFFR_X2 \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.D(_02690_),
    .RN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.mcountinhibit[0] ),
    .QN(_00554_));
 DFFR_X1 \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.D(_02691_),
    .RN(net248),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.mcountinhibit[2] ),
    .QN(_01158_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[0]$_DFFE_PN0P_  (.D(_02692_),
    .RN(net630),
    .CK(clknet_leaf_134_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .QN(_00552_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[10]$_DFFE_PN0P_  (.D(_02693_),
    .RN(net254),
    .CK(clknet_leaf_133_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .QN(_14443_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[11]$_DFFE_PN0P_  (.D(_02694_),
    .RN(net630),
    .CK(clknet_leaf_135_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .QN(_14442_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[12]$_DFFE_PN0P_  (.D(_02695_),
    .RN(net630),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .QN(_14441_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[13]$_DFFE_PN0P_  (.D(_02696_),
    .RN(net630),
    .CK(clknet_leaf_135_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .QN(_14440_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[14]$_DFFE_PN0P_  (.D(_02697_),
    .RN(net630),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .QN(_14439_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[15]$_DFFE_PN0P_  (.D(_02698_),
    .RN(net630),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .QN(_14438_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[16]$_DFFE_PN0P_  (.D(_02699_),
    .RN(net630),
    .CK(clknet_leaf_123_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .QN(_14437_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[17]$_DFFE_PN0P_  (.D(_02700_),
    .RN(net254),
    .CK(clknet_leaf_123_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .QN(_14436_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[18]$_DFFE_PN0P_  (.D(_02701_),
    .RN(net254),
    .CK(clknet_leaf_123_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .QN(_14435_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[19]$_DFFE_PN0P_  (.D(_02702_),
    .RN(net254),
    .CK(clknet_leaf_123_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .QN(_14434_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[1]$_DFFE_PN0P_  (.D(_02703_),
    .RN(net630),
    .CK(clknet_leaf_134_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .QN(_14433_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[20]$_DFFE_PN0P_  (.D(_02704_),
    .RN(net254),
    .CK(clknet_leaf_133_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .QN(_14432_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[21]$_DFFE_PN0P_  (.D(_02705_),
    .RN(net254),
    .CK(clknet_leaf_133_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .QN(_14431_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[22]$_DFFE_PN0P_  (.D(_02706_),
    .RN(net254),
    .CK(clknet_leaf_124_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .QN(_14430_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[23]$_DFFE_PN0P_  (.D(_02707_),
    .RN(net254),
    .CK(clknet_leaf_133_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .QN(_14429_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[24]$_DFFE_PN0P_  (.D(_02708_),
    .RN(net254),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .QN(_14428_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[25]$_DFFE_PN0P_  (.D(_02709_),
    .RN(net253),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .QN(_14427_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[26]$_DFFE_PN0P_  (.D(_02710_),
    .RN(net253),
    .CK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .QN(_14426_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[27]$_DFFE_PN0P_  (.D(_02711_),
    .RN(net254),
    .CK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .QN(_14425_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[28]$_DFFE_PN0P_  (.D(_02712_),
    .RN(net254),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .QN(_14424_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[29]$_DFFE_PN0P_  (.D(_02713_),
    .RN(net254),
    .CK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .QN(_14423_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[2]$_DFFE_PN0P_  (.D(_02714_),
    .RN(net630),
    .CK(clknet_leaf_134_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .QN(_14422_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[30]$_DFFE_PN0P_  (.D(_02715_),
    .RN(net253),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .QN(_14421_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[31]$_DFFE_PN0P_  (.D(_02716_),
    .RN(net630),
    .CK(clknet_leaf_138_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .QN(_14420_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[32]$_DFFE_PN0P_  (.D(_02717_),
    .RN(net254),
    .CK(clknet_leaf_133_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .QN(_14419_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[33]$_DFFE_PN0P_  (.D(_02718_),
    .RN(net630),
    .CK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .QN(_14418_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[34]$_DFFE_PN0P_  (.D(_02719_),
    .RN(net254),
    .CK(clknet_leaf_133_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .QN(_14417_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[35]$_DFFE_PN0P_  (.D(_02720_),
    .RN(net630),
    .CK(clknet_leaf_138_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .QN(_14416_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[36]$_DFFE_PN0P_  (.D(_02721_),
    .RN(net630),
    .CK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .QN(_14415_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[37]$_DFFE_PN0P_  (.D(_02722_),
    .RN(net630),
    .CK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .QN(_14414_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[38]$_DFFE_PN0P_  (.D(_02723_),
    .RN(net630),
    .CK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .QN(_14413_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[39]$_DFFE_PN0P_  (.D(_02724_),
    .RN(net254),
    .CK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .QN(_14412_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[3]$_DFFE_PN0P_  (.D(_02725_),
    .RN(net630),
    .CK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .QN(_14411_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[40]$_DFFE_PN0P_  (.D(_02726_),
    .RN(net254),
    .CK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .QN(_14410_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[41]$_DFFE_PN0P_  (.D(_02727_),
    .RN(net630),
    .CK(clknet_leaf_138_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .QN(_14409_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[42]$_DFFE_PN0P_  (.D(_02728_),
    .RN(net630),
    .CK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .QN(_14408_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[43]$_DFFE_PN0P_  (.D(_02729_),
    .RN(net254),
    .CK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .QN(_14407_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[44]$_DFFE_PN0P_  (.D(_02730_),
    .RN(net254),
    .CK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .QN(_14406_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[45]$_DFFE_PN0P_  (.D(_02731_),
    .RN(net254),
    .CK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .QN(_14405_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[46]$_DFFE_PN0P_  (.D(_02732_),
    .RN(net254),
    .CK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .QN(_14404_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[47]$_DFFE_PN0P_  (.D(_02733_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .QN(_14403_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[48]$_DFFE_PN0P_  (.D(_02734_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .QN(_14402_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[49]$_DFFE_PN0P_  (.D(_02735_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .QN(_14401_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[4]$_DFFE_PN0P_  (.D(_02736_),
    .RN(net630),
    .CK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .QN(_14400_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[50]$_DFFE_PN0P_  (.D(_02737_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .QN(_14399_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[51]$_DFFE_PN0P_  (.D(_02738_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .QN(_14398_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[52]$_DFFE_PN0P_  (.D(_02739_),
    .RN(net254),
    .CK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .QN(_14397_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[53]$_DFFE_PN0P_  (.D(_02740_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .QN(_14396_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[54]$_DFFE_PN0P_  (.D(_02741_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .QN(_14395_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[55]$_DFFE_PN0P_  (.D(_02742_),
    .RN(net254),
    .CK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .QN(_14394_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[56]$_DFFE_PN0P_  (.D(_02743_),
    .RN(net254),
    .CK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .QN(_14393_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[57]$_DFFE_PN0P_  (.D(_02744_),
    .RN(net253),
    .CK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .QN(_14392_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[58]$_DFFE_PN0P_  (.D(_02745_),
    .RN(net254),
    .CK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .QN(_14391_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[59]$_DFFE_PN0P_  (.D(_02746_),
    .RN(net254),
    .CK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .QN(_14390_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[5]$_DFFE_PN0P_  (.D(_02747_),
    .RN(net254),
    .CK(clknet_leaf_133_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .QN(_14389_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[60]$_DFFE_PN0P_  (.D(_02748_),
    .RN(net253),
    .CK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .QN(_14388_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[61]$_DFFE_PN0P_  (.D(_02749_),
    .RN(net254),
    .CK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .QN(_14387_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[62]$_DFFE_PN0P_  (.D(_02750_),
    .RN(net253),
    .CK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .QN(_14386_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[63]$_DFFE_PN0P_  (.D(_02751_),
    .RN(net254),
    .CK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .QN(_14385_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[6]$_DFFE_PN0P_  (.D(_02752_),
    .RN(net630),
    .CK(clknet_leaf_137_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .QN(_14384_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[7]$_DFFE_PN0P_  (.D(_02753_),
    .RN(net630),
    .CK(clknet_leaf_134_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .QN(_14383_));
 DFFR_X1 \cs_registers_i.mcycle_counter_i.counter_q[8]$_DFFE_PN0P_  (.D(_02754_),
    .RN(net630),
    .CK(clknet_leaf_134_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .QN(_14382_));
 DFFR_X2 \cs_registers_i.mcycle_counter_i.counter_q[9]$_DFFE_PN0P_  (.D(_02755_),
    .RN(net630),
    .CK(clknet_leaf_134_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .QN(_14381_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[0]$_DFFE_PN0P_  (.D(_02756_),
    .RN(net253),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mhpmcounter[2][0] ),
    .QN(_00553_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[10]$_DFFE_PN0P_  (.D(_02757_),
    .RN(net254),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mhpmcounter[2][10] ),
    .QN(_14380_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[11]$_DFFE_PN0P_  (.D(_02758_),
    .RN(net248),
    .CK(clknet_leaf_124_clk),
    .Q(\cs_registers_i.mhpmcounter[2][11] ),
    .QN(_14379_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[12]$_DFFE_PN0P_  (.D(_02759_),
    .RN(net254),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mhpmcounter[2][12] ),
    .QN(_14378_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[13]$_DFFE_PN0P_  (.D(_02760_),
    .RN(net630),
    .CK(clknet_leaf_121_clk),
    .Q(\cs_registers_i.mhpmcounter[2][13] ),
    .QN(_14377_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[14]$_DFFE_PN0P_  (.D(_02761_),
    .RN(net254),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.mhpmcounter[2][14] ),
    .QN(_14376_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[15]$_DFFE_PN0P_  (.D(_02762_),
    .RN(net248),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mhpmcounter[2][15] ),
    .QN(_14375_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[16]$_DFFE_PN0P_  (.D(_02763_),
    .RN(net248),
    .CK(clknet_leaf_124_clk),
    .Q(\cs_registers_i.mhpmcounter[2][16] ),
    .QN(_14374_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[17]$_DFFE_PN0P_  (.D(_02764_),
    .RN(net248),
    .CK(clknet_leaf_124_clk),
    .Q(\cs_registers_i.mhpmcounter[2][17] ),
    .QN(_14373_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[18]$_DFFE_PN0P_  (.D(_02765_),
    .RN(net248),
    .CK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mhpmcounter[2][18] ),
    .QN(_14372_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[19]$_DFFE_PN0P_  (.D(_02766_),
    .RN(net248),
    .CK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mhpmcounter[2][19] ),
    .QN(_14371_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[1]$_DFFE_PN0P_  (.D(_02767_),
    .RN(net253),
    .CK(clknet_leaf_126_clk),
    .Q(\cs_registers_i.mhpmcounter[2][1] ),
    .QN(_14370_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[20]$_DFFE_PN0P_  (.D(_02768_),
    .RN(net248),
    .CK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mhpmcounter[2][20] ),
    .QN(_14369_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[21]$_DFFE_PN0P_  (.D(_02769_),
    .RN(net248),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mhpmcounter[2][21] ),
    .QN(_14368_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[22]$_DFFE_PN0P_  (.D(_02770_),
    .RN(net248),
    .CK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mhpmcounter[2][22] ),
    .QN(_14367_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[23]$_DFFE_PN0P_  (.D(_02771_),
    .RN(net248),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mhpmcounter[2][23] ),
    .QN(_14366_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[24]$_DFFE_PN0P_  (.D(_02772_),
    .RN(net248),
    .CK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mhpmcounter[2][24] ),
    .QN(_14365_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[25]$_DFFE_PN0P_  (.D(_02773_),
    .RN(net248),
    .CK(clknet_leaf_124_clk),
    .Q(\cs_registers_i.mhpmcounter[2][25] ),
    .QN(_14364_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[26]$_DFFE_PN0P_  (.D(_02774_),
    .RN(net253),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mhpmcounter[2][26] ),
    .QN(_14363_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[27]$_DFFE_PN0P_  (.D(_02775_),
    .RN(net253),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mhpmcounter[2][27] ),
    .QN(_14362_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[28]$_DFFE_PN0P_  (.D(_02776_),
    .RN(net248),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mhpmcounter[2][28] ),
    .QN(_14361_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[29]$_DFFE_PN0P_  (.D(_02777_),
    .RN(net248),
    .CK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mhpmcounter[2][29] ),
    .QN(_14360_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[2]$_DFFE_PN0P_  (.D(_02778_),
    .RN(net254),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mhpmcounter[2][2] ),
    .QN(_14359_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[30]$_DFFE_PN0P_  (.D(_02779_),
    .RN(net248),
    .CK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mhpmcounter[2][30] ),
    .QN(_14358_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[31]$_DFFE_PN0P_  (.D(_02780_),
    .RN(net253),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mhpmcounter[2][31] ),
    .QN(_14357_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[32]$_DFFE_PN0P_  (.D(_02781_),
    .RN(net253),
    .CK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mhpmcounter[2][32] ),
    .QN(_14356_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[33]$_DFFE_PN0P_  (.D(_02782_),
    .RN(net253),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mhpmcounter[2][33] ),
    .QN(_14355_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[34]$_DFFE_PN0P_  (.D(_02783_),
    .RN(net253),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mhpmcounter[2][34] ),
    .QN(_14354_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[35]$_DFFE_PN0P_  (.D(_02784_),
    .RN(net253),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mhpmcounter[2][35] ),
    .QN(_14353_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[36]$_DFFE_PN0P_  (.D(_02785_),
    .RN(net253),
    .CK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mhpmcounter[2][36] ),
    .QN(_14352_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[37]$_DFFE_PN0P_  (.D(_02786_),
    .RN(net253),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mhpmcounter[2][37] ),
    .QN(_14351_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[38]$_DFFE_PN0P_  (.D(_02787_),
    .RN(net253),
    .CK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mhpmcounter[2][38] ),
    .QN(_14350_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[39]$_DFFE_PN0P_  (.D(_02788_),
    .RN(net253),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mhpmcounter[2][39] ),
    .QN(_14349_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[3]$_DFFE_PN0P_  (.D(_02789_),
    .RN(net254),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mhpmcounter[2][3] ),
    .QN(_14348_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[40]$_DFFE_PN0P_  (.D(_02790_),
    .RN(net253),
    .CK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mhpmcounter[2][40] ),
    .QN(_14347_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[41]$_DFFE_PN0P_  (.D(_02791_),
    .RN(net253),
    .CK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mhpmcounter[2][41] ),
    .QN(_14346_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[42]$_DFFE_PN0P_  (.D(_02792_),
    .RN(net253),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mhpmcounter[2][42] ),
    .QN(_14345_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[43]$_DFFE_PN0P_  (.D(_02793_),
    .RN(net253),
    .CK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mhpmcounter[2][43] ),
    .QN(_14344_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[44]$_DFFE_PN0P_  (.D(_02794_),
    .RN(net253),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mhpmcounter[2][44] ),
    .QN(_14343_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[45]$_DFFE_PN0P_  (.D(_02795_),
    .RN(net253),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mhpmcounter[2][45] ),
    .QN(_14342_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[46]$_DFFE_PN0P_  (.D(_02796_),
    .RN(net253),
    .CK(clknet_leaf_106_clk),
    .Q(\cs_registers_i.mhpmcounter[2][46] ),
    .QN(_14341_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[47]$_DFFE_PN0P_  (.D(_02797_),
    .RN(net253),
    .CK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mhpmcounter[2][47] ),
    .QN(_14340_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[48]$_DFFE_PN0P_  (.D(_02798_),
    .RN(net253),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][48] ),
    .QN(_14339_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[49]$_DFFE_PN0P_  (.D(_02799_),
    .RN(net253),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mhpmcounter[2][49] ),
    .QN(_14338_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[4]$_DFFE_PN0P_  (.D(_02800_),
    .RN(net254),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mhpmcounter[2][4] ),
    .QN(_14337_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[50]$_DFFE_PN0P_  (.D(_02801_),
    .RN(net253),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.mhpmcounter[2][50] ),
    .QN(_14336_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[51]$_DFFE_PN0P_  (.D(_02802_),
    .RN(net253),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mhpmcounter[2][51] ),
    .QN(_14335_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[52]$_DFFE_PN0P_  (.D(_02803_),
    .RN(net253),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.mhpmcounter[2][52] ),
    .QN(_14334_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[53]$_DFFE_PN0P_  (.D(_02804_),
    .RN(net253),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][53] ),
    .QN(_14333_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[54]$_DFFE_PN0P_  (.D(_02805_),
    .RN(net253),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][54] ),
    .QN(_14332_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[55]$_DFFE_PN0P_  (.D(_02806_),
    .RN(net253),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][55] ),
    .QN(_14331_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[56]$_DFFE_PN0P_  (.D(_02807_),
    .RN(net253),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][56] ),
    .QN(_14330_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[57]$_DFFE_PN0P_  (.D(_02808_),
    .RN(net253),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][57] ),
    .QN(_14329_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[58]$_DFFE_PN0P_  (.D(_02809_),
    .RN(net252),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][58] ),
    .QN(_14328_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[59]$_DFFE_PN0P_  (.D(_02810_),
    .RN(net253),
    .CK(clknet_leaf_105_clk),
    .Q(\cs_registers_i.mhpmcounter[2][59] ),
    .QN(_14327_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[5]$_DFFE_PN0P_  (.D(_02811_),
    .RN(net254),
    .CK(clknet_leaf_120_clk),
    .Q(\cs_registers_i.mhpmcounter[2][5] ),
    .QN(_14326_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[60]$_DFFE_PN0P_  (.D(_02812_),
    .RN(net252),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][60] ),
    .QN(_14325_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[61]$_DFFE_PN0P_  (.D(_02813_),
    .RN(net253),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][61] ),
    .QN(_14324_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[62]$_DFFE_PN0P_  (.D(_02814_),
    .RN(net252),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mhpmcounter[2][62] ),
    .QN(_14323_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[63]$_DFFE_PN0P_  (.D(_02815_),
    .RN(net252),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.mhpmcounter[2][63] ),
    .QN(_14322_));
 DFFR_X2 \cs_registers_i.minstret_counter_i.counter_q[6]$_DFFE_PN0P_  (.D(_02816_),
    .RN(net254),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mhpmcounter[2][6] ),
    .QN(_14321_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[7]$_DFFE_PN0P_  (.D(_02817_),
    .RN(net254),
    .CK(clknet_leaf_123_clk),
    .Q(\cs_registers_i.mhpmcounter[2][7] ),
    .QN(_14320_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[8]$_DFFE_PN0P_  (.D(_02818_),
    .RN(net630),
    .CK(clknet_leaf_122_clk),
    .Q(\cs_registers_i.mhpmcounter[2][8] ),
    .QN(_14319_));
 DFFR_X1 \cs_registers_i.minstret_counter_i.counter_q[9]$_DFFE_PN0P_  (.D(_02819_),
    .RN(net254),
    .CK(clknet_leaf_123_clk),
    .Q(\cs_registers_i.mhpmcounter[2][9] ),
    .QN(_14318_));
 DFFS_X1 \cs_registers_i.priv_lvl_q[0]$_DFFE_PN1P_  (.D(_02820_),
    .SN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.priv_lvl_q[0] ),
    .QN(_14317_));
 DFFS_X1 \cs_registers_i.priv_lvl_q[1]$_DFFE_PN1P_  (.D(_02821_),
    .SN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.priv_lvl_q[1] ),
    .QN(_15902_));
 DFFS_X2 \cs_registers_i.u_dcsr_csr.rdata_q[0]$_DFFE_PN1N_  (.D(_02822_),
    .SN(net253),
    .CK(clknet_leaf_112_clk),
    .Q(\cs_registers_i.dcsr_q[0] ),
    .QN(_14316_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02823_),
    .RN(net252),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.dcsr_q[11] ),
    .QN(_14315_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02824_),
    .RN(net253),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.dcsr_q[12] ),
    .QN(_00549_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02825_),
    .RN(net253),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.dcsr_q[13] ),
    .QN(_14314_));
 DFFR_X2 \cs_registers_i.u_dcsr_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02826_),
    .RN(net253),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.dcsr_q[15] ),
    .QN(_00556_));
 DFFS_X2 \cs_registers_i.u_dcsr_csr.rdata_q[1]$_DFFE_PN1N_  (.D(_02827_),
    .SN(net253),
    .CK(clknet_leaf_112_clk),
    .Q(\cs_registers_i.dcsr_q[1] ),
    .QN(_14313_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02828_),
    .RN(net248),
    .CK(clknet_leaf_116_clk),
    .Q(\cs_registers_i.dcsr_q[2] ),
    .QN(_01164_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02829_),
    .RN(net249),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.dcsr_q[6] ),
    .QN(_14312_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02830_),
    .RN(net248),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.dcsr_q[7] ),
    .QN(_14311_));
 DFFR_X1 \cs_registers_i.u_dcsr_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02831_),
    .RN(net249),
    .CK(clknet_leaf_114_clk),
    .Q(\cs_registers_i.dcsr_q[8] ),
    .QN(_14310_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02832_),
    .RN(net250),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.csr_depc_o[10] ),
    .QN(_14309_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02833_),
    .RN(net253),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.csr_depc_o[11] ),
    .QN(_14308_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02834_),
    .RN(net249),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.csr_depc_o[12] ),
    .QN(_14307_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02835_),
    .RN(net249),
    .CK(clknet_leaf_114_clk),
    .Q(\cs_registers_i.csr_depc_o[13] ),
    .QN(_14306_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02836_),
    .RN(net249),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.csr_depc_o[14] ),
    .QN(_14305_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02837_),
    .RN(net249),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.csr_depc_o[15] ),
    .QN(_14304_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02838_),
    .RN(net250),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.csr_depc_o[16] ),
    .QN(_14303_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02839_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.csr_depc_o[17] ),
    .QN(_14302_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02840_),
    .RN(net250),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_depc_o[18] ),
    .QN(_14301_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02841_),
    .RN(net250),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_depc_o[19] ),
    .QN(_14300_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02842_),
    .RN(net249),
    .CK(clknet_leaf_114_clk),
    .Q(\cs_registers_i.csr_depc_o[1] ),
    .QN(_00555_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02843_),
    .RN(net250),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_depc_o[20] ),
    .QN(_14299_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02844_),
    .RN(net250),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.csr_depc_o[21] ),
    .QN(_14298_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02845_),
    .RN(net251),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.csr_depc_o[22] ),
    .QN(_14297_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02846_),
    .RN(net250),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.csr_depc_o[23] ),
    .QN(_14296_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02847_),
    .RN(net251),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.csr_depc_o[24] ),
    .QN(_14295_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_02848_),
    .RN(net250),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.csr_depc_o[25] ),
    .QN(_14294_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_02849_),
    .RN(net251),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.csr_depc_o[26] ),
    .QN(_14293_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_02850_),
    .RN(net250),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.csr_depc_o[27] ),
    .QN(_14292_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02851_),
    .RN(net250),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.csr_depc_o[28] ),
    .QN(_14291_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02852_),
    .RN(net250),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.csr_depc_o[29] ),
    .QN(_14290_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02853_),
    .RN(net250),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.csr_depc_o[2] ),
    .QN(_14289_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02854_),
    .RN(net250),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.csr_depc_o[30] ),
    .QN(_14288_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02855_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.csr_depc_o[31] ),
    .QN(_14287_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02856_),
    .RN(net253),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.csr_depc_o[3] ),
    .QN(_01165_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02857_),
    .RN(net253),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.csr_depc_o[4] ),
    .QN(_01166_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02858_),
    .RN(net249),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.csr_depc_o[5] ),
    .QN(_01167_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02859_),
    .RN(net249),
    .CK(clknet_leaf_114_clk),
    .Q(\cs_registers_i.csr_depc_o[6] ),
    .QN(_01168_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02860_),
    .RN(net249),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.csr_depc_o[7] ),
    .QN(_14286_));
 DFFR_X2 \cs_registers_i.u_depc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02861_),
    .RN(net250),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.csr_depc_o[8] ),
    .QN(_14285_));
 DFFR_X1 \cs_registers_i.u_depc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02862_),
    .RN(net249),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.csr_depc_o[9] ),
    .QN(_14284_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02863_),
    .RN(net252),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.dscratch0_q[0] ),
    .QN(_14283_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02864_),
    .RN(net251),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch0_q[10] ),
    .QN(_14282_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02865_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch0_q[11] ),
    .QN(_14281_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02866_),
    .RN(net252),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.dscratch0_q[12] ),
    .QN(_14280_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02867_),
    .RN(net252),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.dscratch0_q[13] ),
    .QN(_14279_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02868_),
    .RN(net250),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.dscratch0_q[14] ),
    .QN(_14278_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02869_),
    .RN(net253),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.dscratch0_q[15] ),
    .QN(_14277_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02870_),
    .RN(net251),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.dscratch0_q[16] ),
    .QN(_14276_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02871_),
    .RN(net250),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.dscratch0_q[17] ),
    .QN(_14275_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02872_),
    .RN(net252),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.dscratch0_q[18] ),
    .QN(_14274_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02873_),
    .RN(net253),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.dscratch0_q[19] ),
    .QN(_14273_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02874_),
    .RN(net253),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.dscratch0_q[1] ),
    .QN(_14272_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02875_),
    .RN(net252),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.dscratch0_q[20] ),
    .QN(_14271_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02876_),
    .RN(net252),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch0_q[21] ),
    .QN(_14270_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02877_),
    .RN(net252),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch0_q[22] ),
    .QN(_14269_));
 DFFR_X2 \cs_registers_i.u_dscratch0_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02878_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch0_q[23] ),
    .QN(_14268_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02879_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch0_q[24] ),
    .QN(_14267_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_02880_),
    .RN(net251),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch0_q[25] ),
    .QN(_14266_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_02881_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch0_q[26] ),
    .QN(_14265_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_02882_),
    .RN(net251),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch0_q[27] ),
    .QN(_14264_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02883_),
    .RN(net251),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.dscratch0_q[28] ),
    .QN(_14263_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02884_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch0_q[29] ),
    .QN(_14262_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02885_),
    .RN(net252),
    .CK(clknet_leaf_103_clk),
    .Q(\cs_registers_i.dscratch0_q[2] ),
    .QN(_14261_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02886_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch0_q[30] ),
    .QN(_14260_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02887_),
    .RN(net251),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch0_q[31] ),
    .QN(_14259_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02888_),
    .RN(net252),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.dscratch0_q[3] ),
    .QN(_14258_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02889_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch0_q[4] ),
    .QN(_14257_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02890_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch0_q[5] ),
    .QN(_14256_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02891_),
    .RN(net252),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.dscratch0_q[6] ),
    .QN(_14255_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02892_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch0_q[7] ),
    .QN(_14254_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02893_),
    .RN(net252),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.dscratch0_q[8] ),
    .QN(_14253_));
 DFFR_X1 \cs_registers_i.u_dscratch0_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02894_),
    .RN(net252),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.dscratch0_q[9] ),
    .QN(_14252_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02895_),
    .RN(net252),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.dscratch1_q[0] ),
    .QN(_14251_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02896_),
    .RN(net251),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch1_q[10] ),
    .QN(_14250_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02897_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch1_q[11] ),
    .QN(_14249_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02898_),
    .RN(net252),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.dscratch1_q[12] ),
    .QN(_14248_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02899_),
    .RN(net252),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.dscratch1_q[13] ),
    .QN(_14247_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02900_),
    .RN(net253),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.dscratch1_q[14] ),
    .QN(_14246_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02901_),
    .RN(net253),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.dscratch1_q[15] ),
    .QN(_14245_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02902_),
    .RN(net251),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.dscratch1_q[16] ),
    .QN(_14244_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02903_),
    .RN(net250),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.dscratch1_q[17] ),
    .QN(_14243_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02904_),
    .RN(net250),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.dscratch1_q[18] ),
    .QN(_14242_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02905_),
    .RN(net253),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.dscratch1_q[19] ),
    .QN(_14241_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02906_),
    .RN(net252),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.dscratch1_q[1] ),
    .QN(_14240_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02907_),
    .RN(net252),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch1_q[20] ),
    .QN(_14239_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02908_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch1_q[21] ),
    .QN(_14238_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02909_),
    .RN(net252),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch1_q[22] ),
    .QN(_14237_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02910_),
    .RN(net252),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.dscratch1_q[23] ),
    .QN(_14236_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02911_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch1_q[24] ),
    .QN(_14235_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_02912_),
    .RN(net251),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch1_q[25] ),
    .QN(_14234_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_02913_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch1_q[26] ),
    .QN(_14233_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_02914_),
    .RN(net251),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.dscratch1_q[27] ),
    .QN(_14232_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02915_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch1_q[28] ),
    .QN(_14231_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02916_),
    .RN(net251),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.dscratch1_q[29] ),
    .QN(_14230_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02917_),
    .RN(net252),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.dscratch1_q[2] ),
    .QN(_14229_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02918_),
    .RN(net251),
    .CK(clknet_leaf_89_clk),
    .Q(\cs_registers_i.dscratch1_q[30] ),
    .QN(_14228_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02919_),
    .RN(net252),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.dscratch1_q[31] ),
    .QN(_14227_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02920_),
    .RN(net252),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.dscratch1_q[3] ),
    .QN(_14226_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02921_),
    .RN(net252),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.dscratch1_q[4] ),
    .QN(_14225_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02922_),
    .RN(net252),
    .CK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.dscratch1_q[5] ),
    .QN(_14224_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02923_),
    .RN(net251),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.dscratch1_q[6] ),
    .QN(_14223_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02924_),
    .RN(net251),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.dscratch1_q[7] ),
    .QN(_14222_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02925_),
    .RN(net251),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.dscratch1_q[8] ),
    .QN(_14221_));
 DFFR_X1 \cs_registers_i.u_dscratch1_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02926_),
    .RN(net252),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.dscratch1_q[9] ),
    .QN(_14220_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02927_),
    .RN(net249),
    .CK(clknet_leaf_112_clk),
    .Q(\cs_registers_i.mcause_q[0] ),
    .QN(_14219_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02928_),
    .RN(net249),
    .CK(clknet_leaf_113_clk),
    .Q(\cs_registers_i.mcause_q[1] ),
    .QN(_14218_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02929_),
    .RN(net253),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mcause_q[2] ),
    .QN(_14217_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02930_),
    .RN(net253),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mcause_q[3] ),
    .QN(_14216_));
 DFFR_X1 \cs_registers_i.u_mcause_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02931_),
    .RN(net253),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mcause_q[4] ),
    .QN(_14215_));
 DFFR_X2 \cs_registers_i.u_mcause_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02932_),
    .RN(net249),
    .CK(clknet_leaf_113_clk),
    .Q(\cs_registers_i.mcause_q[5] ),
    .QN(_14214_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02933_),
    .RN(net249),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.csr_mepc_o[0] ),
    .QN(_14213_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02934_),
    .RN(net250),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.csr_mepc_o[10] ),
    .QN(_14212_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02935_),
    .RN(net253),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.csr_mepc_o[11] ),
    .QN(_14211_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02936_),
    .RN(net250),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.csr_mepc_o[12] ),
    .QN(_14210_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02937_),
    .RN(net249),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.csr_mepc_o[13] ),
    .QN(_14209_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02938_),
    .RN(net249),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.csr_mepc_o[14] ),
    .QN(_14208_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02939_),
    .RN(net249),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.csr_mepc_o[15] ),
    .QN(_14207_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02940_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.csr_mepc_o[16] ),
    .QN(_14206_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02941_),
    .RN(net250),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.csr_mepc_o[17] ),
    .QN(_14205_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02942_),
    .RN(net250),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mepc_o[18] ),
    .QN(_14204_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02943_),
    .RN(net250),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.csr_mepc_o[19] ),
    .QN(_14203_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02944_),
    .RN(net253),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.csr_mepc_o[1] ),
    .QN(_14202_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02945_),
    .RN(net251),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.csr_mepc_o[20] ),
    .QN(_14201_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02946_),
    .RN(net250),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.csr_mepc_o[21] ),
    .QN(_14200_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02947_),
    .RN(net251),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.csr_mepc_o[22] ),
    .QN(_14199_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02948_),
    .RN(net250),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.csr_mepc_o[23] ),
    .QN(_14198_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02949_),
    .RN(net251),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.csr_mepc_o[24] ),
    .QN(_14197_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_02950_),
    .RN(net251),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.csr_mepc_o[25] ),
    .QN(_14196_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_02951_),
    .RN(net251),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.csr_mepc_o[26] ),
    .QN(_14195_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_02952_),
    .RN(net250),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.csr_mepc_o[27] ),
    .QN(_14194_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_02953_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.csr_mepc_o[28] ),
    .QN(_14193_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_02954_),
    .RN(net250),
    .CK(clknet_leaf_76_clk),
    .Q(\cs_registers_i.csr_mepc_o[29] ),
    .QN(_14192_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02955_),
    .RN(net250),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.csr_mepc_o[2] ),
    .QN(_14191_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_02956_),
    .RN(net251),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.csr_mepc_o[30] ),
    .QN(_14190_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_02957_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.csr_mepc_o[31] ),
    .QN(_14189_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02958_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.csr_mepc_o[3] ),
    .QN(_14188_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02959_),
    .RN(net253),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.csr_mepc_o[4] ),
    .QN(_14187_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02960_),
    .RN(net249),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.csr_mepc_o[5] ),
    .QN(_14186_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02961_),
    .RN(net249),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.csr_mepc_o[6] ),
    .QN(_14185_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02962_),
    .RN(net253),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.csr_mepc_o[7] ),
    .QN(_14184_));
 DFFR_X2 \cs_registers_i.u_mepc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02963_),
    .RN(net250),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.csr_mepc_o[8] ),
    .QN(_14183_));
 DFFR_X1 \cs_registers_i.u_mepc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02964_),
    .RN(net249),
    .CK(clknet_leaf_114_clk),
    .Q(\cs_registers_i.csr_mepc_o[9] ),
    .QN(_14182_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02965_),
    .RN(net251),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mie_q[0] ),
    .QN(_14181_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02966_),
    .RN(net251),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mie_q[10] ),
    .QN(_14180_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02967_),
    .RN(net251),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mie_q[11] ),
    .QN(_14179_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02968_),
    .RN(net252),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mie_q[12] ),
    .QN(_14178_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02969_),
    .RN(net252),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mie_q[13] ),
    .QN(_14177_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02970_),
    .RN(net251),
    .CK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.mie_q[14] ),
    .QN(_14176_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02971_),
    .RN(net252),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mie_q[15] ),
    .QN(_14175_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02972_),
    .RN(net251),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mie_q[16] ),
    .QN(_14174_));
 DFFR_X1 \cs_registers_i.u_mie_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02973_),
    .RN(net252),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mie_q[17] ),
    .QN(_14173_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02974_),
    .RN(net252),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mie_q[1] ),
    .QN(_14172_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_02975_),
    .RN(net251),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mie_q[2] ),
    .QN(_14171_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_02976_),
    .RN(net253),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mie_q[3] ),
    .QN(_14170_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_02977_),
    .RN(net252),
    .CK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mie_q[4] ),
    .QN(_14169_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_02978_),
    .RN(net253),
    .CK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mie_q[5] ),
    .QN(_14168_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_02979_),
    .RN(net252),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mie_q[6] ),
    .QN(_14167_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_02980_),
    .RN(net253),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mie_q[7] ),
    .QN(_14166_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_02981_),
    .RN(net251),
    .CK(clknet_leaf_101_clk),
    .Q(\cs_registers_i.mie_q[8] ),
    .QN(_14165_));
 DFFR_X2 \cs_registers_i.u_mie_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_02982_),
    .RN(net251),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mie_q[9] ),
    .QN(_14164_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_02983_),
    .RN(net249),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mscratch_q[0] ),
    .QN(_14163_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_02984_),
    .RN(net252),
    .CK(clknet_leaf_92_clk),
    .Q(\cs_registers_i.mscratch_q[10] ),
    .QN(_14162_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_02985_),
    .RN(net253),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mscratch_q[11] ),
    .QN(_14161_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_02986_),
    .RN(net250),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[12] ),
    .QN(_14160_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_02987_),
    .RN(net249),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mscratch_q[13] ),
    .QN(_14159_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_02988_),
    .RN(net253),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mscratch_q[14] ),
    .QN(_14158_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_02989_),
    .RN(net253),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.mscratch_q[15] ),
    .QN(_14157_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_02990_),
    .RN(net250),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[16] ),
    .QN(_14156_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_02991_),
    .RN(net250),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mscratch_q[17] ),
    .QN(_14155_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_02992_),
    .RN(net252),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mscratch_q[18] ),
    .QN(_14154_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_02993_),
    .RN(net249),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mscratch_q[19] ),
    .QN(_14153_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_02994_),
    .RN(net249),
    .CK(clknet_leaf_99_clk),
    .Q(\cs_registers_i.mscratch_q[1] ),
    .QN(_14152_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_02995_),
    .RN(net252),
    .CK(clknet_leaf_90_clk),
    .Q(\cs_registers_i.mscratch_q[20] ),
    .QN(_14151_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_02996_),
    .RN(net250),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[21] ),
    .QN(_14150_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_02997_),
    .RN(net252),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[22] ),
    .QN(_14149_));
 DFFR_X2 \cs_registers_i.u_mscratch_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_02998_),
    .RN(net250),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mscratch_q[23] ),
    .QN(_14148_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_02999_),
    .RN(net251),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mscratch_q[24] ),
    .QN(_14147_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_03000_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mscratch_q[25] ),
    .QN(_14146_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_03001_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mscratch_q[26] ),
    .QN(_14145_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_03002_),
    .RN(net251),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mscratch_q[27] ),
    .QN(_14144_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_03003_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mscratch_q[28] ),
    .QN(_14143_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_03004_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mscratch_q[29] ),
    .QN(_14142_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_03005_),
    .RN(net253),
    .CK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mscratch_q[2] ),
    .QN(_14141_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_03006_),
    .RN(net251),
    .CK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mscratch_q[30] ),
    .QN(_14140_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_03007_),
    .RN(net252),
    .CK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[31] ),
    .QN(_14139_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_03008_),
    .RN(net250),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mscratch_q[3] ),
    .QN(_14138_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_03009_),
    .RN(net250),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mscratch_q[4] ),
    .QN(_14137_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_03010_),
    .RN(net250),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mscratch_q[5] ),
    .QN(_14136_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_03011_),
    .RN(net253),
    .CK(clknet_leaf_108_clk),
    .Q(\cs_registers_i.mscratch_q[6] ),
    .QN(_14135_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_03012_),
    .RN(net249),
    .CK(clknet_leaf_112_clk),
    .Q(\cs_registers_i.mscratch_q[7] ),
    .QN(_14134_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_03013_),
    .RN(net249),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mscratch_q[8] ),
    .QN(_14133_));
 DFFR_X1 \cs_registers_i.u_mscratch_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_03014_),
    .RN(net252),
    .CK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mscratch_q[9] ),
    .QN(_14132_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_03015_),
    .RN(net249),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mstack_cause_q[0] ),
    .QN(_14131_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_03016_),
    .RN(net249),
    .CK(clknet_leaf_113_clk),
    .Q(\cs_registers_i.mstack_cause_q[1] ),
    .QN(_14130_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_03017_),
    .RN(net253),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mstack_cause_q[2] ),
    .QN(_14129_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_03018_),
    .RN(net253),
    .CK(clknet_leaf_97_clk),
    .Q(\cs_registers_i.mstack_cause_q[3] ),
    .QN(_14128_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_03019_),
    .RN(net249),
    .CK(clknet_leaf_113_clk),
    .Q(\cs_registers_i.mstack_cause_q[4] ),
    .QN(_14127_));
 DFFR_X1 \cs_registers_i.u_mstack_cause_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_03020_),
    .RN(net249),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mstack_cause_q[5] ),
    .QN(_14126_));
 DFFR_X1 \cs_registers_i.u_mstack_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_03021_),
    .RN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.mstack_q[0] ),
    .QN(_14125_));
 DFFR_X1 \cs_registers_i.u_mstack_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_03022_),
    .RN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.mstack_q[1] ),
    .QN(_14124_));
 DFFS_X1 \cs_registers_i.u_mstack_csr.rdata_q[2]$_DFFE_PN1P_  (.D(_03023_),
    .SN(net249),
    .CK(clknet_leaf_112_clk),
    .Q(\cs_registers_i.mstack_q[2] ),
    .QN(_14123_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_03024_),
    .RN(net249),
    .CK(clknet_leaf_113_clk),
    .Q(\cs_registers_i.mstack_epc_q[0] ),
    .QN(_14122_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_03025_),
    .RN(net250),
    .CK(clknet_leaf_77_clk),
    .Q(\cs_registers_i.mstack_epc_q[10] ),
    .QN(_14121_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_03026_),
    .RN(net253),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.mstack_epc_q[11] ),
    .QN(_14120_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_03027_),
    .RN(net250),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.mstack_epc_q[12] ),
    .QN(_14119_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_03028_),
    .RN(net249),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mstack_epc_q[13] ),
    .QN(_14118_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_03029_),
    .RN(net249),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mstack_epc_q[14] ),
    .QN(_14117_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_03030_),
    .RN(net249),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.mstack_epc_q[15] ),
    .QN(_14116_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_03031_),
    .RN(net250),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mstack_epc_q[16] ),
    .QN(_14115_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_03032_),
    .RN(net250),
    .CK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mstack_epc_q[17] ),
    .QN(_14114_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_03033_),
    .RN(net250),
    .CK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.mstack_epc_q[18] ),
    .QN(_14113_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_03034_),
    .RN(net250),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mstack_epc_q[19] ),
    .QN(_14112_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_03035_),
    .RN(net253),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mstack_epc_q[1] ),
    .QN(_14111_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_03036_),
    .RN(net251),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mstack_epc_q[20] ),
    .QN(_14110_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_03037_),
    .RN(net250),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mstack_epc_q[21] ),
    .QN(_14109_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_03038_),
    .RN(net251),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mstack_epc_q[22] ),
    .QN(_14108_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_03039_),
    .RN(net250),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mstack_epc_q[23] ),
    .QN(_14107_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_03040_),
    .RN(net251),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.mstack_epc_q[24] ),
    .QN(_14106_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_03041_),
    .RN(net251),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.mstack_epc_q[25] ),
    .QN(_14105_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_03042_),
    .RN(net251),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.mstack_epc_q[26] ),
    .QN(_14104_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_03043_),
    .RN(net250),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mstack_epc_q[27] ),
    .QN(_14103_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_03044_),
    .RN(net251),
    .CK(clknet_leaf_86_clk),
    .Q(\cs_registers_i.mstack_epc_q[28] ),
    .QN(_14102_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_03045_),
    .RN(net250),
    .CK(clknet_leaf_75_clk),
    .Q(\cs_registers_i.mstack_epc_q[29] ),
    .QN(_14101_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_03046_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.mstack_epc_q[2] ),
    .QN(_14100_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_03047_),
    .RN(net251),
    .CK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mstack_epc_q[30] ),
    .QN(_14099_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_03048_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.mstack_epc_q[31] ),
    .QN(_14098_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_03049_),
    .RN(net250),
    .CK(clknet_leaf_82_clk),
    .Q(\cs_registers_i.mstack_epc_q[3] ),
    .QN(_14097_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_03050_),
    .RN(net253),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mstack_epc_q[4] ),
    .QN(_14096_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_03051_),
    .RN(net249),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.mstack_epc_q[5] ),
    .QN(_14095_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_03052_),
    .RN(net249),
    .CK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mstack_epc_q[6] ),
    .QN(_14094_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_03053_),
    .RN(net253),
    .CK(clknet_leaf_81_clk),
    .Q(\cs_registers_i.mstack_epc_q[7] ),
    .QN(_14093_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_03054_),
    .RN(net250),
    .CK(clknet_leaf_80_clk),
    .Q(\cs_registers_i.mstack_epc_q[8] ),
    .QN(_14092_));
 DFFR_X1 \cs_registers_i.u_mstack_epc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_03055_),
    .RN(net249),
    .CK(clknet_leaf_114_clk),
    .Q(\cs_registers_i.mstack_epc_q[9] ),
    .QN(_14091_));
 DFFR_X2 \cs_registers_i.u_mstatus_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_03056_),
    .RN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.csr_mstatus_tw_o ),
    .QN(_14090_));
 DFFR_X1 \cs_registers_i.u_mstatus_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_03057_),
    .RN(net249),
    .CK(clknet_leaf_111_clk),
    .Q(\cs_registers_i.mstatus_q[1] ),
    .QN(_14089_));
 DFFR_X1 \cs_registers_i.u_mstatus_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_03058_),
    .RN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.mstack_d[0] ),
    .QN(_14088_));
 DFFR_X1 \cs_registers_i.u_mstatus_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_03059_),
    .RN(net248),
    .CK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.mstack_d[1] ),
    .QN(_14087_));
 DFFS_X2 \cs_registers_i.u_mstatus_csr.rdata_q[4]$_DFFE_PN1P_  (.D(_03060_),
    .SN(net249),
    .CK(clknet_leaf_112_clk),
    .Q(\cs_registers_i.mstack_d[2] ),
    .QN(_14086_));
 DFFR_X2 \cs_registers_i.u_mstatus_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_03061_),
    .RN(net249),
    .CK(clknet_leaf_113_clk),
    .Q(\cs_registers_i.csr_mstatus_mie_o ),
    .QN(_14085_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_03062_),
    .RN(net248),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mtval_q[0] ),
    .QN(_14084_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_03063_),
    .RN(net248),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.mtval_q[10] ),
    .QN(_14083_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_03064_),
    .RN(net249),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mtval_q[11] ),
    .QN(_14082_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_03065_),
    .RN(net248),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.mtval_q[12] ),
    .QN(_14081_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_03066_),
    .RN(net248),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.mtval_q[13] ),
    .QN(_14080_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_03067_),
    .RN(net249),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mtval_q[14] ),
    .QN(_14079_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_03068_),
    .RN(net248),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.mtval_q[15] ),
    .QN(_14078_));
 DFFR_X2 \cs_registers_i.u_mtval_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_03069_),
    .RN(net249),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.mtval_q[16] ),
    .QN(_14077_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_03070_),
    .RN(net249),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mtval_q[17] ),
    .QN(_14076_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_03071_),
    .RN(net248),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mtval_q[18] ),
    .QN(_14075_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_03072_),
    .RN(net248),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.mtval_q[19] ),
    .QN(_14074_));
 DFFR_X2 \cs_registers_i.u_mtval_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_03073_),
    .RN(net248),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.mtval_q[1] ),
    .QN(_14073_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_03074_),
    .RN(net249),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mtval_q[20] ),
    .QN(_14072_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_03075_),
    .RN(net249),
    .CK(clknet_leaf_62_clk),
    .Q(\cs_registers_i.mtval_q[21] ),
    .QN(_14071_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_03076_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[22] ),
    .QN(_14070_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_03077_),
    .RN(net248),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.mtval_q[23] ),
    .QN(_14069_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_03078_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[24] ),
    .QN(_14068_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_03079_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[25] ),
    .QN(_14067_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_03080_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mtval_q[26] ),
    .QN(_14066_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_03081_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mtval_q[27] ),
    .QN(_14065_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_03082_),
    .RN(net251),
    .CK(clknet_leaf_87_clk),
    .Q(\cs_registers_i.mtval_q[28] ),
    .QN(_14064_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_03083_),
    .RN(net249),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mtval_q[29] ),
    .QN(_14063_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_03084_),
    .RN(net248),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mtval_q[2] ),
    .QN(_14062_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_03085_),
    .RN(net250),
    .CK(clknet_leaf_83_clk),
    .Q(\cs_registers_i.mtval_q[30] ),
    .QN(_14061_));
 DFFR_X2 \cs_registers_i.u_mtval_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_03086_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[31] ),
    .QN(_14060_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_03087_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.mtval_q[3] ),
    .QN(_14059_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_03088_),
    .RN(net253),
    .CK(clknet_leaf_96_clk),
    .Q(\cs_registers_i.mtval_q[4] ),
    .QN(_14058_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_03089_),
    .RN(net250),
    .CK(clknet_leaf_94_clk),
    .Q(\cs_registers_i.mtval_q[5] ),
    .QN(_14057_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_03090_),
    .RN(net249),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mtval_q[6] ),
    .QN(_14056_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_03091_),
    .RN(net248),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mtval_q[7] ),
    .QN(_14055_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_03092_),
    .RN(net248),
    .CK(clknet_leaf_115_clk),
    .Q(\cs_registers_i.mtval_q[8] ),
    .QN(_14054_));
 DFFR_X1 \cs_registers_i.u_mtval_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_03093_),
    .RN(net248),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.mtval_q[9] ),
    .QN(_14053_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_03094_),
    .RN(net250),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mtvec_o[10] ),
    .QN(_01171_));
 DFFR_X2 \cs_registers_i.u_mtvec_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_01186_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.csr_mtvec_o[11] ),
    .QN(_00551_));
 DFFR_X2 \cs_registers_i.u_mtvec_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_01187_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.csr_mtvec_o[12] ),
    .QN(_00550_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_01188_),
    .RN(net248),
    .CK(clknet_leaf_60_clk),
    .Q(\cs_registers_i.csr_mtvec_o[13] ),
    .QN(_01172_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_01189_),
    .RN(net249),
    .CK(clknet_leaf_63_clk),
    .Q(\cs_registers_i.csr_mtvec_o[14] ),
    .QN(_01173_));
 DFFR_X2 \cs_registers_i.u_mtvec_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_01190_),
    .RN(net249),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mtvec_o[15] ),
    .QN(_01174_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_01191_),
    .RN(net250),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mtvec_o[16] ),
    .QN(_01175_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_01192_),
    .RN(net250),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.csr_mtvec_o[17] ),
    .QN(_01176_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_01193_),
    .RN(net250),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[18] ),
    .QN(_01177_));
 DFFR_X2 \cs_registers_i.u_mtvec_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_01194_),
    .RN(net250),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_mtvec_o[19] ),
    .QN(_01178_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_01195_),
    .RN(net250),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_mtvec_o[20] ),
    .QN(_01179_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_01196_),
    .RN(net250),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[21] ),
    .QN(_01180_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_01197_),
    .RN(net250),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[22] ),
    .QN(_01181_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_01198_),
    .RN(net250),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[23] ),
    .QN(_01182_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_01199_),
    .RN(net250),
    .CK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[24] ),
    .QN(_01183_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_01200_),
    .RN(net250),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[25] ),
    .QN(_01184_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_01201_),
    .RN(net250),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_mtvec_o[26] ),
    .QN(_01185_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_01202_),
    .RN(net250),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[27] ),
    .QN(_00007_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_01203_),
    .RN(net250),
    .CK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_mtvec_o[28] ),
    .QN(_00008_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_01204_),
    .RN(net250),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[29] ),
    .QN(_00009_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_01205_),
    .RN(net250),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[30] ),
    .QN(_00010_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_01206_),
    .RN(net250),
    .CK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.csr_mtvec_o[31] ),
    .QN(_00011_));
 DFFR_X2 \cs_registers_i.u_mtvec_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_01207_),
    .RN(net250),
    .CK(clknet_leaf_79_clk),
    .Q(\cs_registers_i.csr_mtvec_o[8] ),
    .QN(_01169_));
 DFFR_X1 \cs_registers_i.u_mtvec_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_01208_),
    .RN(net248),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.csr_mtvec_o[9] ),
    .QN(_01170_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.D(_01209_),
    .RN(net246),
    .CK(clknet_leaf_41_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .QN(_14052_));
 DFFR_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.D(_01210_),
    .RN(net246),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .QN(_15940_));
 DFFR_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.D(_01211_),
    .RN(net246),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .QN(_15941_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.D(_01212_),
    .RN(net246),
    .CK(clknet_leaf_38_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .QN(_00066_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.D(_01213_),
    .RN(net246),
    .CK(clknet_leaf_38_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .QN(_00067_));
 DFFR_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.D(_01214_),
    .RN(net246),
    .CK(clknet_leaf_38_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .QN(_01162_));
 DFFS_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.D(_00000_),
    .SN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .QN(_14451_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.D(_00001_),
    .RN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .QN(_01163_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.D(_00002_),
    .RN(net246),
    .CK(clknet_leaf_39_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .QN(_14452_));
 DFFR_X2 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.D(_00003_),
    .RN(net246),
    .CK(clknet_leaf_42_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .QN(_14453_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.D(_00004_),
    .RN(net246),
    .CK(clknet_leaf_39_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .QN(_00178_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.D(_00005_),
    .RN(net246),
    .CK(clknet_leaf_39_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .QN(_14051_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.D(_01215_),
    .RN(net247),
    .CK(clknet_leaf_35_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .QN(_00101_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.D(_01216_),
    .RN(net247),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .QN(_00111_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.D(_01217_),
    .RN(net247),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .QN(_00110_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.D(_01218_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .QN(_00113_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.D(_01219_),
    .RN(net247),
    .CK(clknet_leaf_35_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .QN(_00112_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.D(_01220_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .QN(_00115_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.D(_01221_),
    .RN(net247),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .QN(_00114_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.D(_01222_),
    .RN(net247),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .QN(_00117_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.D(_01223_),
    .RN(net247),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .QN(_00116_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.D(_01224_),
    .RN(net247),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .QN(_00119_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.D(_01225_),
    .RN(net247),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .QN(_00118_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.D(_01226_),
    .RN(net247),
    .CK(clknet_leaf_35_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .QN(_00100_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.D(_01227_),
    .RN(net247),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .QN(_00121_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.D(_01228_),
    .RN(net247),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .QN(_00120_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.D(_01229_),
    .RN(net247),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .QN(_00123_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.D(_01230_),
    .RN(net247),
    .CK(clknet_leaf_34_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .QN(_00122_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.D(_01231_),
    .RN(net247),
    .CK(clknet_leaf_34_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .QN(_00125_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.D(_01232_),
    .RN(net247),
    .CK(clknet_leaf_34_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .QN(_00124_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.D(_01233_),
    .RN(net247),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .QN(_00127_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.D(_01234_),
    .RN(net247),
    .CK(clknet_leaf_34_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .QN(_00126_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.D(_01235_),
    .RN(net246),
    .CK(clknet_leaf_34_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .QN(_00129_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.D(_01236_),
    .RN(net247),
    .CK(clknet_leaf_34_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .QN(_00128_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.D(_01237_),
    .RN(net247),
    .CK(clknet_leaf_35_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .QN(_00103_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.D(_01238_),
    .RN(net246),
    .CK(clknet_leaf_34_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .QN(_00131_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.D(_01239_),
    .RN(net247),
    .CK(clknet_leaf_35_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .QN(_00130_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.D(_01240_),
    .RN(net247),
    .CK(clknet_leaf_35_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .QN(_00102_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.D(_01241_),
    .RN(net246),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .QN(_00105_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.D(_01242_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .QN(_00104_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.D(_01243_),
    .RN(net246),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .QN(_00107_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.D(_01244_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .QN(_00106_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.D(_01245_),
    .RN(net247),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .QN(_00109_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.D(_01246_),
    .RN(net247),
    .CK(clknet_leaf_32_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .QN(_00108_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.D(_01247_),
    .RN(net246),
    .CK(clknet_leaf_43_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .QN(_00068_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.D(_01248_),
    .RN(net246),
    .CK(clknet_leaf_44_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .QN(_00078_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.D(_01249_),
    .RN(net246),
    .CK(clknet_leaf_44_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .QN(_00079_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.D(_01250_),
    .RN(net246),
    .CK(clknet_leaf_43_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .QN(_00080_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.D(_01251_),
    .RN(net246),
    .CK(clknet_leaf_43_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .QN(_00081_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.D(_01252_),
    .RN(net246),
    .CK(clknet_leaf_43_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .QN(_00082_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.D(_01253_),
    .RN(net246),
    .CK(clknet_leaf_44_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .QN(_00083_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.D(_01254_),
    .RN(net246),
    .CK(clknet_leaf_43_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .QN(_00084_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.D(_01255_),
    .RN(net246),
    .CK(clknet_leaf_38_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .QN(_00085_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.D(_01256_),
    .RN(net246),
    .CK(clknet_leaf_38_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .QN(_00086_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.D(_01257_),
    .RN(net246),
    .CK(clknet_leaf_38_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .QN(_00087_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.D(_01258_),
    .RN(net246),
    .CK(clknet_leaf_38_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .QN(_00069_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.D(_01259_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .QN(_00088_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.D(_01260_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .QN(_00089_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.D(_01261_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .QN(_00090_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.D(_01262_),
    .RN(net246),
    .CK(clknet_leaf_39_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .QN(_00091_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.D(_01263_),
    .RN(net246),
    .CK(clknet_leaf_36_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .QN(_00092_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.D(_01264_),
    .RN(net246),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .QN(_00093_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.D(_01265_),
    .RN(net246),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .QN(_00094_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.D(_01266_),
    .RN(net246),
    .CK(clknet_leaf_37_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .QN(_00095_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.D(_01267_),
    .RN(net246),
    .CK(clknet_leaf_42_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .QN(_00096_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.D(_01268_),
    .RN(net246),
    .CK(clknet_leaf_41_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .QN(_00097_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.D(_01269_),
    .RN(net246),
    .CK(clknet_leaf_45_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .QN(_00070_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.D(_01270_),
    .RN(net246),
    .CK(clknet_leaf_42_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .QN(_00098_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.D(_01271_),
    .RN(net246),
    .CK(clknet_leaf_42_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .QN(_00099_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.D(_01272_),
    .RN(net246),
    .CK(clknet_leaf_43_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .QN(_00071_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.D(_01273_),
    .RN(net246),
    .CK(clknet_leaf_42_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .QN(_00072_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.D(_01274_),
    .RN(net246),
    .CK(clknet_leaf_41_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .QN(_00073_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.D(_01275_),
    .RN(net246),
    .CK(clknet_leaf_45_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .QN(_00074_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.D(_01276_),
    .RN(net246),
    .CK(clknet_leaf_45_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .QN(_00075_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.D(_01277_),
    .RN(net246),
    .CK(clknet_leaf_42_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .QN(_00076_));
 DFFR_X1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.D(_01278_),
    .RN(net246),
    .CK(clknet_leaf_42_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .QN(_00077_));
 DFFR_X1 \fetch_enable_q$_DFFE_PN0P_  (.D(_01279_),
    .RN(net144),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(fetch_enable_q),
    .QN(_14050_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[0]$_DFFE_PN0P_  (.D(_01280_),
    .RN(net267),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .QN(_14049_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[100]$_DFFE_PN0P_  (.D(_01281_),
    .RN(net264),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .QN(_00311_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[101]$_DFFE_PN0P_  (.D(_01282_),
    .RN(net267),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .QN(_00341_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[102]$_DFFE_PN0P_  (.D(_01283_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .QN(_00371_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[103]$_DFFE_PN0P_  (.D(_01284_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .QN(_00401_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[104]$_DFFE_PN0P_  (.D(_01285_),
    .RN(net268),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .QN(_00431_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[105]$_DFFE_PN0P_  (.D(_01286_),
    .RN(net267),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .QN(_00461_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[106]$_DFFE_PN0P_  (.D(_01287_),
    .RN(net262),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .QN(_00491_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[107]$_DFFE_PN0P_  (.D(_01288_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .QN(_00521_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[108]$_DFFE_PN0P_  (.D(_01289_),
    .RN(net261),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .QN(_00220_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[109]$_DFFE_PN0P_  (.D(_01290_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .QN(_00571_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[10]$_DFFE_PN0P_  (.D(_01291_),
    .RN(net262),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .QN(_14048_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[110]$_DFFE_PN0P_  (.D(_01292_),
    .RN(net255),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .QN(_00602_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[111]$_DFFE_PN0P_  (.D(_01293_),
    .RN(net255),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .QN(_00633_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[112]$_DFFE_PN0P_  (.D(_01294_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .QN(_00664_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[113]$_DFFE_PN0P_  (.D(_01295_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .QN(_00695_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[114]$_DFFE_PN0P_  (.D(_01296_),
    .RN(net255),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .QN(_00726_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[115]$_DFFE_PN0P_  (.D(_01297_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .QN(_00757_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[116]$_DFFE_PN0P_  (.D(_01298_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .QN(_00788_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[117]$_DFFE_PN0P_  (.D(_01299_),
    .RN(net260),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .QN(_00819_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[118]$_DFFE_PN0P_  (.D(_01300_),
    .RN(net260),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .QN(_00850_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[119]$_DFFE_PN0P_  (.D(_01301_),
    .RN(net261),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .QN(_00881_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[11]$_DFFE_PN0P_  (.D(_01302_),
    .RN(net268),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .QN(_14047_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[120]$_DFFE_PN0P_  (.D(_01303_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .QN(_00912_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[121]$_DFFE_PN0P_  (.D(_01304_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .QN(_00943_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[122]$_DFFE_PN0P_  (.D(_01305_),
    .RN(net257),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .QN(_00974_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[123]$_DFFE_PN0P_  (.D(_01306_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .QN(_01005_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[124]$_DFFE_PN0P_  (.D(_01307_),
    .RN(net258),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .QN(_01036_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[125]$_DFFE_PN0P_  (.D(_01308_),
    .RN(net262),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .QN(_01067_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[126]$_DFFE_PN0P_  (.D(_01309_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .QN(_01098_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[127]$_DFFE_PN0P_  (.D(_01310_),
    .RN(net266),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .QN(_01129_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[128]$_DFFE_PN0P_  (.D(_01311_),
    .RN(net267),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .QN(_00189_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[129]$_DFFE_PN0P_  (.D(_01312_),
    .RN(net266),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .QN(_00144_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[12]$_DFFE_PN0P_  (.D(_01313_),
    .RN(net260),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .QN(_14046_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[130]$_DFFE_PN0P_  (.D(_01314_),
    .RN(net267),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .QN(_00251_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[131]$_DFFE_PN0P_  (.D(_01315_),
    .RN(net267),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .QN(_00282_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[132]$_DFFE_PN0P_  (.D(_01316_),
    .RN(net264),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .QN(_00312_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[133]$_DFFE_PN0P_  (.D(_01317_),
    .RN(net264),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .QN(_00342_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[134]$_DFFE_PN0P_  (.D(_01318_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .QN(_00372_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[135]$_DFFE_PN0P_  (.D(_01319_),
    .RN(net268),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .QN(_00402_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[136]$_DFFE_PN0P_  (.D(_01320_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .QN(_00432_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[137]$_DFFE_PN0P_  (.D(_01321_),
    .RN(net268),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .QN(_00462_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[138]$_DFFE_PN0P_  (.D(_01322_),
    .RN(net262),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .QN(_00492_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[139]$_DFFE_PN0P_  (.D(_01323_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .QN(_00522_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[13]$_DFFE_PN0P_  (.D(_01324_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .QN(_14045_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[140]$_DFFE_PN0P_  (.D(_01325_),
    .RN(net261),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .QN(_00221_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[141]$_DFFE_PN0P_  (.D(_01326_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .QN(_00572_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[142]$_DFFE_PN0P_  (.D(_01327_),
    .RN(net255),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .QN(_00603_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[143]$_DFFE_PN0P_  (.D(_01328_),
    .RN(net255),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .QN(_00634_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[144]$_DFFE_PN0P_  (.D(_01329_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .QN(_00665_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[145]$_DFFE_PN0P_  (.D(_01330_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .QN(_00696_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[146]$_DFFE_PN0P_  (.D(_01331_),
    .RN(net255),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .QN(_00727_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[147]$_DFFE_PN0P_  (.D(_01332_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .QN(_00758_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[148]$_DFFE_PN0P_  (.D(_01333_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .QN(_00789_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[149]$_DFFE_PN0P_  (.D(_01334_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .QN(_00820_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[14]$_DFFE_PN0P_  (.D(_01335_),
    .RN(net261),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .QN(_14044_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[150]$_DFFE_PN0P_  (.D(_01336_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .QN(_00851_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[151]$_DFFE_PN0P_  (.D(_01337_),
    .RN(net259),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .QN(_00882_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[152]$_DFFE_PN0P_  (.D(_01338_),
    .RN(net258),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .QN(_00913_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[153]$_DFFE_PN0P_  (.D(_01339_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .QN(_00944_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[154]$_DFFE_PN0P_  (.D(_01340_),
    .RN(net256),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .QN(_00975_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[155]$_DFFE_PN0P_  (.D(_01341_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .QN(_01006_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[156]$_DFFE_PN0P_  (.D(_01342_),
    .RN(net258),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .QN(_01037_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[157]$_DFFE_PN0P_  (.D(_01343_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .QN(_01068_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[158]$_DFFE_PN0P_  (.D(_01344_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .QN(_01099_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[159]$_DFFE_PN0P_  (.D(_01345_),
    .RN(net262),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .QN(_01130_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[15]$_DFFE_PN0P_  (.D(_01346_),
    .RN(net261),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .QN(_14043_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[160]$_DFFE_PN0P_  (.D(_01347_),
    .RN(net267),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .QN(_00190_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[161]$_DFFE_PN0P_  (.D(_01348_),
    .RN(net266),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .QN(_00145_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[162]$_DFFE_PN0P_  (.D(_01349_),
    .RN(net267),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .QN(_00252_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[163]$_DFFE_PN0P_  (.D(_01350_),
    .RN(net267),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .QN(_00283_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[164]$_DFFE_PN0P_  (.D(_01351_),
    .RN(net267),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .QN(_00313_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[165]$_DFFE_PN0P_  (.D(_01352_),
    .RN(net267),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .QN(_00343_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[166]$_DFFE_PN0P_  (.D(_01353_),
    .RN(net258),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .QN(_00373_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[167]$_DFFE_PN0P_  (.D(_01354_),
    .RN(net268),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .QN(_00403_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[168]$_DFFE_PN0P_  (.D(_01355_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .QN(_00433_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[169]$_DFFE_PN0P_  (.D(_01356_),
    .RN(net267),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .QN(_00463_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[16]$_DFFE_PN0P_  (.D(_01357_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .QN(_14042_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[170]$_DFFE_PN0P_  (.D(_01358_),
    .RN(net262),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .QN(_00493_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[171]$_DFFE_PN0P_  (.D(_01359_),
    .RN(net255),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .QN(_00523_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[172]$_DFFE_PN0P_  (.D(_01360_),
    .RN(net261),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .QN(_00222_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[173]$_DFFE_PN0P_  (.D(_01361_),
    .RN(net255),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .QN(_00573_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[174]$_DFFE_PN0P_  (.D(_01362_),
    .RN(net255),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .QN(_00604_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[175]$_DFFE_PN0P_  (.D(_01363_),
    .RN(net255),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .QN(_00635_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[176]$_DFFE_PN0P_  (.D(_01364_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .QN(_00666_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[177]$_DFFE_PN0P_  (.D(_01365_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .QN(_00697_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[178]$_DFFE_PN0P_  (.D(_01366_),
    .RN(net255),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .QN(_00728_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[179]$_DFFE_PN0P_  (.D(_01367_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .QN(_00759_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[17]$_DFFE_PN0P_  (.D(_01368_),
    .RN(net257),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .QN(_14041_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[180]$_DFFE_PN0P_  (.D(_01369_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .QN(_00790_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[181]$_DFFE_PN0P_  (.D(_01370_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .QN(_00821_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[182]$_DFFE_PN0P_  (.D(_01371_),
    .RN(net260),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .QN(_00852_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[183]$_DFFE_PN0P_  (.D(_01372_),
    .RN(net261),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .QN(_00883_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[184]$_DFFE_PN0P_  (.D(_01373_),
    .RN(net258),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .QN(_00914_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[185]$_DFFE_PN0P_  (.D(_01374_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .QN(_00945_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[186]$_DFFE_PN0P_  (.D(_01375_),
    .RN(net257),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .QN(_00976_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[187]$_DFFE_PN0P_  (.D(_01376_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .QN(_01007_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[188]$_DFFE_PN0P_  (.D(_01377_),
    .RN(net258),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .QN(_01038_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[189]$_DFFE_PN0P_  (.D(_01378_),
    .RN(net262),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .QN(_01069_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[18]$_DFFE_PN0P_  (.D(_01379_),
    .RN(net261),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .QN(_14040_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[190]$_DFFE_PN0P_  (.D(_01380_),
    .RN(net258),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .QN(_01100_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[191]$_DFFE_PN0P_  (.D(_01381_),
    .RN(net262),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .QN(_01131_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[192]$_DFFE_PN0P_  (.D(_01382_),
    .RN(net267),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .QN(_00191_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[193]$_DFFE_PN0P_  (.D(_01383_),
    .RN(net266),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .QN(_00146_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[194]$_DFFE_PN0P_  (.D(_01384_),
    .RN(net267),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .QN(_00253_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[195]$_DFFE_PN0P_  (.D(_01385_),
    .RN(net267),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .QN(_00284_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[196]$_DFFE_PN0P_  (.D(_01386_),
    .RN(net264),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .QN(_00314_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[197]$_DFFE_PN0P_  (.D(_01387_),
    .RN(net264),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .QN(_00344_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[198]$_DFFE_PN0P_  (.D(_01388_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .QN(_00374_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[199]$_DFFE_PN0P_  (.D(_01389_),
    .RN(net262),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .QN(_00404_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[19]$_DFFE_PN0P_  (.D(_01390_),
    .RN(net261),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .QN(_14039_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[1]$_DFFE_PN0P_  (.D(_01391_),
    .RN(net266),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .QN(_14038_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[200]$_DFFE_PN0P_  (.D(_01392_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .QN(_00434_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[201]$_DFFE_PN0P_  (.D(_01393_),
    .RN(net268),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .QN(_00464_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[202]$_DFFE_PN0P_  (.D(_01394_),
    .RN(net262),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .QN(_00494_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[203]$_DFFE_PN0P_  (.D(_01395_),
    .RN(net255),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .QN(_00524_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[204]$_DFFE_PN0P_  (.D(_01396_),
    .RN(net261),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .QN(_00223_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[205]$_DFFE_PN0P_  (.D(_01397_),
    .RN(net255),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .QN(_00574_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[206]$_DFFE_PN0P_  (.D(_01398_),
    .RN(net255),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .QN(_00605_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[207]$_DFFE_PN0P_  (.D(_01399_),
    .RN(net255),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .QN(_00636_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[208]$_DFFE_PN0P_  (.D(_01400_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .QN(_00667_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[209]$_DFFE_PN0P_  (.D(_01401_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .QN(_00698_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[20]$_DFFE_PN0P_  (.D(_01402_),
    .RN(net259),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .QN(_14037_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[210]$_DFFE_PN0P_  (.D(_01403_),
    .RN(net255),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .QN(_00729_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[211]$_DFFE_PN0P_  (.D(_01404_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .QN(_00760_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[212]$_DFFE_PN0P_  (.D(_01405_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .QN(_00791_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[213]$_DFFE_PN0P_  (.D(_01406_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .QN(_00822_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[214]$_DFFE_PN0P_  (.D(_01407_),
    .RN(net260),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .QN(_00853_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[215]$_DFFE_PN0P_  (.D(_01408_),
    .RN(net259),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .QN(_00884_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[216]$_DFFE_PN0P_  (.D(_01409_),
    .RN(net258),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .QN(_00915_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[217]$_DFFE_PN0P_  (.D(_01410_),
    .RN(net260),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .QN(_00946_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[218]$_DFFE_PN0P_  (.D(_01411_),
    .RN(net256),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .QN(_00977_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[219]$_DFFE_PN0P_  (.D(_01412_),
    .RN(net260),
    .CK(clknet_leaf_55_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .QN(_01008_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[21]$_DFFE_PN0P_  (.D(_01413_),
    .RN(net257),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .QN(_14036_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[220]$_DFFE_PN0P_  (.D(_01414_),
    .RN(net258),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .QN(_01039_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[221]$_DFFE_PN0P_  (.D(_01415_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .QN(_01070_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[222]$_DFFE_PN0P_  (.D(_01416_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .QN(_01101_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[223]$_DFFE_PN0P_  (.D(_01417_),
    .RN(net266),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .QN(_01132_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[224]$_DFFE_PN0P_  (.D(_01418_),
    .RN(net267),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .QN(_00192_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[225]$_DFFE_PN0P_  (.D(_01419_),
    .RN(net266),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .QN(_00147_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[226]$_DFFE_PN0P_  (.D(_01420_),
    .RN(net264),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .QN(_00254_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[227]$_DFFE_PN0P_  (.D(_01421_),
    .RN(net267),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .QN(_00285_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[228]$_DFFE_PN0P_  (.D(_01422_),
    .RN(net264),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .QN(_00315_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[229]$_DFFE_PN0P_  (.D(_01423_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .QN(_00345_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[22]$_DFFE_PN0P_  (.D(_01424_),
    .RN(net259),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .QN(_14035_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[230]$_DFFE_PN0P_  (.D(_01425_),
    .RN(net257),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .QN(_00375_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[231]$_DFFE_PN0P_  (.D(_01426_),
    .RN(net262),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .QN(_00405_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[232]$_DFFE_PN0P_  (.D(_01427_),
    .RN(net263),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .QN(_00435_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[233]$_DFFE_PN0P_  (.D(_01428_),
    .RN(net263),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .QN(_00465_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[234]$_DFFE_PN0P_  (.D(_01429_),
    .RN(net262),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .QN(_00495_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[235]$_DFFE_PN0P_  (.D(_01430_),
    .RN(net263),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .QN(_00525_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[236]$_DFFE_PN0P_  (.D(_01431_),
    .RN(net260),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .QN(_00224_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[237]$_DFFE_PN0P_  (.D(_01432_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .QN(_00575_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[238]$_DFFE_PN0P_  (.D(_01433_),
    .RN(net263),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .QN(_00606_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[239]$_DFFE_PN0P_  (.D(_01434_),
    .RN(net261),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .QN(_00637_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[23]$_DFFE_PN0P_  (.D(_01435_),
    .RN(net259),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .QN(_14034_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[240]$_DFFE_PN0P_  (.D(_01436_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .QN(_00668_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[241]$_DFFE_PN0P_  (.D(_01437_),
    .RN(net259),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .QN(_00699_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[242]$_DFFE_PN0P_  (.D(_01438_),
    .RN(net263),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .QN(_00730_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[243]$_DFFE_PN0P_  (.D(_01439_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .QN(_00761_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[244]$_DFFE_PN0P_  (.D(_01440_),
    .RN(net259),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .QN(_00792_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[245]$_DFFE_PN0P_  (.D(_01441_),
    .RN(net259),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .QN(_00823_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[246]$_DFFE_PN0P_  (.D(_01442_),
    .RN(net260),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .QN(_00854_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[247]$_DFFE_PN0P_  (.D(_01443_),
    .RN(net259),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .QN(_00885_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[248]$_DFFE_PN0P_  (.D(_01444_),
    .RN(net258),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .QN(_00916_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[249]$_DFFE_PN0P_  (.D(_01445_),
    .RN(net259),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .QN(_00947_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[24]$_DFFE_PN0P_  (.D(_01446_),
    .RN(net257),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .QN(_14033_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[250]$_DFFE_PN0P_  (.D(_01447_),
    .RN(net257),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .QN(_00978_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[251]$_DFFE_PN0P_  (.D(_01448_),
    .RN(net259),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .QN(_01009_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[252]$_DFFE_PN0P_  (.D(_01449_),
    .RN(net258),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .QN(_01040_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[253]$_DFFE_PN0P_  (.D(_01450_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .QN(_01071_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[254]$_DFFE_PN0P_  (.D(_01451_),
    .RN(net257),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .QN(_01102_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[255]$_DFFE_PN0P_  (.D(_01452_),
    .RN(net266),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .QN(_01133_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[256]$_DFFE_PN0P_  (.D(_01453_),
    .RN(net267),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .QN(_00193_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[257]$_DFFE_PN0P_  (.D(_01454_),
    .RN(net266),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .QN(_00148_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[258]$_DFFE_PN0P_  (.D(_01455_),
    .RN(net264),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .QN(_00255_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[259]$_DFFE_PN0P_  (.D(_01456_),
    .RN(net267),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .QN(_00286_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[25]$_DFFE_PN0P_  (.D(_01457_),
    .RN(net257),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .QN(_14032_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[260]$_DFFE_PN0P_  (.D(_01458_),
    .RN(net267),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .QN(_00316_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[261]$_DFFE_PN0P_  (.D(_01459_),
    .RN(net264),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .QN(_00346_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[262]$_DFFE_PN0P_  (.D(_01460_),
    .RN(net257),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .QN(_00376_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[263]$_DFFE_PN0P_  (.D(_01461_),
    .RN(net268),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .QN(_00406_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[264]$_DFFE_PN0P_  (.D(_01462_),
    .RN(net263),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .QN(_00436_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[265]$_DFFE_PN0P_  (.D(_01463_),
    .RN(net268),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .QN(_00466_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[266]$_DFFE_PN0P_  (.D(_01464_),
    .RN(net262),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .QN(_00496_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[267]$_DFFE_PN0P_  (.D(_01465_),
    .RN(net263),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .QN(_00526_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[268]$_DFFE_PN0P_  (.D(_01466_),
    .RN(net260),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .QN(_00225_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[269]$_DFFE_PN0P_  (.D(_01467_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .QN(_00576_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[26]$_DFFE_PN0P_  (.D(_01468_),
    .RN(net257),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .QN(_14031_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[270]$_DFFE_PN0P_  (.D(_01469_),
    .RN(net263),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .QN(_00607_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[271]$_DFFE_PN0P_  (.D(_01470_),
    .RN(net261),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .QN(_00638_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[272]$_DFFE_PN0P_  (.D(_01471_),
    .RN(net263),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .QN(_00669_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[273]$_DFFE_PN0P_  (.D(_01472_),
    .RN(net259),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .QN(_00700_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[274]$_DFFE_PN0P_  (.D(_01473_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .QN(_00731_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[275]$_DFFE_PN0P_  (.D(_01474_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .QN(_00762_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[276]$_DFFE_PN0P_  (.D(_01475_),
    .RN(net259),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .QN(_00793_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[277]$_DFFE_PN0P_  (.D(_01476_),
    .RN(net259),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .QN(_00824_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[278]$_DFFE_PN0P_  (.D(_01477_),
    .RN(net259),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .QN(_00855_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[279]$_DFFE_PN0P_  (.D(_01478_),
    .RN(net259),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .QN(_00886_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[27]$_DFFE_PN0P_  (.D(_01479_),
    .RN(net259),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .QN(_14030_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[280]$_DFFE_PN0P_  (.D(_01480_),
    .RN(net259),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .QN(_00917_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[281]$_DFFE_PN0P_  (.D(_01481_),
    .RN(net259),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .QN(_00948_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[282]$_DFFE_PN0P_  (.D(_01482_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .QN(_00979_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[283]$_DFFE_PN0P_  (.D(_01483_),
    .RN(net259),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .QN(_01010_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[284]$_DFFE_PN0P_  (.D(_01484_),
    .RN(net259),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .QN(_01041_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[285]$_DFFE_PN0P_  (.D(_01485_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .QN(_01072_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[286]$_DFFE_PN0P_  (.D(_01486_),
    .RN(net257),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .QN(_01103_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[287]$_DFFE_PN0P_  (.D(_01487_),
    .RN(net262),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .QN(_01134_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[288]$_DFFE_PN0P_  (.D(_01488_),
    .RN(net267),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .QN(_00194_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[289]$_DFFE_PN0P_  (.D(_01489_),
    .RN(net266),
    .CK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .QN(_00149_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[28]$_DFFE_PN0P_  (.D(_01490_),
    .RN(net257),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .QN(_14029_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[290]$_DFFE_PN0P_  (.D(_01491_),
    .RN(net264),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .QN(_00256_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[291]$_DFFE_PN0P_  (.D(_01492_),
    .RN(net266),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .QN(_00287_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[292]$_DFFE_PN0P_  (.D(_01493_),
    .RN(net266),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .QN(_00317_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[293]$_DFFE_PN0P_  (.D(_01494_),
    .RN(net264),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .QN(_00347_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[294]$_DFFE_PN0P_  (.D(_01495_),
    .RN(net257),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .QN(_00377_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[295]$_DFFE_PN0P_  (.D(_01496_),
    .RN(net262),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .QN(_00407_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[296]$_DFFE_PN0P_  (.D(_01497_),
    .RN(net255),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .QN(_00437_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[297]$_DFFE_PN0P_  (.D(_01498_),
    .RN(net268),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .QN(_00467_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[298]$_DFFE_PN0P_  (.D(_01499_),
    .RN(net262),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .QN(_00497_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[299]$_DFFE_PN0P_  (.D(_01500_),
    .RN(net263),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .QN(_00527_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[29]$_DFFE_PN0P_  (.D(_01501_),
    .RN(net256),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .QN(_14028_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[2]$_DFFE_PN0P_  (.D(_01502_),
    .RN(net266),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .QN(_14027_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[300]$_DFFE_PN0P_  (.D(_01503_),
    .RN(net260),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .QN(_00226_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[301]$_DFFE_PN0P_  (.D(_01504_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .QN(_00577_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[302]$_DFFE_PN0P_  (.D(_01505_),
    .RN(net263),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .QN(_00608_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[303]$_DFFE_PN0P_  (.D(_01506_),
    .RN(net261),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .QN(_00639_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[304]$_DFFE_PN0P_  (.D(_01507_),
    .RN(net263),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .QN(_00670_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[305]$_DFFE_PN0P_  (.D(_01508_),
    .RN(net259),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .QN(_00701_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[306]$_DFFE_PN0P_  (.D(_01509_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .QN(_00732_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[307]$_DFFE_PN0P_  (.D(_01510_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .QN(_00763_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[308]$_DFFE_PN0P_  (.D(_01511_),
    .RN(net259),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .QN(_00794_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[309]$_DFFE_PN0P_  (.D(_01512_),
    .RN(net260),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .QN(_00825_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[30]$_DFFE_PN0P_  (.D(_01513_),
    .RN(net257),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .QN(_14026_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[310]$_DFFE_PN0P_  (.D(_01514_),
    .RN(net260),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .QN(_00856_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[311]$_DFFE_PN0P_  (.D(_01515_),
    .RN(net259),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .QN(_00887_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[312]$_DFFE_PN0P_  (.D(_01516_),
    .RN(net258),
    .CK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .QN(_00918_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[313]$_DFFE_PN0P_  (.D(_01517_),
    .RN(net259),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .QN(_00949_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[314]$_DFFE_PN0P_  (.D(_01518_),
    .RN(net257),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .QN(_00980_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[315]$_DFFE_PN0P_  (.D(_01519_),
    .RN(net260),
    .CK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .QN(_01011_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[316]$_DFFE_PN0P_  (.D(_01520_),
    .RN(net258),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .QN(_01042_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[317]$_DFFE_PN0P_  (.D(_01521_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .QN(_01073_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[318]$_DFFE_PN0P_  (.D(_01522_),
    .RN(net257),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .QN(_01104_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[319]$_DFFE_PN0P_  (.D(_01523_),
    .RN(net262),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .QN(_01135_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[31]$_DFFE_PN0P_  (.D(_01524_),
    .RN(net266),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .QN(_14025_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[320]$_DFFE_PN0P_  (.D(_01525_),
    .RN(net264),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .QN(_00195_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[321]$_DFFE_PN0P_  (.D(_01526_),
    .RN(net266),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .QN(_00150_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[322]$_DFFE_PN0P_  (.D(_01527_),
    .RN(net264),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .QN(_00257_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[323]$_DFFE_PN0P_  (.D(_01528_),
    .RN(net267),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .QN(_00288_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[324]$_DFFE_PN0P_  (.D(_01529_),
    .RN(net267),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .QN(_00318_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[325]$_DFFE_PN0P_  (.D(_01530_),
    .RN(net264),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .QN(_00348_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[326]$_DFFE_PN0P_  (.D(_01531_),
    .RN(net257),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .QN(_00378_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[327]$_DFFE_PN0P_  (.D(_01532_),
    .RN(net262),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .QN(_00408_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[328]$_DFFE_PN0P_  (.D(_01533_),
    .RN(net263),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .QN(_00438_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[329]$_DFFE_PN0P_  (.D(_01534_),
    .RN(net268),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .QN(_00468_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[32]$_DFFE_PN0P_  (.D(_01535_),
    .RN(net267),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .QN(_00186_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[330]$_DFFE_PN0P_  (.D(_01536_),
    .RN(net262),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .QN(_00498_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[331]$_DFFE_PN0P_  (.D(_01537_),
    .RN(net263),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .QN(_00528_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[332]$_DFFE_PN0P_  (.D(_01538_),
    .RN(net260),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .QN(_00227_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[333]$_DFFE_PN0P_  (.D(_01539_),
    .RN(net262),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .QN(_00578_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[334]$_DFFE_PN0P_  (.D(_01540_),
    .RN(net261),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .QN(_00609_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[335]$_DFFE_PN0P_  (.D(_01541_),
    .RN(net261),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .QN(_00640_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[336]$_DFFE_PN0P_  (.D(_01542_),
    .RN(net263),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .QN(_00671_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[337]$_DFFE_PN0P_  (.D(_01543_),
    .RN(net259),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .QN(_00702_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[338]$_DFFE_PN0P_  (.D(_01544_),
    .RN(net263),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .QN(_00733_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[339]$_DFFE_PN0P_  (.D(_01545_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .QN(_00764_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[33]$_DFFE_PN0P_  (.D(_01546_),
    .RN(net266),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .QN(_00141_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[340]$_DFFE_PN0P_  (.D(_01547_),
    .RN(net259),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .QN(_00795_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[341]$_DFFE_PN0P_  (.D(_01548_),
    .RN(net258),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .QN(_00826_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[342]$_DFFE_PN0P_  (.D(_01549_),
    .RN(net259),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .QN(_00857_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[343]$_DFFE_PN0P_  (.D(_01550_),
    .RN(net261),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .QN(_00888_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[344]$_DFFE_PN0P_  (.D(_01551_),
    .RN(net258),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .QN(_00919_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[345]$_DFFE_PN0P_  (.D(_01552_),
    .RN(net259),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .QN(_00950_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[346]$_DFFE_PN0P_  (.D(_01553_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .QN(_00981_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[347]$_DFFE_PN0P_  (.D(_01554_),
    .RN(net259),
    .CK(clknet_leaf_59_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .QN(_01012_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[348]$_DFFE_PN0P_  (.D(_01555_),
    .RN(net259),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .QN(_01043_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[349]$_DFFE_PN0P_  (.D(_01556_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .QN(_01074_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[34]$_DFFE_PN0P_  (.D(_01557_),
    .RN(net266),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .QN(_00248_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[350]$_DFFE_PN0P_  (.D(_01558_),
    .RN(net257),
    .CK(clknet_leaf_72_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .QN(_01105_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[351]$_DFFE_PN0P_  (.D(_01559_),
    .RN(net266),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .QN(_01136_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[352]$_DFFE_PN0P_  (.D(_01560_),
    .RN(net264),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .QN(_00196_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[353]$_DFFE_PN0P_  (.D(_01561_),
    .RN(net266),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .QN(_00151_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[354]$_DFFE_PN0P_  (.D(_01562_),
    .RN(net264),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .QN(_00258_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[355]$_DFFE_PN0P_  (.D(_01563_),
    .RN(net267),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .QN(_00289_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[356]$_DFFE_PN0P_  (.D(_01564_),
    .RN(net264),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .QN(_00319_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[357]$_DFFE_PN0P_  (.D(_01565_),
    .RN(net264),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .QN(_00349_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[358]$_DFFE_PN0P_  (.D(_01566_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .QN(_00379_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[359]$_DFFE_PN0P_  (.D(_01567_),
    .RN(net262),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .QN(_00409_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[35]$_DFFE_PN0P_  (.D(_01568_),
    .RN(net267),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .QN(_00279_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[360]$_DFFE_PN0P_  (.D(_01569_),
    .RN(net263),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .QN(_00439_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[361]$_DFFE_PN0P_  (.D(_01570_),
    .RN(net268),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .QN(_00469_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[362]$_DFFE_PN0P_  (.D(_01571_),
    .RN(net262),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .QN(_00499_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[363]$_DFFE_PN0P_  (.D(_01572_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .QN(_00529_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[364]$_DFFE_PN0P_  (.D(_01573_),
    .RN(net261),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .QN(_00228_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[365]$_DFFE_PN0P_  (.D(_01574_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .QN(_00579_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[366]$_DFFE_PN0P_  (.D(_01575_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .QN(_00610_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[367]$_DFFE_PN0P_  (.D(_01576_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .QN(_00641_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[368]$_DFFE_PN0P_  (.D(_01577_),
    .RN(net255),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .QN(_00672_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[369]$_DFFE_PN0P_  (.D(_01578_),
    .RN(net260),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .QN(_00703_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[36]$_DFFE_PN0P_  (.D(_01579_),
    .RN(net266),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .QN(_00309_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[370]$_DFFE_PN0P_  (.D(_01580_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .QN(_00734_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[371]$_DFFE_PN0P_  (.D(_01581_),
    .RN(net255),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .QN(_00765_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[372]$_DFFE_PN0P_  (.D(_01582_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .QN(_00796_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[373]$_DFFE_PN0P_  (.D(_01583_),
    .RN(net258),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .QN(_00827_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[374]$_DFFE_PN0P_  (.D(_01584_),
    .RN(net258),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .QN(_00858_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[375]$_DFFE_PN0P_  (.D(_01585_),
    .RN(net261),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .QN(_00889_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[376]$_DFFE_PN0P_  (.D(_01586_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .QN(_00920_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[377]$_DFFE_PN0P_  (.D(_01587_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .QN(_00951_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[378]$_DFFE_PN0P_  (.D(_01588_),
    .RN(net257),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .QN(_00982_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[379]$_DFFE_PN0P_  (.D(_01589_),
    .RN(net260),
    .CK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .QN(_01013_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[37]$_DFFE_PN0P_  (.D(_01590_),
    .RN(net267),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .QN(_00339_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[380]$_DFFE_PN0P_  (.D(_01591_),
    .RN(net258),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .QN(_01044_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[381]$_DFFE_PN0P_  (.D(_01592_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .QN(_01075_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[382]$_DFFE_PN0P_  (.D(_01593_),
    .RN(net258),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .QN(_01106_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[383]$_DFFE_PN0P_  (.D(_01594_),
    .RN(net266),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .QN(_01137_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[384]$_DFFE_PN0P_  (.D(_01595_),
    .RN(net264),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .QN(_00197_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[385]$_DFFE_PN0P_  (.D(_01596_),
    .RN(net266),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .QN(_00152_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[386]$_DFFE_PN0P_  (.D(_01597_),
    .RN(net264),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .QN(_00259_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[387]$_DFFE_PN0P_  (.D(_01598_),
    .RN(net267),
    .CK(clknet_leaf_130_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .QN(_00290_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[388]$_DFFE_PN0P_  (.D(_01599_),
    .RN(net264),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .QN(_00320_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[389]$_DFFE_PN0P_  (.D(_01600_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .QN(_00350_));
 DFFR_X2 \gen_regfile_ff.register_file_i.rf_reg_q[38]$_DFFE_PN0P_  (.D(_01601_),
    .RN(net257),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .QN(_00369_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[390]$_DFFE_PN0P_  (.D(_01602_),
    .RN(net258),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .QN(_00380_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[391]$_DFFE_PN0P_  (.D(_01603_),
    .RN(net268),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .QN(_00410_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[392]$_DFFE_PN0P_  (.D(_01604_),
    .RN(net268),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .QN(_00440_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[393]$_DFFE_PN0P_  (.D(_01605_),
    .RN(net268),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .QN(_00470_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[394]$_DFFE_PN0P_  (.D(_01606_),
    .RN(net262),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .QN(_00500_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[395]$_DFFE_PN0P_  (.D(_01607_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .QN(_00530_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[396]$_DFFE_PN0P_  (.D(_01608_),
    .RN(net261),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .QN(_00229_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[397]$_DFFE_PN0P_  (.D(_01609_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .QN(_00580_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[398]$_DFFE_PN0P_  (.D(_01610_),
    .RN(net255),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .QN(_00611_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[399]$_DFFE_PN0P_  (.D(_01611_),
    .RN(net255),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .QN(_00642_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[39]$_DFFE_PN0P_  (.D(_01612_),
    .RN(net268),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .QN(_00399_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[3]$_DFFE_PN0P_  (.D(_01613_),
    .RN(net268),
    .CK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .QN(_14024_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[400]$_DFFE_PN0P_  (.D(_01614_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .QN(_00673_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[401]$_DFFE_PN0P_  (.D(_01615_),
    .RN(net258),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .QN(_00704_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[402]$_DFFE_PN0P_  (.D(_01616_),
    .RN(net255),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .QN(_00735_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[403]$_DFFE_PN0P_  (.D(_01617_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .QN(_00766_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[404]$_DFFE_PN0P_  (.D(_01618_),
    .RN(net260),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .QN(_00797_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[405]$_DFFE_PN0P_  (.D(_01619_),
    .RN(net259),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .QN(_00828_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[406]$_DFFE_PN0P_  (.D(_01620_),
    .RN(net260),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .QN(_00859_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[407]$_DFFE_PN0P_  (.D(_01621_),
    .RN(net261),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .QN(_00890_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[408]$_DFFE_PN0P_  (.D(_01622_),
    .RN(net258),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .QN(_00921_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[409]$_DFFE_PN0P_  (.D(_01623_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .QN(_00952_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[40]$_DFFE_PN0P_  (.D(_01624_),
    .RN(net268),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .QN(_00429_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[410]$_DFFE_PN0P_  (.D(_01625_),
    .RN(net257),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .QN(_00983_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[411]$_DFFE_PN0P_  (.D(_01626_),
    .RN(net260),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .QN(_01014_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[412]$_DFFE_PN0P_  (.D(_01627_),
    .RN(net259),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .QN(_01045_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[413]$_DFFE_PN0P_  (.D(_01628_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .QN(_01076_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[414]$_DFFE_PN0P_  (.D(_01629_),
    .RN(net259),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .QN(_01107_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[415]$_DFFE_PN0P_  (.D(_01630_),
    .RN(net262),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .QN(_01138_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[416]$_DFFE_PN0P_  (.D(_01631_),
    .RN(net264),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .QN(_00198_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[417]$_DFFE_PN0P_  (.D(_01632_),
    .RN(net266),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .QN(_00153_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[418]$_DFFE_PN0P_  (.D(_01633_),
    .RN(net264),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .QN(_00260_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[419]$_DFFE_PN0P_  (.D(_01634_),
    .RN(net266),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .QN(_00291_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[41]$_DFFE_PN0P_  (.D(_01635_),
    .RN(net268),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .QN(_00459_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[420]$_DFFE_PN0P_  (.D(_01636_),
    .RN(net264),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .QN(_00321_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[421]$_DFFE_PN0P_  (.D(_01637_),
    .RN(net264),
    .CK(clknet_leaf_131_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .QN(_00351_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[422]$_DFFE_PN0P_  (.D(_01638_),
    .RN(net258),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .QN(_00381_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[423]$_DFFE_PN0P_  (.D(_01639_),
    .RN(net262),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .QN(_00411_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[424]$_DFFE_PN0P_  (.D(_01640_),
    .RN(net268),
    .CK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .QN(_00441_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[425]$_DFFE_PN0P_  (.D(_01641_),
    .RN(net268),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .QN(_00471_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[426]$_DFFE_PN0P_  (.D(_01642_),
    .RN(net262),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .QN(_00501_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[427]$_DFFE_PN0P_  (.D(_01643_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .QN(_00531_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[428]$_DFFE_PN0P_  (.D(_01644_),
    .RN(net261),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .QN(_00230_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[429]$_DFFE_PN0P_  (.D(_01645_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .QN(_00581_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[42]$_DFFE_PN0P_  (.D(_01646_),
    .RN(net262),
    .CK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .QN(_00489_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[430]$_DFFE_PN0P_  (.D(_01647_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .QN(_00612_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[431]$_DFFE_PN0P_  (.D(_01648_),
    .RN(net255),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .QN(_00643_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[432]$_DFFE_PN0P_  (.D(_01649_),
    .RN(net255),
    .CK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .QN(_00674_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[433]$_DFFE_PN0P_  (.D(_01650_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .QN(_00705_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[434]$_DFFE_PN0P_  (.D(_01651_),
    .RN(net255),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .QN(_00736_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[435]$_DFFE_PN0P_  (.D(_01652_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .QN(_00767_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[436]$_DFFE_PN0P_  (.D(_01653_),
    .RN(net260),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .QN(_00798_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[437]$_DFFE_PN0P_  (.D(_01654_),
    .RN(net258),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .QN(_00829_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[438]$_DFFE_PN0P_  (.D(_01655_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .QN(_00860_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[439]$_DFFE_PN0P_  (.D(_01656_),
    .RN(net261),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .QN(_00891_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[43]$_DFFE_PN0P_  (.D(_01657_),
    .RN(net268),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .QN(_00519_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[440]$_DFFE_PN0P_  (.D(_01658_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .QN(_00922_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[441]$_DFFE_PN0P_  (.D(_01659_),
    .RN(net258),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .QN(_00953_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[442]$_DFFE_PN0P_  (.D(_01660_),
    .RN(net257),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .QN(_00984_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[443]$_DFFE_PN0P_  (.D(_01661_),
    .RN(net258),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .QN(_01015_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[444]$_DFFE_PN0P_  (.D(_01662_),
    .RN(net259),
    .CK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .QN(_01046_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[445]$_DFFE_PN0P_  (.D(_01663_),
    .RN(net256),
    .CK(clknet_leaf_70_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .QN(_01077_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[446]$_DFFE_PN0P_  (.D(_01664_),
    .RN(net259),
    .CK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .QN(_01108_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[447]$_DFFE_PN0P_  (.D(_01665_),
    .RN(net266),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .QN(_01139_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[448]$_DFFE_PN0P_  (.D(_01666_),
    .RN(net264),
    .CK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .QN(_00199_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[449]$_DFFE_PN0P_  (.D(_01667_),
    .RN(net267),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .QN(_00154_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[44]$_DFFE_PN0P_  (.D(_01668_),
    .RN(net260),
    .CK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .QN(_00218_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[450]$_DFFE_PN0P_  (.D(_01669_),
    .RN(net264),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .QN(_00261_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[451]$_DFFE_PN0P_  (.D(_01670_),
    .RN(net267),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .QN(_00292_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[452]$_DFFE_PN0P_  (.D(_01671_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .QN(_00322_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[453]$_DFFE_PN0P_  (.D(_01672_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .QN(_00352_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[454]$_DFFE_PN0P_  (.D(_01673_),
    .RN(net258),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .QN(_00382_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[455]$_DFFE_PN0P_  (.D(_01674_),
    .RN(net262),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .QN(_00412_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[456]$_DFFE_PN0P_  (.D(_01675_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .QN(_00442_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[457]$_DFFE_PN0P_  (.D(_01676_),
    .RN(net268),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .QN(_00472_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[458]$_DFFE_PN0P_  (.D(_01677_),
    .RN(net262),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .QN(_00502_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[459]$_DFFE_PN0P_  (.D(_01678_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .QN(_00532_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[45]$_DFFE_PN0P_  (.D(_01679_),
    .RN(net261),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .QN(_00569_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[460]$_DFFE_PN0P_  (.D(_01680_),
    .RN(net261),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .QN(_00231_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[461]$_DFFE_PN0P_  (.D(_01681_),
    .RN(net255),
    .CK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .QN(_00582_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[462]$_DFFE_PN0P_  (.D(_01682_),
    .RN(net255),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .QN(_00613_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[463]$_DFFE_PN0P_  (.D(_01683_),
    .RN(net255),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .QN(_00644_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[464]$_DFFE_PN0P_  (.D(_01684_),
    .RN(net255),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .QN(_00675_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[465]$_DFFE_PN0P_  (.D(_01685_),
    .RN(net258),
    .CK(clknet_leaf_81_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .QN(_00706_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[466]$_DFFE_PN0P_  (.D(_01686_),
    .RN(net255),
    .CK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .QN(_00737_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[467]$_DFFE_PN0P_  (.D(_01687_),
    .RN(net255),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .QN(_00768_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[468]$_DFFE_PN0P_  (.D(_01688_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .QN(_00799_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[469]$_DFFE_PN0P_  (.D(_01689_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .QN(_00830_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[46]$_DFFE_PN0P_  (.D(_01690_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .QN(_00600_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[470]$_DFFE_PN0P_  (.D(_01691_),
    .RN(net260),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .QN(_00861_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[471]$_DFFE_PN0P_  (.D(_01692_),
    .RN(net261),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .QN(_00892_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[472]$_DFFE_PN0P_  (.D(_01693_),
    .RN(net258),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .QN(_00923_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[473]$_DFFE_PN0P_  (.D(_01694_),
    .RN(net258),
    .CK(clknet_leaf_83_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .QN(_00954_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[474]$_DFFE_PN0P_  (.D(_01695_),
    .RN(net257),
    .CK(clknet_leaf_66_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .QN(_00985_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[475]$_DFFE_PN0P_  (.D(_01696_),
    .RN(net260),
    .CK(clknet_leaf_82_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .QN(_01016_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[476]$_DFFE_PN0P_  (.D(_01697_),
    .RN(net259),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .QN(_01047_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[477]$_DFFE_PN0P_  (.D(_01698_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .QN(_01078_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[478]$_DFFE_PN0P_  (.D(_01699_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .QN(_01109_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[479]$_DFFE_PN0P_  (.D(_01700_),
    .RN(net266),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .QN(_01140_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[47]$_DFFE_PN0P_  (.D(_01701_),
    .RN(net261),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .QN(_00631_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[480]$_DFFE_PN0P_  (.D(_01702_),
    .RN(net267),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .QN(_00200_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[481]$_DFFE_PN0P_  (.D(_01703_),
    .RN(net266),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .QN(_00155_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[482]$_DFFE_PN0P_  (.D(_01704_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .QN(_00262_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[483]$_DFFE_PN0P_  (.D(_01705_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .QN(_00293_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[484]$_DFFE_PN0P_  (.D(_01706_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .QN(_00323_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[485]$_DFFE_PN0P_  (.D(_01707_),
    .RN(net264),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .QN(_00353_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[486]$_DFFE_PN0P_  (.D(_01708_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .QN(_00383_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[487]$_DFFE_PN0P_  (.D(_01709_),
    .RN(net261),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .QN(_00413_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[488]$_DFFE_PN0P_  (.D(_01710_),
    .RN(net267),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .QN(_00443_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[489]$_DFFE_PN0P_  (.D(_01711_),
    .RN(net267),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .QN(_00473_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[48]$_DFFE_PN0P_  (.D(_01712_),
    .RN(net261),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .QN(_00662_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[490]$_DFFE_PN0P_  (.D(_01713_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .QN(_00503_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[491]$_DFFE_PN0P_  (.D(_01714_),
    .RN(net263),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .QN(_00533_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[492]$_DFFE_PN0P_  (.D(_01715_),
    .RN(net261),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .QN(_00232_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[493]$_DFFE_PN0P_  (.D(_01716_),
    .RN(net262),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .QN(_00583_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[494]$_DFFE_PN0P_  (.D(_01717_),
    .RN(net261),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .QN(_00614_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[495]$_DFFE_PN0P_  (.D(_01718_),
    .RN(net261),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .QN(_00645_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[496]$_DFFE_PN0P_  (.D(_01719_),
    .RN(net261),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .QN(_00676_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[497]$_DFFE_PN0P_  (.D(_01720_),
    .RN(net257),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .QN(_00707_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[498]$_DFFE_PN0P_  (.D(_01721_),
    .RN(net261),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .QN(_00738_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[499]$_DFFE_PN0P_  (.D(_01722_),
    .RN(net261),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .QN(_00769_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[49]$_DFFE_PN0P_  (.D(_01723_),
    .RN(net257),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .QN(_00693_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[4]$_DFFE_PN0P_  (.D(_01724_),
    .RN(net266),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .QN(_14023_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[500]$_DFFE_PN0P_  (.D(_01725_),
    .RN(net260),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .QN(_00800_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[501]$_DFFE_PN0P_  (.D(_01726_),
    .RN(net257),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .QN(_00831_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[502]$_DFFE_PN0P_  (.D(_01727_),
    .RN(net258),
    .CK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .QN(_00862_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[503]$_DFFE_PN0P_  (.D(_01728_),
    .RN(net261),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .QN(_00893_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[504]$_DFFE_PN0P_  (.D(_01729_),
    .RN(net257),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .QN(_00924_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[505]$_DFFE_PN0P_  (.D(_01730_),
    .RN(net258),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .QN(_00955_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[506]$_DFFE_PN0P_  (.D(_01731_),
    .RN(net256),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .QN(_00986_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[507]$_DFFE_PN0P_  (.D(_01732_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .QN(_01017_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[508]$_DFFE_PN0P_  (.D(_01733_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .QN(_01048_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[509]$_DFFE_PN0P_  (.D(_01734_),
    .RN(net262),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .QN(_01079_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[50]$_DFFE_PN0P_  (.D(_01735_),
    .RN(net261),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .QN(_00724_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[510]$_DFFE_PN0P_  (.D(_01736_),
    .RN(net256),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .QN(_01110_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[511]$_DFFE_PN0P_  (.D(_01737_),
    .RN(net266),
    .CK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .QN(_01141_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[512]$_DFFE_PN0P_  (.D(_01738_),
    .RN(net267),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .QN(_00201_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[513]$_DFFE_PN0P_  (.D(_01739_),
    .RN(net266),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .QN(_00156_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[514]$_DFFE_PN0P_  (.D(_01740_),
    .RN(net264),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .QN(_00263_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[515]$_DFFE_PN0P_  (.D(_01741_),
    .RN(net267),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .QN(_00294_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[516]$_DFFE_PN0P_  (.D(_01742_),
    .RN(net264),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .QN(_00324_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[517]$_DFFE_PN0P_  (.D(_01743_),
    .RN(net264),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .QN(_00354_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[518]$_DFFE_PN0P_  (.D(_01744_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .QN(_00384_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[519]$_DFFE_PN0P_  (.D(_01745_),
    .RN(net262),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .QN(_00414_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[51]$_DFFE_PN0P_  (.D(_01746_),
    .RN(net261),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .QN(_00755_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[520]$_DFFE_PN0P_  (.D(_01747_),
    .RN(net267),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .QN(_00444_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[521]$_DFFE_PN0P_  (.D(_01748_),
    .RN(net267),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .QN(_00474_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[522]$_DFFE_PN0P_  (.D(_01749_),
    .RN(net262),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .QN(_00504_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[523]$_DFFE_PN0P_  (.D(_01750_),
    .RN(net262),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .QN(_00534_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[524]$_DFFE_PN0P_  (.D(_01751_),
    .RN(net261),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .QN(_00233_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[525]$_DFFE_PN0P_  (.D(_01752_),
    .RN(net262),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .QN(_00584_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[526]$_DFFE_PN0P_  (.D(_01753_),
    .RN(net260),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .QN(_00615_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[527]$_DFFE_PN0P_  (.D(_01754_),
    .RN(net261),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .QN(_00646_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[528]$_DFFE_PN0P_  (.D(_01755_),
    .RN(net261),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .QN(_00677_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[529]$_DFFE_PN0P_  (.D(_01756_),
    .RN(net257),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .QN(_00708_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[52]$_DFFE_PN0P_  (.D(_01757_),
    .RN(net259),
    .CK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .QN(_00786_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[530]$_DFFE_PN0P_  (.D(_01758_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .QN(_00739_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[531]$_DFFE_PN0P_  (.D(_01759_),
    .RN(net261),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .QN(_00770_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[532]$_DFFE_PN0P_  (.D(_01760_),
    .RN(net260),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .QN(_00801_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[533]$_DFFE_PN0P_  (.D(_01761_),
    .RN(net257),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .QN(_00832_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[534]$_DFFE_PN0P_  (.D(_01762_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .QN(_00863_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[535]$_DFFE_PN0P_  (.D(_01763_),
    .RN(net261),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .QN(_00894_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[536]$_DFFE_PN0P_  (.D(_01764_),
    .RN(net257),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .QN(_00925_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[537]$_DFFE_PN0P_  (.D(_01765_),
    .RN(net258),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .QN(_00956_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[538]$_DFFE_PN0P_  (.D(_01766_),
    .RN(net262),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .QN(_00987_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[539]$_DFFE_PN0P_  (.D(_01767_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .QN(_01018_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[53]$_DFFE_PN0P_  (.D(_01768_),
    .RN(net259),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .QN(_00817_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[540]$_DFFE_PN0P_  (.D(_01769_),
    .RN(net256),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .QN(_01049_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[541]$_DFFE_PN0P_  (.D(_01770_),
    .RN(net262),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .QN(_01080_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[542]$_DFFE_PN0P_  (.D(_01771_),
    .RN(net262),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .QN(_01111_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[543]$_DFFE_PN0P_  (.D(_01772_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .QN(_01142_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[544]$_DFFE_PN0P_  (.D(_01773_),
    .RN(net267),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .QN(_00202_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[545]$_DFFE_PN0P_  (.D(_01774_),
    .RN(net266),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .QN(_00157_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[546]$_DFFE_PN0P_  (.D(_01775_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .QN(_00264_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[547]$_DFFE_PN0P_  (.D(_01776_),
    .RN(net267),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .QN(_00295_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[548]$_DFFE_PN0P_  (.D(_01777_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .QN(_00325_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[549]$_DFFE_PN0P_  (.D(_01778_),
    .RN(net267),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .QN(_00355_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[54]$_DFFE_PN0P_  (.D(_01779_),
    .RN(net259),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .QN(_00848_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[550]$_DFFE_PN0P_  (.D(_01780_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .QN(_00385_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[551]$_DFFE_PN0P_  (.D(_01781_),
    .RN(net268),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .QN(_00415_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[552]$_DFFE_PN0P_  (.D(_01782_),
    .RN(net267),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .QN(_00445_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[553]$_DFFE_PN0P_  (.D(_01783_),
    .RN(net267),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .QN(_00475_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[554]$_DFFE_PN0P_  (.D(_01784_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .QN(_00505_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[555]$_DFFE_PN0P_  (.D(_01785_),
    .RN(net263),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .QN(_00535_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[556]$_DFFE_PN0P_  (.D(_01786_),
    .RN(net260),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .QN(_00234_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[557]$_DFFE_PN0P_  (.D(_01787_),
    .RN(net262),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .QN(_00585_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[558]$_DFFE_PN0P_  (.D(_01788_),
    .RN(net261),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .QN(_00616_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[559]$_DFFE_PN0P_  (.D(_01789_),
    .RN(net261),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .QN(_00647_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[55]$_DFFE_PN0P_  (.D(_01790_),
    .RN(net259),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .QN(_00879_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[560]$_DFFE_PN0P_  (.D(_01791_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .QN(_00678_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[561]$_DFFE_PN0P_  (.D(_01792_),
    .RN(net257),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .QN(_00709_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[562]$_DFFE_PN0P_  (.D(_01793_),
    .RN(net261),
    .CK(clknet_leaf_41_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .QN(_00740_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[563]$_DFFE_PN0P_  (.D(_01794_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .QN(_00771_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[564]$_DFFE_PN0P_  (.D(_01795_),
    .RN(net260),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .QN(_00802_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[565]$_DFFE_PN0P_  (.D(_01796_),
    .RN(net257),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .QN(_00833_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[566]$_DFFE_PN0P_  (.D(_01797_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .QN(_00864_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[567]$_DFFE_PN0P_  (.D(_01798_),
    .RN(net261),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .QN(_00895_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[568]$_DFFE_PN0P_  (.D(_01799_),
    .RN(net257),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .QN(_00926_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[569]$_DFFE_PN0P_  (.D(_01800_),
    .RN(net258),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .QN(_00957_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[56]$_DFFE_PN0P_  (.D(_01801_),
    .RN(net259),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .QN(_00910_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[570]$_DFFE_PN0P_  (.D(_01802_),
    .RN(net256),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .QN(_00988_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[571]$_DFFE_PN0P_  (.D(_01803_),
    .RN(net258),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .QN(_01019_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[572]$_DFFE_PN0P_  (.D(_01804_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .QN(_01050_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[573]$_DFFE_PN0P_  (.D(_01805_),
    .RN(net266),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .QN(_01081_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[574]$_DFFE_PN0P_  (.D(_01806_),
    .RN(net256),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .QN(_01112_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[575]$_DFFE_PN0P_  (.D(_01807_),
    .RN(net266),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .QN(_01143_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[576]$_DFFE_PN0P_  (.D(_01808_),
    .RN(net267),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .QN(_00203_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[577]$_DFFE_PN0P_  (.D(_01809_),
    .RN(net266),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .QN(_00158_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[578]$_DFFE_PN0P_  (.D(_01810_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .QN(_00265_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[579]$_DFFE_PN0P_  (.D(_01811_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .QN(_00296_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[57]$_DFFE_PN0P_  (.D(_01812_),
    .RN(net259),
    .CK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .QN(_00941_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[580]$_DFFE_PN0P_  (.D(_01813_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .QN(_00326_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[581]$_DFFE_PN0P_  (.D(_01814_),
    .RN(net264),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .QN(_00356_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[582]$_DFFE_PN0P_  (.D(_01815_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .QN(_00386_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[583]$_DFFE_PN0P_  (.D(_01816_),
    .RN(net261),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .QN(_00416_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[584]$_DFFE_PN0P_  (.D(_01817_),
    .RN(net267),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .QN(_00446_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[585]$_DFFE_PN0P_  (.D(_01818_),
    .RN(net267),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .QN(_00476_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[586]$_DFFE_PN0P_  (.D(_01819_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .QN(_00506_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[587]$_DFFE_PN0P_  (.D(_01820_),
    .RN(net262),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .QN(_00536_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[588]$_DFFE_PN0P_  (.D(_01821_),
    .RN(net260),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .QN(_00235_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[589]$_DFFE_PN0P_  (.D(_01822_),
    .RN(net262),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .QN(_00586_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[58]$_DFFE_PN0P_  (.D(_01823_),
    .RN(net257),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .QN(_00972_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[590]$_DFFE_PN0P_  (.D(_01824_),
    .RN(net260),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .QN(_00617_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[591]$_DFFE_PN0P_  (.D(_01825_),
    .RN(net261),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .QN(_00648_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[592]$_DFFE_PN0P_  (.D(_01826_),
    .RN(net261),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .QN(_00679_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[593]$_DFFE_PN0P_  (.D(_01827_),
    .RN(net257),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .QN(_00710_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[594]$_DFFE_PN0P_  (.D(_01828_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .QN(_00741_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[595]$_DFFE_PN0P_  (.D(_01829_),
    .RN(net261),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .QN(_00772_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[596]$_DFFE_PN0P_  (.D(_01830_),
    .RN(net260),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .QN(_00803_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[597]$_DFFE_PN0P_  (.D(_01831_),
    .RN(net259),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .QN(_00834_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[598]$_DFFE_PN0P_  (.D(_01832_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .QN(_00865_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[599]$_DFFE_PN0P_  (.D(_01833_),
    .RN(net261),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .QN(_00896_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[59]$_DFFE_PN0P_  (.D(_01834_),
    .RN(net259),
    .CK(clknet_leaf_78_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .QN(_01003_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[5]$_DFFE_PN0P_  (.D(_01835_),
    .RN(net267),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .QN(_14022_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[600]$_DFFE_PN0P_  (.D(_01836_),
    .RN(net257),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .QN(_00927_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[601]$_DFFE_PN0P_  (.D(_01837_),
    .RN(net258),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .QN(_00958_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[602]$_DFFE_PN0P_  (.D(_01838_),
    .RN(net262),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .QN(_00989_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[603]$_DFFE_PN0P_  (.D(_01839_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .QN(_01020_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[604]$_DFFE_PN0P_  (.D(_01840_),
    .RN(net256),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .QN(_01051_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[605]$_DFFE_PN0P_  (.D(_01841_),
    .RN(net266),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .QN(_01082_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[606]$_DFFE_PN0P_  (.D(_01842_),
    .RN(net256),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .QN(_01113_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[607]$_DFFE_PN0P_  (.D(_01843_),
    .RN(net266),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .QN(_01144_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[608]$_DFFE_PN0P_  (.D(_01844_),
    .RN(net264),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .QN(_00204_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[609]$_DFFE_PN0P_  (.D(_01845_),
    .RN(net266),
    .CK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .QN(_00159_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[60]$_DFFE_PN0P_  (.D(_01846_),
    .RN(net257),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .QN(_01034_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[610]$_DFFE_PN0P_  (.D(_01847_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .QN(_00266_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[611]$_DFFE_PN0P_  (.D(_01848_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .QN(_00297_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[612]$_DFFE_PN0P_  (.D(_01849_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .QN(_00327_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[613]$_DFFE_PN0P_  (.D(_01850_),
    .RN(net264),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .QN(_00357_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[614]$_DFFE_PN0P_  (.D(_01851_),
    .RN(net258),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .QN(_00387_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[615]$_DFFE_PN0P_  (.D(_01852_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .QN(_00417_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[616]$_DFFE_PN0P_  (.D(_01853_),
    .RN(net267),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .QN(_00447_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[617]$_DFFE_PN0P_  (.D(_01854_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .QN(_00477_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[618]$_DFFE_PN0P_  (.D(_01855_),
    .RN(net262),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .QN(_00507_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[619]$_DFFE_PN0P_  (.D(_01856_),
    .RN(net263),
    .CK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .QN(_00537_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[61]$_DFFE_PN0P_  (.D(_01857_),
    .RN(net256),
    .CK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .QN(_01065_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[620]$_DFFE_PN0P_  (.D(_01858_),
    .RN(net261),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .QN(_00236_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[621]$_DFFE_PN0P_  (.D(_01859_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .QN(_00587_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[622]$_DFFE_PN0P_  (.D(_01860_),
    .RN(net263),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .QN(_00618_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[623]$_DFFE_PN0P_  (.D(_01861_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .QN(_00649_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[624]$_DFFE_PN0P_  (.D(_01862_),
    .RN(net263),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .QN(_00680_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[625]$_DFFE_PN0P_  (.D(_01863_),
    .RN(net257),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .QN(_00711_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[626]$_DFFE_PN0P_  (.D(_01864_),
    .RN(net255),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .QN(_00742_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[627]$_DFFE_PN0P_  (.D(_01865_),
    .RN(net255),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .QN(_00773_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[628]$_DFFE_PN0P_  (.D(_01866_),
    .RN(net260),
    .CK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .QN(_00804_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[629]$_DFFE_PN0P_  (.D(_01867_),
    .RN(net259),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .QN(_00835_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[62]$_DFFE_PN0P_  (.D(_01868_),
    .RN(net257),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .QN(_01096_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[630]$_DFFE_PN0P_  (.D(_01869_),
    .RN(net257),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .QN(_00866_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[631]$_DFFE_PN0P_  (.D(_01870_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .QN(_00897_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[632]$_DFFE_PN0P_  (.D(_01871_),
    .RN(net257),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .QN(_00928_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[633]$_DFFE_PN0P_  (.D(_01872_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .QN(_00959_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[634]$_DFFE_PN0P_  (.D(_01873_),
    .RN(net262),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .QN(_00990_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[635]$_DFFE_PN0P_  (.D(_01874_),
    .RN(net257),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .QN(_01021_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[636]$_DFFE_PN0P_  (.D(_01875_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .QN(_01052_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[637]$_DFFE_PN0P_  (.D(_01876_),
    .RN(net266),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .QN(_01083_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[638]$_DFFE_PN0P_  (.D(_01877_),
    .RN(net262),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .QN(_01114_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[639]$_DFFE_PN0P_  (.D(_01878_),
    .RN(net266),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .QN(_01145_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[63]$_DFFE_PN0P_  (.D(_01879_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .QN(_01127_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[640]$_DFFE_PN0P_  (.D(_01880_),
    .RN(net264),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .QN(_00205_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[641]$_DFFE_PN0P_  (.D(_01881_),
    .RN(net265),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .QN(_00160_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[642]$_DFFE_PN0P_  (.D(_01882_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .QN(_00267_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[643]$_DFFE_PN0P_  (.D(_01883_),
    .RN(net267),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .QN(_00298_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[644]$_DFFE_PN0P_  (.D(_01884_),
    .RN(net264),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .QN(_00328_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[645]$_DFFE_PN0P_  (.D(_01885_),
    .RN(net264),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .QN(_00358_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[646]$_DFFE_PN0P_  (.D(_01886_),
    .RN(net258),
    .CK(clknet_leaf_85_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .QN(_00388_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[647]$_DFFE_PN0P_  (.D(_01887_),
    .RN(net262),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .QN(_00418_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[648]$_DFFE_PN0P_  (.D(_01888_),
    .RN(net267),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .QN(_00448_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[649]$_DFFE_PN0P_  (.D(_01889_),
    .RN(net267),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .QN(_00478_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[64]$_DFFE_PN0P_  (.D(_01890_),
    .RN(net267),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .QN(_00187_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[650]$_DFFE_PN0P_  (.D(_01891_),
    .RN(net262),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .QN(_00508_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[651]$_DFFE_PN0P_  (.D(_01892_),
    .RN(net263),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .QN(_00538_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[652]$_DFFE_PN0P_  (.D(_01893_),
    .RN(net261),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .QN(_00237_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[653]$_DFFE_PN0P_  (.D(_01894_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .QN(_00588_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[654]$_DFFE_PN0P_  (.D(_01895_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .QN(_00619_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[655]$_DFFE_PN0P_  (.D(_01896_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .QN(_00650_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[656]$_DFFE_PN0P_  (.D(_01897_),
    .RN(net263),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .QN(_00681_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[657]$_DFFE_PN0P_  (.D(_01898_),
    .RN(net257),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .QN(_00712_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[658]$_DFFE_PN0P_  (.D(_01899_),
    .RN(net255),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .QN(_00743_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[659]$_DFFE_PN0P_  (.D(_01900_),
    .RN(net255),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .QN(_00774_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[65]$_DFFE_PN0P_  (.D(_01901_),
    .RN(net266),
    .CK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .QN(_00142_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[660]$_DFFE_PN0P_  (.D(_01902_),
    .RN(net260),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .QN(_00805_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[661]$_DFFE_PN0P_  (.D(_01903_),
    .RN(net259),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .QN(_00836_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[662]$_DFFE_PN0P_  (.D(_01904_),
    .RN(net257),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .QN(_00867_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[663]$_DFFE_PN0P_  (.D(_01905_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .QN(_00898_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[664]$_DFFE_PN0P_  (.D(_01906_),
    .RN(net256),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .QN(_00929_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[665]$_DFFE_PN0P_  (.D(_01907_),
    .RN(net259),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .QN(_00960_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[666]$_DFFE_PN0P_  (.D(_01908_),
    .RN(net262),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .QN(_00991_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[667]$_DFFE_PN0P_  (.D(_01909_),
    .RN(net257),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .QN(_01022_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[668]$_DFFE_PN0P_  (.D(_01910_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .QN(_01053_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[669]$_DFFE_PN0P_  (.D(_01911_),
    .RN(net266),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .QN(_01084_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[66]$_DFFE_PN0P_  (.D(_01912_),
    .RN(net264),
    .CK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .QN(_00249_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[670]$_DFFE_PN0P_  (.D(_01913_),
    .RN(net262),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .QN(_01115_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[671]$_DFFE_PN0P_  (.D(_01914_),
    .RN(net262),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .QN(_01146_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[672]$_DFFE_PN0P_  (.D(_01915_),
    .RN(net264),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .QN(_00206_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[673]$_DFFE_PN0P_  (.D(_01916_),
    .RN(net266),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .QN(_00161_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[674]$_DFFE_PN0P_  (.D(_01917_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .QN(_00268_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[675]$_DFFE_PN0P_  (.D(_01918_),
    .RN(net267),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .QN(_00299_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[676]$_DFFE_PN0P_  (.D(_01919_),
    .RN(net264),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .QN(_00329_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[677]$_DFFE_PN0P_  (.D(_01920_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .QN(_00359_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[678]$_DFFE_PN0P_  (.D(_01921_),
    .RN(net258),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .QN(_00389_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[679]$_DFFE_PN0P_  (.D(_01922_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .QN(_00419_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[67]$_DFFE_PN0P_  (.D(_01923_),
    .RN(net268),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .QN(_00280_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[680]$_DFFE_PN0P_  (.D(_01924_),
    .RN(net267),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .QN(_00449_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[681]$_DFFE_PN0P_  (.D(_01925_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .QN(_00479_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[682]$_DFFE_PN0P_  (.D(_01926_),
    .RN(net266),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .QN(_00509_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[683]$_DFFE_PN0P_  (.D(_01927_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .QN(_00539_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[684]$_DFFE_PN0P_  (.D(_01928_),
    .RN(net261),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .QN(_00238_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[685]$_DFFE_PN0P_  (.D(_01929_),
    .RN(net263),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .QN(_00589_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[686]$_DFFE_PN0P_  (.D(_01930_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .QN(_00620_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[687]$_DFFE_PN0P_  (.D(_01931_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .QN(_00651_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[688]$_DFFE_PN0P_  (.D(_01932_),
    .RN(net263),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .QN(_00682_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[689]$_DFFE_PN0P_  (.D(_01933_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .QN(_00713_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[68]$_DFFE_PN0P_  (.D(_01934_),
    .RN(net264),
    .CK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .QN(_00310_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[690]$_DFFE_PN0P_  (.D(_01935_),
    .RN(net255),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .QN(_00744_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[691]$_DFFE_PN0P_  (.D(_01936_),
    .RN(net255),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .QN(_00775_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[692]$_DFFE_PN0P_  (.D(_01937_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .QN(_00806_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[693]$_DFFE_PN0P_  (.D(_01938_),
    .RN(net257),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .QN(_00837_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[694]$_DFFE_PN0P_  (.D(_01939_),
    .RN(net257),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .QN(_00868_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[695]$_DFFE_PN0P_  (.D(_01940_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .QN(_00899_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[696]$_DFFE_PN0P_  (.D(_01941_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .QN(_00930_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[697]$_DFFE_PN0P_  (.D(_01942_),
    .RN(net257),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .QN(_00961_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[698]$_DFFE_PN0P_  (.D(_01943_),
    .RN(net262),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .QN(_00992_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[699]$_DFFE_PN0P_  (.D(_01944_),
    .RN(net257),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .QN(_01023_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[69]$_DFFE_PN0P_  (.D(_01945_),
    .RN(net264),
    .CK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .QN(_00340_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[6]$_DFFE_PN0P_  (.D(_01946_),
    .RN(net262),
    .CK(clknet_leaf_69_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .QN(_14021_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[700]$_DFFE_PN0P_  (.D(_01947_),
    .RN(net256),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .QN(_01054_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[701]$_DFFE_PN0P_  (.D(_01948_),
    .RN(net266),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .QN(_01085_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[702]$_DFFE_PN0P_  (.D(_01949_),
    .RN(net262),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .QN(_01116_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[703]$_DFFE_PN0P_  (.D(_01950_),
    .RN(net265),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .QN(_01147_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[704]$_DFFE_PN0P_  (.D(_01951_),
    .RN(net264),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .QN(_00207_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[705]$_DFFE_PN0P_  (.D(_01952_),
    .RN(net265),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .QN(_00162_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[706]$_DFFE_PN0P_  (.D(_01953_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .QN(_00269_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[707]$_DFFE_PN0P_  (.D(_01954_),
    .RN(net267),
    .CK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .QN(_00300_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[708]$_DFFE_PN0P_  (.D(_01955_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .QN(_00330_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[709]$_DFFE_PN0P_  (.D(_01956_),
    .RN(net264),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .QN(_00360_));
 DFFR_X2 \gen_regfile_ff.register_file_i.rf_reg_q[70]$_DFFE_PN0P_  (.D(_01957_),
    .RN(net256),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .QN(_00370_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[710]$_DFFE_PN0P_  (.D(_01958_),
    .RN(net258),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .QN(_00390_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[711]$_DFFE_PN0P_  (.D(_01959_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .QN(_00420_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[712]$_DFFE_PN0P_  (.D(_01960_),
    .RN(net267),
    .CK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .QN(_00450_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[713]$_DFFE_PN0P_  (.D(_01961_),
    .RN(net267),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .QN(_00480_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[714]$_DFFE_PN0P_  (.D(_01962_),
    .RN(net262),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .QN(_00510_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[715]$_DFFE_PN0P_  (.D(_01963_),
    .RN(net268),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .QN(_00540_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[716]$_DFFE_PN0P_  (.D(_01964_),
    .RN(net261),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .QN(_00239_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[717]$_DFFE_PN0P_  (.D(_01965_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .QN(_00590_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[718]$_DFFE_PN0P_  (.D(_01966_),
    .RN(net263),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .QN(_00621_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[719]$_DFFE_PN0P_  (.D(_01967_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .QN(_00652_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[71]$_DFFE_PN0P_  (.D(_01968_),
    .RN(net262),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .QN(_00400_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[720]$_DFFE_PN0P_  (.D(_01969_),
    .RN(net263),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .QN(_00683_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[721]$_DFFE_PN0P_  (.D(_01970_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .QN(_00714_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[722]$_DFFE_PN0P_  (.D(_01971_),
    .RN(net255),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .QN(_00745_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[723]$_DFFE_PN0P_  (.D(_01972_),
    .RN(net255),
    .CK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .QN(_00776_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[724]$_DFFE_PN0P_  (.D(_01973_),
    .RN(net260),
    .CK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .QN(_00807_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[725]$_DFFE_PN0P_  (.D(_01974_),
    .RN(net257),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .QN(_00838_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[726]$_DFFE_PN0P_  (.D(_01975_),
    .RN(net257),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .QN(_00869_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[727]$_DFFE_PN0P_  (.D(_01976_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .QN(_00900_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[728]$_DFFE_PN0P_  (.D(_01977_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .QN(_00931_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[729]$_DFFE_PN0P_  (.D(_01978_),
    .RN(net257),
    .CK(clknet_leaf_93_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .QN(_00962_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[72]$_DFFE_PN0P_  (.D(_01979_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .QN(_00430_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[730]$_DFFE_PN0P_  (.D(_01980_),
    .RN(net262),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .QN(_00993_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[731]$_DFFE_PN0P_  (.D(_01981_),
    .RN(net257),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .QN(_01024_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[732]$_DFFE_PN0P_  (.D(_01982_),
    .RN(net256),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .QN(_01055_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[733]$_DFFE_PN0P_  (.D(_01983_),
    .RN(net266),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .QN(_01086_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[734]$_DFFE_PN0P_  (.D(_01984_),
    .RN(net262),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .QN(_01117_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[735]$_DFFE_PN0P_  (.D(_01985_),
    .RN(net265),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .QN(_01148_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[736]$_DFFE_PN0P_  (.D(_01986_),
    .RN(net267),
    .CK(clknet_leaf_121_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .QN(_00208_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[737]$_DFFE_PN0P_  (.D(_01987_),
    .RN(net266),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .QN(_00163_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[738]$_DFFE_PN0P_  (.D(_01988_),
    .RN(net264),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .QN(_00270_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[739]$_DFFE_PN0P_  (.D(_01989_),
    .RN(net267),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .QN(_00301_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[73]$_DFFE_PN0P_  (.D(_01990_),
    .RN(net267),
    .CK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .QN(_00460_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[740]$_DFFE_PN0P_  (.D(_01991_),
    .RN(net264),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .QN(_00331_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[741]$_DFFE_PN0P_  (.D(_01992_),
    .RN(net264),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .QN(_00361_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[742]$_DFFE_PN0P_  (.D(_01993_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .QN(_00391_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[743]$_DFFE_PN0P_  (.D(_01994_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .QN(_00421_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[744]$_DFFE_PN0P_  (.D(_01995_),
    .RN(net268),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .QN(_00451_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[745]$_DFFE_PN0P_  (.D(_01996_),
    .RN(net268),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .QN(_00481_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[746]$_DFFE_PN0P_  (.D(_01997_),
    .RN(net266),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .QN(_00511_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[747]$_DFFE_PN0P_  (.D(_01998_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .QN(_00541_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[748]$_DFFE_PN0P_  (.D(_01999_),
    .RN(net261),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .QN(_00240_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[749]$_DFFE_PN0P_  (.D(_02000_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .QN(_00591_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[74]$_DFFE_PN0P_  (.D(_02001_),
    .RN(net262),
    .CK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .QN(_00490_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[750]$_DFFE_PN0P_  (.D(_02002_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .QN(_00622_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[751]$_DFFE_PN0P_  (.D(_02003_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .QN(_00653_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[752]$_DFFE_PN0P_  (.D(_02004_),
    .RN(net263),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .QN(_00684_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[753]$_DFFE_PN0P_  (.D(_02005_),
    .RN(net257),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .QN(_00715_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[754]$_DFFE_PN0P_  (.D(_02006_),
    .RN(net263),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .QN(_00746_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[755]$_DFFE_PN0P_  (.D(_02007_),
    .RN(net255),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .QN(_00777_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[756]$_DFFE_PN0P_  (.D(_02008_),
    .RN(net260),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .QN(_00808_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[757]$_DFFE_PN0P_  (.D(_02009_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .QN(_00839_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[758]$_DFFE_PN0P_  (.D(_02010_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .QN(_00870_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[759]$_DFFE_PN0P_  (.D(_02011_),
    .RN(net261),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .QN(_00901_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[75]$_DFFE_PN0P_  (.D(_02012_),
    .RN(net268),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .QN(_00520_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[760]$_DFFE_PN0P_  (.D(_02013_),
    .RN(net257),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .QN(_00932_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[761]$_DFFE_PN0P_  (.D(_02014_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .QN(_00963_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[762]$_DFFE_PN0P_  (.D(_02015_),
    .RN(net256),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .QN(_00994_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[763]$_DFFE_PN0P_  (.D(_02016_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .QN(_01025_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[764]$_DFFE_PN0P_  (.D(_02017_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .QN(_01056_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[765]$_DFFE_PN0P_  (.D(_02018_),
    .RN(net262),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .QN(_01087_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[766]$_DFFE_PN0P_  (.D(_02019_),
    .RN(net256),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .QN(_01118_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[767]$_DFFE_PN0P_  (.D(_02020_),
    .RN(net265),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .QN(_01149_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[768]$_DFFE_PN0P_  (.D(_02021_),
    .RN(net267),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .QN(_00209_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[769]$_DFFE_PN0P_  (.D(_02022_),
    .RN(net266),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .QN(_00164_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[76]$_DFFE_PN0P_  (.D(_02023_),
    .RN(net261),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .QN(_00219_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[770]$_DFFE_PN0P_  (.D(_02024_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .QN(_00271_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[771]$_DFFE_PN0P_  (.D(_02025_),
    .RN(net267),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .QN(_00302_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[772]$_DFFE_PN0P_  (.D(_02026_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .QN(_00332_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[773]$_DFFE_PN0P_  (.D(_02027_),
    .RN(net264),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .QN(_00362_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[774]$_DFFE_PN0P_  (.D(_02028_),
    .RN(net259),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .QN(_00392_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[775]$_DFFE_PN0P_  (.D(_02029_),
    .RN(net268),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .QN(_00422_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[776]$_DFFE_PN0P_  (.D(_02030_),
    .RN(net268),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .QN(_00452_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[777]$_DFFE_PN0P_  (.D(_02031_),
    .RN(net268),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .QN(_00482_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[778]$_DFFE_PN0P_  (.D(_02032_),
    .RN(net266),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .QN(_00512_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[779]$_DFFE_PN0P_  (.D(_02033_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .QN(_00542_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[77]$_DFFE_PN0P_  (.D(_02034_),
    .RN(net261),
    .CK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .QN(_00570_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[780]$_DFFE_PN0P_  (.D(_02035_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .QN(_00241_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[781]$_DFFE_PN0P_  (.D(_02036_),
    .RN(net263),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .QN(_00592_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[782]$_DFFE_PN0P_  (.D(_02037_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .QN(_00623_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[783]$_DFFE_PN0P_  (.D(_02038_),
    .RN(net255),
    .CK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .QN(_00654_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[784]$_DFFE_PN0P_  (.D(_02039_),
    .RN(net263),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .QN(_00685_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[785]$_DFFE_PN0P_  (.D(_02040_),
    .RN(net257),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .QN(_00716_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[786]$_DFFE_PN0P_  (.D(_02041_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .QN(_00747_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[787]$_DFFE_PN0P_  (.D(_02042_),
    .RN(net255),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .QN(_00778_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[788]$_DFFE_PN0P_  (.D(_02043_),
    .RN(net260),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .QN(_00809_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[789]$_DFFE_PN0P_  (.D(_02044_),
    .RN(net259),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .QN(_00840_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[78]$_DFFE_PN0P_  (.D(_02045_),
    .RN(net261),
    .CK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .QN(_00601_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[790]$_DFFE_PN0P_  (.D(_02046_),
    .RN(net259),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .QN(_00871_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[791]$_DFFE_PN0P_  (.D(_02047_),
    .RN(net262),
    .CK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .QN(_00902_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[792]$_DFFE_PN0P_  (.D(_02048_),
    .RN(net257),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .QN(_00933_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[793]$_DFFE_PN0P_  (.D(_02049_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .QN(_00964_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[794]$_DFFE_PN0P_  (.D(_02050_),
    .RN(net256),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .QN(_00995_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[795]$_DFFE_PN0P_  (.D(_02051_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .QN(_01026_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[796]$_DFFE_PN0P_  (.D(_02052_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .QN(_01057_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[797]$_DFFE_PN0P_  (.D(_02053_),
    .RN(net262),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .QN(_01088_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[798]$_DFFE_PN0P_  (.D(_02054_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .QN(_01119_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[799]$_DFFE_PN0P_  (.D(_02055_),
    .RN(net265),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .QN(_01150_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[79]$_DFFE_PN0P_  (.D(_02056_),
    .RN(net261),
    .CK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .QN(_00632_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[7]$_DFFE_PN0P_  (.D(_02057_),
    .RN(net268),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .QN(_14020_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[800]$_DFFE_PN0P_  (.D(_02058_),
    .RN(net267),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .QN(_00210_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[801]$_DFFE_PN0P_  (.D(_02059_),
    .RN(net266),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .QN(_00165_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[802]$_DFFE_PN0P_  (.D(_02060_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .QN(_00272_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[803]$_DFFE_PN0P_  (.D(_02061_),
    .RN(net267),
    .CK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .QN(_00303_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[804]$_DFFE_PN0P_  (.D(_02062_),
    .RN(net264),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .QN(_00333_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[805]$_DFFE_PN0P_  (.D(_02063_),
    .RN(net264),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .QN(_00363_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[806]$_DFFE_PN0P_  (.D(_02064_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .QN(_00393_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[807]$_DFFE_PN0P_  (.D(_02065_),
    .RN(net268),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .QN(_00423_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[808]$_DFFE_PN0P_  (.D(_02066_),
    .RN(net268),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .QN(_00453_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[809]$_DFFE_PN0P_  (.D(_02067_),
    .RN(net255),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .QN(_00483_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[80]$_DFFE_PN0P_  (.D(_02068_),
    .RN(net261),
    .CK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .QN(_00663_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[810]$_DFFE_PN0P_  (.D(_02069_),
    .RN(net266),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .QN(_00513_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[811]$_DFFE_PN0P_  (.D(_02070_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .QN(_00543_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[812]$_DFFE_PN0P_  (.D(_02071_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .QN(_00242_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[813]$_DFFE_PN0P_  (.D(_02072_),
    .RN(net263),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .QN(_00593_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[814]$_DFFE_PN0P_  (.D(_02073_),
    .RN(net263),
    .CK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .QN(_00624_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[815]$_DFFE_PN0P_  (.D(_02074_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .QN(_00655_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[816]$_DFFE_PN0P_  (.D(_02075_),
    .RN(net263),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .QN(_00686_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[817]$_DFFE_PN0P_  (.D(_02076_),
    .RN(net256),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .QN(_00717_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[818]$_DFFE_PN0P_  (.D(_02077_),
    .RN(net263),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .QN(_00748_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[819]$_DFFE_PN0P_  (.D(_02078_),
    .RN(net255),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .QN(_00779_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[81]$_DFFE_PN0P_  (.D(_02079_),
    .RN(net257),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .QN(_00694_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[820]$_DFFE_PN0P_  (.D(_02080_),
    .RN(net259),
    .CK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .QN(_00810_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[821]$_DFFE_PN0P_  (.D(_02081_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .QN(_00841_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[822]$_DFFE_PN0P_  (.D(_02082_),
    .RN(net259),
    .CK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .QN(_00872_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[823]$_DFFE_PN0P_  (.D(_02083_),
    .RN(net262),
    .CK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .QN(_00903_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[824]$_DFFE_PN0P_  (.D(_02084_),
    .RN(net257),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .QN(_00934_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[825]$_DFFE_PN0P_  (.D(_02085_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .QN(_00965_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[826]$_DFFE_PN0P_  (.D(_02086_),
    .RN(net256),
    .CK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .QN(_00996_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[827]$_DFFE_PN0P_  (.D(_02087_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .QN(_01027_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[828]$_DFFE_PN0P_  (.D(_02088_),
    .RN(net256),
    .CK(clknet_leaf_99_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .QN(_01058_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[829]$_DFFE_PN0P_  (.D(_02089_),
    .RN(net262),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .QN(_01089_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[82]$_DFFE_PN0P_  (.D(_02090_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .QN(_00725_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[830]$_DFFE_PN0P_  (.D(_02091_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .QN(_01120_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[831]$_DFFE_PN0P_  (.D(_02092_),
    .RN(net266),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .QN(_01151_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[832]$_DFFE_PN0P_  (.D(_02093_),
    .RN(net264),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .QN(_00211_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[833]$_DFFE_PN0P_  (.D(_02094_),
    .RN(net266),
    .CK(clknet_leaf_116_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .QN(_00166_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[834]$_DFFE_PN0P_  (.D(_02095_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .QN(_00273_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[835]$_DFFE_PN0P_  (.D(_02096_),
    .RN(net268),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .QN(_00304_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[836]$_DFFE_PN0P_  (.D(_02097_),
    .RN(net264),
    .CK(clknet_leaf_135_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .QN(_00334_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[837]$_DFFE_PN0P_  (.D(_02098_),
    .RN(net264),
    .CK(clknet_leaf_132_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .QN(_00364_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[838]$_DFFE_PN0P_  (.D(_02099_),
    .RN(net259),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .QN(_00394_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[839]$_DFFE_PN0P_  (.D(_02100_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .QN(_00424_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[83]$_DFFE_PN0P_  (.D(_02101_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .QN(_00756_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[840]$_DFFE_PN0P_  (.D(_02102_),
    .RN(net267),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .QN(_00454_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[841]$_DFFE_PN0P_  (.D(_02103_),
    .RN(net268),
    .CK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .QN(_00484_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[842]$_DFFE_PN0P_  (.D(_02104_),
    .RN(net266),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .QN(_00514_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[843]$_DFFE_PN0P_  (.D(_02105_),
    .RN(net255),
    .CK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .QN(_00544_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[844]$_DFFE_PN0P_  (.D(_02106_),
    .RN(net261),
    .CK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .QN(_00243_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[845]$_DFFE_PN0P_  (.D(_02107_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .QN(_00594_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[846]$_DFFE_PN0P_  (.D(_02108_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .QN(_00625_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[847]$_DFFE_PN0P_  (.D(_02109_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .QN(_00656_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[848]$_DFFE_PN0P_  (.D(_02110_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .QN(_00687_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[849]$_DFFE_PN0P_  (.D(_02111_),
    .RN(net256),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .QN(_00718_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[84]$_DFFE_PN0P_  (.D(_02112_),
    .RN(net259),
    .CK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .QN(_00787_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[850]$_DFFE_PN0P_  (.D(_02113_),
    .RN(net263),
    .CK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .QN(_00749_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[851]$_DFFE_PN0P_  (.D(_02114_),
    .RN(net255),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .QN(_00780_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[852]$_DFFE_PN0P_  (.D(_02115_),
    .RN(net260),
    .CK(clknet_leaf_61_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .QN(_00811_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[853]$_DFFE_PN0P_  (.D(_02116_),
    .RN(net257),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .QN(_00842_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[854]$_DFFE_PN0P_  (.D(_02117_),
    .RN(net259),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .QN(_00873_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[855]$_DFFE_PN0P_  (.D(_02118_),
    .RN(net261),
    .CK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .QN(_00904_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[856]$_DFFE_PN0P_  (.D(_02119_),
    .RN(net257),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .QN(_00935_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[857]$_DFFE_PN0P_  (.D(_02120_),
    .RN(net259),
    .CK(clknet_leaf_92_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .QN(_00966_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[858]$_DFFE_PN0P_  (.D(_02121_),
    .RN(net256),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .QN(_00997_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[859]$_DFFE_PN0P_  (.D(_02122_),
    .RN(net259),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .QN(_01028_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[85]$_DFFE_PN0P_  (.D(_02123_),
    .RN(net257),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .QN(_00818_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[860]$_DFFE_PN0P_  (.D(_02124_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .QN(_01059_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[861]$_DFFE_PN0P_  (.D(_02125_),
    .RN(net262),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .QN(_01090_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[862]$_DFFE_PN0P_  (.D(_02126_),
    .RN(net256),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .QN(_01121_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[863]$_DFFE_PN0P_  (.D(_02127_),
    .RN(net265),
    .CK(clknet_leaf_114_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .QN(_01152_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[864]$_DFFE_PN0P_  (.D(_02128_),
    .RN(net267),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .QN(_00212_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[865]$_DFFE_PN0P_  (.D(_02129_),
    .RN(net265),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .QN(_00167_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[866]$_DFFE_PN0P_  (.D(_02130_),
    .RN(net264),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .QN(_00274_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[867]$_DFFE_PN0P_  (.D(_02131_),
    .RN(net268),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .QN(_00305_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[868]$_DFFE_PN0P_  (.D(_02132_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .QN(_00335_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[869]$_DFFE_PN0P_  (.D(_02133_),
    .RN(net264),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .QN(_00365_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[86]$_DFFE_PN0P_  (.D(_02134_),
    .RN(net257),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .QN(_00849_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[870]$_DFFE_PN0P_  (.D(_02135_),
    .RN(net257),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .QN(_00395_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[871]$_DFFE_PN0P_  (.D(_02136_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .QN(_00425_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[872]$_DFFE_PN0P_  (.D(_02137_),
    .RN(net267),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .QN(_00455_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[873]$_DFFE_PN0P_  (.D(_02138_),
    .RN(net268),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .QN(_00485_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[874]$_DFFE_PN0P_  (.D(_02139_),
    .RN(net266),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .QN(_00515_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[875]$_DFFE_PN0P_  (.D(_02140_),
    .RN(net263),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .QN(_00545_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[876]$_DFFE_PN0P_  (.D(_02141_),
    .RN(net261),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .QN(_00244_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[877]$_DFFE_PN0P_  (.D(_02142_),
    .RN(net263),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .QN(_00595_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[878]$_DFFE_PN0P_  (.D(_02143_),
    .RN(net263),
    .CK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .QN(_00626_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[879]$_DFFE_PN0P_  (.D(_02144_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .QN(_00657_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[87]$_DFFE_PN0P_  (.D(_02145_),
    .RN(net261),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .QN(_00880_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[880]$_DFFE_PN0P_  (.D(_02146_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .QN(_00688_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[881]$_DFFE_PN0P_  (.D(_02147_),
    .RN(net256),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .QN(_00719_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[882]$_DFFE_PN0P_  (.D(_02148_),
    .RN(net255),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .QN(_00750_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[883]$_DFFE_PN0P_  (.D(_02149_),
    .RN(net255),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .QN(_00781_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[884]$_DFFE_PN0P_  (.D(_02150_),
    .RN(net260),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .QN(_00812_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[885]$_DFFE_PN0P_  (.D(_02151_),
    .RN(net257),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .QN(_00843_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[886]$_DFFE_PN0P_  (.D(_02152_),
    .RN(net257),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .QN(_00874_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[887]$_DFFE_PN0P_  (.D(_02153_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .QN(_00905_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[888]$_DFFE_PN0P_  (.D(_02154_),
    .RN(net257),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .QN(_00936_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[889]$_DFFE_PN0P_  (.D(_02155_),
    .RN(net257),
    .CK(clknet_leaf_91_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .QN(_00967_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[88]$_DFFE_PN0P_  (.D(_02156_),
    .RN(net257),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .QN(_00911_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[890]$_DFFE_PN0P_  (.D(_02157_),
    .RN(net256),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .QN(_00998_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[891]$_DFFE_PN0P_  (.D(_02158_),
    .RN(net257),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .QN(_01029_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[892]$_DFFE_PN0P_  (.D(_02159_),
    .RN(net256),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .QN(_01060_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[893]$_DFFE_PN0P_  (.D(_02160_),
    .RN(net262),
    .CK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .QN(_01091_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[894]$_DFFE_PN0P_  (.D(_02161_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .QN(_01122_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[895]$_DFFE_PN0P_  (.D(_02162_),
    .RN(net265),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .QN(_01153_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[896]$_DFFE_PN0P_  (.D(_02163_),
    .RN(net267),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .QN(_00213_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[897]$_DFFE_PN0P_  (.D(_02164_),
    .RN(net265),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .QN(_00168_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[898]$_DFFE_PN0P_  (.D(_02165_),
    .RN(net264),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .QN(_00275_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[899]$_DFFE_PN0P_  (.D(_02166_),
    .RN(net268),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .QN(_00306_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[89]$_DFFE_PN0P_  (.D(_02167_),
    .RN(net257),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .QN(_00942_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[8]$_DFFE_PN0P_  (.D(_02168_),
    .RN(net268),
    .CK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .QN(_14019_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[900]$_DFFE_PN0P_  (.D(_02169_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .QN(_00336_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[901]$_DFFE_PN0P_  (.D(_02170_),
    .RN(net264),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .QN(_00366_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[902]$_DFFE_PN0P_  (.D(_02171_),
    .RN(net257),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .QN(_00396_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[903]$_DFFE_PN0P_  (.D(_02172_),
    .RN(net262),
    .CK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .QN(_00426_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[904]$_DFFE_PN0P_  (.D(_02173_),
    .RN(net268),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .QN(_00456_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[905]$_DFFE_PN0P_  (.D(_02174_),
    .RN(net268),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .QN(_00486_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[906]$_DFFE_PN0P_  (.D(_02175_),
    .RN(net266),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .QN(_00516_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[907]$_DFFE_PN0P_  (.D(_02176_),
    .RN(net263),
    .CK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .QN(_00546_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[908]$_DFFE_PN0P_  (.D(_02177_),
    .RN(net261),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .QN(_00245_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[909]$_DFFE_PN0P_  (.D(_02178_),
    .RN(net263),
    .CK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .QN(_00596_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[90]$_DFFE_PN0P_  (.D(_02179_),
    .RN(net257),
    .CK(clknet_leaf_73_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .QN(_00973_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[910]$_DFFE_PN0P_  (.D(_02180_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .QN(_00627_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[911]$_DFFE_PN0P_  (.D(_02181_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .QN(_00658_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[912]$_DFFE_PN0P_  (.D(_02182_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .QN(_00689_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[913]$_DFFE_PN0P_  (.D(_02183_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .QN(_00720_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[914]$_DFFE_PN0P_  (.D(_02184_),
    .RN(net255),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .QN(_00751_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[915]$_DFFE_PN0P_  (.D(_02185_),
    .RN(net255),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .QN(_00782_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[916]$_DFFE_PN0P_  (.D(_02186_),
    .RN(net260),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .QN(_00813_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[917]$_DFFE_PN0P_  (.D(_02187_),
    .RN(net257),
    .CK(clknet_leaf_88_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .QN(_00844_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[918]$_DFFE_PN0P_  (.D(_02188_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .QN(_00875_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[919]$_DFFE_PN0P_  (.D(_02189_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .QN(_00906_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[91]$_DFFE_PN0P_  (.D(_02190_),
    .RN(net257),
    .CK(clknet_leaf_76_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .QN(_01004_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[920]$_DFFE_PN0P_  (.D(_02191_),
    .RN(net256),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .QN(_00937_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[921]$_DFFE_PN0P_  (.D(_02192_),
    .RN(net257),
    .CK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .QN(_00968_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[922]$_DFFE_PN0P_  (.D(_02193_),
    .RN(net256),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .QN(_00999_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[923]$_DFFE_PN0P_  (.D(_02194_),
    .RN(net256),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .QN(_01030_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[924]$_DFFE_PN0P_  (.D(_02195_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .QN(_01061_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[925]$_DFFE_PN0P_  (.D(_02196_),
    .RN(net265),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .QN(_01092_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[926]$_DFFE_PN0P_  (.D(_02197_),
    .RN(net256),
    .CK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .QN(_01123_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[927]$_DFFE_PN0P_  (.D(_02198_),
    .RN(net266),
    .CK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .QN(_01154_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[928]$_DFFE_PN0P_  (.D(_02199_),
    .RN(net264),
    .CK(clknet_leaf_120_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .QN(_00214_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[929]$_DFFE_PN0P_  (.D(_02200_),
    .RN(net265),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .QN(_00169_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[92]$_DFFE_PN0P_  (.D(_02201_),
    .RN(net257),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .QN(_01035_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[930]$_DFFE_PN0P_  (.D(_02202_),
    .RN(net264),
    .CK(clknet_leaf_118_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .QN(_00276_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[931]$_DFFE_PN0P_  (.D(_02203_),
    .RN(net268),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .QN(_00307_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[932]$_DFFE_PN0P_  (.D(_02204_),
    .RN(net264),
    .CK(clknet_leaf_133_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .QN(_00337_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[933]$_DFFE_PN0P_  (.D(_02205_),
    .RN(net264),
    .CK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .QN(_00367_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[934]$_DFFE_PN0P_  (.D(_02206_),
    .RN(net259),
    .CK(clknet_leaf_86_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .QN(_00397_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[935]$_DFFE_PN0P_  (.D(_02207_),
    .RN(net268),
    .CK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .QN(_00427_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[936]$_DFFE_PN0P_  (.D(_02208_),
    .RN(net267),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .QN(_00457_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[937]$_DFFE_PN0P_  (.D(_02209_),
    .RN(net268),
    .CK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .QN(_00487_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[938]$_DFFE_PN0P_  (.D(_02210_),
    .RN(net266),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .QN(_00517_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[939]$_DFFE_PN0P_  (.D(_02211_),
    .RN(net263),
    .CK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .QN(_00547_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[93]$_DFFE_PN0P_  (.D(_02212_),
    .RN(net256),
    .CK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .QN(_01066_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[940]$_DFFE_PN0P_  (.D(_02213_),
    .RN(net261),
    .CK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .QN(_00246_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[941]$_DFFE_PN0P_  (.D(_02214_),
    .RN(net263),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .QN(_00597_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[942]$_DFFE_PN0P_  (.D(_02215_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .QN(_00628_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[943]$_DFFE_PN0P_  (.D(_02216_),
    .RN(net263),
    .CK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .QN(_00659_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[944]$_DFFE_PN0P_  (.D(_02217_),
    .RN(net263),
    .CK(clknet_leaf_37_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .QN(_00690_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[945]$_DFFE_PN0P_  (.D(_02218_),
    .RN(net256),
    .CK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .QN(_00721_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[946]$_DFFE_PN0P_  (.D(_02219_),
    .RN(net255),
    .CK(clknet_leaf_45_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .QN(_00752_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[947]$_DFFE_PN0P_  (.D(_02220_),
    .RN(net255),
    .CK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .QN(_00783_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[948]$_DFFE_PN0P_  (.D(_02221_),
    .RN(net260),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .QN(_00814_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[949]$_DFFE_PN0P_  (.D(_02222_),
    .RN(net257),
    .CK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .QN(_00845_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[94]$_DFFE_PN0P_  (.D(_02223_),
    .RN(net256),
    .CK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .QN(_01097_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[950]$_DFFE_PN0P_  (.D(_02224_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .QN(_00876_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[951]$_DFFE_PN0P_  (.D(_02225_),
    .RN(net261),
    .CK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .QN(_00907_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[952]$_DFFE_PN0P_  (.D(_02226_),
    .RN(net257),
    .CK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .QN(_00938_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[953]$_DFFE_PN0P_  (.D(_02227_),
    .RN(net257),
    .CK(clknet_leaf_94_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .QN(_00969_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[954]$_DFFE_PN0P_  (.D(_02228_),
    .RN(net256),
    .CK(clknet_leaf_107_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .QN(_01000_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[955]$_DFFE_PN0P_  (.D(_02229_),
    .RN(net257),
    .CK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .QN(_01031_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[956]$_DFFE_PN0P_  (.D(_02230_),
    .RN(net256),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .QN(_01062_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[957]$_DFFE_PN0P_  (.D(_02231_),
    .RN(net265),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .QN(_01093_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[958]$_DFFE_PN0P_  (.D(_02232_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .QN(_01124_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[959]$_DFFE_PN0P_  (.D(_02233_),
    .RN(net265),
    .CK(clknet_leaf_115_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .QN(_01155_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[95]$_DFFE_PN0P_  (.D(_02234_),
    .RN(net266),
    .CK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .QN(_01128_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[960]$_DFFE_PN0P_  (.D(_02235_),
    .RN(net267),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .QN(_00215_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[961]$_DFFE_PN0P_  (.D(_02236_),
    .RN(net265),
    .CK(clknet_leaf_117_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .QN(_00170_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[962]$_DFFE_PN0P_  (.D(_02237_),
    .RN(net264),
    .CK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .QN(_00277_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[963]$_DFFE_PN0P_  (.D(_02238_),
    .RN(net268),
    .CK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .QN(_00308_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[964]$_DFFE_PN0P_  (.D(_02239_),
    .RN(net264),
    .CK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .QN(_00338_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[965]$_DFFE_PN0P_  (.D(_02240_),
    .RN(net264),
    .CK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .QN(_00368_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[966]$_DFFE_PN0P_  (.D(_02241_),
    .RN(net256),
    .CK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .QN(_00398_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[967]$_DFFE_PN0P_  (.D(_02242_),
    .RN(net262),
    .CK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .QN(_00428_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[968]$_DFFE_PN0P_  (.D(_02243_),
    .RN(net268),
    .CK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .QN(_00458_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[969]$_DFFE_PN0P_  (.D(_02244_),
    .RN(net268),
    .CK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .QN(_00488_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[96]$_DFFE_PN0P_  (.D(_02245_),
    .RN(net267),
    .CK(clknet_leaf_123_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .QN(_00188_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[970]$_DFFE_PN0P_  (.D(_02246_),
    .RN(net266),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .QN(_00518_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[971]$_DFFE_PN0P_  (.D(_02247_),
    .RN(net263),
    .CK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .QN(_00548_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[972]$_DFFE_PN0P_  (.D(_02248_),
    .RN(net261),
    .CK(clknet_leaf_50_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .QN(_00247_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[973]$_DFFE_PN0P_  (.D(_02249_),
    .RN(net262),
    .CK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .QN(_00598_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[974]$_DFFE_PN0P_  (.D(_02250_),
    .RN(net263),
    .CK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .QN(_00629_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[975]$_DFFE_PN0P_  (.D(_02251_),
    .RN(net263),
    .CK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .QN(_00660_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[976]$_DFFE_PN0P_  (.D(_02252_),
    .RN(net263),
    .CK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .QN(_00691_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[977]$_DFFE_PN0P_  (.D(_02253_),
    .RN(net256),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .QN(_00722_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[978]$_DFFE_PN0P_  (.D(_02254_),
    .RN(net255),
    .CK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .QN(_00753_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[979]$_DFFE_PN0P_  (.D(_02255_),
    .RN(net255),
    .CK(clknet_leaf_46_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .QN(_00784_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[97]$_DFFE_PN0P_  (.D(_02256_),
    .RN(net266),
    .CK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .QN(_00143_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[980]$_DFFE_PN0P_  (.D(_02257_),
    .RN(net260),
    .CK(clknet_leaf_52_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .QN(_00815_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[981]$_DFFE_PN0P_  (.D(_02258_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .QN(_00846_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[982]$_DFFE_PN0P_  (.D(_02259_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .QN(_00877_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[983]$_DFFE_PN0P_  (.D(_02260_),
    .RN(net261),
    .CK(clknet_leaf_64_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .QN(_00908_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[984]$_DFFE_PN0P_  (.D(_02261_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .QN(_00939_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[985]$_DFFE_PN0P_  (.D(_02262_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .QN(_00970_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[986]$_DFFE_PN0P_  (.D(_02263_),
    .RN(net256),
    .CK(clknet_leaf_105_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .QN(_01001_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[987]$_DFFE_PN0P_  (.D(_02264_),
    .RN(net256),
    .CK(clknet_leaf_96_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .QN(_01032_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[988]$_DFFE_PN0P_  (.D(_02265_),
    .RN(net256),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .QN(_01063_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[989]$_DFFE_PN0P_  (.D(_02266_),
    .RN(net265),
    .CK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .QN(_01094_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[98]$_DFFE_PN0P_  (.D(_02267_),
    .RN(net267),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .QN(_00250_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[990]$_DFFE_PN0P_  (.D(_02268_),
    .RN(net265),
    .CK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .QN(_01125_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[991]$_DFFE_PN0P_  (.D(_02269_),
    .RN(net265),
    .CK(clknet_leaf_103_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .QN(_01156_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[99]$_DFFE_PN0P_  (.D(_02270_),
    .RN(net266),
    .CK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .QN(_00281_));
 DFFR_X1 \gen_regfile_ff.register_file_i.rf_reg_q[9]$_DFFE_PN0P_  (.D(_02271_),
    .RN(net268),
    .CK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .QN(_14018_));
 DFFR_X1 \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.D(_02272_),
    .RN(net248),
    .CK(clknet_leaf_116_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .QN(_14017_));
 DFFR_X1 \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.D(_02273_),
    .RN(net248),
    .CK(clknet_leaf_117_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .QN(_14016_));
 DFFR_X1 \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.D(_02274_),
    .RN(net248),
    .CK(clknet_leaf_116_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .QN(_14015_));
 DFFR_X2 \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.D(_02275_),
    .RN(net248),
    .CK(clknet_leaf_117_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .QN(_14014_));
 DFFR_X1 \id_stage_i.controller_i.debug_mode_q$_DFFE_PN0P_  (.D(_02276_),
    .RN(net248),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.debug_mode_i ),
    .QN(_01160_));
 DFFR_X1 \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.exc_req_d ),
    .RN(net248),
    .CK(clknet_leaf_55_clk),
    .Q(\id_stage_i.controller_i.exc_req_q ),
    .QN(_14454_));
 DFFR_X1 \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.illegal_insn_d ),
    .RN(net248),
    .CK(clknet_leaf_55_clk),
    .Q(\id_stage_i.controller_i.illegal_insn_q ),
    .QN(_00557_));
 DFFR_X2 \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.load_err_d ),
    .RN(net248),
    .CK(clknet_leaf_117_clk),
    .Q(\id_stage_i.controller_i.load_err_q ),
    .QN(_14013_));
 DFFR_X2 \id_stage_i.controller_i.nmi_mode_q$_DFFE_PN0P_  (.D(_02277_),
    .RN(net249),
    .CK(clknet_leaf_113_clk),
    .Q(\cs_registers_i.nmi_mode_i ),
    .QN(_14455_));
 DFFR_X2 \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.store_err_d ),
    .RN(net248),
    .CK(clknet_leaf_117_clk),
    .Q(\id_stage_i.controller_i.store_err_q ),
    .QN(_14456_));
 DFFR_X1 \id_stage_i.g_branch_set_flop.branch_set_q$_DFF_PN0_  (.D(\id_stage_i.branch_set_d ),
    .RN(net248),
    .CK(clknet_leaf_118_clk),
    .Q(\id_stage_i.branch_set ),
    .QN(_14012_));
 DFFR_X1 \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.D(_02278_),
    .RN(net248),
    .CK(clknet_leaf_13_clk),
    .Q(\id_stage_i.id_fsm_q ),
    .QN(_14011_));
 DFFR_X1 \id_stage_i.imd_val_q[0]$_DFFE_PN0P_  (.D(_02279_),
    .RN(net265),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .QN(_14010_));
 DFFR_X1 \id_stage_i.imd_val_q[10]$_DFFE_PN0P_  (.D(_02280_),
    .RN(net265),
    .CK(clknet_leaf_21_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .QN(_14009_));
 DFFR_X1 \id_stage_i.imd_val_q[11]$_DFFE_PN0P_  (.D(_02281_),
    .RN(net265),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .QN(_14008_));
 DFFR_X1 \id_stage_i.imd_val_q[12]$_DFFE_PN0P_  (.D(_02282_),
    .RN(net265),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .QN(_14007_));
 DFFR_X1 \id_stage_i.imd_val_q[13]$_DFFE_PN0P_  (.D(_02283_),
    .RN(net265),
    .CK(clknet_leaf_21_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .QN(_14006_));
 DFFR_X1 \id_stage_i.imd_val_q[14]$_DFFE_PN0P_  (.D(_02284_),
    .RN(net265),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .QN(_14005_));
 DFFR_X1 \id_stage_i.imd_val_q[15]$_DFFE_PN0P_  (.D(_02285_),
    .RN(net265),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .QN(_14004_));
 DFFR_X1 \id_stage_i.imd_val_q[16]$_DFFE_PN0P_  (.D(_02286_),
    .RN(net265),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .QN(_14003_));
 DFFR_X1 \id_stage_i.imd_val_q[17]$_DFFE_PN0P_  (.D(_02287_),
    .RN(net246),
    .CK(clknet_leaf_41_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .QN(_14002_));
 DFFR_X1 \id_stage_i.imd_val_q[18]$_DFFE_PN0P_  (.D(_02288_),
    .RN(net265),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .QN(_14001_));
 DFFR_X1 \id_stage_i.imd_val_q[19]$_DFFE_PN0P_  (.D(_02289_),
    .RN(net265),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .QN(_14000_));
 DFFR_X1 \id_stage_i.imd_val_q[1]$_DFFE_PN0P_  (.D(_02290_),
    .RN(net265),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .QN(_13999_));
 DFFR_X1 \id_stage_i.imd_val_q[20]$_DFFE_PN0P_  (.D(_02291_),
    .RN(net265),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .QN(_13998_));
 DFFR_X1 \id_stage_i.imd_val_q[21]$_DFFE_PN0P_  (.D(_02292_),
    .RN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .QN(_13997_));
 DFFR_X1 \id_stage_i.imd_val_q[22]$_DFFE_PN0P_  (.D(_02293_),
    .RN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .QN(_13996_));
 DFFR_X1 \id_stage_i.imd_val_q[23]$_DFFE_PN0P_  (.D(_02294_),
    .RN(net265),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .QN(_13995_));
 DFFR_X1 \id_stage_i.imd_val_q[24]$_DFFE_PN0P_  (.D(_02295_),
    .RN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .QN(_13994_));
 DFFR_X1 \id_stage_i.imd_val_q[25]$_DFFE_PN0P_  (.D(_02296_),
    .RN(net265),
    .CK(clknet_leaf_24_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .QN(_13993_));
 DFFR_X1 \id_stage_i.imd_val_q[26]$_DFFE_PN0P_  (.D(_02297_),
    .RN(net265),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .QN(_13992_));
 DFFR_X1 \id_stage_i.imd_val_q[27]$_DFFE_PN0P_  (.D(_02298_),
    .RN(net265),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .QN(_13991_));
 DFFR_X1 \id_stage_i.imd_val_q[28]$_DFFE_PN0P_  (.D(_02299_),
    .RN(net265),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .QN(_13990_));
 DFFR_X1 \id_stage_i.imd_val_q[29]$_DFFE_PN0P_  (.D(_02300_),
    .RN(net265),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .QN(_13989_));
 DFFR_X1 \id_stage_i.imd_val_q[2]$_DFFE_PN0P_  (.D(_02301_),
    .RN(net265),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .QN(_13988_));
 DFFR_X1 \id_stage_i.imd_val_q[30]$_DFFE_PN0P_  (.D(_02302_),
    .RN(net265),
    .CK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .QN(_13987_));
 DFFR_X1 \id_stage_i.imd_val_q[31]$_DFFE_PN0P_  (.D(_02303_),
    .RN(net246),
    .CK(clknet_leaf_41_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .QN(_13986_));
 DFFR_X2 \id_stage_i.imd_val_q[34]$_DFFE_PN0P_  (.D(_02304_),
    .RN(net246),
    .CK(clknet_leaf_40_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .QN(_00217_));
 DFFR_X2 \id_stage_i.imd_val_q[35]$_DFFE_PN0P_  (.D(_02305_),
    .RN(net265),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .QN(_00185_));
 DFFR_X2 \id_stage_i.imd_val_q[36]$_DFFE_PN0P_  (.D(_02306_),
    .RN(net246),
    .CK(clknet_leaf_40_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .QN(_00558_));
 DFFR_X2 \id_stage_i.imd_val_q[37]$_DFFE_PN0P_  (.D(_02307_),
    .RN(net247),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .QN(_00559_));
 DFFR_X2 \id_stage_i.imd_val_q[38]$_DFFE_PN0P_  (.D(_02308_),
    .RN(net246),
    .CK(clknet_leaf_40_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .QN(_00560_));
 DFFR_X2 \id_stage_i.imd_val_q[39]$_DFFE_PN0P_  (.D(_02309_),
    .RN(net247),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .QN(_00561_));
 DFFR_X1 \id_stage_i.imd_val_q[3]$_DFFE_PN0P_  (.D(_02310_),
    .RN(net265),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .QN(_13985_));
 DFFR_X2 \id_stage_i.imd_val_q[40]$_DFFE_PN0P_  (.D(_02311_),
    .RN(net247),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .QN(_00562_));
 DFFR_X2 \id_stage_i.imd_val_q[41]$_DFFE_PN0P_  (.D(_02312_),
    .RN(net246),
    .CK(clknet_leaf_40_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .QN(_00563_));
 DFFR_X2 \id_stage_i.imd_val_q[42]$_DFFE_PN0P_  (.D(_02313_),
    .RN(net247),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .QN(_00564_));
 DFFR_X2 \id_stage_i.imd_val_q[43]$_DFFE_PN0P_  (.D(_02314_),
    .RN(net246),
    .CK(clknet_leaf_40_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .QN(_00565_));
 DFFR_X2 \id_stage_i.imd_val_q[44]$_DFFE_PN0P_  (.D(_02315_),
    .RN(net247),
    .CK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .QN(_00566_));
 DFFR_X2 \id_stage_i.imd_val_q[45]$_DFFE_PN0P_  (.D(_02316_),
    .RN(net246),
    .CK(clknet_leaf_40_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .QN(_00567_));
 DFFR_X2 \id_stage_i.imd_val_q[46]$_DFFE_PN0P_  (.D(_02317_),
    .RN(net246),
    .CK(clknet_leaf_40_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .QN(_00568_));
 DFFR_X1 \id_stage_i.imd_val_q[47]$_DFFE_PN0P_  (.D(_02318_),
    .RN(net246),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .QN(_00599_));
 DFFR_X2 \id_stage_i.imd_val_q[48]$_DFFE_PN0P_  (.D(_02319_),
    .RN(net247),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .QN(_00630_));
 DFFR_X2 \id_stage_i.imd_val_q[49]$_DFFE_PN0P_  (.D(_02320_),
    .RN(net247),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .QN(_00661_));
 DFFR_X1 \id_stage_i.imd_val_q[4]$_DFFE_PN0P_  (.D(_02321_),
    .RN(net265),
    .CK(clknet_leaf_21_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .QN(_13984_));
 DFFR_X2 \id_stage_i.imd_val_q[50]$_DFFE_PN0P_  (.D(_02322_),
    .RN(net247),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .QN(_00692_));
 DFFR_X2 \id_stage_i.imd_val_q[51]$_DFFE_PN0P_  (.D(_02323_),
    .RN(net247),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .QN(_00723_));
 DFFR_X2 \id_stage_i.imd_val_q[52]$_DFFE_PN0P_  (.D(_02324_),
    .RN(net247),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .QN(_00754_));
 DFFR_X2 \id_stage_i.imd_val_q[53]$_DFFE_PN0P_  (.D(_02325_),
    .RN(net247),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .QN(_00785_));
 DFFR_X2 \id_stage_i.imd_val_q[54]$_DFFE_PN0P_  (.D(_02326_),
    .RN(net247),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .QN(_00816_));
 DFFR_X2 \id_stage_i.imd_val_q[55]$_DFFE_PN0P_  (.D(_02327_),
    .RN(net247),
    .CK(clknet_leaf_33_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .QN(_00847_));
 DFFR_X2 \id_stage_i.imd_val_q[56]$_DFFE_PN0P_  (.D(_02328_),
    .RN(net247),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .QN(_00878_));
 DFFR_X2 \id_stage_i.imd_val_q[57]$_DFFE_PN0P_  (.D(_02329_),
    .RN(net247),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .QN(_00909_));
 DFFR_X2 \id_stage_i.imd_val_q[58]$_DFFE_PN0P_  (.D(_02330_),
    .RN(net265),
    .CK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .QN(_00940_));
 DFFR_X2 \id_stage_i.imd_val_q[59]$_DFFE_PN0P_  (.D(_02331_),
    .RN(net247),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .QN(_00971_));
 DFFR_X1 \id_stage_i.imd_val_q[5]$_DFFE_PN0P_  (.D(_02332_),
    .RN(net247),
    .CK(clknet_leaf_21_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .QN(_13983_));
 DFFR_X2 \id_stage_i.imd_val_q[60]$_DFFE_PN0P_  (.D(_02333_),
    .RN(net247),
    .CK(clknet_leaf_29_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .QN(_01002_));
 DFFR_X2 \id_stage_i.imd_val_q[61]$_DFFE_PN0P_  (.D(_02334_),
    .RN(net247),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .QN(_01033_));
 DFFR_X2 \id_stage_i.imd_val_q[62]$_DFFE_PN0P_  (.D(_02335_),
    .RN(net247),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .QN(_01064_));
 DFFR_X2 \id_stage_i.imd_val_q[63]$_DFFE_PN0P_  (.D(_02336_),
    .RN(net265),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .QN(_01095_));
 DFFR_X2 \id_stage_i.imd_val_q[64]$_DFFE_PN0P_  (.D(_02337_),
    .RN(net265),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .QN(_01126_));
 DFFR_X1 \id_stage_i.imd_val_q[65]$_DFFE_PN0P_  (.D(_02338_),
    .RN(net247),
    .CK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .QN(_01157_));
 DFFR_X1 \id_stage_i.imd_val_q[66]$_DFFE_PN0P_  (.D(_02339_),
    .RN(net265),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .QN(_13982_));
 DFFR_X1 \id_stage_i.imd_val_q[67]$_DFFE_PN0P_  (.D(_02340_),
    .RN(net265),
    .CK(clknet_leaf_23_clk),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .QN(_00132_));
 DFFR_X1 \id_stage_i.imd_val_q[6]$_DFFE_PN0P_  (.D(_02341_),
    .RN(net265),
    .CK(clknet_leaf_27_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .QN(_13981_));
 DFFR_X1 \id_stage_i.imd_val_q[7]$_DFFE_PN0P_  (.D(_02342_),
    .RN(net247),
    .CK(clknet_leaf_53_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .QN(_13980_));
 DFFR_X1 \id_stage_i.imd_val_q[8]$_DFFE_PN0P_  (.D(_02343_),
    .RN(net265),
    .CK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .QN(_13979_));
 DFFR_X1 \id_stage_i.imd_val_q[9]$_DFFE_PN0P_  (.D(_02344_),
    .RN(net265),
    .CK(clknet_leaf_21_clk),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .QN(_14457_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .RN(net254),
    .CK(clknet_leaf_120_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .QN(_14458_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .RN(net254),
    .CK(clknet_leaf_120_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .QN(_14459_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .RN(net254),
    .CK(clknet_leaf_120_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .QN(_13978_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.D(_02345_),
    .CK(clknet_leaf_68_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .QN(_13977_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.D(_02346_),
    .CK(clknet_leaf_71_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .QN(_13976_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.D(_02347_),
    .CK(clknet_leaf_68_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .QN(_13975_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.D(_02348_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .QN(_13974_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.D(_02349_),
    .CK(clknet_leaf_69_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .QN(_13973_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.D(_02350_),
    .CK(clknet_leaf_69_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .QN(_13972_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.D(_02351_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .QN(_13971_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.D(_02352_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .QN(_13970_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.D(_02353_),
    .CK(clknet_leaf_47_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .QN(_13969_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.D(_02354_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .QN(_13968_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.D(_02355_),
    .CK(clknet_leaf_45_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .QN(_13967_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.D(_02356_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .QN(_13966_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.D(_02357_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .QN(_13965_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.D(_02358_),
    .CK(clknet_leaf_45_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .QN(_13964_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.D(_02359_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .QN(_13963_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.D(_02360_),
    .CK(clknet_leaf_47_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .QN(_13962_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.D(_02361_),
    .CK(clknet_leaf_48_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .QN(_13961_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.D(_02362_),
    .CK(clknet_leaf_48_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .QN(_13960_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.D(_02363_),
    .CK(clknet_leaf_48_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .QN(_13959_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.D(_02364_),
    .CK(clknet_leaf_47_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .QN(_13958_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.D(_02365_),
    .CK(clknet_leaf_72_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .QN(_13957_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.D(_02366_),
    .CK(clknet_leaf_48_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .QN(_13956_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.D(_02367_),
    .CK(clknet_leaf_48_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .QN(_13955_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.D(_02368_),
    .CK(clknet_leaf_73_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .QN(_13954_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.D(_02369_),
    .CK(clknet_leaf_73_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .QN(_13953_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.D(_02370_),
    .CK(clknet_leaf_72_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .QN(_13952_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.D(_02371_),
    .CK(clknet_leaf_72_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .QN(_13951_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.D(_02372_),
    .CK(clknet_leaf_71_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .QN(_13950_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.D(_02373_),
    .CK(clknet_leaf_72_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .QN(_13949_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.D(_02374_),
    .CK(clknet_leaf_71_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .QN(_13948_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.D(_02375_),
    .CK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .QN(_13947_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.D(_02376_),
    .CK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .QN(_13946_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.D(_02377_),
    .CK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .QN(_13945_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.D(_02378_),
    .CK(clknet_leaf_119_clk),
    .Q(\cs_registers_i.pc_if_i[1] ),
    .QN(_00137_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.D(_02379_),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.pc_if_i[11] ),
    .QN(_13944_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.D(_02380_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_if_i[12] ),
    .QN(_13943_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.D(_02381_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_if_i[13] ),
    .QN(_13942_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.D(_02382_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_if_i[14] ),
    .QN(_13941_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.D(_02383_),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.pc_if_i[15] ),
    .QN(_13940_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.D(_02384_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_if_i[16] ),
    .QN(_13939_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.D(_02385_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[17] ),
    .QN(_13938_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.D(_02386_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_if_i[18] ),
    .QN(_13937_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.D(_02387_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_if_i[19] ),
    .QN(_13936_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.D(_02388_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_if_i[20] ),
    .QN(_13935_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.D(_02389_),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.pc_if_i[2] ),
    .QN(_15754_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.D(_02390_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[21] ),
    .QN(_13934_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.D(_02391_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[22] ),
    .QN(_13933_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.D(_02392_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_if_i[23] ),
    .QN(_13932_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.D(_02393_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[24] ),
    .QN(_13931_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.D(_02394_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[25] ),
    .QN(_13930_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.D(_02395_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[26] ),
    .QN(_13929_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.D(_02396_),
    .CK(clknet_leaf_49_clk),
    .Q(\cs_registers_i.pc_if_i[27] ),
    .QN(_13928_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.D(_02397_),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.pc_if_i[28] ),
    .QN(_13927_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.D(_02398_),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.pc_if_i[29] ),
    .QN(_13926_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.D(_02399_),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.pc_if_i[30] ),
    .QN(_13925_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.D(_02400_),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.pc_if_i[3] ),
    .QN(_13924_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.D(_02401_),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.pc_if_i[31] ),
    .QN(_13923_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.D(_02402_),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.pc_if_i[4] ),
    .QN(_13922_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.D(_02403_),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.pc_if_i[5] ),
    .QN(_13921_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.D(_02404_),
    .CK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.pc_if_i[6] ),
    .QN(_13920_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.D(_02405_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_if_i[7] ),
    .QN(_13919_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.D(_02406_),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.pc_if_i[8] ),
    .QN(_13918_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.D(_02407_),
    .CK(clknet_leaf_68_clk),
    .Q(\cs_registers_i.pc_if_i[9] ),
    .QN(_13917_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.D(_02408_),
    .CK(clknet_leaf_69_clk),
    .Q(\cs_registers_i.pc_if_i[10] ),
    .QN(_13916_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.D(_02409_),
    .CK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .QN(_13915_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.D(_02410_),
    .CK(clknet_leaf_142_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .QN(_13914_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.D(_02411_),
    .CK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .QN(_13913_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.D(_02412_),
    .CK(clknet_leaf_141_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .QN(_13912_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.D(_02413_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .QN(_13911_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.D(_02414_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .QN(_13910_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.D(_02415_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .QN(_13909_));
 DFF_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.D(_02416_),
    .CK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .QN(_13908_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.D(_02417_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .QN(_13907_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.D(_02418_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .QN(_13906_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.D(_02419_),
    .CK(clknet_leaf_4_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .QN(_13905_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.D(_02420_),
    .CK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .QN(_13904_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.D(_02421_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .QN(_13903_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.D(_02422_),
    .CK(clknet_leaf_5_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .QN(_13902_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.D(_02423_),
    .CK(clknet_leaf_141_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .QN(_13901_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.D(_02424_),
    .CK(clknet_leaf_5_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .QN(_13900_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.D(_02425_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .QN(_13899_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.D(_02426_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .QN(_13898_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.D(_02427_),
    .CK(clknet_leaf_142_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .QN(_13897_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.D(_02428_),
    .CK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .QN(_13896_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.D(_02429_),
    .CK(clknet_leaf_142_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .QN(_13895_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.D(_02430_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .QN(_13894_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.D(_02431_),
    .CK(clknet_leaf_5_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .QN(_13893_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.D(_02432_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .QN(_13892_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.D(_02433_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .QN(_13891_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.D(_02434_),
    .CK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .QN(_13890_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.D(_02435_),
    .CK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .QN(_13889_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.D(_02436_),
    .CK(clknet_leaf_5_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .QN(_13888_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.D(_02437_),
    .CK(clknet_leaf_4_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .QN(_13887_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.D(_02438_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .QN(_13886_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.D(_02439_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .QN(_13885_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.D(_02440_),
    .CK(clknet_leaf_7_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .QN(_13884_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.D(_02441_),
    .CK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .QN(_13883_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.D(_02442_),
    .CK(clknet_leaf_4_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .QN(_13882_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.D(_02443_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .QN(_13881_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.D(_02444_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .QN(_13880_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.D(_02445_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .QN(_13879_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.D(_02446_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .QN(_13878_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.D(_02447_),
    .CK(clknet_leaf_142_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .QN(_13877_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.D(_02448_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .QN(_13876_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.D(_02449_),
    .CK(clknet_leaf_137_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .QN(_13875_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.D(_02450_),
    .CK(clknet_leaf_137_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .QN(_13874_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.D(_02451_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .QN(_13873_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.D(_02452_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .QN(_13872_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.D(_02453_),
    .CK(clknet_leaf_7_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .QN(_13871_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.D(_02454_),
    .CK(clknet_leaf_139_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .QN(_13870_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.D(_02455_),
    .CK(clknet_leaf_5_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .QN(_13869_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.D(_02456_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .QN(_13868_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.D(_02457_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .QN(_13867_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.D(_02458_),
    .CK(clknet_leaf_141_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .QN(_13866_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.D(_02459_),
    .CK(clknet_leaf_141_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .QN(_13865_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.D(_02460_),
    .CK(clknet_leaf_139_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .QN(_13864_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.D(_02461_),
    .CK(clknet_leaf_142_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .QN(_13863_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.D(_02462_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .QN(_13862_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.D(_02463_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .QN(_13861_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.D(_02464_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .QN(_13860_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.D(_02465_),
    .CK(clknet_leaf_142_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .QN(_13859_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.D(_02466_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .QN(_13858_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.D(_02467_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .QN(_13857_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.D(_02468_),
    .CK(clknet_leaf_121_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .QN(_13856_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.D(_02469_),
    .CK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .QN(_13855_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.D(_02470_),
    .CK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .QN(_13854_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.D(_02471_),
    .CK(clknet_leaf_5_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .QN(_13853_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.D(_02472_),
    .CK(clknet_leaf_5_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .QN(_13852_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.D(_02473_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .QN(_13851_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.D(_02474_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .QN(_13850_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.D(_02475_),
    .CK(clknet_leaf_4_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .QN(_13849_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.D(_02476_),
    .CK(clknet_leaf_7_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .QN(_13848_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.D(_02477_),
    .CK(clknet_leaf_4_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .QN(_13847_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.D(_02478_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .QN(_13846_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.D(_02479_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .QN(_13845_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.D(_02480_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .QN(_13844_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.D(_02481_),
    .CK(clknet_leaf_137_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .QN(_13843_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.D(_02482_),
    .CK(clknet_leaf_139_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .QN(_13842_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.D(_02483_),
    .CK(clknet_leaf_137_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .QN(_13841_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.D(_02484_),
    .CK(clknet_leaf_137_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .QN(_13840_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.D(_02485_),
    .CK(clknet_leaf_137_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .QN(_13839_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.D(_02486_),
    .CK(clknet_leaf_4_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .QN(_13838_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.D(_02487_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .QN(_13837_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.D(_02488_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .QN(_13836_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.D(_02489_),
    .CK(clknet_leaf_139_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .QN(_13835_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.D(_02490_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .QN(_13834_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.D(_02491_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .QN(_13833_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.D(_02492_),
    .CK(clknet_leaf_140_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .QN(_13832_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.D(_02493_),
    .CK(clknet_leaf_141_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .QN(_13831_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.D(_02494_),
    .CK(clknet_leaf_139_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .QN(_13830_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.D(_02495_),
    .CK(clknet_leaf_139_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .QN(_13829_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.D(_02496_),
    .CK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .QN(_13828_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.D(_02497_),
    .CK(clknet_leaf_6_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .QN(_13827_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.D(_02498_),
    .CK(clknet_leaf_142_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .QN(_13826_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.D(_02499_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .QN(_13825_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.D(_02500_),
    .CK(clknet_leaf_141_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .QN(_13824_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.D(_02501_),
    .CK(clknet_leaf_135_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .QN(_13823_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.D(_02502_),
    .CK(clknet_leaf_136_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .QN(_13822_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.D(_02503_),
    .CK(clknet_leaf_121_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .QN(_13821_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.D(_02504_),
    .CK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .QN(_14460_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .RN(net630),
    .CK(clknet_leaf_122_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .QN(_00136_));
 DFFR_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .RN(net630),
    .CK(clknet_leaf_121_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .QN(_00135_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .RN(net630),
    .CK(clknet_leaf_121_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .QN(_14461_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .RN(net254),
    .CK(clknet_leaf_120_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .QN(_14462_));
 DFFR_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .RN(net254),
    .CK(clknet_leaf_120_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .QN(_00134_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.D(_02505_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .QN(_13820_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.D(_02506_),
    .CK(clknet_leaf_71_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .QN(_13819_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.D(_02507_),
    .CK(clknet_leaf_71_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .QN(_13818_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.D(_02508_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .QN(_13817_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.D(_02509_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .QN(_13816_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.D(_02510_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .QN(_13815_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.D(_02511_),
    .CK(clknet_leaf_47_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .QN(_13814_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.D(_02512_),
    .CK(clknet_leaf_47_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .QN(_13813_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.D(_02513_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .QN(_13812_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.D(_02514_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .QN(_13811_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.D(_02515_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .QN(_13810_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.D(_02516_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .QN(_13809_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.D(_02517_),
    .CK(clknet_leaf_45_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .QN(_13808_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.D(_02518_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .QN(_13807_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.D(_02519_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .QN(_13806_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.D(_02520_),
    .CK(clknet_leaf_46_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .QN(_13805_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.D(_02521_),
    .CK(clknet_leaf_47_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .QN(_13804_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.D(_02522_),
    .CK(clknet_leaf_48_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .QN(_13803_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.D(_02523_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .QN(_13802_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.D(_02524_),
    .CK(clknet_leaf_44_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .QN(_13801_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.D(_02525_),
    .CK(clknet_leaf_74_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .QN(_13800_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.D(_02526_),
    .CK(clknet_leaf_47_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .QN(_13799_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.D(_02527_),
    .CK(clknet_leaf_48_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .QN(_13798_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.D(_02528_),
    .CK(clknet_leaf_74_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .QN(_13797_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.D(_02529_),
    .CK(clknet_leaf_74_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .QN(_13796_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.D(_02530_),
    .CK(clknet_leaf_71_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .QN(_13795_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.D(_02531_),
    .CK(clknet_leaf_74_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .QN(_13794_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.D(_02532_),
    .CK(clknet_leaf_74_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .QN(_13793_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.D(_02533_),
    .CK(clknet_leaf_70_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .QN(_13792_));
 DFF_X1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.D(_02534_),
    .CK(clknet_leaf_71_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .QN(_14463_));
 DFFR_X2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .RN(net254),
    .CK(clknet_leaf_119_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .QN(_00133_));
 DFF_X1 \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.D(_02535_),
    .CK(clknet_leaf_10_clk),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .QN(_13791_));
 DFF_X1 \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.D(_02536_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ),
    .QN(_13790_));
 DFF_X1 \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.D(_02537_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .QN(_13789_));
 DFF_X1 \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.D(_02538_),
    .CK(clknet_leaf_11_clk),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ),
    .QN(_00278_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[0]$_DFFE_PN_  (.D(_02539_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_i[0] ),
    .QN(_13788_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[10]$_DFFE_PN_  (.D(_02540_),
    .CK(clknet_leaf_10_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .QN(_00036_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[11]$_DFFE_PN_  (.D(_02541_),
    .CK(clknet_leaf_14_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .QN(_00039_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[12]$_DFFE_PN_  (.D(_02542_),
    .CK(clknet_leaf_14_clk),
    .Q(\id_stage_i.controller_i.instr_i[12] ),
    .QN(_00176_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[13]$_DFFE_PN_  (.D(_02543_),
    .CK(clknet_leaf_13_clk),
    .Q(\id_stage_i.controller_i.instr_i[13] ),
    .QN(_00175_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[14]$_DFFE_PN_  (.D(_02544_),
    .CK(clknet_leaf_13_clk),
    .Q(\id_stage_i.controller_i.instr_i[14] ),
    .QN(_00173_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[15]$_DFFE_PN_  (.D(_02545_),
    .CK(clknet_leaf_10_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .QN(_00184_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[16]$_DFFE_PN_  (.D(_02546_),
    .CK(clknet_leaf_14_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .QN(_00183_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[17]$_DFFE_PN_  (.D(_02547_),
    .CK(clknet_leaf_14_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .QN(_00182_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[18]$_DFFE_PN_  (.D(_02548_),
    .CK(clknet_leaf_14_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .QN(_00181_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[19]$_DFFE_PN_  (.D(_02549_),
    .CK(clknet_leaf_15_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .QN(_00180_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[1]$_DFFE_PN_  (.D(_02550_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_i[1] ),
    .QN(_00013_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[20]$_DFFE_PN_  (.D(_02551_),
    .CK(clknet_leaf_15_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .QN(_00140_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[21]$_DFFE_PN_  (.D(_02552_),
    .CK(clknet_leaf_8_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .QN(_13787_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[22]$_DFFE_PN_  (.D(_02553_),
    .CK(clknet_leaf_14_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .QN(_13786_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[23]$_DFFE_PN_  (.D(_02554_),
    .CK(clknet_leaf_15_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .QN(_00139_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[24]$_DFFE_PN_  (.D(_02555_),
    .CK(clknet_leaf_14_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .QN(_00138_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[25]$_DFFE_PN_  (.D(_02556_),
    .CK(clknet_leaf_10_clk),
    .Q(\id_stage_i.controller_i.instr_i[25] ),
    .QN(_13785_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[26]$_DFFE_PN_  (.D(_02557_),
    .CK(clknet_leaf_13_clk),
    .Q(\id_stage_i.controller_i.instr_i[26] ),
    .QN(_00177_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[27]$_DFFE_PN_  (.D(_02558_),
    .CK(clknet_leaf_10_clk),
    .Q(\id_stage_i.controller_i.instr_i[27] ),
    .QN(_13784_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[28]$_DFFE_PN_  (.D(_02559_),
    .CK(clknet_leaf_118_clk),
    .Q(\id_stage_i.controller_i.instr_i[28] ),
    .QN(_13783_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[29]$_DFFE_PN_  (.D(_02560_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_i[29] ),
    .QN(_13782_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[2]$_DFFE_PN_  (.D(_02561_),
    .CK(clknet_leaf_11_clk),
    .Q(\id_stage_i.controller_i.instr_i[2] ),
    .QN(_00015_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[30]$_DFFE_PN_  (.D(_02562_),
    .CK(clknet_leaf_13_clk),
    .Q(\id_stage_i.controller_i.instr_i[30] ),
    .QN(_13781_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[31]$_DFFE_PN_  (.D(_02563_),
    .CK(clknet_leaf_13_clk),
    .Q(\id_stage_i.controller_i.instr_i[31] ),
    .QN(_00174_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[3]$_DFFE_PN_  (.D(_02564_),
    .CK(clknet_leaf_11_clk),
    .Q(\id_stage_i.controller_i.instr_i[3] ),
    .QN(_00017_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[4]$_DFFE_PN_  (.D(_02565_),
    .CK(clknet_leaf_12_clk),
    .Q(\id_stage_i.controller_i.instr_i[4] ),
    .QN(_00020_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[5]$_DFFE_PN_  (.D(_02566_),
    .CK(clknet_leaf_12_clk),
    .Q(\id_stage_i.controller_i.instr_i[5] ),
    .QN(_00023_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[6]$_DFFE_PN_  (.D(_02567_),
    .CK(clknet_leaf_12_clk),
    .Q(\id_stage_i.controller_i.instr_i[6] ),
    .QN(_00172_));
 DFF_X2 \if_stage_i.instr_rdata_alu_id_o[7]$_DFFE_PN_  (.D(_02568_),
    .CK(clknet_leaf_11_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .QN(_00216_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[8]$_DFFE_PN_  (.D(_02569_),
    .CK(clknet_leaf_10_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .QN(_00030_));
 DFF_X1 \if_stage_i.instr_rdata_alu_id_o[9]$_DFFE_PN_  (.D(_02570_),
    .CK(clknet_leaf_9_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .QN(_00033_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.D(_02571_),
    .CK(clknet_leaf_11_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .QN(_13780_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.D(_02572_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .QN(_00037_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.D(_02573_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .QN(_00040_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.D(_02574_),
    .CK(clknet_leaf_11_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .QN(_00042_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.D(_02575_),
    .CK(clknet_leaf_12_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .QN(_00044_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.D(_02576_),
    .CK(clknet_leaf_119_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .QN(_00046_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.D(_02577_),
    .CK(clknet_leaf_119_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .QN(_00048_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.D(_02578_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .QN(_00014_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.D(_02579_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .QN(_00016_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.D(_02580_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .QN(_00018_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.D(_02581_),
    .CK(clknet_leaf_119_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .QN(_00021_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.D(_02582_),
    .CK(clknet_leaf_118_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .QN(_00024_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.D(_02583_),
    .CK(clknet_leaf_119_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .QN(_00026_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.D(_02584_),
    .CK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .QN(_00028_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.D(_02585_),
    .CK(clknet_leaf_10_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .QN(_00031_));
 DFF_X1 \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.D(_02586_),
    .CK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .QN(_00034_));
 DFFR_X2 \if_stage_i.instr_valid_id_q$_DFF_PN0_  (.D(\if_stage_i.instr_valid_id_d ),
    .RN(net248),
    .CK(clknet_leaf_118_clk),
    .Q(\id_stage_i.controller_i.instr_valid_i ),
    .QN(_01161_));
 DFF_X1 \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.D(_02587_),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.pc_id_i[10] ),
    .QN(_00038_));
 DFF_X1 \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.D(_02588_),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.pc_id_i[11] ),
    .QN(_00041_));
 DFF_X1 \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.D(_02589_),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.pc_id_i[12] ),
    .QN(_00043_));
 DFF_X1 \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.D(_02590_),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.pc_id_i[13] ),
    .QN(_00045_));
 DFF_X1 \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.D(_02591_),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.pc_id_i[14] ),
    .QN(_00047_));
 DFF_X1 \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.D(_02592_),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.pc_id_i[15] ),
    .QN(_00049_));
 DFF_X1 \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.D(_02593_),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.pc_id_i[16] ),
    .QN(_00050_));
 DFF_X1 \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.D(_02594_),
    .CK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.pc_id_i[17] ),
    .QN(_00051_));
 DFF_X1 \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.D(_02595_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[18] ),
    .QN(_00052_));
 DFF_X2 \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.D(_02596_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[19] ),
    .QN(_00053_));
 DFF_X1 \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.D(_02597_),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.pc_id_i[1] ),
    .QN(_13779_));
 DFF_X1 \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.D(_02598_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[20] ),
    .QN(_00054_));
 DFF_X1 \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.D(_02599_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[21] ),
    .QN(_00055_));
 DFF_X1 \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.D(_02600_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[22] ),
    .QN(_00056_));
 DFF_X1 \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.D(_02601_),
    .CK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.pc_id_i[23] ),
    .QN(_00057_));
 DFF_X2 \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.D(_02602_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[24] ),
    .QN(_00058_));
 DFF_X1 \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.D(_02603_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[25] ),
    .QN(_00059_));
 DFF_X1 \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.D(_02604_),
    .CK(clknet_leaf_51_clk),
    .Q(\cs_registers_i.pc_id_i[26] ),
    .QN(_00060_));
 DFF_X1 \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.D(_02605_),
    .CK(clknet_leaf_50_clk),
    .Q(\cs_registers_i.pc_id_i[27] ),
    .QN(_00061_));
 DFF_X1 \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.D(_02606_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_id_i[28] ),
    .QN(_00062_));
 DFF_X1 \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.D(_02607_),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.pc_id_i[29] ),
    .QN(_00063_));
 DFF_X2 \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.D(_02608_),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.pc_id_i[2] ),
    .QN(_00012_));
 DFF_X2 \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.D(_02609_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_id_i[30] ),
    .QN(_00064_));
 DFF_X1 \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.D(_02610_),
    .CK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.pc_id_i[31] ),
    .QN(_00065_));
 DFF_X1 \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.D(_02611_),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.pc_id_i[3] ),
    .QN(_00019_));
 DFF_X1 \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.D(_02612_),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.pc_id_i[4] ),
    .QN(_00022_));
 DFF_X1 \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.D(_02613_),
    .CK(clknet_leaf_65_clk),
    .Q(\cs_registers_i.pc_id_i[5] ),
    .QN(_00025_));
 DFF_X1 \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.D(_02614_),
    .CK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.pc_id_i[6] ),
    .QN(_00027_));
 DFF_X1 \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.D(_02615_),
    .CK(clknet_leaf_59_clk),
    .Q(\cs_registers_i.pc_id_i[7] ),
    .QN(_00029_));
 DFF_X1 \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.D(_02616_),
    .CK(clknet_leaf_67_clk),
    .Q(\cs_registers_i.pc_id_i[8] ),
    .QN(_00032_));
 DFF_X1 \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.D(_02617_),
    .CK(clknet_leaf_57_clk),
    .Q(\cs_registers_i.pc_id_i[9] ),
    .QN(_00035_));
 DFFR_X1 \load_store_unit_i.addr_last_q[0]$_DFFE_PN0P_  (.D(_02618_),
    .RN(net248),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .QN(_13778_));
 DFFR_X1 \load_store_unit_i.addr_last_q[10]$_DFFE_PN0P_  (.D(_02619_),
    .RN(net247),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .QN(_13777_));
 DFFR_X1 \load_store_unit_i.addr_last_q[11]$_DFFE_PN0P_  (.D(_02620_),
    .RN(net247),
    .CK(clknet_leaf_55_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .QN(_13776_));
 DFFR_X1 \load_store_unit_i.addr_last_q[12]$_DFFE_PN0P_  (.D(_02621_),
    .RN(net247),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .QN(_13775_));
 DFFR_X1 \load_store_unit_i.addr_last_q[13]$_DFFE_PN0P_  (.D(_02622_),
    .RN(net247),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .QN(_13774_));
 DFFR_X1 \load_store_unit_i.addr_last_q[14]$_DFFE_PN0P_  (.D(_02623_),
    .RN(net247),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .QN(_13773_));
 DFFR_X1 \load_store_unit_i.addr_last_q[15]$_DFFE_PN0P_  (.D(_02624_),
    .RN(net247),
    .CK(clknet_leaf_55_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .QN(_13772_));
 DFFR_X1 \load_store_unit_i.addr_last_q[16]$_DFFE_PN0P_  (.D(_02625_),
    .RN(net247),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .QN(_13771_));
 DFFR_X1 \load_store_unit_i.addr_last_q[17]$_DFFE_PN0P_  (.D(_02626_),
    .RN(net247),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .QN(_13770_));
 DFFR_X1 \load_store_unit_i.addr_last_q[18]$_DFFE_PN0P_  (.D(_02627_),
    .RN(net247),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .QN(_13769_));
 DFFR_X1 \load_store_unit_i.addr_last_q[19]$_DFFE_PN0P_  (.D(_02628_),
    .RN(net247),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .QN(_13768_));
 DFFR_X2 \load_store_unit_i.addr_last_q[1]$_DFFE_PN0P_  (.D(_02629_),
    .RN(net247),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .QN(_13767_));
 DFFR_X1 \load_store_unit_i.addr_last_q[20]$_DFFE_PN0P_  (.D(_02630_),
    .RN(net247),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .QN(_13766_));
 DFFR_X1 \load_store_unit_i.addr_last_q[21]$_DFFE_PN0P_  (.D(_02631_),
    .RN(net247),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .QN(_13765_));
 DFFR_X1 \load_store_unit_i.addr_last_q[22]$_DFFE_PN0P_  (.D(_02632_),
    .RN(net247),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .QN(_13764_));
 DFFR_X1 \load_store_unit_i.addr_last_q[23]$_DFFE_PN0P_  (.D(_02633_),
    .RN(net247),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .QN(_13763_));
 DFFR_X1 \load_store_unit_i.addr_last_q[24]$_DFFE_PN0P_  (.D(_02634_),
    .RN(net247),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .QN(_13762_));
 DFFR_X1 \load_store_unit_i.addr_last_q[25]$_DFFE_PN0P_  (.D(_02635_),
    .RN(net247),
    .CK(clknet_leaf_54_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .QN(_13761_));
 DFFR_X1 \load_store_unit_i.addr_last_q[26]$_DFFE_PN0P_  (.D(_02636_),
    .RN(net247),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .QN(_13760_));
 DFFR_X1 \load_store_unit_i.addr_last_q[27]$_DFFE_PN0P_  (.D(_02637_),
    .RN(net247),
    .CK(clknet_leaf_52_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .QN(_13759_));
 DFFR_X1 \load_store_unit_i.addr_last_q[28]$_DFFE_PN0P_  (.D(_02638_),
    .RN(net247),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .QN(_13758_));
 DFFR_X1 \load_store_unit_i.addr_last_q[29]$_DFFE_PN0P_  (.D(_02639_),
    .RN(net247),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .QN(_13757_));
 DFFR_X1 \load_store_unit_i.addr_last_q[2]$_DFFE_PN0P_  (.D(_02640_),
    .RN(net248),
    .CK(clknet_leaf_55_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .QN(_13756_));
 DFFR_X1 \load_store_unit_i.addr_last_q[30]$_DFFE_PN0P_  (.D(_02641_),
    .RN(net247),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .QN(_13755_));
 DFFR_X2 \load_store_unit_i.addr_last_q[31]$_DFFE_PN0P_  (.D(_02642_),
    .RN(net247),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .QN(_13754_));
 DFFR_X1 \load_store_unit_i.addr_last_q[3]$_DFFE_PN0P_  (.D(_02643_),
    .RN(net248),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .QN(_13753_));
 DFFR_X1 \load_store_unit_i.addr_last_q[4]$_DFFE_PN0P_  (.D(_02644_),
    .RN(net247),
    .CK(clknet_leaf_66_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .QN(_13752_));
 DFFR_X1 \load_store_unit_i.addr_last_q[5]$_DFFE_PN0P_  (.D(_02645_),
    .RN(net247),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .QN(_13751_));
 DFFR_X1 \load_store_unit_i.addr_last_q[6]$_DFFE_PN0P_  (.D(_02646_),
    .RN(net247),
    .CK(clknet_leaf_57_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .QN(_13750_));
 DFFR_X1 \load_store_unit_i.addr_last_q[7]$_DFFE_PN0P_  (.D(_02647_),
    .RN(net248),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .QN(_13749_));
 DFFR_X1 \load_store_unit_i.addr_last_q[8]$_DFFE_PN0P_  (.D(_02648_),
    .RN(net247),
    .CK(clknet_leaf_53_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .QN(_13748_));
 DFFR_X1 \load_store_unit_i.addr_last_q[9]$_DFFE_PN0P_  (.D(_02649_),
    .RN(net247),
    .CK(clknet_leaf_56_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .QN(_13747_));
 DFFR_X2 \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.D(_02650_),
    .RN(net265),
    .CK(clknet_leaf_19_clk),
    .Q(\load_store_unit_i.data_sign_ext_q ),
    .QN(_13746_));
 DFFR_X1 \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.D(_02651_),
    .RN(net265),
    .CK(clknet_leaf_20_clk),
    .Q(\load_store_unit_i.data_we_q ),
    .QN(_01159_));
 DFFR_X2 \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.D(_02652_),
    .RN(net265),
    .CK(clknet_leaf_19_clk),
    .Q(\load_store_unit_i.handle_misaligned_q ),
    .QN(_16486_));
 DFFR_X1 \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.D(_02653_),
    .RN(net265),
    .CK(clknet_leaf_19_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[0] ),
    .QN(_13745_));
 DFFR_X1 \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.D(_02654_),
    .RN(net265),
    .CK(clknet_leaf_20_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[1] ),
    .QN(_13744_));
 DFFR_X1 \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.D(_02655_),
    .RN(net265),
    .CK(clknet_leaf_20_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[2] ),
    .QN(_00171_));
 DFFR_X1 \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.D(_02656_),
    .RN(net265),
    .CK(clknet_leaf_20_clk),
    .Q(\load_store_unit_i.lsu_err_q ),
    .QN(_13743_));
 DFFR_X1 \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.D(_02657_),
    .RN(net265),
    .CK(clknet_leaf_18_clk),
    .Q(\load_store_unit_i.rdata_offset_q[0] ),
    .QN(_13742_));
 DFFR_X1 \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.D(_02658_),
    .RN(net265),
    .CK(clknet_leaf_19_clk),
    .Q(\load_store_unit_i.rdata_offset_q[1] ),
    .QN(_13741_));
 DFFR_X1 \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.D(_02659_),
    .RN(net265),
    .CK(clknet_leaf_17_clk),
    .Q(\load_store_unit_i.rdata_q[8] ),
    .QN(_13740_));
 DFFR_X1 \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.D(_02660_),
    .RN(net256),
    .CK(clknet_leaf_22_clk),
    .Q(\load_store_unit_i.rdata_q[18] ),
    .QN(_13739_));
 DFFR_X1 \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.D(_02661_),
    .RN(net265),
    .CK(clknet_leaf_22_clk),
    .Q(\load_store_unit_i.rdata_q[19] ),
    .QN(_13738_));
 DFFR_X1 \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.D(_02662_),
    .RN(net256),
    .CK(clknet_leaf_22_clk),
    .Q(\load_store_unit_i.rdata_q[20] ),
    .QN(_13737_));
 DFFR_X1 \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.D(_02663_),
    .RN(net256),
    .CK(clknet_leaf_16_clk),
    .Q(\load_store_unit_i.rdata_q[21] ),
    .QN(_13736_));
 DFFR_X1 \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.D(_02664_),
    .RN(net256),
    .CK(clknet_leaf_16_clk),
    .Q(\load_store_unit_i.rdata_q[22] ),
    .QN(_13735_));
 DFFR_X1 \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.D(_02665_),
    .RN(net265),
    .CK(clknet_leaf_18_clk),
    .Q(\load_store_unit_i.rdata_q[23] ),
    .QN(_13734_));
 DFFR_X1 \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.D(_02666_),
    .RN(net265),
    .CK(clknet_leaf_17_clk),
    .Q(\load_store_unit_i.rdata_q[24] ),
    .QN(_13733_));
 DFFR_X1 \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.D(_02667_),
    .RN(net265),
    .CK(clknet_leaf_17_clk),
    .Q(\load_store_unit_i.rdata_q[25] ),
    .QN(_13732_));
 DFFR_X1 \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.D(_02668_),
    .RN(net265),
    .CK(clknet_leaf_22_clk),
    .Q(\load_store_unit_i.rdata_q[26] ),
    .QN(_13731_));
 DFFR_X1 \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.D(_02669_),
    .RN(net265),
    .CK(clknet_leaf_22_clk),
    .Q(\load_store_unit_i.rdata_q[27] ),
    .QN(_13730_));
 DFFR_X1 \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.D(_02670_),
    .RN(net265),
    .CK(clknet_leaf_16_clk),
    .Q(\load_store_unit_i.rdata_q[9] ),
    .QN(_13729_));
 DFFR_X1 \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.D(_02671_),
    .RN(net256),
    .CK(clknet_leaf_23_clk),
    .Q(\load_store_unit_i.rdata_q[28] ),
    .QN(_13728_));
 DFFR_X1 \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.D(_02672_),
    .RN(net256),
    .CK(clknet_leaf_17_clk),
    .Q(\load_store_unit_i.rdata_q[29] ),
    .QN(_13727_));
 DFFR_X1 \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.D(_02673_),
    .RN(net256),
    .CK(clknet_leaf_16_clk),
    .Q(\load_store_unit_i.rdata_q[30] ),
    .QN(_13726_));
 DFFR_X1 \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.D(_02674_),
    .RN(net265),
    .CK(clknet_leaf_18_clk),
    .Q(\load_store_unit_i.rdata_q[31] ),
    .QN(_13725_));
 DFFR_X1 \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.D(_02675_),
    .RN(net256),
    .CK(clknet_leaf_22_clk),
    .Q(\load_store_unit_i.rdata_q[10] ),
    .QN(_13724_));
 DFFR_X1 \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.D(_02676_),
    .RN(net265),
    .CK(clknet_leaf_17_clk),
    .Q(\load_store_unit_i.rdata_q[11] ),
    .QN(_13723_));
 DFFR_X1 \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.D(_02677_),
    .RN(net256),
    .CK(clknet_leaf_23_clk),
    .Q(\load_store_unit_i.rdata_q[12] ),
    .QN(_13722_));
 DFFR_X1 \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.D(_02678_),
    .RN(net256),
    .CK(clknet_leaf_16_clk),
    .Q(\load_store_unit_i.rdata_q[13] ),
    .QN(_13721_));
 DFFR_X1 \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.D(_02679_),
    .RN(net256),
    .CK(clknet_leaf_16_clk),
    .Q(\load_store_unit_i.rdata_q[14] ),
    .QN(_13720_));
 DFFR_X1 \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.D(_02680_),
    .RN(net265),
    .CK(clknet_leaf_18_clk),
    .Q(\load_store_unit_i.rdata_q[15] ),
    .QN(_13719_));
 DFFR_X1 \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.D(_02681_),
    .RN(net265),
    .CK(clknet_leaf_18_clk),
    .Q(\load_store_unit_i.rdata_q[16] ),
    .QN(_13718_));
 DFFR_X1 \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.D(_02682_),
    .RN(net256),
    .CK(clknet_leaf_16_clk),
    .Q(\load_store_unit_i.rdata_q[17] ),
    .QN(_13717_));
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_425 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_426 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_427 ();
 CLKBUF_X3 max_cap7 (.A(\alu_adder_result_ex[14] ),
    .Z(net7));
 BUF_X4 max_cap8 (.A(\alu_adder_result_ex[6] ),
    .Z(net8));
 CLKBUF_X3 wire9 (.A(_11923_),
    .Z(net9));
 BUF_X4 wire10 (.A(_11571_),
    .Z(net10));
 BUF_X1 max_cap11 (.A(net13),
    .Z(net11));
 CLKBUF_X3 max_cap12 (.A(_04490_),
    .Z(net12));
 CLKBUF_X2 wire13 (.A(_03568_),
    .Z(net13));
 CLKBUF_X2 wire14 (.A(_03545_),
    .Z(net14));
 BUF_X1 input1 (.A(boot_addr_i[10]),
    .Z(net1));
 BUF_X2 input2 (.A(boot_addr_i[11]),
    .Z(net2));
 BUF_X1 input3 (.A(boot_addr_i[12]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(boot_addr_i[13]),
    .Z(net4));
 BUF_X1 input5 (.A(boot_addr_i[14]),
    .Z(net5));
 BUF_X2 input6 (.A(boot_addr_i[15]),
    .Z(net6));
 BUF_X1 input7 (.A(boot_addr_i[16]),
    .Z(net15));
 BUF_X1 input8 (.A(boot_addr_i[17]),
    .Z(net16));
 BUF_X1 input9 (.A(boot_addr_i[18]),
    .Z(net17));
 BUF_X1 input10 (.A(boot_addr_i[19]),
    .Z(net18));
 BUF_X1 input11 (.A(boot_addr_i[20]),
    .Z(net19));
 BUF_X1 input12 (.A(boot_addr_i[21]),
    .Z(net20));
 BUF_X1 input13 (.A(boot_addr_i[22]),
    .Z(net21));
 BUF_X1 input14 (.A(boot_addr_i[23]),
    .Z(net22));
 BUF_X1 input15 (.A(boot_addr_i[24]),
    .Z(net23));
 BUF_X1 input16 (.A(boot_addr_i[25]),
    .Z(net24));
 CLKBUF_X2 input17 (.A(boot_addr_i[26]),
    .Z(net25));
 BUF_X1 input18 (.A(boot_addr_i[27]),
    .Z(net26));
 BUF_X1 input19 (.A(boot_addr_i[28]),
    .Z(net27));
 BUF_X1 input20 (.A(boot_addr_i[29]),
    .Z(net28));
 BUF_X1 input21 (.A(boot_addr_i[30]),
    .Z(net29));
 BUF_X1 input22 (.A(boot_addr_i[31]),
    .Z(net30));
 BUF_X1 input23 (.A(boot_addr_i[8]),
    .Z(net31));
 CLKBUF_X2 input24 (.A(boot_addr_i[9]),
    .Z(net32));
 CLKBUF_X3 input25 (.A(data_err_i),
    .Z(net33));
 CLKBUF_X2 input26 (.A(data_rdata_i[0]),
    .Z(net34));
 BUF_X2 input27 (.A(data_rdata_i[14]),
    .Z(net35));
 BUF_X2 input28 (.A(data_rdata_i[16]),
    .Z(net36));
 BUF_X2 input29 (.A(data_rdata_i[17]),
    .Z(net37));
 BUF_X2 input30 (.A(data_rdata_i[18]),
    .Z(net38));
 BUF_X2 input31 (.A(data_rdata_i[19]),
    .Z(net39));
 CLKBUF_X2 input32 (.A(data_rdata_i[1]),
    .Z(net40));
 BUF_X2 input33 (.A(data_rdata_i[20]),
    .Z(net41));
 CLKBUF_X2 input34 (.A(data_rdata_i[21]),
    .Z(net42));
 BUF_X1 input35 (.A(data_rdata_i[22]),
    .Z(net43));
 BUF_X2 input36 (.A(data_rdata_i[23]),
    .Z(net44));
 CLKBUF_X2 input37 (.A(data_rdata_i[24]),
    .Z(net45));
 BUF_X2 input38 (.A(data_rdata_i[25]),
    .Z(net46));
 BUF_X2 input39 (.A(data_rdata_i[26]),
    .Z(net47));
 BUF_X2 input40 (.A(data_rdata_i[27]),
    .Z(net48));
 BUF_X2 input41 (.A(data_rdata_i[28]),
    .Z(net49));
 BUF_X2 input42 (.A(data_rdata_i[29]),
    .Z(net50));
 BUF_X2 input43 (.A(data_rdata_i[2]),
    .Z(net51));
 BUF_X2 input44 (.A(data_rdata_i[30]),
    .Z(net52));
 BUF_X2 input45 (.A(data_rdata_i[31]),
    .Z(net53));
 BUF_X2 input46 (.A(data_rdata_i[3]),
    .Z(net54));
 BUF_X2 input47 (.A(data_rdata_i[4]),
    .Z(net55));
 CLKBUF_X2 input48 (.A(data_rdata_i[5]),
    .Z(net56));
 BUF_X1 input49 (.A(data_rdata_i[6]),
    .Z(net57));
 BUF_X2 input50 (.A(data_rdata_i[7]),
    .Z(net58));
 CLKBUF_X3 input51 (.A(data_rvalid_i),
    .Z(net59));
 BUF_X1 input52 (.A(fetch_enable_i),
    .Z(net60));
 BUF_X1 input53 (.A(hart_id_i[0]),
    .Z(net61));
 BUF_X1 input54 (.A(hart_id_i[10]),
    .Z(net62));
 CLKBUF_X2 input55 (.A(hart_id_i[11]),
    .Z(net63));
 BUF_X1 input56 (.A(hart_id_i[12]),
    .Z(net64));
 BUF_X1 input57 (.A(hart_id_i[13]),
    .Z(net65));
 BUF_X1 input58 (.A(hart_id_i[14]),
    .Z(net66));
 BUF_X1 input59 (.A(hart_id_i[15]),
    .Z(net67));
 BUF_X1 input60 (.A(hart_id_i[16]),
    .Z(net68));
 BUF_X1 input61 (.A(hart_id_i[17]),
    .Z(net69));
 BUF_X1 input62 (.A(hart_id_i[18]),
    .Z(net70));
 BUF_X1 input63 (.A(hart_id_i[19]),
    .Z(net71));
 BUF_X1 input64 (.A(hart_id_i[1]),
    .Z(net72));
 BUF_X1 input65 (.A(hart_id_i[20]),
    .Z(net73));
 BUF_X1 input66 (.A(hart_id_i[21]),
    .Z(net74));
 BUF_X1 input67 (.A(hart_id_i[22]),
    .Z(net75));
 BUF_X1 input68 (.A(hart_id_i[23]),
    .Z(net76));
 BUF_X1 input69 (.A(hart_id_i[24]),
    .Z(net77));
 BUF_X1 input70 (.A(hart_id_i[25]),
    .Z(net78));
 BUF_X1 input71 (.A(hart_id_i[26]),
    .Z(net79));
 BUF_X1 input72 (.A(hart_id_i[27]),
    .Z(net80));
 BUF_X1 input73 (.A(hart_id_i[28]),
    .Z(net81));
 BUF_X1 input74 (.A(hart_id_i[29]),
    .Z(net82));
 BUF_X1 input75 (.A(hart_id_i[2]),
    .Z(net83));
 BUF_X1 input76 (.A(hart_id_i[30]),
    .Z(net84));
 CLKBUF_X2 input77 (.A(hart_id_i[31]),
    .Z(net85));
 BUF_X1 input78 (.A(hart_id_i[3]),
    .Z(net86));
 BUF_X1 input79 (.A(hart_id_i[4]),
    .Z(net87));
 BUF_X1 input80 (.A(hart_id_i[5]),
    .Z(net88));
 BUF_X1 input81 (.A(hart_id_i[6]),
    .Z(net89));
 BUF_X1 input82 (.A(hart_id_i[7]),
    .Z(net90));
 BUF_X1 input83 (.A(hart_id_i[8]),
    .Z(net91));
 BUF_X1 input84 (.A(hart_id_i[9]),
    .Z(net92));
 CLKBUF_X3 input85 (.A(instr_gnt_i),
    .Z(net93));
 BUF_X2 input86 (.A(instr_rdata_i[0]),
    .Z(net94));
 CLKBUF_X2 input87 (.A(instr_rdata_i[10]),
    .Z(net95));
 BUF_X1 input88 (.A(instr_rdata_i[11]),
    .Z(net96));
 CLKBUF_X2 input89 (.A(instr_rdata_i[12]),
    .Z(net97));
 BUF_X1 input90 (.A(instr_rdata_i[13]),
    .Z(net98));
 BUF_X1 input91 (.A(instr_rdata_i[14]),
    .Z(net99));
 BUF_X1 input92 (.A(instr_rdata_i[15]),
    .Z(net100));
 BUF_X2 input93 (.A(instr_rdata_i[18]),
    .Z(net101));
 BUF_X2 input94 (.A(instr_rdata_i[19]),
    .Z(net102));
 BUF_X2 input95 (.A(instr_rdata_i[1]),
    .Z(net103));
 BUF_X2 input96 (.A(instr_rdata_i[20]),
    .Z(net104));
 BUF_X2 input97 (.A(instr_rdata_i[21]),
    .Z(net105));
 BUF_X2 input98 (.A(instr_rdata_i[22]),
    .Z(net106));
 BUF_X2 input99 (.A(instr_rdata_i[23]),
    .Z(net107));
 BUF_X2 input100 (.A(instr_rdata_i[24]),
    .Z(net108));
 CLKBUF_X2 input101 (.A(instr_rdata_i[25]),
    .Z(net109));
 BUF_X2 input102 (.A(instr_rdata_i[26]),
    .Z(net110));
 CLKBUF_X2 input103 (.A(instr_rdata_i[27]),
    .Z(net111));
 BUF_X2 input104 (.A(instr_rdata_i[28]),
    .Z(net112));
 CLKBUF_X2 input105 (.A(instr_rdata_i[29]),
    .Z(net113));
 CLKBUF_X2 input106 (.A(instr_rdata_i[2]),
    .Z(net114));
 CLKBUF_X2 input107 (.A(instr_rdata_i[30]),
    .Z(net115));
 CLKBUF_X2 input108 (.A(instr_rdata_i[31]),
    .Z(net116));
 CLKBUF_X2 input109 (.A(instr_rdata_i[3]),
    .Z(net117));
 BUF_X2 input110 (.A(instr_rdata_i[4]),
    .Z(net118));
 CLKBUF_X2 input111 (.A(instr_rdata_i[5]),
    .Z(net119));
 BUF_X2 input112 (.A(instr_rdata_i[6]),
    .Z(net120));
 CLKBUF_X2 input113 (.A(instr_rdata_i[7]),
    .Z(net121));
 CLKBUF_X2 input114 (.A(instr_rdata_i[8]),
    .Z(net122));
 CLKBUF_X2 input115 (.A(instr_rdata_i[9]),
    .Z(net123));
 CLKBUF_X2 input116 (.A(instr_rvalid_i),
    .Z(net124));
 BUF_X2 input117 (.A(irq_external_i),
    .Z(net125));
 CLKBUF_X2 input118 (.A(irq_fast_i[0]),
    .Z(net126));
 BUF_X2 input119 (.A(irq_fast_i[10]),
    .Z(net127));
 BUF_X2 input120 (.A(irq_fast_i[11]),
    .Z(net128));
 BUF_X2 input121 (.A(irq_fast_i[12]),
    .Z(net129));
 BUF_X2 input122 (.A(irq_fast_i[13]),
    .Z(net130));
 CLKBUF_X2 input123 (.A(irq_fast_i[14]),
    .Z(net131));
 CLKBUF_X2 input124 (.A(irq_fast_i[1]),
    .Z(net132));
 BUF_X1 input125 (.A(irq_fast_i[2]),
    .Z(net133));
 BUF_X1 input126 (.A(irq_fast_i[3]),
    .Z(net134));
 BUF_X2 input127 (.A(irq_fast_i[4]),
    .Z(net135));
 BUF_X2 input128 (.A(irq_fast_i[5]),
    .Z(net136));
 BUF_X2 input129 (.A(irq_fast_i[6]),
    .Z(net137));
 CLKBUF_X3 input130 (.A(irq_fast_i[7]),
    .Z(net138));
 BUF_X2 input131 (.A(irq_fast_i[8]),
    .Z(net139));
 BUF_X2 input132 (.A(irq_fast_i[9]),
    .Z(net140));
 BUF_X2 input133 (.A(irq_nm_i),
    .Z(net141));
 CLKBUF_X2 input134 (.A(irq_software_i),
    .Z(net142));
 CLKBUF_X2 input135 (.A(irq_timer_i),
    .Z(net143));
 BUF_X4 input136 (.A(net629),
    .Z(net144));
 BUF_X1 input137 (.A(test_en_i),
    .Z(net145));
 BUF_X1 output138 (.A(net146),
    .Z(core_sleep_o));
 BUF_X1 output139 (.A(net147),
    .Z(data_addr_o[10]));
 BUF_X1 output140 (.A(net148),
    .Z(data_addr_o[11]));
 BUF_X1 output141 (.A(net149),
    .Z(data_addr_o[12]));
 BUF_X1 output142 (.A(net150),
    .Z(data_addr_o[13]));
 BUF_X1 output143 (.A(net151),
    .Z(data_addr_o[14]));
 BUF_X1 output144 (.A(net152),
    .Z(data_addr_o[15]));
 BUF_X1 output145 (.A(net153),
    .Z(data_addr_o[16]));
 BUF_X1 output146 (.A(net154),
    .Z(data_addr_o[17]));
 BUF_X1 output147 (.A(net155),
    .Z(data_addr_o[18]));
 BUF_X1 output148 (.A(net156),
    .Z(data_addr_o[19]));
 BUF_X1 output149 (.A(net157),
    .Z(data_addr_o[20]));
 BUF_X1 output150 (.A(net158),
    .Z(data_addr_o[21]));
 BUF_X1 output151 (.A(net159),
    .Z(data_addr_o[22]));
 BUF_X1 output152 (.A(net160),
    .Z(data_addr_o[23]));
 BUF_X1 output153 (.A(net161),
    .Z(data_addr_o[24]));
 BUF_X1 output154 (.A(net162),
    .Z(data_addr_o[25]));
 BUF_X1 output155 (.A(net163),
    .Z(data_addr_o[26]));
 BUF_X1 output156 (.A(net164),
    .Z(data_addr_o[27]));
 BUF_X1 output157 (.A(net165),
    .Z(data_addr_o[28]));
 BUF_X1 output158 (.A(net166),
    .Z(data_addr_o[29]));
 BUF_X1 output159 (.A(net167),
    .Z(data_addr_o[2]));
 BUF_X1 output160 (.A(net168),
    .Z(data_addr_o[30]));
 BUF_X1 output161 (.A(net169),
    .Z(data_addr_o[31]));
 BUF_X1 output162 (.A(net170),
    .Z(data_addr_o[3]));
 BUF_X1 output163 (.A(net171),
    .Z(data_addr_o[4]));
 BUF_X1 output164 (.A(net172),
    .Z(data_addr_o[5]));
 BUF_X1 output165 (.A(net173),
    .Z(data_addr_o[6]));
 BUF_X1 output166 (.A(net174),
    .Z(data_addr_o[7]));
 BUF_X1 output167 (.A(net175),
    .Z(data_addr_o[8]));
 BUF_X1 output168 (.A(net176),
    .Z(data_addr_o[9]));
 BUF_X1 output169 (.A(net177),
    .Z(data_be_o[0]));
 BUF_X1 output170 (.A(net178),
    .Z(data_be_o[1]));
 BUF_X1 output171 (.A(net179),
    .Z(data_be_o[2]));
 BUF_X1 output172 (.A(net180),
    .Z(data_be_o[3]));
 BUF_X1 output173 (.A(net181),
    .Z(data_req_o));
 BUF_X1 output174 (.A(net182),
    .Z(data_wdata_o[0]));
 BUF_X1 output175 (.A(net183),
    .Z(data_wdata_o[10]));
 BUF_X1 output176 (.A(net184),
    .Z(data_wdata_o[11]));
 BUF_X1 output177 (.A(net185),
    .Z(data_wdata_o[12]));
 BUF_X1 output178 (.A(net186),
    .Z(data_wdata_o[13]));
 BUF_X1 output179 (.A(net187),
    .Z(data_wdata_o[14]));
 BUF_X1 output180 (.A(net188),
    .Z(data_wdata_o[15]));
 BUF_X1 output181 (.A(net189),
    .Z(data_wdata_o[16]));
 BUF_X1 output182 (.A(net190),
    .Z(data_wdata_o[17]));
 BUF_X1 output183 (.A(net191),
    .Z(data_wdata_o[18]));
 BUF_X1 output184 (.A(net192),
    .Z(data_wdata_o[19]));
 BUF_X1 output185 (.A(net193),
    .Z(data_wdata_o[1]));
 BUF_X1 output186 (.A(net194),
    .Z(data_wdata_o[20]));
 BUF_X1 output187 (.A(net195),
    .Z(data_wdata_o[21]));
 BUF_X1 output188 (.A(net196),
    .Z(data_wdata_o[22]));
 BUF_X1 output189 (.A(net197),
    .Z(data_wdata_o[23]));
 BUF_X1 output190 (.A(net198),
    .Z(data_wdata_o[24]));
 BUF_X1 output191 (.A(net199),
    .Z(data_wdata_o[25]));
 BUF_X1 output192 (.A(net200),
    .Z(data_wdata_o[26]));
 BUF_X1 output193 (.A(net201),
    .Z(data_wdata_o[27]));
 BUF_X1 output194 (.A(net202),
    .Z(data_wdata_o[28]));
 BUF_X1 output195 (.A(net203),
    .Z(data_wdata_o[29]));
 BUF_X1 output196 (.A(net204),
    .Z(data_wdata_o[2]));
 BUF_X1 output197 (.A(net205),
    .Z(data_wdata_o[30]));
 BUF_X1 output198 (.A(net206),
    .Z(data_wdata_o[31]));
 BUF_X1 output199 (.A(net207),
    .Z(data_wdata_o[3]));
 BUF_X1 output200 (.A(net208),
    .Z(data_wdata_o[4]));
 BUF_X1 output201 (.A(net209),
    .Z(data_wdata_o[5]));
 BUF_X1 output202 (.A(net210),
    .Z(data_wdata_o[6]));
 BUF_X1 output203 (.A(net211),
    .Z(data_wdata_o[7]));
 BUF_X1 output204 (.A(net212),
    .Z(data_wdata_o[8]));
 BUF_X1 output205 (.A(net213),
    .Z(data_wdata_o[9]));
 BUF_X1 output206 (.A(net214),
    .Z(data_we_o));
 BUF_X1 output207 (.A(net215),
    .Z(instr_addr_o[10]));
 BUF_X1 output208 (.A(net216),
    .Z(instr_addr_o[11]));
 BUF_X1 output209 (.A(net217),
    .Z(instr_addr_o[12]));
 BUF_X1 output210 (.A(net218),
    .Z(instr_addr_o[13]));
 BUF_X1 output211 (.A(net219),
    .Z(instr_addr_o[14]));
 BUF_X1 output212 (.A(net220),
    .Z(instr_addr_o[15]));
 BUF_X1 output213 (.A(net221),
    .Z(instr_addr_o[16]));
 BUF_X1 output214 (.A(net222),
    .Z(instr_addr_o[17]));
 BUF_X1 output215 (.A(net223),
    .Z(instr_addr_o[18]));
 BUF_X1 output216 (.A(net224),
    .Z(instr_addr_o[19]));
 BUF_X1 output217 (.A(net225),
    .Z(instr_addr_o[20]));
 BUF_X1 output218 (.A(net226),
    .Z(instr_addr_o[21]));
 BUF_X1 output219 (.A(net227),
    .Z(instr_addr_o[22]));
 BUF_X1 output220 (.A(net228),
    .Z(instr_addr_o[23]));
 BUF_X1 output221 (.A(net229),
    .Z(instr_addr_o[24]));
 BUF_X1 output222 (.A(net230),
    .Z(instr_addr_o[25]));
 BUF_X1 output223 (.A(net231),
    .Z(instr_addr_o[26]));
 BUF_X1 output224 (.A(net232),
    .Z(instr_addr_o[27]));
 BUF_X1 output225 (.A(net233),
    .Z(instr_addr_o[28]));
 BUF_X1 output226 (.A(net234),
    .Z(instr_addr_o[29]));
 BUF_X1 output227 (.A(net235),
    .Z(instr_addr_o[2]));
 BUF_X1 output228 (.A(net236),
    .Z(instr_addr_o[30]));
 BUF_X1 output229 (.A(net237),
    .Z(instr_addr_o[31]));
 BUF_X1 output230 (.A(net238),
    .Z(instr_addr_o[3]));
 BUF_X1 output231 (.A(net239),
    .Z(instr_addr_o[4]));
 BUF_X1 output232 (.A(net240),
    .Z(instr_addr_o[5]));
 BUF_X1 output233 (.A(net241),
    .Z(instr_addr_o[6]));
 BUF_X1 output234 (.A(net242),
    .Z(instr_addr_o[7]));
 BUF_X1 output235 (.A(net243),
    .Z(instr_addr_o[8]));
 BUF_X1 output236 (.A(net244),
    .Z(instr_addr_o[9]));
 BUF_X1 output237 (.A(net245),
    .Z(instr_req_o));
 BUF_X4 max_cap238 (.A(net247),
    .Z(net246));
 BUF_X4 max_cap239 (.A(net248),
    .Z(net247));
 BUF_X4 max_cap240 (.A(net254),
    .Z(net248));
 BUF_X4 max_cap241 (.A(net253),
    .Z(net249));
 BUF_X4 max_cap242 (.A(net252),
    .Z(net250));
 BUF_X4 max_cap243 (.A(net252),
    .Z(net251));
 BUF_X4 max_cap244 (.A(net253),
    .Z(net252));
 BUF_X4 max_cap245 (.A(net254),
    .Z(net253));
 BUF_X4 max_cap246 (.A(net144),
    .Z(net254));
 BUF_X4 max_cap247 (.A(net268),
    .Z(net255));
 BUF_X4 wire248 (.A(net257),
    .Z(net256));
 BUF_X4 max_cap249 (.A(net262),
    .Z(net257));
 BUF_X4 max_cap250 (.A(net259),
    .Z(net258));
 BUF_X4 max_cap251 (.A(net260),
    .Z(net259));
 BUF_X4 max_cap252 (.A(net261),
    .Z(net260));
 BUF_X4 max_cap253 (.A(net262),
    .Z(net261));
 BUF_X4 max_cap254 (.A(net268),
    .Z(net262));
 BUF_X4 max_cap255 (.A(net268),
    .Z(net263));
 BUF_X4 max_cap256 (.A(net267),
    .Z(net264));
 BUF_X4 max_cap257 (.A(net266),
    .Z(net265));
 BUF_X4 max_cap258 (.A(net267),
    .Z(net266));
 BUF_X4 max_cap259 (.A(net268),
    .Z(net267));
 BUF_X4 max_cap260 (.A(net144),
    .Z(net268));
 LOGIC0_X1 _30653__261 (.Z(net269));
 LOGIC0_X1 _30654__262 (.Z(net270));
 LOGIC0_X1 _30655__263 (.Z(net271));
 LOGIC0_X1 _30656__264 (.Z(net272));
 LOGIC0_X1 _30687__265 (.Z(net273));
 LOGIC0_X1 _30688__266 (.Z(net274));
 CLKBUF_X3 clkbuf_0_clk_i (.A(clk_i),
    .Z(clknet_0_clk_i));
 CLKBUF_X3 clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_1_0__leaf_clk_i));
 CLKBUF_X3 clkbuf_leaf_0_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_0_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_1_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_1_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_2_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_2_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_3_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_3_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_4_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_4_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_5_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_5_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_6_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_6_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_7_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_7_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_8_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_8_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_9_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_9_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_10_clk_i_regs (.A(clknet_4_0_0_clk_i_regs),
    .Z(clknet_leaf_10_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_11_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_11_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_12_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_12_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_13_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_13_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_14_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_14_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_15_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_15_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_16_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_16_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_17_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_17_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_18_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_18_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_19_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_19_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_20_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_20_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_21_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_21_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_22_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_22_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_23_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_23_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_24_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_24_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_25_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_25_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_26_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_26_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_27_clk_i_regs (.A(clknet_4_3_0_clk_i_regs),
    .Z(clknet_leaf_27_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_28_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_28_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_29_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_29_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_30_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_30_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_31_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_31_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_32_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_32_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_33_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_33_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_34_clk_i_regs (.A(clknet_4_2_0_clk_i_regs),
    .Z(clknet_leaf_34_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_35_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_35_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_36_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_36_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_37_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_37_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_38_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_38_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_39_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_39_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_40_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_40_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_41_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_41_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_42_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_42_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_43_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_43_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_44_clk_i_regs (.A(clknet_4_8_0_clk_i_regs),
    .Z(clknet_leaf_44_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_45_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_45_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_46_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_46_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_47_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_47_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_48_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_48_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_49_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_49_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_50_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_50_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_51_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_51_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_52_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_52_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_53_clk_i_regs (.A(clknet_4_10_0_clk_i_regs),
    .Z(clknet_leaf_53_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_54_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_54_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_55_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_55_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_56_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_56_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_57_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_57_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_58_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_58_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_59_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_59_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_60_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_60_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_61_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_61_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_62_clk_i_regs (.A(clknet_4_11_0_clk_i_regs),
    .Z(clknet_leaf_62_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_63_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_63_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_64_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_64_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_65_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_65_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_66_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_66_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_67_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_67_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_68_clk_i_regs (.A(clknet_4_9_0_clk_i_regs),
    .Z(clknet_leaf_68_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_69_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_69_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_70_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_70_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_71_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_71_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_72_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_72_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_73_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_73_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_74_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_74_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_75_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_75_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_76_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_76_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_77_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_77_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_78_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_78_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_79_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_79_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_80_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_80_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_81_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_81_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_82_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_82_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_83_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_83_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_84_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_84_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_85_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_85_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_86_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_86_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_87_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_87_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_88_clk_i_regs (.A(clknet_4_14_0_clk_i_regs),
    .Z(clknet_leaf_88_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_89_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_89_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_90_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_90_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_91_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_91_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_92_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_92_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_93_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_93_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_94_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_94_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_95_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_95_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_96_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_96_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_97_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_97_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_98_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_98_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_99_clk_i_regs (.A(clknet_4_15_0_clk_i_regs),
    .Z(clknet_leaf_99_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_100_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_100_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_101_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_101_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_102_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_102_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_103_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_103_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_104_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_104_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_105_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_105_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_106_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_106_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_107_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_107_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_108_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_108_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_109_clk_i_regs (.A(clknet_4_13_0_clk_i_regs),
    .Z(clknet_leaf_109_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_110_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_110_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_111_clk_i_regs (.A(clknet_4_12_0_clk_i_regs),
    .Z(clknet_leaf_111_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_112_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_112_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_113_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_113_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_114_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_114_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_115_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_115_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_116_clk_i_regs (.A(clknet_4_7_0_clk_i_regs),
    .Z(clknet_leaf_116_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_117_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_117_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_118_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_118_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_119_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_119_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_120_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_120_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_121_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_121_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_122_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_122_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_123_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_123_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_124_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_124_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_125_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_125_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_126_clk_i_regs (.A(clknet_4_6_0_clk_i_regs),
    .Z(clknet_leaf_126_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_127_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_127_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_128_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_128_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_129_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_129_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_130_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_130_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_131_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_131_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_132_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_132_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_133_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_133_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_134_clk_i_regs (.A(clknet_4_4_0_clk_i_regs),
    .Z(clknet_leaf_134_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_135_clk_i_regs (.A(clknet_4_5_0_clk_i_regs),
    .Z(clknet_leaf_135_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_136_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_136_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_137_clk_i_regs (.A(clknet_4_1_0_clk_i_regs),
    .Z(clknet_leaf_137_clk_i_regs));
 CLKBUF_X3 clkbuf_0_clk_i_regs (.A(clk_i_regs),
    .Z(clknet_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_0_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_0_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_1_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_1_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_2_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_2_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_3_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_3_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_4_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_4_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_5_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_5_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_6_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_6_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_7_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_7_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_8_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_8_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_9_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_9_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_10_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_10_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_11_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_11_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_12_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_12_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_13_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_13_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_14_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_14_0_clk_i_regs));
 CLKBUF_X3 clkbuf_4_15_0_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Z(clknet_4_15_0_clk_i_regs));
 INV_X4 clkload0 (.A(clknet_4_0_0_clk_i_regs));
 INV_X4 clkload1 (.A(clknet_4_1_0_clk_i_regs));
 INV_X4 clkload2 (.A(clknet_4_2_0_clk_i_regs));
 INV_X4 clkload3 (.A(clknet_4_3_0_clk_i_regs));
 INV_X2 clkload4 (.A(clknet_4_4_0_clk_i_regs));
 INV_X4 clkload5 (.A(clknet_4_5_0_clk_i_regs));
 INV_X4 clkload6 (.A(clknet_4_6_0_clk_i_regs));
 INV_X4 clkload7 (.A(clknet_4_7_0_clk_i_regs));
 INV_X2 clkload8 (.A(clknet_4_8_0_clk_i_regs));
 INV_X4 clkload9 (.A(clknet_4_9_0_clk_i_regs));
 INV_X2 clkload10 (.A(clknet_4_10_0_clk_i_regs));
 INV_X2 clkload11 (.A(clknet_4_11_0_clk_i_regs));
 CLKBUF_X3 clkload12 (.A(clknet_4_12_0_clk_i_regs));
 INV_X4 clkload13 (.A(clknet_4_13_0_clk_i_regs));
 CLKBUF_X3 clkload14 (.A(clknet_4_15_0_clk_i_regs));
 CLKBUF_X1 clkload15 (.A(clknet_leaf_2_clk_i_regs));
 INV_X1 clkload16 (.A(clknet_leaf_3_clk_i_regs));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_4_clk_i_regs));
 CLKBUF_X1 clkload18 (.A(clknet_leaf_6_clk_i_regs));
 INV_X1 clkload19 (.A(clknet_leaf_7_clk_i_regs));
 INV_X1 clkload20 (.A(clknet_leaf_8_clk_i_regs));
 INV_X2 clkload21 (.A(clknet_leaf_10_clk_i_regs));
 CLKBUF_X1 clkload22 (.A(clknet_leaf_0_clk_i_regs));
 CLKBUF_X1 clkload23 (.A(clknet_leaf_1_clk_i_regs));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_12_clk_i_regs));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_16_clk_i_regs));
 INV_X2 clkload26 (.A(clknet_leaf_136_clk_i_regs));
 INV_X1 clkload27 (.A(clknet_leaf_9_clk_i_regs));
 INV_X1 clkload28 (.A(clknet_leaf_28_clk_i_regs));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_29_clk_i_regs));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_30_clk_i_regs));
 INV_X1 clkload31 (.A(clknet_leaf_31_clk_i_regs));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_32_clk_i_regs));
 INV_X1 clkload33 (.A(clknet_leaf_33_clk_i_regs));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_15_clk_i_regs));
 INV_X1 clkload35 (.A(clknet_leaf_19_clk_i_regs));
 INV_X1 clkload36 (.A(clknet_leaf_20_clk_i_regs));
 CLKBUF_X1 clkload37 (.A(clknet_leaf_21_clk_i_regs));
 INV_X1 clkload38 (.A(clknet_leaf_22_clk_i_regs));
 CLKBUF_X1 clkload39 (.A(clknet_leaf_23_clk_i_regs));
 INV_X1 clkload40 (.A(clknet_leaf_27_clk_i_regs));
 INV_X1 clkload41 (.A(clknet_leaf_13_clk_i_regs));
 INV_X2 clkload42 (.A(clknet_leaf_127_clk_i_regs));
 CLKBUF_X1 clkload43 (.A(clknet_leaf_129_clk_i_regs));
 INV_X1 clkload44 (.A(clknet_leaf_130_clk_i_regs));
 INV_X2 clkload45 (.A(clknet_leaf_131_clk_i_regs));
 INV_X1 clkload46 (.A(clknet_leaf_133_clk_i_regs));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_134_clk_i_regs));
 INV_X4 clkload48 (.A(clknet_leaf_117_clk_i_regs));
 INV_X2 clkload49 (.A(clknet_leaf_118_clk_i_regs));
 INV_X2 clkload50 (.A(clknet_leaf_119_clk_i_regs));
 CLKBUF_X1 clkload51 (.A(clknet_leaf_121_clk_i_regs));
 CLKBUF_X1 clkload52 (.A(clknet_leaf_14_clk_i_regs));
 INV_X2 clkload53 (.A(clknet_leaf_17_clk_i_regs));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_18_clk_i_regs));
 INV_X1 clkload55 (.A(clknet_leaf_124_clk_i_regs));
 CLKBUF_X1 clkload56 (.A(clknet_leaf_125_clk_i_regs));
 INV_X1 clkload57 (.A(clknet_leaf_126_clk_i_regs));
 CLKBUF_X1 clkload58 (.A(clknet_leaf_112_clk_i_regs));
 INV_X1 clkload59 (.A(clknet_leaf_113_clk_i_regs));
 CLKBUF_X1 clkload60 (.A(clknet_leaf_114_clk_i_regs));
 INV_X1 clkload61 (.A(clknet_leaf_115_clk_i_regs));
 INV_X1 clkload62 (.A(clknet_leaf_116_clk_i_regs));
 INV_X1 clkload63 (.A(clknet_leaf_39_clk_i_regs));
 CLKBUF_X1 clkload64 (.A(clknet_leaf_40_clk_i_regs));
 INV_X1 clkload65 (.A(clknet_leaf_41_clk_i_regs));
 CLKBUF_X1 clkload66 (.A(clknet_leaf_44_clk_i_regs));
 CLKBUF_X1 clkload67 (.A(clknet_leaf_24_clk_i_regs));
 CLKBUF_X1 clkload68 (.A(clknet_leaf_63_clk_i_regs));
 CLKBUF_X1 clkload69 (.A(clknet_leaf_66_clk_i_regs));
 CLKBUF_X1 clkload70 (.A(clknet_leaf_68_clk_i_regs));
 CLKBUF_X1 clkload71 (.A(clknet_leaf_46_clk_i_regs));
 INV_X2 clkload72 (.A(clknet_leaf_47_clk_i_regs));
 CLKBUF_X1 clkload73 (.A(clknet_leaf_48_clk_i_regs));
 INV_X1 clkload74 (.A(clknet_leaf_49_clk_i_regs));
 CLKBUF_X1 clkload75 (.A(clknet_leaf_51_clk_i_regs));
 CLKBUF_X1 clkload76 (.A(clknet_leaf_53_clk_i_regs));
 CLKBUF_X1 clkload77 (.A(clknet_leaf_56_clk_i_regs));
 CLKBUF_X1 clkload78 (.A(clknet_leaf_58_clk_i_regs));
 CLKBUF_X1 clkload79 (.A(clknet_leaf_59_clk_i_regs));
 INV_X1 clkload80 (.A(clknet_leaf_60_clk_i_regs));
 CLKBUF_X1 clkload81 (.A(clknet_leaf_61_clk_i_regs));
 CLKBUF_X1 clkload82 (.A(clknet_leaf_62_clk_i_regs));
 CLKBUF_X1 clkload83 (.A(clknet_leaf_69_clk_i_regs));
 CLKBUF_X1 clkload84 (.A(clknet_leaf_70_clk_i_regs));
 CLKBUF_X1 clkload85 (.A(clknet_leaf_71_clk_i_regs));
 INV_X1 clkload86 (.A(clknet_leaf_73_clk_i_regs));
 INV_X1 clkload87 (.A(clknet_leaf_74_clk_i_regs));
 CLKBUF_X1 clkload88 (.A(clknet_leaf_76_clk_i_regs));
 CLKBUF_X1 clkload89 (.A(clknet_leaf_100_clk_i_regs));
 INV_X1 clkload90 (.A(clknet_leaf_101_clk_i_regs));
 INV_X1 clkload91 (.A(clknet_leaf_102_clk_i_regs));
 CLKBUF_X1 clkload92 (.A(clknet_leaf_104_clk_i_regs));
 CLKBUF_X1 clkload93 (.A(clknet_leaf_105_clk_i_regs));
 CLKBUF_X1 clkload94 (.A(clknet_leaf_106_clk_i_regs));
 INV_X1 clkload95 (.A(clknet_leaf_109_clk_i_regs));
 INV_X1 clkload96 (.A(clknet_leaf_77_clk_i_regs));
 CLKBUF_X1 clkload97 (.A(clknet_leaf_78_clk_i_regs));
 CLKBUF_X1 clkload98 (.A(clknet_leaf_82_clk_i_regs));
 CLKBUF_X1 clkload99 (.A(clknet_leaf_88_clk_i_regs));
 CLKBUF_X1 clkload100 (.A(clknet_leaf_89_clk_i_regs));
 INV_X1 clkload101 (.A(clknet_leaf_90_clk_i_regs));
 CLKBUF_X1 clkload102 (.A(clknet_leaf_91_clk_i_regs));
 CLKBUF_X1 clkload103 (.A(clknet_leaf_92_clk_i_regs));
 INV_X1 clkload104 (.A(clknet_leaf_93_clk_i_regs));
 INV_X2 clkload105 (.A(clknet_leaf_94_clk_i_regs));
 INV_X1 clkload106 (.A(clknet_leaf_95_clk_i_regs));
 INV_X2 clkload107 (.A(clknet_leaf_97_clk_i_regs));
 INV_X2 clkload108 (.A(clknet_leaf_98_clk_i_regs));
 CLKBUF_X1 clkload109 (.A(clknet_leaf_99_clk_i_regs));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_leaf_83_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_83_clk));
 CLKBUF_X3 clkbuf_leaf_84_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_84_clk));
 CLKBUF_X3 clkbuf_leaf_85_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_85_clk));
 CLKBUF_X3 clkbuf_leaf_86_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_86_clk));
 CLKBUF_X3 clkbuf_leaf_87_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_87_clk));
 CLKBUF_X3 clkbuf_leaf_88_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_88_clk));
 CLKBUF_X3 clkbuf_leaf_89_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_89_clk));
 CLKBUF_X3 clkbuf_leaf_90_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_90_clk));
 CLKBUF_X3 clkbuf_leaf_91_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_91_clk));
 CLKBUF_X3 clkbuf_leaf_92_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_92_clk));
 CLKBUF_X3 clkbuf_leaf_93_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_93_clk));
 CLKBUF_X3 clkbuf_leaf_94_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_94_clk));
 CLKBUF_X3 clkbuf_leaf_95_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_95_clk));
 CLKBUF_X3 clkbuf_leaf_96_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_96_clk));
 CLKBUF_X3 clkbuf_leaf_97_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_97_clk));
 CLKBUF_X3 clkbuf_leaf_98_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_98_clk));
 CLKBUF_X3 clkbuf_leaf_99_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_99_clk));
 CLKBUF_X3 clkbuf_leaf_100_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_100_clk));
 CLKBUF_X3 clkbuf_leaf_101_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_101_clk));
 CLKBUF_X3 clkbuf_leaf_102_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_102_clk));
 CLKBUF_X3 clkbuf_leaf_103_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_103_clk));
 CLKBUF_X3 clkbuf_leaf_104_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_104_clk));
 CLKBUF_X3 clkbuf_leaf_105_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_105_clk));
 CLKBUF_X3 clkbuf_leaf_106_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_106_clk));
 CLKBUF_X3 clkbuf_leaf_107_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_107_clk));
 CLKBUF_X3 clkbuf_leaf_108_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_108_clk));
 CLKBUF_X3 clkbuf_leaf_109_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_109_clk));
 CLKBUF_X3 clkbuf_leaf_110_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_110_clk));
 CLKBUF_X3 clkbuf_leaf_111_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_111_clk));
 CLKBUF_X3 clkbuf_leaf_112_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_112_clk));
 CLKBUF_X3 clkbuf_leaf_113_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_113_clk));
 CLKBUF_X3 clkbuf_leaf_114_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_114_clk));
 CLKBUF_X3 clkbuf_leaf_115_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_115_clk));
 CLKBUF_X3 clkbuf_leaf_116_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_116_clk));
 CLKBUF_X3 clkbuf_leaf_117_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_117_clk));
 CLKBUF_X3 clkbuf_leaf_118_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_118_clk));
 CLKBUF_X3 clkbuf_leaf_119_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_119_clk));
 CLKBUF_X3 clkbuf_leaf_120_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_120_clk));
 CLKBUF_X3 clkbuf_leaf_121_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_121_clk));
 CLKBUF_X3 clkbuf_leaf_122_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_122_clk));
 CLKBUF_X3 clkbuf_leaf_123_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_123_clk));
 CLKBUF_X3 clkbuf_leaf_124_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_124_clk));
 CLKBUF_X3 clkbuf_leaf_125_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_125_clk));
 CLKBUF_X3 clkbuf_leaf_126_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_126_clk));
 CLKBUF_X3 clkbuf_leaf_127_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_127_clk));
 CLKBUF_X3 clkbuf_leaf_128_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_128_clk));
 CLKBUF_X3 clkbuf_leaf_129_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_129_clk));
 CLKBUF_X3 clkbuf_leaf_130_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_130_clk));
 CLKBUF_X3 clkbuf_leaf_131_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_131_clk));
 CLKBUF_X3 clkbuf_leaf_132_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_132_clk));
 CLKBUF_X3 clkbuf_leaf_133_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_133_clk));
 CLKBUF_X3 clkbuf_leaf_134_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_134_clk));
 CLKBUF_X3 clkbuf_leaf_135_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_135_clk));
 CLKBUF_X3 clkbuf_leaf_136_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_136_clk));
 CLKBUF_X3 clkbuf_leaf_137_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_137_clk));
 CLKBUF_X3 clkbuf_leaf_138_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_138_clk));
 CLKBUF_X3 clkbuf_leaf_139_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_139_clk));
 CLKBUF_X3 clkbuf_leaf_140_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_140_clk));
 CLKBUF_X3 clkbuf_leaf_141_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_141_clk));
 CLKBUF_X3 clkbuf_leaf_142_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_142_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X4 clkload110 (.A(clknet_4_0_0_clk));
 INV_X2 clkload111 (.A(clknet_4_1_0_clk));
 INV_X4 clkload112 (.A(clknet_4_2_0_clk));
 INV_X8 clkload113 (.A(clknet_4_3_0_clk));
 INV_X8 clkload114 (.A(clknet_4_4_0_clk));
 INV_X8 clkload115 (.A(clknet_4_5_0_clk));
 INV_X4 clkload116 (.A(clknet_4_6_0_clk));
 INV_X8 clkload117 (.A(clknet_4_7_0_clk));
 INV_X2 clkload118 (.A(clknet_4_8_0_clk));
 INV_X8 clkload119 (.A(clknet_4_9_0_clk));
 CLKBUF_X3 clkload120 (.A(clknet_4_10_0_clk));
 INV_X8 clkload121 (.A(clknet_4_12_0_clk));
 INV_X4 clkload122 (.A(clknet_4_13_0_clk));
 INV_X2 clkload123 (.A(clknet_4_14_0_clk));
 INV_X2 clkload124 (.A(clknet_4_15_0_clk));
 CLKBUF_X1 clkload125 (.A(clknet_leaf_0_clk));
 CLKBUF_X1 clkload126 (.A(clknet_leaf_132_clk));
 INV_X1 clkload127 (.A(clknet_leaf_134_clk));
 CLKBUF_X1 clkload128 (.A(clknet_leaf_135_clk));
 CLKBUF_X2 clkload129 (.A(clknet_leaf_136_clk));
 CLKBUF_X1 clkload130 (.A(clknet_leaf_137_clk));
 INV_X4 clkload131 (.A(clknet_leaf_138_clk));
 CLKBUF_X1 clkload132 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload133 (.A(clknet_leaf_2_clk));
 INV_X1 clkload134 (.A(clknet_leaf_3_clk));
 INV_X1 clkload135 (.A(clknet_leaf_4_clk));
 CLKBUF_X1 clkload136 (.A(clknet_leaf_5_clk));
 INV_X2 clkload137 (.A(clknet_leaf_7_clk));
 INV_X1 clkload138 (.A(clknet_leaf_139_clk));
 INV_X1 clkload139 (.A(clknet_leaf_141_clk));
 CLKBUF_X1 clkload140 (.A(clknet_leaf_142_clk));
 INV_X1 clkload141 (.A(clknet_leaf_105_clk));
 INV_X1 clkload142 (.A(clknet_leaf_106_clk));
 INV_X1 clkload143 (.A(clknet_leaf_126_clk));
 INV_X1 clkload144 (.A(clknet_leaf_127_clk));
 INV_X1 clkload145 (.A(clknet_leaf_128_clk));
 INV_X1 clkload146 (.A(clknet_leaf_129_clk));
 INV_X1 clkload147 (.A(clknet_leaf_131_clk));
 CLKBUF_X1 clkload148 (.A(clknet_leaf_133_clk));
 INV_X2 clkload149 (.A(clknet_leaf_107_clk));
 INV_X1 clkload150 (.A(clknet_leaf_108_clk));
 CLKBUF_X1 clkload151 (.A(clknet_leaf_109_clk));
 CLKBUF_X1 clkload152 (.A(clknet_leaf_122_clk));
 INV_X1 clkload153 (.A(clknet_leaf_123_clk));
 INV_X2 clkload154 (.A(clknet_leaf_12_clk));
 CLKBUF_X1 clkload155 (.A(clknet_leaf_13_clk));
 CLKBUF_X1 clkload156 (.A(clknet_leaf_14_clk));
 INV_X2 clkload157 (.A(clknet_leaf_15_clk));
 INV_X1 clkload158 (.A(clknet_leaf_17_clk));
 CLKBUF_X1 clkload159 (.A(clknet_leaf_18_clk));
 INV_X1 clkload160 (.A(clknet_leaf_19_clk));
 INV_X2 clkload161 (.A(clknet_leaf_20_clk));
 INV_X1 clkload162 (.A(clknet_leaf_8_clk));
 INV_X1 clkload163 (.A(clknet_leaf_11_clk));
 INV_X2 clkload164 (.A(clknet_leaf_118_clk));
 CLKBUF_X1 clkload165 (.A(clknet_leaf_119_clk));
 CLKBUF_X1 clkload166 (.A(clknet_leaf_120_clk));
 INV_X2 clkload167 (.A(clknet_leaf_124_clk));
 INV_X1 clkload168 (.A(clknet_leaf_125_clk));
 INV_X2 clkload169 (.A(clknet_leaf_55_clk));
 CLKBUF_X1 clkload170 (.A(clknet_leaf_59_clk));
 CLKBUF_X1 clkload171 (.A(clknet_leaf_115_clk));
 INV_X2 clkload172 (.A(clknet_leaf_116_clk));
 INV_X2 clkload173 (.A(clknet_leaf_117_clk));
 CLKBUF_X1 clkload174 (.A(clknet_leaf_92_clk));
 CLKBUF_X1 clkload175 (.A(clknet_leaf_93_clk));
 CLKBUF_X1 clkload176 (.A(clknet_leaf_94_clk));
 CLKBUF_X1 clkload177 (.A(clknet_leaf_96_clk));
 CLKBUF_X1 clkload178 (.A(clknet_leaf_98_clk));
 CLKBUF_X1 clkload179 (.A(clknet_leaf_100_clk));
 CLKBUF_X1 clkload180 (.A(clknet_leaf_101_clk));
 CLKBUF_X1 clkload181 (.A(clknet_leaf_102_clk));
 INV_X1 clkload182 (.A(clknet_leaf_103_clk));
 CLKBUF_X1 clkload183 (.A(clknet_leaf_104_clk));
 CLKBUF_X1 clkload184 (.A(clknet_leaf_111_clk));
 CLKBUF_X1 clkload185 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload186 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload187 (.A(clknet_leaf_97_clk));
 CLKBUF_X1 clkload188 (.A(clknet_leaf_112_clk));
 CLKBUF_X1 clkload189 (.A(clknet_leaf_113_clk));
 CLKBUF_X1 clkload190 (.A(clknet_leaf_114_clk));
 CLKBUF_X1 clkload191 (.A(clknet_leaf_80_clk));
 CLKBUF_X1 clkload192 (.A(clknet_leaf_81_clk));
 CLKBUF_X1 clkload193 (.A(clknet_leaf_82_clk));
 CLKBUF_X1 clkload194 (.A(clknet_leaf_83_clk));
 INV_X1 clkload195 (.A(clknet_leaf_84_clk));
 CLKBUF_X1 clkload196 (.A(clknet_leaf_85_clk));
 INV_X1 clkload197 (.A(clknet_leaf_86_clk));
 CLKBUF_X1 clkload198 (.A(clknet_leaf_87_clk));
 CLKBUF_X1 clkload199 (.A(clknet_leaf_88_clk));
 CLKBUF_X1 clkload200 (.A(clknet_leaf_90_clk));
 CLKBUF_X1 clkload201 (.A(clknet_leaf_91_clk));
 CLKBUF_X1 clkload202 (.A(clknet_leaf_95_clk));
 CLKBUF_X1 clkload203 (.A(clknet_leaf_62_clk));
 INV_X1 clkload204 (.A(clknet_leaf_64_clk));
 CLKBUF_X1 clkload205 (.A(clknet_leaf_65_clk));
 CLKBUF_X2 clkload206 (.A(clknet_leaf_68_clk));
 CLKBUF_X2 clkload207 (.A(clknet_leaf_71_clk));
 CLKBUF_X1 clkload208 (.A(clknet_leaf_72_clk));
 INV_X1 clkload209 (.A(clknet_leaf_73_clk));
 INV_X1 clkload210 (.A(clknet_leaf_74_clk));
 CLKBUF_X1 clkload211 (.A(clknet_leaf_75_clk));
 INV_X1 clkload212 (.A(clknet_leaf_76_clk));
 INV_X2 clkload213 (.A(clknet_leaf_77_clk));
 CLKBUF_X1 clkload214 (.A(clknet_leaf_78_clk));
 INV_X1 clkload215 (.A(clknet_leaf_79_clk));
 INV_X1 clkload216 (.A(clknet_leaf_21_clk));
 CLKBUF_X1 clkload217 (.A(clknet_leaf_28_clk));
 CLKBUF_X1 clkload218 (.A(clknet_leaf_52_clk));
 INV_X1 clkload219 (.A(clknet_leaf_53_clk));
 CLKBUF_X1 clkload220 (.A(clknet_leaf_54_clk));
 CLKBUF_X1 clkload221 (.A(clknet_leaf_66_clk));
 INV_X1 clkload222 (.A(clknet_leaf_22_clk));
 INV_X1 clkload223 (.A(clknet_leaf_23_clk));
 INV_X2 clkload224 (.A(clknet_leaf_25_clk));
 INV_X1 clkload225 (.A(clknet_leaf_26_clk));
 CLKBUF_X1 clkload226 (.A(clknet_leaf_27_clk));
 INV_X1 clkload227 (.A(clknet_leaf_29_clk));
 INV_X2 clkload228 (.A(clknet_leaf_30_clk));
 CLKBUF_X1 clkload229 (.A(clknet_leaf_40_clk));
 INV_X1 clkload230 (.A(clknet_leaf_45_clk));
 CLKBUF_X1 clkload231 (.A(clknet_leaf_46_clk));
 CLKBUF_X1 clkload232 (.A(clknet_leaf_47_clk));
 CLKBUF_X1 clkload233 (.A(clknet_leaf_48_clk));
 CLKBUF_X1 clkload234 (.A(clknet_leaf_49_clk));
 CLKBUF_X1 clkload235 (.A(clknet_leaf_50_clk));
 INV_X1 clkload236 (.A(clknet_leaf_51_clk));
 CLKBUF_X1 clkload237 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload238 (.A(clknet_leaf_69_clk));
 CLKBUF_X1 clkload239 (.A(clknet_leaf_70_clk));
 CLKBUF_X1 clkload240 (.A(clknet_leaf_31_clk));
 CLKBUF_X1 clkload241 (.A(clknet_leaf_32_clk));
 CLKBUF_X1 clkload242 (.A(clknet_leaf_33_clk));
 CLKBUF_X1 clkload243 (.A(clknet_leaf_34_clk));
 INV_X1 clkload244 (.A(clknet_leaf_35_clk));
 CLKBUF_X1 clkload245 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload246 (.A(clknet_leaf_38_clk));
 INV_X1 clkload247 (.A(clknet_leaf_39_clk));
 INV_X1 clkload248 (.A(clknet_leaf_41_clk));
 CLKBUF_X1 clkload249 (.A(clknet_leaf_42_clk));
 INV_X1 clkload250 (.A(clknet_leaf_43_clk));
 CLKBUF_X3 delaybuf_0_core_clock (.A(delaynet_0_core_clock),
    .Z(delaynet_1_core_clock));
 CLKBUF_X3 delaybuf_1_core_clock (.A(delaynet_1_core_clock),
    .Z(clk_i_regs));
 BUF_X4 rebuffer1 (.A(_12527_),
    .Z(net275));
 BUF_X1 rebuffer2 (.A(_11166_),
    .Z(net276));
 BUF_X1 rebuffer3 (.A(net276),
    .Z(net277));
 BUF_X1 rebuffer4 (.A(net276),
    .Z(net278));
 BUF_X1 rebuffer5 (.A(_16102_),
    .Z(net279));
 BUF_X1 rebuffer6 (.A(_16109_),
    .Z(net280));
 BUF_X4 rebuffer7 (.A(_12752_),
    .Z(net281));
 BUF_X1 rebuffer8 (.A(net281),
    .Z(net282));
 BUF_X4 rebuffer9 (.A(_13012_),
    .Z(net283));
 BUF_X1 rebuffer10 (.A(net283),
    .Z(net284));
 BUF_X1 rebuffer11 (.A(net283),
    .Z(net285));
 BUF_X8 rebuffer12 (.A(_12936_),
    .Z(net286));
 BUF_X1 rebuffer13 (.A(net286),
    .Z(net287));
 XOR2_X1 clone15 (.A(_03511_),
    .B(_03516_),
    .Z(net289));
 BUF_X4 clone16 (.A(_03508_),
    .Z(net290));
 BUF_X2 rebuffer18 (.A(\id_stage_i.controller_i.instr_i[14] ),
    .Z(net292));
 BUF_X2 rebuffer19 (.A(net292),
    .Z(net293));
 BUF_X1 rebuffer20 (.A(_10901_),
    .Z(net294));
 BUF_X1 rebuffer21 (.A(_10901_),
    .Z(net295));
 BUF_X1 rebuffer22 (.A(_10901_),
    .Z(net296));
 BUF_X4 rebuffer23 (.A(_10870_),
    .Z(net297));
 BUF_X1 rebuffer24 (.A(net297),
    .Z(net298));
 BUF_X1 rebuffer26 (.A(_10879_),
    .Z(net300));
 BUF_X2 rebuffer27 (.A(_10765_),
    .Z(net301));
 BUF_X1 rebuffer28 (.A(net301),
    .Z(net302));
 BUF_X4 clone29 (.A(net304),
    .Z(net303));
 BUF_X1 rebuffer30 (.A(\id_stage_i.controller_i.instr_i[14] ),
    .Z(net304));
 BUF_X1 rebuffer31 (.A(_10950_),
    .Z(net305));
 BUF_X8 clone33 (.A(net414),
    .Z(net307));
 BUF_X1 rebuffer35 (.A(net308),
    .Z(net309));
 BUF_X4 rebuffer36 (.A(_10786_),
    .Z(net310));
 BUF_X1 rebuffer37 (.A(net310),
    .Z(net311));
 BUF_X2 rebuffer38 (.A(_13118_),
    .Z(net312));
 BUF_X16 clone40 (.A(net372),
    .Z(net314));
 NOR2_X2 clone41 (.A1(_03931_),
    .A2(_03791_),
    .ZN(net315));
 BUF_X4 clone42 (.A(_03850_),
    .Z(net316));
 MUX2_X1 clone43 (.A(_03849_),
    .B(_13384_),
    .S(_03789_),
    .Z(net317));
 BUF_X1 rebuffer44 (.A(_12656_),
    .Z(net318));
 AOI21_X2 clone45 (.A(_13368_),
    .B1(_13117_),
    .B2(net320),
    .ZN(net319));
 BUF_X1 rebuffer46 (.A(_13383_),
    .Z(net320));
 BUF_X4 clone47 (.A(_03840_),
    .Z(net321));
 MUX2_X1 clone48 (.A(net363),
    .B(_13307_),
    .S(_03788_),
    .Z(net322));
 AOI21_X2 clone49 (.A(_13288_),
    .B1(_13117_),
    .B2(net324),
    .ZN(net323));
 BUF_X1 rebuffer50 (.A(_13306_),
    .Z(net324));
 BUF_X1 rebuffer51 (.A(_12473_),
    .Z(net325));
 BUF_X2 rebuffer52 (.A(_14983_),
    .Z(net326));
 BUF_X1 rebuffer53 (.A(net326),
    .Z(net327));
 BUF_X16 clone84 (.A(net372),
    .Z(net358));
 BUF_X16 clone97 (.A(net372),
    .Z(net371));
 BUF_X8 rebuffer98 (.A(_06476_),
    .Z(net372));
 BUF_X4 clone99 (.A(_03832_),
    .Z(net373));
 BUF_X32 clone100 (.A(_10750_),
    .Z(net374));
 BUF_X8 clone101 (.A(_10699_),
    .Z(net375));
 BUF_X1 rebuffer102 (.A(_16074_),
    .Z(net376));
 BUF_X16 clone103 (.A(net380),
    .Z(net377));
 BUF_X16 clone104 (.A(_10703_),
    .Z(net378));
 BUF_X16 clone105 (.A(_10704_),
    .Z(net379));
 BUF_X16 clone106 (.A(net342),
    .Z(net380));
 BUF_X4 clone325 (.A(_06422_),
    .Z(net599));
 CLKBUF_X1 hold355 (.A(net631),
    .Z(net629));
 CLKBUF_X3 hold356 (.A(net144),
    .Z(net630));
 CLKBUF_X1 hold357 (.A(rst_ni),
    .Z(net631));
 BUF_X1 rebuffer15 (.A(_03517_),
    .Z(net313));
 BUF_X1 rebuffer16 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .Z(net328));
 BUF_X1 rebuffer29 (.A(net332),
    .Z(net329));
 BUF_X2 rebuffer33 (.A(_11470_),
    .Z(net330));
 BUF_X1 rebuffer39 (.A(net330),
    .Z(net331));
 BUF_X1 rebuffer40 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .Z(net332));
 BUF_X1 rebuffer41 (.A(_10909_),
    .Z(net333));
 BUF_X16 clone53 (.A(_10704_),
    .Z(net341));
 BUF_X16 clone54 (.A(_10700_),
    .Z(net342));
 BUF_X16 clone55 (.A(net374),
    .Z(net343));
 BUF_X16 clone56 (.A(net374),
    .Z(net344));
 BUF_X1 rebuffer57 (.A(\alu_adder_result_ex[30] ),
    .Z(net345));
 BUF_X1 rebuffer58 (.A(net345),
    .Z(net346));
 BUF_X2 rebuffer59 (.A(_15788_),
    .Z(net347));
 BUF_X1 rebuffer60 (.A(net347),
    .Z(net348));
 BUF_X1 rebuffer61 (.A(_15812_),
    .Z(net349));
 BUF_X4 rebuffer62 (.A(_13384_),
    .Z(net350));
 BUF_X1 rebuffer69 (.A(net356),
    .Z(net357));
 BUF_X1 rebuffer70 (.A(\alu_adder_result_ex[23] ),
    .Z(net359));
 BUF_X1 rebuffer71 (.A(_11929_),
    .Z(net360));
 BUF_X1 rebuffer72 (.A(_11570_),
    .Z(net361));
 BUF_X1 rebuffer73 (.A(net361),
    .Z(net362));
 BUF_X1 rebuffer74 (.A(net361),
    .Z(net363));
 BUF_X2 rebuffer75 (.A(_11375_),
    .Z(net364));
 BUF_X1 rebuffer76 (.A(net364),
    .Z(net365));
 BUF_X1 rebuffer77 (.A(_10840_),
    .Z(net366));
 BUF_X1 rebuffer78 (.A(_10840_),
    .Z(net367));
 BUF_X8 rebuffer79 (.A(_13118_),
    .Z(net368));
 BUF_X1 rebuffer80 (.A(net368),
    .Z(net369));
 XNOR2_X1 clone87 (.A(_03336_),
    .B(_03321_),
    .ZN(net386));
 BUF_X1 rebuffer89 (.A(\alu_adder_result_ex[25] ),
    .Z(net388));
 BUF_X1 rebuffer90 (.A(net388),
    .Z(net389));
 BUF_X1 rebuffer91 (.A(\alu_adder_result_ex[25] ),
    .Z(net390));
 BUF_X1 rebuffer92 (.A(_03162_),
    .Z(net391));
 BUF_X1 rebuffer93 (.A(_03162_),
    .Z(net392));
 AOI21_X2 clone120 (.A(_03327_),
    .B1(_03332_),
    .B2(_03329_),
    .ZN(net411));
 BUF_X4 rebuffer121 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .Z(net412));
 BUF_X1 rebuffer122 (.A(_10903_),
    .Z(net413));
 BUF_X8 clone123 (.A(_10776_),
    .Z(net414));
 BUF_X1 rebuffer144 (.A(_13266_),
    .Z(net435));
 BUF_X1 rebuffer147 (.A(net437),
    .Z(net438));
 BUF_X1 rebuffer148 (.A(net437),
    .Z(net439));
 BUF_X4 clone159 (.A(_06422_),
    .Z(net450));
 BUF_X16 clone165 (.A(_06456_),
    .Z(net456));
 BUF_X16 clone166 (.A(_06456_),
    .Z(net457));
 BUF_X4 clone167 (.A(_06422_),
    .Z(net458));
 BUF_X16 clone168 (.A(_06456_),
    .Z(net459));
 BUF_X4 clone169 (.A(net461),
    .Z(net460));
 BUF_X4 rebuffer170 (.A(_06255_),
    .Z(net461));
 BUF_X4 clone192 (.A(_06328_),
    .Z(net483));
 BUF_X4 clone193 (.A(_06328_),
    .Z(net484));
 BUF_X4 clone194 (.A(_06328_),
    .Z(net485));
 XNOR2_X1 clone195 (.A(_12333_),
    .B(_12325_),
    .ZN(net486));
 BUF_X8 clone196 (.A(_06309_),
    .Z(net487));
 BUF_X8 clone197 (.A(_06309_),
    .Z(net488));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_17 ();
 FILLCELL_X4 FILLER_0_25 ();
 FILLCELL_X2 FILLER_0_29 ();
 FILLCELL_X1 FILLER_0_31 ();
 FILLCELL_X4 FILLER_0_35 ();
 FILLCELL_X8 FILLER_0_42 ();
 FILLCELL_X2 FILLER_0_50 ();
 FILLCELL_X1 FILLER_0_52 ();
 FILLCELL_X32 FILLER_0_60 ();
 FILLCELL_X32 FILLER_0_92 ();
 FILLCELL_X32 FILLER_0_124 ();
 FILLCELL_X32 FILLER_0_156 ();
 FILLCELL_X32 FILLER_0_188 ();
 FILLCELL_X32 FILLER_0_220 ();
 FILLCELL_X32 FILLER_0_252 ();
 FILLCELL_X32 FILLER_0_284 ();
 FILLCELL_X32 FILLER_0_316 ();
 FILLCELL_X8 FILLER_0_348 ();
 FILLCELL_X4 FILLER_0_356 ();
 FILLCELL_X2 FILLER_0_360 ();
 FILLCELL_X2 FILLER_0_366 ();
 FILLCELL_X4 FILLER_0_372 ();
 FILLCELL_X4 FILLER_0_384 ();
 FILLCELL_X2 FILLER_0_388 ();
 FILLCELL_X4 FILLER_0_394 ();
 FILLCELL_X1 FILLER_0_398 ();
 FILLCELL_X16 FILLER_0_407 ();
 FILLCELL_X2 FILLER_0_423 ();
 FILLCELL_X8 FILLER_0_433 ();
 FILLCELL_X2 FILLER_0_441 ();
 FILLCELL_X1 FILLER_0_443 ();
 FILLCELL_X1 FILLER_0_448 ();
 FILLCELL_X4 FILLER_0_453 ();
 FILLCELL_X2 FILLER_0_457 ();
 FILLCELL_X2 FILLER_0_471 ();
 FILLCELL_X1 FILLER_0_473 ();
 FILLCELL_X4 FILLER_0_478 ();
 FILLCELL_X1 FILLER_0_482 ();
 FILLCELL_X8 FILLER_0_491 ();
 FILLCELL_X4 FILLER_0_503 ();
 FILLCELL_X2 FILLER_0_507 ();
 FILLCELL_X1 FILLER_0_509 ();
 FILLCELL_X4 FILLER_0_527 ();
 FILLCELL_X8 FILLER_0_535 ();
 FILLCELL_X4 FILLER_0_546 ();
 FILLCELL_X1 FILLER_0_570 ();
 FILLCELL_X2 FILLER_0_584 ();
 FILLCELL_X1 FILLER_0_613 ();
 FILLCELL_X1 FILLER_0_621 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X16 FILLER_0_654 ();
 FILLCELL_X8 FILLER_0_670 ();
 FILLCELL_X1 FILLER_0_678 ();
 FILLCELL_X4 FILLER_0_706 ();
 FILLCELL_X2 FILLER_0_710 ();
 FILLCELL_X1 FILLER_0_716 ();
 FILLCELL_X4 FILLER_0_737 ();
 FILLCELL_X1 FILLER_0_745 ();
 FILLCELL_X1 FILLER_0_749 ();
 FILLCELL_X4 FILLER_0_754 ();
 FILLCELL_X1 FILLER_0_758 ();
 FILLCELL_X1 FILLER_0_802 ();
 FILLCELL_X1 FILLER_0_831 ();
 FILLCELL_X2 FILLER_0_855 ();
 FILLCELL_X2 FILLER_0_912 ();
 FILLCELL_X4 FILLER_0_949 ();
 FILLCELL_X1 FILLER_0_961 ();
 FILLCELL_X4 FILLER_0_973 ();
 FILLCELL_X1 FILLER_0_977 ();
 FILLCELL_X4 FILLER_0_1017 ();
 FILLCELL_X1 FILLER_0_1021 ();
 FILLCELL_X8 FILLER_0_1029 ();
 FILLCELL_X4 FILLER_0_1037 ();
 FILLCELL_X32 FILLER_0_1063 ();
 FILLCELL_X32 FILLER_0_1095 ();
 FILLCELL_X32 FILLER_0_1127 ();
 FILLCELL_X32 FILLER_0_1159 ();
 FILLCELL_X32 FILLER_0_1191 ();
 FILLCELL_X32 FILLER_0_1223 ();
 FILLCELL_X4 FILLER_0_1255 ();
 FILLCELL_X1 FILLER_0_1259 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X16 FILLER_1_321 ();
 FILLCELL_X8 FILLER_1_337 ();
 FILLCELL_X4 FILLER_1_345 ();
 FILLCELL_X2 FILLER_1_349 ();
 FILLCELL_X1 FILLER_1_351 ();
 FILLCELL_X16 FILLER_1_356 ();
 FILLCELL_X1 FILLER_1_372 ();
 FILLCELL_X32 FILLER_1_377 ();
 FILLCELL_X32 FILLER_1_409 ();
 FILLCELL_X32 FILLER_1_441 ();
 FILLCELL_X8 FILLER_1_473 ();
 FILLCELL_X4 FILLER_1_481 ();
 FILLCELL_X2 FILLER_1_485 ();
 FILLCELL_X8 FILLER_1_495 ();
 FILLCELL_X2 FILLER_1_503 ();
 FILLCELL_X16 FILLER_1_525 ();
 FILLCELL_X4 FILLER_1_541 ();
 FILLCELL_X1 FILLER_1_545 ();
 FILLCELL_X1 FILLER_1_568 ();
 FILLCELL_X8 FILLER_1_638 ();
 FILLCELL_X2 FILLER_1_646 ();
 FILLCELL_X1 FILLER_1_648 ();
 FILLCELL_X16 FILLER_1_673 ();
 FILLCELL_X8 FILLER_1_689 ();
 FILLCELL_X2 FILLER_1_697 ();
 FILLCELL_X1 FILLER_1_699 ();
 FILLCELL_X1 FILLER_1_719 ();
 FILLCELL_X1 FILLER_1_723 ();
 FILLCELL_X4 FILLER_1_728 ();
 FILLCELL_X1 FILLER_1_732 ();
 FILLCELL_X8 FILLER_1_783 ();
 FILLCELL_X2 FILLER_1_791 ();
 FILLCELL_X2 FILLER_1_800 ();
 FILLCELL_X1 FILLER_1_802 ();
 FILLCELL_X1 FILLER_1_806 ();
 FILLCELL_X2 FILLER_1_811 ();
 FILLCELL_X1 FILLER_1_820 ();
 FILLCELL_X1 FILLER_1_824 ();
 FILLCELL_X1 FILLER_1_834 ();
 FILLCELL_X1 FILLER_1_838 ();
 FILLCELL_X4 FILLER_1_846 ();
 FILLCELL_X2 FILLER_1_872 ();
 FILLCELL_X1 FILLER_1_884 ();
 FILLCELL_X1 FILLER_1_906 ();
 FILLCELL_X2 FILLER_1_936 ();
 FILLCELL_X1 FILLER_1_967 ();
 FILLCELL_X2 FILLER_1_993 ();
 FILLCELL_X1 FILLER_1_995 ();
 FILLCELL_X8 FILLER_1_1003 ();
 FILLCELL_X4 FILLER_1_1011 ();
 FILLCELL_X1 FILLER_1_1015 ();
 FILLCELL_X16 FILLER_1_1019 ();
 FILLCELL_X2 FILLER_1_1035 ();
 FILLCELL_X1 FILLER_1_1037 ();
 FILLCELL_X32 FILLER_1_1065 ();
 FILLCELL_X32 FILLER_1_1097 ();
 FILLCELL_X32 FILLER_1_1129 ();
 FILLCELL_X32 FILLER_1_1161 ();
 FILLCELL_X32 FILLER_1_1193 ();
 FILLCELL_X32 FILLER_1_1225 ();
 FILLCELL_X2 FILLER_1_1257 ();
 FILLCELL_X1 FILLER_1_1259 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X16 FILLER_2_449 ();
 FILLCELL_X4 FILLER_2_465 ();
 FILLCELL_X2 FILLER_2_518 ();
 FILLCELL_X2 FILLER_2_544 ();
 FILLCELL_X1 FILLER_2_546 ();
 FILLCELL_X4 FILLER_2_569 ();
 FILLCELL_X2 FILLER_2_573 ();
 FILLCELL_X8 FILLER_2_595 ();
 FILLCELL_X2 FILLER_2_603 ();
 FILLCELL_X1 FILLER_2_605 ();
 FILLCELL_X8 FILLER_2_610 ();
 FILLCELL_X4 FILLER_2_618 ();
 FILLCELL_X1 FILLER_2_622 ();
 FILLCELL_X16 FILLER_2_659 ();
 FILLCELL_X8 FILLER_2_695 ();
 FILLCELL_X4 FILLER_2_703 ();
 FILLCELL_X1 FILLER_2_707 ();
 FILLCELL_X2 FILLER_2_714 ();
 FILLCELL_X16 FILLER_2_738 ();
 FILLCELL_X2 FILLER_2_754 ();
 FILLCELL_X2 FILLER_2_760 ();
 FILLCELL_X1 FILLER_2_762 ();
 FILLCELL_X2 FILLER_2_772 ();
 FILLCELL_X1 FILLER_2_774 ();
 FILLCELL_X2 FILLER_2_780 ();
 FILLCELL_X4 FILLER_2_800 ();
 FILLCELL_X1 FILLER_2_804 ();
 FILLCELL_X1 FILLER_2_871 ();
 FILLCELL_X1 FILLER_2_877 ();
 FILLCELL_X1 FILLER_2_888 ();
 FILLCELL_X2 FILLER_2_913 ();
 FILLCELL_X1 FILLER_2_928 ();
 FILLCELL_X4 FILLER_2_946 ();
 FILLCELL_X1 FILLER_2_959 ();
 FILLCELL_X2 FILLER_2_973 ();
 FILLCELL_X1 FILLER_2_975 ();
 FILLCELL_X2 FILLER_2_1032 ();
 FILLCELL_X4 FILLER_2_1039 ();
 FILLCELL_X1 FILLER_2_1043 ();
 FILLCELL_X8 FILLER_2_1051 ();
 FILLCELL_X4 FILLER_2_1059 ();
 FILLCELL_X32 FILLER_2_1070 ();
 FILLCELL_X32 FILLER_2_1102 ();
 FILLCELL_X32 FILLER_2_1134 ();
 FILLCELL_X32 FILLER_2_1166 ();
 FILLCELL_X32 FILLER_2_1198 ();
 FILLCELL_X16 FILLER_2_1230 ();
 FILLCELL_X8 FILLER_2_1246 ();
 FILLCELL_X4 FILLER_2_1254 ();
 FILLCELL_X2 FILLER_2_1258 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X4 FILLER_3_481 ();
 FILLCELL_X2 FILLER_3_485 ();
 FILLCELL_X2 FILLER_3_491 ();
 FILLCELL_X2 FILLER_3_497 ();
 FILLCELL_X2 FILLER_3_510 ();
 FILLCELL_X2 FILLER_3_538 ();
 FILLCELL_X1 FILLER_3_540 ();
 FILLCELL_X8 FILLER_3_545 ();
 FILLCELL_X2 FILLER_3_553 ();
 FILLCELL_X2 FILLER_3_558 ();
 FILLCELL_X1 FILLER_3_560 ();
 FILLCELL_X4 FILLER_3_583 ();
 FILLCELL_X2 FILLER_3_587 ();
 FILLCELL_X4 FILLER_3_598 ();
 FILLCELL_X2 FILLER_3_606 ();
 FILLCELL_X1 FILLER_3_608 ();
 FILLCELL_X2 FILLER_3_613 ();
 FILLCELL_X2 FILLER_3_630 ();
 FILLCELL_X1 FILLER_3_644 ();
 FILLCELL_X2 FILLER_3_652 ();
 FILLCELL_X1 FILLER_3_654 ();
 FILLCELL_X8 FILLER_3_672 ();
 FILLCELL_X2 FILLER_3_689 ();
 FILLCELL_X2 FILLER_3_696 ();
 FILLCELL_X1 FILLER_3_702 ();
 FILLCELL_X2 FILLER_3_707 ();
 FILLCELL_X2 FILLER_3_714 ();
 FILLCELL_X1 FILLER_3_731 ();
 FILLCELL_X1 FILLER_3_736 ();
 FILLCELL_X4 FILLER_3_740 ();
 FILLCELL_X2 FILLER_3_744 ();
 FILLCELL_X1 FILLER_3_748 ();
 FILLCELL_X2 FILLER_3_753 ();
 FILLCELL_X1 FILLER_3_768 ();
 FILLCELL_X4 FILLER_3_778 ();
 FILLCELL_X2 FILLER_3_782 ();
 FILLCELL_X4 FILLER_3_795 ();
 FILLCELL_X1 FILLER_3_799 ();
 FILLCELL_X16 FILLER_3_805 ();
 FILLCELL_X2 FILLER_3_821 ();
 FILLCELL_X1 FILLER_3_827 ();
 FILLCELL_X2 FILLER_3_832 ();
 FILLCELL_X8 FILLER_3_839 ();
 FILLCELL_X1 FILLER_3_852 ();
 FILLCELL_X2 FILLER_3_856 ();
 FILLCELL_X1 FILLER_3_858 ();
 FILLCELL_X1 FILLER_3_863 ();
 FILLCELL_X1 FILLER_3_868 ();
 FILLCELL_X2 FILLER_3_872 ();
 FILLCELL_X4 FILLER_3_899 ();
 FILLCELL_X8 FILLER_3_907 ();
 FILLCELL_X2 FILLER_3_915 ();
 FILLCELL_X1 FILLER_3_917 ();
 FILLCELL_X2 FILLER_3_920 ();
 FILLCELL_X1 FILLER_3_948 ();
 FILLCELL_X16 FILLER_3_1003 ();
 FILLCELL_X2 FILLER_3_1019 ();
 FILLCELL_X1 FILLER_3_1041 ();
 FILLCELL_X8 FILLER_3_1049 ();
 FILLCELL_X2 FILLER_3_1057 ();
 FILLCELL_X1 FILLER_3_1059 ();
 FILLCELL_X8 FILLER_3_1087 ();
 FILLCELL_X2 FILLER_3_1099 ();
 FILLCELL_X8 FILLER_3_1132 ();
 FILLCELL_X32 FILLER_3_1147 ();
 FILLCELL_X32 FILLER_3_1179 ();
 FILLCELL_X32 FILLER_3_1211 ();
 FILLCELL_X16 FILLER_3_1243 ();
 FILLCELL_X1 FILLER_3_1259 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X16 FILLER_4_65 ();
 FILLCELL_X1 FILLER_4_81 ();
 FILLCELL_X32 FILLER_4_89 ();
 FILLCELL_X32 FILLER_4_121 ();
 FILLCELL_X32 FILLER_4_153 ();
 FILLCELL_X32 FILLER_4_185 ();
 FILLCELL_X32 FILLER_4_217 ();
 FILLCELL_X32 FILLER_4_249 ();
 FILLCELL_X32 FILLER_4_281 ();
 FILLCELL_X32 FILLER_4_313 ();
 FILLCELL_X32 FILLER_4_345 ();
 FILLCELL_X32 FILLER_4_377 ();
 FILLCELL_X32 FILLER_4_409 ();
 FILLCELL_X32 FILLER_4_441 ();
 FILLCELL_X4 FILLER_4_473 ();
 FILLCELL_X2 FILLER_4_477 ();
 FILLCELL_X2 FILLER_4_486 ();
 FILLCELL_X2 FILLER_4_491 ();
 FILLCELL_X1 FILLER_4_493 ();
 FILLCELL_X1 FILLER_4_497 ();
 FILLCELL_X1 FILLER_4_505 ();
 FILLCELL_X2 FILLER_4_511 ();
 FILLCELL_X1 FILLER_4_513 ();
 FILLCELL_X1 FILLER_4_525 ();
 FILLCELL_X1 FILLER_4_534 ();
 FILLCELL_X2 FILLER_4_545 ();
 FILLCELL_X1 FILLER_4_547 ();
 FILLCELL_X2 FILLER_4_564 ();
 FILLCELL_X8 FILLER_4_575 ();
 FILLCELL_X2 FILLER_4_583 ();
 FILLCELL_X2 FILLER_4_595 ();
 FILLCELL_X1 FILLER_4_597 ();
 FILLCELL_X2 FILLER_4_607 ();
 FILLCELL_X1 FILLER_4_609 ();
 FILLCELL_X2 FILLER_4_628 ();
 FILLCELL_X1 FILLER_4_630 ();
 FILLCELL_X2 FILLER_4_640 ();
 FILLCELL_X1 FILLER_4_642 ();
 FILLCELL_X2 FILLER_4_665 ();
 FILLCELL_X1 FILLER_4_667 ();
 FILLCELL_X8 FILLER_4_685 ();
 FILLCELL_X4 FILLER_4_695 ();
 FILLCELL_X1 FILLER_4_702 ();
 FILLCELL_X2 FILLER_4_706 ();
 FILLCELL_X2 FILLER_4_713 ();
 FILLCELL_X4 FILLER_4_733 ();
 FILLCELL_X2 FILLER_4_737 ();
 FILLCELL_X1 FILLER_4_744 ();
 FILLCELL_X2 FILLER_4_752 ();
 FILLCELL_X1 FILLER_4_758 ();
 FILLCELL_X8 FILLER_4_775 ();
 FILLCELL_X2 FILLER_4_783 ();
 FILLCELL_X8 FILLER_4_811 ();
 FILLCELL_X2 FILLER_4_819 ();
 FILLCELL_X1 FILLER_4_821 ();
 FILLCELL_X2 FILLER_4_830 ();
 FILLCELL_X1 FILLER_4_832 ();
 FILLCELL_X2 FILLER_4_845 ();
 FILLCELL_X1 FILLER_4_852 ();
 FILLCELL_X2 FILLER_4_871 ();
 FILLCELL_X4 FILLER_4_877 ();
 FILLCELL_X2 FILLER_4_891 ();
 FILLCELL_X2 FILLER_4_896 ();
 FILLCELL_X1 FILLER_4_898 ();
 FILLCELL_X4 FILLER_4_919 ();
 FILLCELL_X2 FILLER_4_923 ();
 FILLCELL_X1 FILLER_4_925 ();
 FILLCELL_X1 FILLER_4_964 ();
 FILLCELL_X4 FILLER_4_968 ();
 FILLCELL_X2 FILLER_4_972 ();
 FILLCELL_X2 FILLER_4_1061 ();
 FILLCELL_X2 FILLER_4_1087 ();
 FILLCELL_X1 FILLER_4_1089 ();
 FILLCELL_X16 FILLER_4_1113 ();
 FILLCELL_X4 FILLER_4_1129 ();
 FILLCELL_X2 FILLER_4_1133 ();
 FILLCELL_X1 FILLER_4_1135 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X16 FILLER_4_1240 ();
 FILLCELL_X4 FILLER_4_1256 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X8 FILLER_5_449 ();
 FILLCELL_X4 FILLER_5_457 ();
 FILLCELL_X2 FILLER_5_461 ();
 FILLCELL_X1 FILLER_5_463 ();
 FILLCELL_X1 FILLER_5_488 ();
 FILLCELL_X4 FILLER_5_494 ();
 FILLCELL_X2 FILLER_5_498 ();
 FILLCELL_X1 FILLER_5_500 ();
 FILLCELL_X1 FILLER_5_511 ();
 FILLCELL_X1 FILLER_5_539 ();
 FILLCELL_X1 FILLER_5_544 ();
 FILLCELL_X1 FILLER_5_549 ();
 FILLCELL_X1 FILLER_5_562 ();
 FILLCELL_X4 FILLER_5_567 ();
 FILLCELL_X1 FILLER_5_598 ();
 FILLCELL_X1 FILLER_5_604 ();
 FILLCELL_X4 FILLER_5_614 ();
 FILLCELL_X2 FILLER_5_618 ();
 FILLCELL_X1 FILLER_5_623 ();
 FILLCELL_X1 FILLER_5_626 ();
 FILLCELL_X4 FILLER_5_645 ();
 FILLCELL_X2 FILLER_5_649 ();
 FILLCELL_X8 FILLER_5_664 ();
 FILLCELL_X4 FILLER_5_672 ();
 FILLCELL_X1 FILLER_5_676 ();
 FILLCELL_X1 FILLER_5_743 ();
 FILLCELL_X1 FILLER_5_750 ();
 FILLCELL_X1 FILLER_5_758 ();
 FILLCELL_X1 FILLER_5_779 ();
 FILLCELL_X1 FILLER_5_790 ();
 FILLCELL_X2 FILLER_5_828 ();
 FILLCELL_X1 FILLER_5_830 ();
 FILLCELL_X4 FILLER_5_835 ();
 FILLCELL_X2 FILLER_5_842 ();
 FILLCELL_X2 FILLER_5_847 ();
 FILLCELL_X1 FILLER_5_849 ();
 FILLCELL_X8 FILLER_5_860 ();
 FILLCELL_X1 FILLER_5_868 ();
 FILLCELL_X1 FILLER_5_877 ();
 FILLCELL_X1 FILLER_5_892 ();
 FILLCELL_X8 FILLER_5_900 ();
 FILLCELL_X1 FILLER_5_908 ();
 FILLCELL_X16 FILLER_5_913 ();
 FILLCELL_X2 FILLER_5_933 ();
 FILLCELL_X2 FILLER_5_966 ();
 FILLCELL_X1 FILLER_5_983 ();
 FILLCELL_X8 FILLER_5_996 ();
 FILLCELL_X4 FILLER_5_1004 ();
 FILLCELL_X2 FILLER_5_1008 ();
 FILLCELL_X1 FILLER_5_1010 ();
 FILLCELL_X1 FILLER_5_1015 ();
 FILLCELL_X16 FILLER_5_1024 ();
 FILLCELL_X4 FILLER_5_1040 ();
 FILLCELL_X2 FILLER_5_1044 ();
 FILLCELL_X2 FILLER_5_1051 ();
 FILLCELL_X1 FILLER_5_1053 ();
 FILLCELL_X1 FILLER_5_1071 ();
 FILLCELL_X2 FILLER_5_1110 ();
 FILLCELL_X1 FILLER_5_1112 ();
 FILLCELL_X2 FILLER_5_1117 ();
 FILLCELL_X1 FILLER_5_1119 ();
 FILLCELL_X1 FILLER_5_1140 ();
 FILLCELL_X4 FILLER_5_1145 ();
 FILLCELL_X2 FILLER_5_1149 ();
 FILLCELL_X2 FILLER_5_1164 ();
 FILLCELL_X32 FILLER_5_1169 ();
 FILLCELL_X32 FILLER_5_1201 ();
 FILLCELL_X16 FILLER_5_1233 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X2 FILLER_5_1257 ();
 FILLCELL_X1 FILLER_5_1259 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X4 FILLER_6_449 ();
 FILLCELL_X2 FILLER_6_453 ();
 FILLCELL_X1 FILLER_6_455 ();
 FILLCELL_X4 FILLER_6_476 ();
 FILLCELL_X2 FILLER_6_480 ();
 FILLCELL_X1 FILLER_6_482 ();
 FILLCELL_X4 FILLER_6_504 ();
 FILLCELL_X1 FILLER_6_508 ();
 FILLCELL_X2 FILLER_6_521 ();
 FILLCELL_X1 FILLER_6_528 ();
 FILLCELL_X1 FILLER_6_549 ();
 FILLCELL_X2 FILLER_6_555 ();
 FILLCELL_X1 FILLER_6_557 ();
 FILLCELL_X1 FILLER_6_582 ();
 FILLCELL_X2 FILLER_6_587 ();
 FILLCELL_X2 FILLER_6_593 ();
 FILLCELL_X1 FILLER_6_600 ();
 FILLCELL_X1 FILLER_6_605 ();
 FILLCELL_X1 FILLER_6_610 ();
 FILLCELL_X2 FILLER_6_615 ();
 FILLCELL_X1 FILLER_6_623 ();
 FILLCELL_X1 FILLER_6_626 ();
 FILLCELL_X1 FILLER_6_630 ();
 FILLCELL_X1 FILLER_6_632 ();
 FILLCELL_X4 FILLER_6_641 ();
 FILLCELL_X2 FILLER_6_645 ();
 FILLCELL_X1 FILLER_6_647 ();
 FILLCELL_X1 FILLER_6_682 ();
 FILLCELL_X8 FILLER_6_718 ();
 FILLCELL_X8 FILLER_6_740 ();
 FILLCELL_X8 FILLER_6_760 ();
 FILLCELL_X4 FILLER_6_768 ();
 FILLCELL_X1 FILLER_6_772 ();
 FILLCELL_X2 FILLER_6_782 ();
 FILLCELL_X1 FILLER_6_810 ();
 FILLCELL_X2 FILLER_6_814 ();
 FILLCELL_X1 FILLER_6_816 ();
 FILLCELL_X1 FILLER_6_823 ();
 FILLCELL_X1 FILLER_6_829 ();
 FILLCELL_X2 FILLER_6_843 ();
 FILLCELL_X2 FILLER_6_849 ();
 FILLCELL_X1 FILLER_6_865 ();
 FILLCELL_X1 FILLER_6_870 ();
 FILLCELL_X1 FILLER_6_876 ();
 FILLCELL_X1 FILLER_6_882 ();
 FILLCELL_X4 FILLER_6_903 ();
 FILLCELL_X2 FILLER_6_907 ();
 FILLCELL_X1 FILLER_6_909 ();
 FILLCELL_X4 FILLER_6_952 ();
 FILLCELL_X2 FILLER_6_967 ();
 FILLCELL_X4 FILLER_6_991 ();
 FILLCELL_X4 FILLER_6_1002 ();
 FILLCELL_X1 FILLER_6_1006 ();
 FILLCELL_X4 FILLER_6_1011 ();
 FILLCELL_X1 FILLER_6_1015 ();
 FILLCELL_X4 FILLER_6_1022 ();
 FILLCELL_X2 FILLER_6_1026 ();
 FILLCELL_X2 FILLER_6_1032 ();
 FILLCELL_X2 FILLER_6_1037 ();
 FILLCELL_X1 FILLER_6_1044 ();
 FILLCELL_X16 FILLER_6_1050 ();
 FILLCELL_X8 FILLER_6_1066 ();
 FILLCELL_X2 FILLER_6_1074 ();
 FILLCELL_X4 FILLER_6_1085 ();
 FILLCELL_X2 FILLER_6_1089 ();
 FILLCELL_X4 FILLER_6_1134 ();
 FILLCELL_X1 FILLER_6_1138 ();
 FILLCELL_X32 FILLER_6_1162 ();
 FILLCELL_X32 FILLER_6_1194 ();
 FILLCELL_X32 FILLER_6_1226 ();
 FILLCELL_X2 FILLER_6_1258 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X1 FILLER_7_5 ();
 FILLCELL_X2 FILLER_7_9 ();
 FILLCELL_X1 FILLER_7_11 ();
 FILLCELL_X1 FILLER_7_14 ();
 FILLCELL_X32 FILLER_7_20 ();
 FILLCELL_X32 FILLER_7_52 ();
 FILLCELL_X32 FILLER_7_84 ();
 FILLCELL_X32 FILLER_7_116 ();
 FILLCELL_X32 FILLER_7_148 ();
 FILLCELL_X32 FILLER_7_180 ();
 FILLCELL_X32 FILLER_7_212 ();
 FILLCELL_X32 FILLER_7_244 ();
 FILLCELL_X32 FILLER_7_276 ();
 FILLCELL_X32 FILLER_7_308 ();
 FILLCELL_X32 FILLER_7_340 ();
 FILLCELL_X32 FILLER_7_372 ();
 FILLCELL_X32 FILLER_7_404 ();
 FILLCELL_X16 FILLER_7_436 ();
 FILLCELL_X8 FILLER_7_452 ();
 FILLCELL_X4 FILLER_7_460 ();
 FILLCELL_X2 FILLER_7_464 ();
 FILLCELL_X1 FILLER_7_466 ();
 FILLCELL_X1 FILLER_7_493 ();
 FILLCELL_X4 FILLER_7_502 ();
 FILLCELL_X2 FILLER_7_506 ();
 FILLCELL_X1 FILLER_7_508 ();
 FILLCELL_X4 FILLER_7_523 ();
 FILLCELL_X2 FILLER_7_527 ();
 FILLCELL_X1 FILLER_7_529 ();
 FILLCELL_X2 FILLER_7_539 ();
 FILLCELL_X2 FILLER_7_545 ();
 FILLCELL_X1 FILLER_7_547 ();
 FILLCELL_X1 FILLER_7_556 ();
 FILLCELL_X1 FILLER_7_577 ();
 FILLCELL_X4 FILLER_7_580 ();
 FILLCELL_X2 FILLER_7_584 ();
 FILLCELL_X4 FILLER_7_599 ();
 FILLCELL_X1 FILLER_7_603 ();
 FILLCELL_X1 FILLER_7_628 ();
 FILLCELL_X1 FILLER_7_632 ();
 FILLCELL_X1 FILLER_7_641 ();
 FILLCELL_X8 FILLER_7_664 ();
 FILLCELL_X4 FILLER_7_672 ();
 FILLCELL_X1 FILLER_7_676 ();
 FILLCELL_X2 FILLER_7_694 ();
 FILLCELL_X4 FILLER_7_703 ();
 FILLCELL_X4 FILLER_7_714 ();
 FILLCELL_X1 FILLER_7_718 ();
 FILLCELL_X1 FILLER_7_722 ();
 FILLCELL_X1 FILLER_7_725 ();
 FILLCELL_X2 FILLER_7_761 ();
 FILLCELL_X1 FILLER_7_763 ();
 FILLCELL_X8 FILLER_7_773 ();
 FILLCELL_X1 FILLER_7_781 ();
 FILLCELL_X16 FILLER_7_791 ();
 FILLCELL_X4 FILLER_7_835 ();
 FILLCELL_X2 FILLER_7_839 ();
 FILLCELL_X1 FILLER_7_864 ();
 FILLCELL_X8 FILLER_7_869 ();
 FILLCELL_X4 FILLER_7_877 ();
 FILLCELL_X8 FILLER_7_918 ();
 FILLCELL_X2 FILLER_7_926 ();
 FILLCELL_X1 FILLER_7_928 ();
 FILLCELL_X8 FILLER_7_934 ();
 FILLCELL_X4 FILLER_7_942 ();
 FILLCELL_X2 FILLER_7_946 ();
 FILLCELL_X32 FILLER_7_955 ();
 FILLCELL_X4 FILLER_7_1047 ();
 FILLCELL_X1 FILLER_7_1051 ();
 FILLCELL_X4 FILLER_7_1079 ();
 FILLCELL_X4 FILLER_7_1103 ();
 FILLCELL_X2 FILLER_7_1107 ();
 FILLCELL_X1 FILLER_7_1109 ();
 FILLCELL_X4 FILLER_7_1120 ();
 FILLCELL_X1 FILLER_7_1124 ();
 FILLCELL_X1 FILLER_7_1129 ();
 FILLCELL_X1 FILLER_7_1135 ();
 FILLCELL_X1 FILLER_7_1140 ();
 FILLCELL_X2 FILLER_7_1157 ();
 FILLCELL_X32 FILLER_7_1183 ();
 FILLCELL_X32 FILLER_7_1215 ();
 FILLCELL_X8 FILLER_7_1247 ();
 FILLCELL_X4 FILLER_7_1255 ();
 FILLCELL_X1 FILLER_7_1259 ();
 FILLCELL_X1 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_5 ();
 FILLCELL_X1 FILLER_8_8 ();
 FILLCELL_X1 FILLER_8_12 ();
 FILLCELL_X8 FILLER_8_15 ();
 FILLCELL_X1 FILLER_8_23 ();
 FILLCELL_X4 FILLER_8_29 ();
 FILLCELL_X1 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_39 ();
 FILLCELL_X32 FILLER_8_71 ();
 FILLCELL_X32 FILLER_8_103 ();
 FILLCELL_X32 FILLER_8_135 ();
 FILLCELL_X32 FILLER_8_167 ();
 FILLCELL_X32 FILLER_8_199 ();
 FILLCELL_X32 FILLER_8_231 ();
 FILLCELL_X32 FILLER_8_263 ();
 FILLCELL_X32 FILLER_8_295 ();
 FILLCELL_X32 FILLER_8_327 ();
 FILLCELL_X32 FILLER_8_359 ();
 FILLCELL_X32 FILLER_8_391 ();
 FILLCELL_X32 FILLER_8_423 ();
 FILLCELL_X8 FILLER_8_455 ();
 FILLCELL_X1 FILLER_8_463 ();
 FILLCELL_X4 FILLER_8_486 ();
 FILLCELL_X2 FILLER_8_490 ();
 FILLCELL_X1 FILLER_8_492 ();
 FILLCELL_X2 FILLER_8_497 ();
 FILLCELL_X1 FILLER_8_499 ();
 FILLCELL_X8 FILLER_8_503 ();
 FILLCELL_X2 FILLER_8_511 ();
 FILLCELL_X1 FILLER_8_513 ();
 FILLCELL_X4 FILLER_8_522 ();
 FILLCELL_X2 FILLER_8_526 ();
 FILLCELL_X1 FILLER_8_528 ();
 FILLCELL_X8 FILLER_8_534 ();
 FILLCELL_X2 FILLER_8_542 ();
 FILLCELL_X1 FILLER_8_553 ();
 FILLCELL_X4 FILLER_8_556 ();
 FILLCELL_X1 FILLER_8_560 ();
 FILLCELL_X1 FILLER_8_565 ();
 FILLCELL_X1 FILLER_8_570 ();
 FILLCELL_X1 FILLER_8_575 ();
 FILLCELL_X1 FILLER_8_580 ();
 FILLCELL_X4 FILLER_8_583 ();
 FILLCELL_X2 FILLER_8_598 ();
 FILLCELL_X4 FILLER_8_603 ();
 FILLCELL_X1 FILLER_8_630 ();
 FILLCELL_X16 FILLER_8_638 ();
 FILLCELL_X8 FILLER_8_671 ();
 FILLCELL_X4 FILLER_8_679 ();
 FILLCELL_X1 FILLER_8_683 ();
 FILLCELL_X2 FILLER_8_693 ();
 FILLCELL_X2 FILLER_8_736 ();
 FILLCELL_X4 FILLER_8_748 ();
 FILLCELL_X1 FILLER_8_752 ();
 FILLCELL_X8 FILLER_8_760 ();
 FILLCELL_X2 FILLER_8_768 ();
 FILLCELL_X1 FILLER_8_770 ();
 FILLCELL_X4 FILLER_8_794 ();
 FILLCELL_X2 FILLER_8_802 ();
 FILLCELL_X1 FILLER_8_804 ();
 FILLCELL_X2 FILLER_8_812 ();
 FILLCELL_X8 FILLER_8_838 ();
 FILLCELL_X4 FILLER_8_846 ();
 FILLCELL_X2 FILLER_8_850 ();
 FILLCELL_X2 FILLER_8_883 ();
 FILLCELL_X2 FILLER_8_889 ();
 FILLCELL_X4 FILLER_8_939 ();
 FILLCELL_X4 FILLER_8_963 ();
 FILLCELL_X8 FILLER_8_987 ();
 FILLCELL_X4 FILLER_8_995 ();
 FILLCELL_X1 FILLER_8_1003 ();
 FILLCELL_X2 FILLER_8_1007 ();
 FILLCELL_X1 FILLER_8_1021 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X4 FILLER_8_1080 ();
 FILLCELL_X1 FILLER_8_1088 ();
 FILLCELL_X1 FILLER_8_1093 ();
 FILLCELL_X8 FILLER_8_1097 ();
 FILLCELL_X1 FILLER_8_1105 ();
 FILLCELL_X2 FILLER_8_1126 ();
 FILLCELL_X1 FILLER_8_1128 ();
 FILLCELL_X4 FILLER_8_1149 ();
 FILLCELL_X32 FILLER_8_1173 ();
 FILLCELL_X32 FILLER_8_1205 ();
 FILLCELL_X16 FILLER_8_1237 ();
 FILLCELL_X4 FILLER_8_1253 ();
 FILLCELL_X2 FILLER_8_1257 ();
 FILLCELL_X1 FILLER_8_1259 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X8 FILLER_9_449 ();
 FILLCELL_X4 FILLER_9_457 ();
 FILLCELL_X2 FILLER_9_461 ();
 FILLCELL_X1 FILLER_9_500 ();
 FILLCELL_X1 FILLER_9_508 ();
 FILLCELL_X16 FILLER_9_514 ();
 FILLCELL_X8 FILLER_9_530 ();
 FILLCELL_X4 FILLER_9_538 ();
 FILLCELL_X1 FILLER_9_542 ();
 FILLCELL_X4 FILLER_9_549 ();
 FILLCELL_X2 FILLER_9_553 ();
 FILLCELL_X1 FILLER_9_555 ();
 FILLCELL_X2 FILLER_9_560 ();
 FILLCELL_X1 FILLER_9_562 ();
 FILLCELL_X8 FILLER_9_612 ();
 FILLCELL_X2 FILLER_9_620 ();
 FILLCELL_X1 FILLER_9_622 ();
 FILLCELL_X8 FILLER_9_626 ();
 FILLCELL_X4 FILLER_9_634 ();
 FILLCELL_X8 FILLER_9_641 ();
 FILLCELL_X4 FILLER_9_649 ();
 FILLCELL_X2 FILLER_9_666 ();
 FILLCELL_X8 FILLER_9_711 ();
 FILLCELL_X4 FILLER_9_719 ();
 FILLCELL_X2 FILLER_9_725 ();
 FILLCELL_X1 FILLER_9_727 ();
 FILLCELL_X1 FILLER_9_735 ();
 FILLCELL_X1 FILLER_9_741 ();
 FILLCELL_X4 FILLER_9_779 ();
 FILLCELL_X1 FILLER_9_783 ();
 FILLCELL_X1 FILLER_9_799 ();
 FILLCELL_X2 FILLER_9_842 ();
 FILLCELL_X4 FILLER_9_855 ();
 FILLCELL_X2 FILLER_9_859 ();
 FILLCELL_X1 FILLER_9_861 ();
 FILLCELL_X8 FILLER_9_870 ();
 FILLCELL_X4 FILLER_9_878 ();
 FILLCELL_X2 FILLER_9_882 ();
 FILLCELL_X8 FILLER_9_887 ();
 FILLCELL_X1 FILLER_9_895 ();
 FILLCELL_X4 FILLER_9_903 ();
 FILLCELL_X1 FILLER_9_907 ();
 FILLCELL_X4 FILLER_9_928 ();
 FILLCELL_X1 FILLER_9_959 ();
 FILLCELL_X8 FILLER_9_963 ();
 FILLCELL_X4 FILLER_9_971 ();
 FILLCELL_X1 FILLER_9_982 ();
 FILLCELL_X1 FILLER_9_986 ();
 FILLCELL_X1 FILLER_9_990 ();
 FILLCELL_X2 FILLER_9_1031 ();
 FILLCELL_X1 FILLER_9_1033 ();
 FILLCELL_X2 FILLER_9_1037 ();
 FILLCELL_X32 FILLER_9_1047 ();
 FILLCELL_X1 FILLER_9_1079 ();
 FILLCELL_X8 FILLER_9_1100 ();
 FILLCELL_X2 FILLER_9_1108 ();
 FILLCELL_X1 FILLER_9_1110 ();
 FILLCELL_X16 FILLER_9_1118 ();
 FILLCELL_X2 FILLER_9_1134 ();
 FILLCELL_X2 FILLER_9_1140 ();
 FILLCELL_X1 FILLER_9_1142 ();
 FILLCELL_X4 FILLER_9_1146 ();
 FILLCELL_X1 FILLER_9_1150 ();
 FILLCELL_X1 FILLER_9_1156 ();
 FILLCELL_X1 FILLER_9_1161 ();
 FILLCELL_X32 FILLER_9_1169 ();
 FILLCELL_X32 FILLER_9_1201 ();
 FILLCELL_X16 FILLER_9_1233 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X2 FILLER_9_1257 ();
 FILLCELL_X1 FILLER_9_1259 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X4 FILLER_10_449 ();
 FILLCELL_X2 FILLER_10_463 ();
 FILLCELL_X1 FILLER_10_465 ();
 FILLCELL_X8 FILLER_10_474 ();
 FILLCELL_X1 FILLER_10_496 ();
 FILLCELL_X8 FILLER_10_522 ();
 FILLCELL_X2 FILLER_10_530 ();
 FILLCELL_X1 FILLER_10_532 ();
 FILLCELL_X8 FILLER_10_555 ();
 FILLCELL_X4 FILLER_10_563 ();
 FILLCELL_X1 FILLER_10_567 ();
 FILLCELL_X2 FILLER_10_571 ();
 FILLCELL_X2 FILLER_10_575 ();
 FILLCELL_X2 FILLER_10_581 ();
 FILLCELL_X8 FILLER_10_586 ();
 FILLCELL_X2 FILLER_10_594 ();
 FILLCELL_X1 FILLER_10_596 ();
 FILLCELL_X1 FILLER_10_600 ();
 FILLCELL_X4 FILLER_10_604 ();
 FILLCELL_X1 FILLER_10_608 ();
 FILLCELL_X2 FILLER_10_615 ();
 FILLCELL_X2 FILLER_10_626 ();
 FILLCELL_X2 FILLER_10_632 ();
 FILLCELL_X16 FILLER_10_645 ();
 FILLCELL_X4 FILLER_10_661 ();
 FILLCELL_X1 FILLER_10_691 ();
 FILLCELL_X2 FILLER_10_709 ();
 FILLCELL_X8 FILLER_10_720 ();
 FILLCELL_X2 FILLER_10_751 ();
 FILLCELL_X4 FILLER_10_758 ();
 FILLCELL_X1 FILLER_10_766 ();
 FILLCELL_X4 FILLER_10_773 ();
 FILLCELL_X1 FILLER_10_777 ();
 FILLCELL_X2 FILLER_10_786 ();
 FILLCELL_X4 FILLER_10_792 ();
 FILLCELL_X1 FILLER_10_796 ();
 FILLCELL_X4 FILLER_10_801 ();
 FILLCELL_X2 FILLER_10_805 ();
 FILLCELL_X2 FILLER_10_814 ();
 FILLCELL_X1 FILLER_10_816 ();
 FILLCELL_X2 FILLER_10_828 ();
 FILLCELL_X2 FILLER_10_856 ();
 FILLCELL_X2 FILLER_10_862 ();
 FILLCELL_X1 FILLER_10_868 ();
 FILLCELL_X8 FILLER_10_894 ();
 FILLCELL_X1 FILLER_10_909 ();
 FILLCELL_X4 FILLER_10_917 ();
 FILLCELL_X2 FILLER_10_921 ();
 FILLCELL_X4 FILLER_10_927 ();
 FILLCELL_X2 FILLER_10_935 ();
 FILLCELL_X4 FILLER_10_940 ();
 FILLCELL_X2 FILLER_10_944 ();
 FILLCELL_X1 FILLER_10_974 ();
 FILLCELL_X2 FILLER_10_1024 ();
 FILLCELL_X2 FILLER_10_1046 ();
 FILLCELL_X4 FILLER_10_1080 ();
 FILLCELL_X1 FILLER_10_1084 ();
 FILLCELL_X4 FILLER_10_1092 ();
 FILLCELL_X2 FILLER_10_1104 ();
 FILLCELL_X4 FILLER_10_1126 ();
 FILLCELL_X1 FILLER_10_1130 ();
 FILLCELL_X2 FILLER_10_1151 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X16 FILLER_10_1240 ();
 FILLCELL_X4 FILLER_10_1256 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X8 FILLER_11_449 ();
 FILLCELL_X1 FILLER_11_457 ();
 FILLCELL_X4 FILLER_11_480 ();
 FILLCELL_X1 FILLER_11_503 ();
 FILLCELL_X1 FILLER_11_506 ();
 FILLCELL_X4 FILLER_11_534 ();
 FILLCELL_X8 FILLER_11_543 ();
 FILLCELL_X2 FILLER_11_551 ();
 FILLCELL_X8 FILLER_11_558 ();
 FILLCELL_X2 FILLER_11_575 ();
 FILLCELL_X1 FILLER_11_577 ();
 FILLCELL_X4 FILLER_11_589 ();
 FILLCELL_X1 FILLER_11_593 ();
 FILLCELL_X2 FILLER_11_624 ();
 FILLCELL_X1 FILLER_11_630 ();
 FILLCELL_X8 FILLER_11_657 ();
 FILLCELL_X2 FILLER_11_665 ();
 FILLCELL_X1 FILLER_11_667 ();
 FILLCELL_X4 FILLER_11_681 ();
 FILLCELL_X2 FILLER_11_685 ();
 FILLCELL_X1 FILLER_11_687 ();
 FILLCELL_X4 FILLER_11_726 ();
 FILLCELL_X2 FILLER_11_734 ();
 FILLCELL_X8 FILLER_11_739 ();
 FILLCELL_X2 FILLER_11_747 ();
 FILLCELL_X1 FILLER_11_749 ();
 FILLCELL_X8 FILLER_11_759 ();
 FILLCELL_X1 FILLER_11_767 ();
 FILLCELL_X1 FILLER_11_776 ();
 FILLCELL_X1 FILLER_11_786 ();
 FILLCELL_X2 FILLER_11_805 ();
 FILLCELL_X1 FILLER_11_807 ();
 FILLCELL_X4 FILLER_11_815 ();
 FILLCELL_X1 FILLER_11_819 ();
 FILLCELL_X8 FILLER_11_829 ();
 FILLCELL_X8 FILLER_11_844 ();
 FILLCELL_X2 FILLER_11_856 ();
 FILLCELL_X1 FILLER_11_858 ();
 FILLCELL_X4 FILLER_11_870 ();
 FILLCELL_X1 FILLER_11_874 ();
 FILLCELL_X8 FILLER_11_879 ();
 FILLCELL_X8 FILLER_11_915 ();
 FILLCELL_X2 FILLER_11_923 ();
 FILLCELL_X1 FILLER_11_925 ();
 FILLCELL_X1 FILLER_11_946 ();
 FILLCELL_X16 FILLER_11_969 ();
 FILLCELL_X16 FILLER_11_990 ();
 FILLCELL_X4 FILLER_11_1006 ();
 FILLCELL_X1 FILLER_11_1010 ();
 FILLCELL_X2 FILLER_11_1018 ();
 FILLCELL_X1 FILLER_11_1064 ();
 FILLCELL_X1 FILLER_11_1069 ();
 FILLCELL_X1 FILLER_11_1077 ();
 FILLCELL_X16 FILLER_11_1112 ();
 FILLCELL_X8 FILLER_11_1135 ();
 FILLCELL_X4 FILLER_11_1143 ();
 FILLCELL_X2 FILLER_11_1149 ();
 FILLCELL_X1 FILLER_11_1151 ();
 FILLCELL_X4 FILLER_11_1157 ();
 FILLCELL_X2 FILLER_11_1161 ();
 FILLCELL_X32 FILLER_11_1194 ();
 FILLCELL_X32 FILLER_11_1226 ();
 FILLCELL_X2 FILLER_11_1258 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X4 FILLER_12_449 ();
 FILLCELL_X2 FILLER_12_453 ();
 FILLCELL_X8 FILLER_12_479 ();
 FILLCELL_X2 FILLER_12_493 ();
 FILLCELL_X1 FILLER_12_499 ();
 FILLCELL_X1 FILLER_12_503 ();
 FILLCELL_X2 FILLER_12_517 ();
 FILLCELL_X8 FILLER_12_533 ();
 FILLCELL_X2 FILLER_12_541 ();
 FILLCELL_X1 FILLER_12_543 ();
 FILLCELL_X4 FILLER_12_547 ();
 FILLCELL_X1 FILLER_12_551 ();
 FILLCELL_X4 FILLER_12_557 ();
 FILLCELL_X1 FILLER_12_609 ();
 FILLCELL_X1 FILLER_12_614 ();
 FILLCELL_X1 FILLER_12_619 ();
 FILLCELL_X1 FILLER_12_622 ();
 FILLCELL_X4 FILLER_12_635 ();
 FILLCELL_X2 FILLER_12_639 ();
 FILLCELL_X1 FILLER_12_641 ();
 FILLCELL_X8 FILLER_12_666 ();
 FILLCELL_X4 FILLER_12_679 ();
 FILLCELL_X2 FILLER_12_683 ();
 FILLCELL_X1 FILLER_12_685 ();
 FILLCELL_X2 FILLER_12_693 ();
 FILLCELL_X1 FILLER_12_730 ();
 FILLCELL_X1 FILLER_12_740 ();
 FILLCELL_X2 FILLER_12_745 ();
 FILLCELL_X1 FILLER_12_758 ();
 FILLCELL_X1 FILLER_12_783 ();
 FILLCELL_X2 FILLER_12_814 ();
 FILLCELL_X1 FILLER_12_823 ();
 FILLCELL_X4 FILLER_12_828 ();
 FILLCELL_X2 FILLER_12_841 ();
 FILLCELL_X1 FILLER_12_843 ();
 FILLCELL_X4 FILLER_12_905 ();
 FILLCELL_X1 FILLER_12_909 ();
 FILLCELL_X4 FILLER_12_950 ();
 FILLCELL_X2 FILLER_12_954 ();
 FILLCELL_X1 FILLER_12_956 ();
 FILLCELL_X8 FILLER_12_960 ();
 FILLCELL_X2 FILLER_12_968 ();
 FILLCELL_X1 FILLER_12_970 ();
 FILLCELL_X1 FILLER_12_978 ();
 FILLCELL_X4 FILLER_12_999 ();
 FILLCELL_X1 FILLER_12_1023 ();
 FILLCELL_X4 FILLER_12_1060 ();
 FILLCELL_X2 FILLER_12_1064 ();
 FILLCELL_X1 FILLER_12_1098 ();
 FILLCELL_X8 FILLER_12_1102 ();
 FILLCELL_X4 FILLER_12_1110 ();
 FILLCELL_X4 FILLER_12_1119 ();
 FILLCELL_X1 FILLER_12_1123 ();
 FILLCELL_X2 FILLER_12_1151 ();
 FILLCELL_X1 FILLER_12_1153 ();
 FILLCELL_X4 FILLER_12_1163 ();
 FILLCELL_X1 FILLER_12_1167 ();
 FILLCELL_X32 FILLER_12_1170 ();
 FILLCELL_X32 FILLER_12_1202 ();
 FILLCELL_X16 FILLER_12_1234 ();
 FILLCELL_X8 FILLER_12_1250 ();
 FILLCELL_X2 FILLER_12_1258 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X16 FILLER_13_449 ();
 FILLCELL_X1 FILLER_13_465 ();
 FILLCELL_X1 FILLER_13_486 ();
 FILLCELL_X1 FILLER_13_502 ();
 FILLCELL_X1 FILLER_13_507 ();
 FILLCELL_X1 FILLER_13_510 ();
 FILLCELL_X1 FILLER_13_519 ();
 FILLCELL_X2 FILLER_13_547 ();
 FILLCELL_X1 FILLER_13_549 ();
 FILLCELL_X2 FILLER_13_560 ();
 FILLCELL_X1 FILLER_13_562 ();
 FILLCELL_X4 FILLER_13_578 ();
 FILLCELL_X1 FILLER_13_582 ();
 FILLCELL_X4 FILLER_13_586 ();
 FILLCELL_X2 FILLER_13_614 ();
 FILLCELL_X1 FILLER_13_616 ();
 FILLCELL_X2 FILLER_13_625 ();
 FILLCELL_X1 FILLER_13_627 ();
 FILLCELL_X16 FILLER_13_632 ();
 FILLCELL_X8 FILLER_13_648 ();
 FILLCELL_X4 FILLER_13_656 ();
 FILLCELL_X2 FILLER_13_660 ();
 FILLCELL_X1 FILLER_13_662 ();
 FILLCELL_X8 FILLER_13_710 ();
 FILLCELL_X1 FILLER_13_718 ();
 FILLCELL_X4 FILLER_13_728 ();
 FILLCELL_X1 FILLER_13_741 ();
 FILLCELL_X4 FILLER_13_749 ();
 FILLCELL_X2 FILLER_13_753 ();
 FILLCELL_X4 FILLER_13_794 ();
 FILLCELL_X2 FILLER_13_817 ();
 FILLCELL_X8 FILLER_13_827 ();
 FILLCELL_X4 FILLER_13_835 ();
 FILLCELL_X8 FILLER_13_845 ();
 FILLCELL_X1 FILLER_13_853 ();
 FILLCELL_X4 FILLER_13_858 ();
 FILLCELL_X8 FILLER_13_870 ();
 FILLCELL_X4 FILLER_13_878 ();
 FILLCELL_X8 FILLER_13_889 ();
 FILLCELL_X1 FILLER_13_924 ();
 FILLCELL_X2 FILLER_13_929 ();
 FILLCELL_X1 FILLER_13_938 ();
 FILLCELL_X4 FILLER_13_942 ();
 FILLCELL_X2 FILLER_13_946 ();
 FILLCELL_X1 FILLER_13_955 ();
 FILLCELL_X8 FILLER_13_987 ();
 FILLCELL_X4 FILLER_13_995 ();
 FILLCELL_X2 FILLER_13_999 ();
 FILLCELL_X16 FILLER_13_1004 ();
 FILLCELL_X1 FILLER_13_1043 ();
 FILLCELL_X2 FILLER_13_1051 ();
 FILLCELL_X2 FILLER_13_1060 ();
 FILLCELL_X1 FILLER_13_1067 ();
 FILLCELL_X8 FILLER_13_1073 ();
 FILLCELL_X4 FILLER_13_1081 ();
 FILLCELL_X1 FILLER_13_1085 ();
 FILLCELL_X1 FILLER_13_1116 ();
 FILLCELL_X4 FILLER_13_1159 ();
 FILLCELL_X2 FILLER_13_1163 ();
 FILLCELL_X32 FILLER_13_1194 ();
 FILLCELL_X32 FILLER_13_1226 ();
 FILLCELL_X2 FILLER_13_1258 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X8 FILLER_14_449 ();
 FILLCELL_X4 FILLER_14_457 ();
 FILLCELL_X1 FILLER_14_461 ();
 FILLCELL_X4 FILLER_14_482 ();
 FILLCELL_X2 FILLER_14_490 ();
 FILLCELL_X8 FILLER_14_496 ();
 FILLCELL_X2 FILLER_14_504 ();
 FILLCELL_X1 FILLER_14_509 ();
 FILLCELL_X16 FILLER_14_513 ();
 FILLCELL_X2 FILLER_14_529 ();
 FILLCELL_X1 FILLER_14_531 ();
 FILLCELL_X2 FILLER_14_535 ();
 FILLCELL_X2 FILLER_14_540 ();
 FILLCELL_X2 FILLER_14_567 ();
 FILLCELL_X1 FILLER_14_571 ();
 FILLCELL_X1 FILLER_14_575 ();
 FILLCELL_X16 FILLER_14_579 ();
 FILLCELL_X2 FILLER_14_595 ();
 FILLCELL_X2 FILLER_14_606 ();
 FILLCELL_X4 FILLER_14_658 ();
 FILLCELL_X1 FILLER_14_662 ();
 FILLCELL_X8 FILLER_14_680 ();
 FILLCELL_X1 FILLER_14_688 ();
 FILLCELL_X8 FILLER_14_719 ();
 FILLCELL_X4 FILLER_14_727 ();
 FILLCELL_X1 FILLER_14_731 ();
 FILLCELL_X8 FILLER_14_768 ();
 FILLCELL_X2 FILLER_14_776 ();
 FILLCELL_X16 FILLER_14_781 ();
 FILLCELL_X2 FILLER_14_797 ();
 FILLCELL_X1 FILLER_14_799 ();
 FILLCELL_X1 FILLER_14_838 ();
 FILLCELL_X16 FILLER_14_887 ();
 FILLCELL_X2 FILLER_14_907 ();
 FILLCELL_X2 FILLER_14_917 ();
 FILLCELL_X1 FILLER_14_919 ();
 FILLCELL_X4 FILLER_14_940 ();
 FILLCELL_X1 FILLER_14_944 ();
 FILLCELL_X1 FILLER_14_965 ();
 FILLCELL_X8 FILLER_14_975 ();
 FILLCELL_X4 FILLER_14_983 ();
 FILLCELL_X2 FILLER_14_987 ();
 FILLCELL_X1 FILLER_14_989 ();
 FILLCELL_X4 FILLER_14_1027 ();
 FILLCELL_X2 FILLER_14_1031 ();
 FILLCELL_X4 FILLER_14_1062 ();
 FILLCELL_X2 FILLER_14_1070 ();
 FILLCELL_X4 FILLER_14_1079 ();
 FILLCELL_X2 FILLER_14_1083 ();
 FILLCELL_X1 FILLER_14_1085 ();
 FILLCELL_X16 FILLER_14_1096 ();
 FILLCELL_X2 FILLER_14_1119 ();
 FILLCELL_X1 FILLER_14_1121 ();
 FILLCELL_X8 FILLER_14_1129 ();
 FILLCELL_X2 FILLER_14_1137 ();
 FILLCELL_X4 FILLER_14_1149 ();
 FILLCELL_X1 FILLER_14_1153 ();
 FILLCELL_X1 FILLER_14_1161 ();
 FILLCELL_X32 FILLER_14_1194 ();
 FILLCELL_X32 FILLER_14_1226 ();
 FILLCELL_X2 FILLER_14_1258 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X1 FILLER_15_488 ();
 FILLCELL_X4 FILLER_15_515 ();
 FILLCELL_X4 FILLER_15_549 ();
 FILLCELL_X2 FILLER_15_553 ();
 FILLCELL_X2 FILLER_15_567 ();
 FILLCELL_X1 FILLER_15_569 ();
 FILLCELL_X1 FILLER_15_574 ();
 FILLCELL_X1 FILLER_15_578 ();
 FILLCELL_X2 FILLER_15_591 ();
 FILLCELL_X4 FILLER_15_610 ();
 FILLCELL_X4 FILLER_15_633 ();
 FILLCELL_X4 FILLER_15_640 ();
 FILLCELL_X1 FILLER_15_644 ();
 FILLCELL_X8 FILLER_15_650 ();
 FILLCELL_X1 FILLER_15_658 ();
 FILLCELL_X1 FILLER_15_693 ();
 FILLCELL_X4 FILLER_15_722 ();
 FILLCELL_X1 FILLER_15_726 ();
 FILLCELL_X16 FILLER_15_747 ();
 FILLCELL_X8 FILLER_15_763 ();
 FILLCELL_X4 FILLER_15_771 ();
 FILLCELL_X4 FILLER_15_788 ();
 FILLCELL_X2 FILLER_15_792 ();
 FILLCELL_X4 FILLER_15_811 ();
 FILLCELL_X8 FILLER_15_827 ();
 FILLCELL_X2 FILLER_15_835 ();
 FILLCELL_X8 FILLER_15_849 ();
 FILLCELL_X1 FILLER_15_857 ();
 FILLCELL_X2 FILLER_15_867 ();
 FILLCELL_X2 FILLER_15_882 ();
 FILLCELL_X1 FILLER_15_884 ();
 FILLCELL_X2 FILLER_15_905 ();
 FILLCELL_X4 FILLER_15_912 ();
 FILLCELL_X2 FILLER_15_920 ();
 FILLCELL_X4 FILLER_15_925 ();
 FILLCELL_X8 FILLER_15_933 ();
 FILLCELL_X16 FILLER_15_946 ();
 FILLCELL_X4 FILLER_15_971 ();
 FILLCELL_X2 FILLER_15_975 ();
 FILLCELL_X1 FILLER_15_977 ();
 FILLCELL_X4 FILLER_15_1007 ();
 FILLCELL_X2 FILLER_15_1011 ();
 FILLCELL_X2 FILLER_15_1023 ();
 FILLCELL_X2 FILLER_15_1044 ();
 FILLCELL_X1 FILLER_15_1046 ();
 FILLCELL_X2 FILLER_15_1054 ();
 FILLCELL_X1 FILLER_15_1086 ();
 FILLCELL_X8 FILLER_15_1118 ();
 FILLCELL_X2 FILLER_15_1140 ();
 FILLCELL_X4 FILLER_15_1145 ();
 FILLCELL_X2 FILLER_15_1149 ();
 FILLCELL_X4 FILLER_15_1168 ();
 FILLCELL_X2 FILLER_15_1172 ();
 FILLCELL_X32 FILLER_15_1198 ();
 FILLCELL_X16 FILLER_15_1230 ();
 FILLCELL_X8 FILLER_15_1246 ();
 FILLCELL_X4 FILLER_15_1254 ();
 FILLCELL_X2 FILLER_15_1258 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X16 FILLER_16_449 ();
 FILLCELL_X2 FILLER_16_465 ();
 FILLCELL_X2 FILLER_16_497 ();
 FILLCELL_X1 FILLER_16_504 ();
 FILLCELL_X4 FILLER_16_513 ();
 FILLCELL_X2 FILLER_16_534 ();
 FILLCELL_X4 FILLER_16_548 ();
 FILLCELL_X2 FILLER_16_552 ();
 FILLCELL_X1 FILLER_16_554 ();
 FILLCELL_X1 FILLER_16_558 ();
 FILLCELL_X2 FILLER_16_599 ();
 FILLCELL_X2 FILLER_16_623 ();
 FILLCELL_X1 FILLER_16_630 ();
 FILLCELL_X1 FILLER_16_661 ();
 FILLCELL_X2 FILLER_16_679 ();
 FILLCELL_X4 FILLER_16_690 ();
 FILLCELL_X1 FILLER_16_694 ();
 FILLCELL_X4 FILLER_16_704 ();
 FILLCELL_X1 FILLER_16_708 ();
 FILLCELL_X4 FILLER_16_713 ();
 FILLCELL_X2 FILLER_16_717 ();
 FILLCELL_X8 FILLER_16_732 ();
 FILLCELL_X1 FILLER_16_740 ();
 FILLCELL_X4 FILLER_16_774 ();
 FILLCELL_X16 FILLER_16_787 ();
 FILLCELL_X4 FILLER_16_807 ();
 FILLCELL_X2 FILLER_16_811 ();
 FILLCELL_X2 FILLER_16_820 ();
 FILLCELL_X1 FILLER_16_822 ();
 FILLCELL_X2 FILLER_16_847 ();
 FILLCELL_X1 FILLER_16_849 ();
 FILLCELL_X4 FILLER_16_855 ();
 FILLCELL_X2 FILLER_16_859 ();
 FILLCELL_X4 FILLER_16_868 ();
 FILLCELL_X2 FILLER_16_872 ();
 FILLCELL_X2 FILLER_16_895 ();
 FILLCELL_X1 FILLER_16_897 ();
 FILLCELL_X2 FILLER_16_905 ();
 FILLCELL_X4 FILLER_16_927 ();
 FILLCELL_X2 FILLER_16_953 ();
 FILLCELL_X4 FILLER_16_1006 ();
 FILLCELL_X1 FILLER_16_1015 ();
 FILLCELL_X1 FILLER_16_1025 ();
 FILLCELL_X2 FILLER_16_1029 ();
 FILLCELL_X1 FILLER_16_1053 ();
 FILLCELL_X4 FILLER_16_1061 ();
 FILLCELL_X2 FILLER_16_1065 ();
 FILLCELL_X1 FILLER_16_1067 ();
 FILLCELL_X2 FILLER_16_1071 ();
 FILLCELL_X1 FILLER_16_1073 ();
 FILLCELL_X2 FILLER_16_1081 ();
 FILLCELL_X2 FILLER_16_1092 ();
 FILLCELL_X2 FILLER_16_1103 ();
 FILLCELL_X4 FILLER_16_1112 ();
 FILLCELL_X2 FILLER_16_1116 ();
 FILLCELL_X8 FILLER_16_1125 ();
 FILLCELL_X1 FILLER_16_1133 ();
 FILLCELL_X1 FILLER_16_1141 ();
 FILLCELL_X2 FILLER_16_1146 ();
 FILLCELL_X1 FILLER_16_1162 ();
 FILLCELL_X1 FILLER_16_1166 ();
 FILLCELL_X1 FILLER_16_1171 ();
 FILLCELL_X1 FILLER_16_1192 ();
 FILLCELL_X32 FILLER_16_1196 ();
 FILLCELL_X32 FILLER_16_1228 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X16 FILLER_17_289 ();
 FILLCELL_X2 FILLER_17_305 ();
 FILLCELL_X32 FILLER_17_312 ();
 FILLCELL_X32 FILLER_17_344 ();
 FILLCELL_X32 FILLER_17_376 ();
 FILLCELL_X32 FILLER_17_408 ();
 FILLCELL_X16 FILLER_17_440 ();
 FILLCELL_X8 FILLER_17_456 ();
 FILLCELL_X4 FILLER_17_464 ();
 FILLCELL_X2 FILLER_17_468 ();
 FILLCELL_X1 FILLER_17_470 ();
 FILLCELL_X1 FILLER_17_475 ();
 FILLCELL_X1 FILLER_17_496 ();
 FILLCELL_X4 FILLER_17_520 ();
 FILLCELL_X1 FILLER_17_524 ();
 FILLCELL_X8 FILLER_17_532 ();
 FILLCELL_X1 FILLER_17_560 ();
 FILLCELL_X1 FILLER_17_569 ();
 FILLCELL_X1 FILLER_17_574 ();
 FILLCELL_X2 FILLER_17_579 ();
 FILLCELL_X1 FILLER_17_581 ();
 FILLCELL_X1 FILLER_17_588 ();
 FILLCELL_X4 FILLER_17_616 ();
 FILLCELL_X2 FILLER_17_620 ();
 FILLCELL_X16 FILLER_17_639 ();
 FILLCELL_X2 FILLER_17_660 ();
 FILLCELL_X8 FILLER_17_735 ();
 FILLCELL_X2 FILLER_17_743 ();
 FILLCELL_X1 FILLER_17_745 ();
 FILLCELL_X4 FILLER_17_748 ();
 FILLCELL_X2 FILLER_17_752 ();
 FILLCELL_X1 FILLER_17_754 ();
 FILLCELL_X1 FILLER_17_764 ();
 FILLCELL_X2 FILLER_17_774 ();
 FILLCELL_X2 FILLER_17_787 ();
 FILLCELL_X2 FILLER_17_800 ();
 FILLCELL_X8 FILLER_17_827 ();
 FILLCELL_X2 FILLER_17_835 ();
 FILLCELL_X2 FILLER_17_846 ();
 FILLCELL_X4 FILLER_17_868 ();
 FILLCELL_X2 FILLER_17_872 ();
 FILLCELL_X1 FILLER_17_874 ();
 FILLCELL_X4 FILLER_17_882 ();
 FILLCELL_X2 FILLER_17_886 ();
 FILLCELL_X16 FILLER_17_902 ();
 FILLCELL_X2 FILLER_17_922 ();
 FILLCELL_X8 FILLER_17_933 ();
 FILLCELL_X1 FILLER_17_946 ();
 FILLCELL_X4 FILLER_17_956 ();
 FILLCELL_X2 FILLER_17_960 ();
 FILLCELL_X4 FILLER_17_989 ();
 FILLCELL_X8 FILLER_17_1041 ();
 FILLCELL_X4 FILLER_17_1049 ();
 FILLCELL_X2 FILLER_17_1053 ();
 FILLCELL_X1 FILLER_17_1055 ();
 FILLCELL_X4 FILLER_17_1067 ();
 FILLCELL_X1 FILLER_17_1071 ();
 FILLCELL_X8 FILLER_17_1079 ();
 FILLCELL_X4 FILLER_17_1087 ();
 FILLCELL_X1 FILLER_17_1109 ();
 FILLCELL_X1 FILLER_17_1114 ();
 FILLCELL_X4 FILLER_17_1132 ();
 FILLCELL_X2 FILLER_17_1136 ();
 FILLCELL_X8 FILLER_17_1154 ();
 FILLCELL_X16 FILLER_17_1176 ();
 FILLCELL_X32 FILLER_17_1196 ();
 FILLCELL_X32 FILLER_17_1228 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X16 FILLER_18_385 ();
 FILLCELL_X8 FILLER_18_401 ();
 FILLCELL_X2 FILLER_18_409 ();
 FILLCELL_X32 FILLER_18_416 ();
 FILLCELL_X8 FILLER_18_448 ();
 FILLCELL_X4 FILLER_18_456 ();
 FILLCELL_X2 FILLER_18_460 ();
 FILLCELL_X1 FILLER_18_462 ();
 FILLCELL_X1 FILLER_18_485 ();
 FILLCELL_X1 FILLER_18_501 ();
 FILLCELL_X1 FILLER_18_505 ();
 FILLCELL_X1 FILLER_18_513 ();
 FILLCELL_X4 FILLER_18_552 ();
 FILLCELL_X2 FILLER_18_556 ();
 FILLCELL_X1 FILLER_18_558 ();
 FILLCELL_X2 FILLER_18_563 ();
 FILLCELL_X1 FILLER_18_565 ();
 FILLCELL_X16 FILLER_18_588 ();
 FILLCELL_X8 FILLER_18_604 ();
 FILLCELL_X2 FILLER_18_612 ();
 FILLCELL_X2 FILLER_18_632 ();
 FILLCELL_X1 FILLER_18_634 ();
 FILLCELL_X8 FILLER_18_676 ();
 FILLCELL_X2 FILLER_18_684 ();
 FILLCELL_X4 FILLER_18_703 ();
 FILLCELL_X2 FILLER_18_736 ();
 FILLCELL_X2 FILLER_18_757 ();
 FILLCELL_X1 FILLER_18_759 ();
 FILLCELL_X4 FILLER_18_771 ();
 FILLCELL_X2 FILLER_18_775 ();
 FILLCELL_X2 FILLER_18_788 ();
 FILLCELL_X1 FILLER_18_807 ();
 FILLCELL_X2 FILLER_18_815 ();
 FILLCELL_X1 FILLER_18_817 ();
 FILLCELL_X2 FILLER_18_825 ();
 FILLCELL_X1 FILLER_18_827 ();
 FILLCELL_X1 FILLER_18_841 ();
 FILLCELL_X2 FILLER_18_862 ();
 FILLCELL_X2 FILLER_18_868 ();
 FILLCELL_X8 FILLER_18_890 ();
 FILLCELL_X1 FILLER_18_898 ();
 FILLCELL_X2 FILLER_18_903 ();
 FILLCELL_X1 FILLER_18_905 ();
 FILLCELL_X4 FILLER_18_909 ();
 FILLCELL_X4 FILLER_18_936 ();
 FILLCELL_X2 FILLER_18_940 ();
 FILLCELL_X1 FILLER_18_942 ();
 FILLCELL_X2 FILLER_18_947 ();
 FILLCELL_X2 FILLER_18_958 ();
 FILLCELL_X1 FILLER_18_960 ();
 FILLCELL_X1 FILLER_18_972 ();
 FILLCELL_X8 FILLER_18_985 ();
 FILLCELL_X2 FILLER_18_993 ();
 FILLCELL_X1 FILLER_18_995 ();
 FILLCELL_X4 FILLER_18_999 ();
 FILLCELL_X2 FILLER_18_1003 ();
 FILLCELL_X1 FILLER_18_1005 ();
 FILLCELL_X4 FILLER_18_1018 ();
 FILLCELL_X1 FILLER_18_1022 ();
 FILLCELL_X2 FILLER_18_1030 ();
 FILLCELL_X1 FILLER_18_1032 ();
 FILLCELL_X2 FILLER_18_1038 ();
 FILLCELL_X4 FILLER_18_1081 ();
 FILLCELL_X1 FILLER_18_1085 ();
 FILLCELL_X8 FILLER_18_1095 ();
 FILLCELL_X4 FILLER_18_1103 ();
 FILLCELL_X1 FILLER_18_1107 ();
 FILLCELL_X16 FILLER_18_1114 ();
 FILLCELL_X1 FILLER_18_1130 ();
 FILLCELL_X1 FILLER_18_1152 ();
 FILLCELL_X2 FILLER_18_1160 ();
 FILLCELL_X2 FILLER_18_1169 ();
 FILLCELL_X2 FILLER_18_1191 ();
 FILLCELL_X32 FILLER_18_1213 ();
 FILLCELL_X8 FILLER_18_1245 ();
 FILLCELL_X4 FILLER_18_1253 ();
 FILLCELL_X2 FILLER_18_1257 ();
 FILLCELL_X1 FILLER_18_1259 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X8 FILLER_19_353 ();
 FILLCELL_X2 FILLER_19_361 ();
 FILLCELL_X4 FILLER_19_383 ();
 FILLCELL_X2 FILLER_19_387 ();
 FILLCELL_X1 FILLER_19_389 ();
 FILLCELL_X32 FILLER_19_394 ();
 FILLCELL_X16 FILLER_19_426 ();
 FILLCELL_X8 FILLER_19_442 ();
 FILLCELL_X2 FILLER_19_450 ();
 FILLCELL_X1 FILLER_19_452 ();
 FILLCELL_X8 FILLER_19_473 ();
 FILLCELL_X8 FILLER_19_485 ();
 FILLCELL_X2 FILLER_19_497 ();
 FILLCELL_X1 FILLER_19_499 ();
 FILLCELL_X4 FILLER_19_505 ();
 FILLCELL_X2 FILLER_19_509 ();
 FILLCELL_X1 FILLER_19_518 ();
 FILLCELL_X16 FILLER_19_526 ();
 FILLCELL_X4 FILLER_19_542 ();
 FILLCELL_X2 FILLER_19_546 ();
 FILLCELL_X4 FILLER_19_551 ();
 FILLCELL_X1 FILLER_19_555 ();
 FILLCELL_X1 FILLER_19_572 ();
 FILLCELL_X2 FILLER_19_577 ();
 FILLCELL_X1 FILLER_19_579 ();
 FILLCELL_X32 FILLER_19_586 ();
 FILLCELL_X1 FILLER_19_618 ();
 FILLCELL_X8 FILLER_19_628 ();
 FILLCELL_X4 FILLER_19_636 ();
 FILLCELL_X2 FILLER_19_640 ();
 FILLCELL_X1 FILLER_19_642 ();
 FILLCELL_X16 FILLER_19_651 ();
 FILLCELL_X8 FILLER_19_667 ();
 FILLCELL_X2 FILLER_19_675 ();
 FILLCELL_X1 FILLER_19_677 ();
 FILLCELL_X1 FILLER_19_683 ();
 FILLCELL_X1 FILLER_19_689 ();
 FILLCELL_X1 FILLER_19_714 ();
 FILLCELL_X8 FILLER_19_724 ();
 FILLCELL_X2 FILLER_19_732 ();
 FILLCELL_X4 FILLER_19_743 ();
 FILLCELL_X8 FILLER_19_750 ();
 FILLCELL_X1 FILLER_19_758 ();
 FILLCELL_X1 FILLER_19_765 ();
 FILLCELL_X1 FILLER_19_771 ();
 FILLCELL_X16 FILLER_19_779 ();
 FILLCELL_X1 FILLER_19_795 ();
 FILLCELL_X8 FILLER_19_807 ();
 FILLCELL_X4 FILLER_19_815 ();
 FILLCELL_X2 FILLER_19_819 ();
 FILLCELL_X1 FILLER_19_821 ();
 FILLCELL_X4 FILLER_19_831 ();
 FILLCELL_X2 FILLER_19_835 ();
 FILLCELL_X1 FILLER_19_837 ();
 FILLCELL_X4 FILLER_19_845 ();
 FILLCELL_X2 FILLER_19_849 ();
 FILLCELL_X32 FILLER_19_866 ();
 FILLCELL_X2 FILLER_19_898 ();
 FILLCELL_X2 FILLER_19_920 ();
 FILLCELL_X4 FILLER_19_960 ();
 FILLCELL_X1 FILLER_19_964 ();
 FILLCELL_X1 FILLER_19_982 ();
 FILLCELL_X2 FILLER_19_995 ();
 FILLCELL_X4 FILLER_19_1009 ();
 FILLCELL_X1 FILLER_19_1013 ();
 FILLCELL_X2 FILLER_19_1041 ();
 FILLCELL_X8 FILLER_19_1046 ();
 FILLCELL_X4 FILLER_19_1054 ();
 FILLCELL_X2 FILLER_19_1058 ();
 FILLCELL_X8 FILLER_19_1089 ();
 FILLCELL_X1 FILLER_19_1097 ();
 FILLCELL_X1 FILLER_19_1121 ();
 FILLCELL_X2 FILLER_19_1127 ();
 FILLCELL_X2 FILLER_19_1133 ();
 FILLCELL_X2 FILLER_19_1140 ();
 FILLCELL_X1 FILLER_19_1142 ();
 FILLCELL_X2 FILLER_19_1155 ();
 FILLCELL_X1 FILLER_19_1157 ();
 FILLCELL_X1 FILLER_19_1192 ();
 FILLCELL_X32 FILLER_19_1196 ();
 FILLCELL_X32 FILLER_19_1228 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X16 FILLER_20_353 ();
 FILLCELL_X2 FILLER_20_369 ();
 FILLCELL_X4 FILLER_20_375 ();
 FILLCELL_X1 FILLER_20_379 ();
 FILLCELL_X1 FILLER_20_392 ();
 FILLCELL_X32 FILLER_20_405 ();
 FILLCELL_X16 FILLER_20_437 ();
 FILLCELL_X8 FILLER_20_453 ();
 FILLCELL_X4 FILLER_20_461 ();
 FILLCELL_X1 FILLER_20_522 ();
 FILLCELL_X2 FILLER_20_527 ();
 FILLCELL_X1 FILLER_20_529 ();
 FILLCELL_X2 FILLER_20_542 ();
 FILLCELL_X1 FILLER_20_544 ();
 FILLCELL_X2 FILLER_20_548 ();
 FILLCELL_X1 FILLER_20_559 ();
 FILLCELL_X4 FILLER_20_567 ();
 FILLCELL_X2 FILLER_20_571 ();
 FILLCELL_X2 FILLER_20_595 ();
 FILLCELL_X2 FILLER_20_601 ();
 FILLCELL_X2 FILLER_20_612 ();
 FILLCELL_X8 FILLER_20_632 ();
 FILLCELL_X4 FILLER_20_640 ();
 FILLCELL_X2 FILLER_20_644 ();
 FILLCELL_X1 FILLER_20_646 ();
 FILLCELL_X1 FILLER_20_654 ();
 FILLCELL_X1 FILLER_20_681 ();
 FILLCELL_X4 FILLER_20_696 ();
 FILLCELL_X2 FILLER_20_700 ();
 FILLCELL_X2 FILLER_20_732 ();
 FILLCELL_X1 FILLER_20_734 ();
 FILLCELL_X2 FILLER_20_745 ();
 FILLCELL_X2 FILLER_20_750 ();
 FILLCELL_X1 FILLER_20_752 ();
 FILLCELL_X1 FILLER_20_760 ();
 FILLCELL_X2 FILLER_20_768 ();
 FILLCELL_X4 FILLER_20_792 ();
 FILLCELL_X2 FILLER_20_796 ();
 FILLCELL_X1 FILLER_20_798 ();
 FILLCELL_X8 FILLER_20_833 ();
 FILLCELL_X1 FILLER_20_841 ();
 FILLCELL_X1 FILLER_20_862 ();
 FILLCELL_X1 FILLER_20_866 ();
 FILLCELL_X1 FILLER_20_887 ();
 FILLCELL_X1 FILLER_20_906 ();
 FILLCELL_X8 FILLER_20_924 ();
 FILLCELL_X4 FILLER_20_932 ();
 FILLCELL_X1 FILLER_20_936 ();
 FILLCELL_X8 FILLER_20_965 ();
 FILLCELL_X1 FILLER_20_973 ();
 FILLCELL_X4 FILLER_20_978 ();
 FILLCELL_X2 FILLER_20_982 ();
 FILLCELL_X1 FILLER_20_1000 ();
 FILLCELL_X2 FILLER_20_1004 ();
 FILLCELL_X2 FILLER_20_1020 ();
 FILLCELL_X4 FILLER_20_1024 ();
 FILLCELL_X2 FILLER_20_1028 ();
 FILLCELL_X1 FILLER_20_1030 ();
 FILLCELL_X4 FILLER_20_1051 ();
 FILLCELL_X4 FILLER_20_1059 ();
 FILLCELL_X2 FILLER_20_1063 ();
 FILLCELL_X1 FILLER_20_1065 ();
 FILLCELL_X1 FILLER_20_1073 ();
 FILLCELL_X1 FILLER_20_1089 ();
 FILLCELL_X16 FILLER_20_1103 ();
 FILLCELL_X2 FILLER_20_1119 ();
 FILLCELL_X1 FILLER_20_1121 ();
 FILLCELL_X8 FILLER_20_1129 ();
 FILLCELL_X4 FILLER_20_1137 ();
 FILLCELL_X1 FILLER_20_1141 ();
 FILLCELL_X1 FILLER_20_1154 ();
 FILLCELL_X8 FILLER_20_1160 ();
 FILLCELL_X1 FILLER_20_1168 ();
 FILLCELL_X8 FILLER_20_1176 ();
 FILLCELL_X1 FILLER_20_1184 ();
 FILLCELL_X2 FILLER_20_1192 ();
 FILLCELL_X32 FILLER_20_1214 ();
 FILLCELL_X8 FILLER_20_1246 ();
 FILLCELL_X4 FILLER_20_1254 ();
 FILLCELL_X2 FILLER_20_1258 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X8 FILLER_21_289 ();
 FILLCELL_X4 FILLER_21_297 ();
 FILLCELL_X2 FILLER_21_301 ();
 FILLCELL_X16 FILLER_21_310 ();
 FILLCELL_X2 FILLER_21_326 ();
 FILLCELL_X1 FILLER_21_328 ();
 FILLCELL_X1 FILLER_21_336 ();
 FILLCELL_X8 FILLER_21_368 ();
 FILLCELL_X4 FILLER_21_376 ();
 FILLCELL_X1 FILLER_21_380 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X16 FILLER_21_417 ();
 FILLCELL_X16 FILLER_21_450 ();
 FILLCELL_X2 FILLER_21_466 ();
 FILLCELL_X1 FILLER_21_497 ();
 FILLCELL_X1 FILLER_21_507 ();
 FILLCELL_X4 FILLER_21_513 ();
 FILLCELL_X8 FILLER_21_521 ();
 FILLCELL_X1 FILLER_21_529 ();
 FILLCELL_X4 FILLER_21_544 ();
 FILLCELL_X2 FILLER_21_548 ();
 FILLCELL_X2 FILLER_21_554 ();
 FILLCELL_X1 FILLER_21_561 ();
 FILLCELL_X1 FILLER_21_570 ();
 FILLCELL_X1 FILLER_21_575 ();
 FILLCELL_X4 FILLER_21_583 ();
 FILLCELL_X8 FILLER_21_592 ();
 FILLCELL_X2 FILLER_21_600 ();
 FILLCELL_X8 FILLER_21_619 ();
 FILLCELL_X2 FILLER_21_627 ();
 FILLCELL_X4 FILLER_21_670 ();
 FILLCELL_X1 FILLER_21_691 ();
 FILLCELL_X4 FILLER_21_705 ();
 FILLCELL_X8 FILLER_21_736 ();
 FILLCELL_X1 FILLER_21_744 ();
 FILLCELL_X2 FILLER_21_762 ();
 FILLCELL_X8 FILLER_21_792 ();
 FILLCELL_X1 FILLER_21_800 ();
 FILLCELL_X4 FILLER_21_834 ();
 FILLCELL_X2 FILLER_21_838 ();
 FILLCELL_X1 FILLER_21_840 ();
 FILLCELL_X4 FILLER_21_854 ();
 FILLCELL_X4 FILLER_21_876 ();
 FILLCELL_X2 FILLER_21_880 ();
 FILLCELL_X8 FILLER_21_921 ();
 FILLCELL_X4 FILLER_21_929 ();
 FILLCELL_X2 FILLER_21_948 ();
 FILLCELL_X8 FILLER_21_970 ();
 FILLCELL_X4 FILLER_21_978 ();
 FILLCELL_X2 FILLER_21_982 ();
 FILLCELL_X2 FILLER_21_995 ();
 FILLCELL_X4 FILLER_21_1037 ();
 FILLCELL_X1 FILLER_21_1041 ();
 FILLCELL_X1 FILLER_21_1060 ();
 FILLCELL_X4 FILLER_21_1097 ();
 FILLCELL_X2 FILLER_21_1101 ();
 FILLCELL_X2 FILLER_21_1107 ();
 FILLCELL_X2 FILLER_21_1114 ();
 FILLCELL_X1 FILLER_21_1116 ();
 FILLCELL_X8 FILLER_21_1146 ();
 FILLCELL_X4 FILLER_21_1168 ();
 FILLCELL_X1 FILLER_21_1172 ();
 FILLCELL_X8 FILLER_21_1177 ();
 FILLCELL_X2 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1216 ();
 FILLCELL_X8 FILLER_21_1248 ();
 FILLCELL_X4 FILLER_21_1256 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X1 FILLER_22_257 ();
 FILLCELL_X8 FILLER_22_282 ();
 FILLCELL_X1 FILLER_22_290 ();
 FILLCELL_X4 FILLER_22_315 ();
 FILLCELL_X1 FILLER_22_319 ();
 FILLCELL_X2 FILLER_22_344 ();
 FILLCELL_X8 FILLER_22_353 ();
 FILLCELL_X16 FILLER_22_368 ();
 FILLCELL_X8 FILLER_22_384 ();
 FILLCELL_X2 FILLER_22_392 ();
 FILLCELL_X2 FILLER_22_401 ();
 FILLCELL_X1 FILLER_22_403 ();
 FILLCELL_X4 FILLER_22_428 ();
 FILLCELL_X2 FILLER_22_432 ();
 FILLCELL_X2 FILLER_22_441 ();
 FILLCELL_X16 FILLER_22_450 ();
 FILLCELL_X8 FILLER_22_466 ();
 FILLCELL_X2 FILLER_22_474 ();
 FILLCELL_X1 FILLER_22_476 ();
 FILLCELL_X4 FILLER_22_484 ();
 FILLCELL_X2 FILLER_22_488 ();
 FILLCELL_X1 FILLER_22_490 ();
 FILLCELL_X1 FILLER_22_501 ();
 FILLCELL_X1 FILLER_22_512 ();
 FILLCELL_X8 FILLER_22_527 ();
 FILLCELL_X4 FILLER_22_542 ();
 FILLCELL_X1 FILLER_22_550 ();
 FILLCELL_X1 FILLER_22_556 ();
 FILLCELL_X2 FILLER_22_560 ();
 FILLCELL_X2 FILLER_22_569 ();
 FILLCELL_X1 FILLER_22_571 ();
 FILLCELL_X8 FILLER_22_598 ();
 FILLCELL_X2 FILLER_22_606 ();
 FILLCELL_X1 FILLER_22_608 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X8 FILLER_22_636 ();
 FILLCELL_X4 FILLER_22_644 ();
 FILLCELL_X2 FILLER_22_648 ();
 FILLCELL_X1 FILLER_22_650 ();
 FILLCELL_X4 FILLER_22_660 ();
 FILLCELL_X1 FILLER_22_664 ();
 FILLCELL_X1 FILLER_22_714 ();
 FILLCELL_X2 FILLER_22_724 ();
 FILLCELL_X1 FILLER_22_726 ();
 FILLCELL_X16 FILLER_22_740 ();
 FILLCELL_X2 FILLER_22_780 ();
 FILLCELL_X8 FILLER_22_786 ();
 FILLCELL_X1 FILLER_22_794 ();
 FILLCELL_X16 FILLER_22_804 ();
 FILLCELL_X4 FILLER_22_820 ();
 FILLCELL_X8 FILLER_22_842 ();
 FILLCELL_X2 FILLER_22_850 ();
 FILLCELL_X1 FILLER_22_852 ();
 FILLCELL_X4 FILLER_22_857 ();
 FILLCELL_X2 FILLER_22_888 ();
 FILLCELL_X1 FILLER_22_890 ();
 FILLCELL_X1 FILLER_22_898 ();
 FILLCELL_X2 FILLER_22_903 ();
 FILLCELL_X2 FILLER_22_908 ();
 FILLCELL_X1 FILLER_22_915 ();
 FILLCELL_X8 FILLER_22_928 ();
 FILLCELL_X2 FILLER_22_936 ();
 FILLCELL_X1 FILLER_22_950 ();
 FILLCELL_X2 FILLER_22_958 ();
 FILLCELL_X2 FILLER_22_974 ();
 FILLCELL_X1 FILLER_22_976 ();
 FILLCELL_X8 FILLER_22_988 ();
 FILLCELL_X4 FILLER_22_999 ();
 FILLCELL_X8 FILLER_22_1035 ();
 FILLCELL_X4 FILLER_22_1043 ();
 FILLCELL_X1 FILLER_22_1067 ();
 FILLCELL_X8 FILLER_22_1071 ();
 FILLCELL_X2 FILLER_22_1079 ();
 FILLCELL_X1 FILLER_22_1081 ();
 FILLCELL_X1 FILLER_22_1085 ();
 FILLCELL_X8 FILLER_22_1107 ();
 FILLCELL_X1 FILLER_22_1115 ();
 FILLCELL_X1 FILLER_22_1120 ();
 FILLCELL_X1 FILLER_22_1124 ();
 FILLCELL_X2 FILLER_22_1130 ();
 FILLCELL_X2 FILLER_22_1152 ();
 FILLCELL_X2 FILLER_22_1174 ();
 FILLCELL_X8 FILLER_22_1179 ();
 FILLCELL_X2 FILLER_22_1187 ();
 FILLCELL_X1 FILLER_22_1189 ();
 FILLCELL_X4 FILLER_22_1193 ();
 FILLCELL_X32 FILLER_22_1200 ();
 FILLCELL_X16 FILLER_22_1232 ();
 FILLCELL_X8 FILLER_22_1248 ();
 FILLCELL_X4 FILLER_22_1256 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X16 FILLER_23_225 ();
 FILLCELL_X4 FILLER_23_241 ();
 FILLCELL_X2 FILLER_23_245 ();
 FILLCELL_X2 FILLER_23_278 ();
 FILLCELL_X1 FILLER_23_280 ();
 FILLCELL_X2 FILLER_23_319 ();
 FILLCELL_X1 FILLER_23_321 ();
 FILLCELL_X16 FILLER_23_364 ();
 FILLCELL_X4 FILLER_23_380 ();
 FILLCELL_X2 FILLER_23_384 ();
 FILLCELL_X1 FILLER_23_403 ();
 FILLCELL_X2 FILLER_23_428 ();
 FILLCELL_X8 FILLER_23_438 ();
 FILLCELL_X1 FILLER_23_446 ();
 FILLCELL_X16 FILLER_23_454 ();
 FILLCELL_X2 FILLER_23_470 ();
 FILLCELL_X1 FILLER_23_472 ();
 FILLCELL_X1 FILLER_23_495 ();
 FILLCELL_X1 FILLER_23_501 ();
 FILLCELL_X4 FILLER_23_504 ();
 FILLCELL_X2 FILLER_23_508 ();
 FILLCELL_X2 FILLER_23_519 ();
 FILLCELL_X1 FILLER_23_533 ();
 FILLCELL_X2 FILLER_23_559 ();
 FILLCELL_X2 FILLER_23_568 ();
 FILLCELL_X1 FILLER_23_574 ();
 FILLCELL_X16 FILLER_23_584 ();
 FILLCELL_X4 FILLER_23_600 ();
 FILLCELL_X2 FILLER_23_604 ();
 FILLCELL_X1 FILLER_23_606 ();
 FILLCELL_X2 FILLER_23_614 ();
 FILLCELL_X1 FILLER_23_616 ();
 FILLCELL_X2 FILLER_23_630 ();
 FILLCELL_X1 FILLER_23_642 ();
 FILLCELL_X1 FILLER_23_647 ();
 FILLCELL_X8 FILLER_23_652 ();
 FILLCELL_X1 FILLER_23_680 ();
 FILLCELL_X1 FILLER_23_698 ();
 FILLCELL_X1 FILLER_23_712 ();
 FILLCELL_X1 FILLER_23_722 ();
 FILLCELL_X8 FILLER_23_746 ();
 FILLCELL_X1 FILLER_23_754 ();
 FILLCELL_X1 FILLER_23_759 ();
 FILLCELL_X8 FILLER_23_768 ();
 FILLCELL_X4 FILLER_23_776 ();
 FILLCELL_X1 FILLER_23_780 ();
 FILLCELL_X4 FILLER_23_784 ();
 FILLCELL_X2 FILLER_23_788 ();
 FILLCELL_X1 FILLER_23_790 ();
 FILLCELL_X8 FILLER_23_806 ();
 FILLCELL_X4 FILLER_23_814 ();
 FILLCELL_X2 FILLER_23_818 ();
 FILLCELL_X8 FILLER_23_838 ();
 FILLCELL_X1 FILLER_23_882 ();
 FILLCELL_X8 FILLER_23_925 ();
 FILLCELL_X4 FILLER_23_933 ();
 FILLCELL_X2 FILLER_23_941 ();
 FILLCELL_X1 FILLER_23_943 ();
 FILLCELL_X2 FILLER_23_958 ();
 FILLCELL_X1 FILLER_23_980 ();
 FILLCELL_X16 FILLER_23_1001 ();
 FILLCELL_X8 FILLER_23_1017 ();
 FILLCELL_X2 FILLER_23_1025 ();
 FILLCELL_X1 FILLER_23_1027 ();
 FILLCELL_X4 FILLER_23_1053 ();
 FILLCELL_X1 FILLER_23_1057 ();
 FILLCELL_X2 FILLER_23_1072 ();
 FILLCELL_X16 FILLER_23_1085 ();
 FILLCELL_X8 FILLER_23_1101 ();
 FILLCELL_X4 FILLER_23_1109 ();
 FILLCELL_X4 FILLER_23_1147 ();
 FILLCELL_X8 FILLER_23_1158 ();
 FILLCELL_X4 FILLER_23_1166 ();
 FILLCELL_X8 FILLER_23_1190 ();
 FILLCELL_X1 FILLER_23_1198 ();
 FILLCELL_X2 FILLER_23_1206 ();
 FILLCELL_X16 FILLER_23_1230 ();
 FILLCELL_X8 FILLER_23_1246 ();
 FILLCELL_X4 FILLER_23_1254 ();
 FILLCELL_X2 FILLER_23_1258 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X16 FILLER_24_264 ();
 FILLCELL_X4 FILLER_24_297 ();
 FILLCELL_X2 FILLER_24_301 ();
 FILLCELL_X4 FILLER_24_320 ();
 FILLCELL_X2 FILLER_24_348 ();
 FILLCELL_X1 FILLER_24_350 ();
 FILLCELL_X4 FILLER_24_356 ();
 FILLCELL_X1 FILLER_24_360 ();
 FILLCELL_X4 FILLER_24_385 ();
 FILLCELL_X1 FILLER_24_394 ();
 FILLCELL_X1 FILLER_24_402 ();
 FILLCELL_X4 FILLER_24_410 ();
 FILLCELL_X2 FILLER_24_414 ();
 FILLCELL_X1 FILLER_24_416 ();
 FILLCELL_X1 FILLER_24_429 ();
 FILLCELL_X1 FILLER_24_447 ();
 FILLCELL_X2 FILLER_24_472 ();
 FILLCELL_X8 FILLER_24_481 ();
 FILLCELL_X1 FILLER_24_509 ();
 FILLCELL_X2 FILLER_24_517 ();
 FILLCELL_X2 FILLER_24_523 ();
 FILLCELL_X2 FILLER_24_533 ();
 FILLCELL_X1 FILLER_24_535 ();
 FILLCELL_X8 FILLER_24_543 ();
 FILLCELL_X4 FILLER_24_551 ();
 FILLCELL_X1 FILLER_24_555 ();
 FILLCELL_X1 FILLER_24_567 ();
 FILLCELL_X2 FILLER_24_572 ();
 FILLCELL_X1 FILLER_24_574 ();
 FILLCELL_X4 FILLER_24_582 ();
 FILLCELL_X2 FILLER_24_606 ();
 FILLCELL_X1 FILLER_24_608 ();
 FILLCELL_X1 FILLER_24_623 ();
 FILLCELL_X2 FILLER_24_628 ();
 FILLCELL_X1 FILLER_24_630 ();
 FILLCELL_X2 FILLER_24_638 ();
 FILLCELL_X1 FILLER_24_640 ();
 FILLCELL_X16 FILLER_24_646 ();
 FILLCELL_X2 FILLER_24_662 ();
 FILLCELL_X2 FILLER_24_683 ();
 FILLCELL_X2 FILLER_24_688 ();
 FILLCELL_X4 FILLER_24_699 ();
 FILLCELL_X4 FILLER_24_710 ();
 FILLCELL_X4 FILLER_24_727 ();
 FILLCELL_X1 FILLER_24_742 ();
 FILLCELL_X4 FILLER_24_748 ();
 FILLCELL_X2 FILLER_24_752 ();
 FILLCELL_X1 FILLER_24_754 ();
 FILLCELL_X1 FILLER_24_759 ();
 FILLCELL_X2 FILLER_24_787 ();
 FILLCELL_X16 FILLER_24_807 ();
 FILLCELL_X4 FILLER_24_825 ();
 FILLCELL_X2 FILLER_24_829 ();
 FILLCELL_X8 FILLER_24_903 ();
 FILLCELL_X1 FILLER_24_911 ();
 FILLCELL_X8 FILLER_24_921 ();
 FILLCELL_X1 FILLER_24_952 ();
 FILLCELL_X8 FILLER_24_957 ();
 FILLCELL_X2 FILLER_24_965 ();
 FILLCELL_X1 FILLER_24_967 ();
 FILLCELL_X2 FILLER_24_972 ();
 FILLCELL_X2 FILLER_24_977 ();
 FILLCELL_X1 FILLER_24_979 ();
 FILLCELL_X1 FILLER_24_984 ();
 FILLCELL_X4 FILLER_24_996 ();
 FILLCELL_X1 FILLER_24_1000 ();
 FILLCELL_X4 FILLER_24_1015 ();
 FILLCELL_X2 FILLER_24_1019 ();
 FILLCELL_X8 FILLER_24_1044 ();
 FILLCELL_X1 FILLER_24_1052 ();
 FILLCELL_X4 FILLER_24_1075 ();
 FILLCELL_X1 FILLER_24_1079 ();
 FILLCELL_X8 FILLER_24_1101 ();
 FILLCELL_X4 FILLER_24_1109 ();
 FILLCELL_X2 FILLER_24_1113 ();
 FILLCELL_X1 FILLER_24_1115 ();
 FILLCELL_X4 FILLER_24_1130 ();
 FILLCELL_X2 FILLER_24_1134 ();
 FILLCELL_X1 FILLER_24_1136 ();
 FILLCELL_X16 FILLER_24_1172 ();
 FILLCELL_X4 FILLER_24_1188 ();
 FILLCELL_X2 FILLER_24_1192 ();
 FILLCELL_X32 FILLER_24_1216 ();
 FILLCELL_X8 FILLER_24_1248 ();
 FILLCELL_X4 FILLER_24_1256 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X16 FILLER_25_225 ();
 FILLCELL_X1 FILLER_25_265 ();
 FILLCELL_X8 FILLER_25_280 ();
 FILLCELL_X1 FILLER_25_288 ();
 FILLCELL_X16 FILLER_25_320 ();
 FILLCELL_X1 FILLER_25_336 ();
 FILLCELL_X8 FILLER_25_344 ();
 FILLCELL_X2 FILLER_25_352 ();
 FILLCELL_X4 FILLER_25_368 ();
 FILLCELL_X16 FILLER_25_379 ();
 FILLCELL_X1 FILLER_25_395 ();
 FILLCELL_X2 FILLER_25_417 ();
 FILLCELL_X1 FILLER_25_419 ();
 FILLCELL_X1 FILLER_25_434 ();
 FILLCELL_X4 FILLER_25_456 ();
 FILLCELL_X2 FILLER_25_460 ();
 FILLCELL_X2 FILLER_25_479 ();
 FILLCELL_X8 FILLER_25_488 ();
 FILLCELL_X1 FILLER_25_496 ();
 FILLCELL_X4 FILLER_25_504 ();
 FILLCELL_X2 FILLER_25_508 ();
 FILLCELL_X1 FILLER_25_510 ();
 FILLCELL_X1 FILLER_25_535 ();
 FILLCELL_X4 FILLER_25_544 ();
 FILLCELL_X2 FILLER_25_548 ();
 FILLCELL_X1 FILLER_25_550 ();
 FILLCELL_X4 FILLER_25_562 ();
 FILLCELL_X2 FILLER_25_612 ();
 FILLCELL_X1 FILLER_25_681 ();
 FILLCELL_X4 FILLER_25_695 ();
 FILLCELL_X1 FILLER_25_704 ();
 FILLCELL_X1 FILLER_25_708 ();
 FILLCELL_X1 FILLER_25_715 ();
 FILLCELL_X1 FILLER_25_719 ();
 FILLCELL_X4 FILLER_25_722 ();
 FILLCELL_X2 FILLER_25_726 ();
 FILLCELL_X1 FILLER_25_728 ();
 FILLCELL_X4 FILLER_25_759 ();
 FILLCELL_X4 FILLER_25_766 ();
 FILLCELL_X2 FILLER_25_775 ();
 FILLCELL_X1 FILLER_25_777 ();
 FILLCELL_X8 FILLER_25_802 ();
 FILLCELL_X4 FILLER_25_824 ();
 FILLCELL_X1 FILLER_25_828 ();
 FILLCELL_X8 FILLER_25_838 ();
 FILLCELL_X8 FILLER_25_853 ();
 FILLCELL_X4 FILLER_25_861 ();
 FILLCELL_X2 FILLER_25_865 ();
 FILLCELL_X2 FILLER_25_870 ();
 FILLCELL_X1 FILLER_25_872 ();
 FILLCELL_X8 FILLER_25_880 ();
 FILLCELL_X4 FILLER_25_888 ();
 FILLCELL_X1 FILLER_25_892 ();
 FILLCELL_X4 FILLER_25_907 ();
 FILLCELL_X2 FILLER_25_911 ();
 FILLCELL_X8 FILLER_25_920 ();
 FILLCELL_X4 FILLER_25_928 ();
 FILLCELL_X1 FILLER_25_932 ();
 FILLCELL_X1 FILLER_25_950 ();
 FILLCELL_X1 FILLER_25_954 ();
 FILLCELL_X1 FILLER_25_975 ();
 FILLCELL_X2 FILLER_25_983 ();
 FILLCELL_X1 FILLER_25_988 ();
 FILLCELL_X2 FILLER_25_996 ();
 FILLCELL_X8 FILLER_25_1007 ();
 FILLCELL_X4 FILLER_25_1015 ();
 FILLCELL_X2 FILLER_25_1019 ();
 FILLCELL_X2 FILLER_25_1059 ();
 FILLCELL_X16 FILLER_25_1065 ();
 FILLCELL_X2 FILLER_25_1081 ();
 FILLCELL_X2 FILLER_25_1117 ();
 FILLCELL_X16 FILLER_25_1148 ();
 FILLCELL_X2 FILLER_25_1186 ();
 FILLCELL_X8 FILLER_25_1195 ();
 FILLCELL_X4 FILLER_25_1203 ();
 FILLCELL_X2 FILLER_25_1207 ();
 FILLCELL_X16 FILLER_25_1231 ();
 FILLCELL_X8 FILLER_25_1247 ();
 FILLCELL_X4 FILLER_25_1255 ();
 FILLCELL_X1 FILLER_25_1259 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X16 FILLER_26_193 ();
 FILLCELL_X8 FILLER_26_209 ();
 FILLCELL_X1 FILLER_26_217 ();
 FILLCELL_X2 FILLER_26_225 ();
 FILLCELL_X2 FILLER_26_253 ();
 FILLCELL_X1 FILLER_26_272 ();
 FILLCELL_X2 FILLER_26_297 ();
 FILLCELL_X1 FILLER_26_299 ();
 FILLCELL_X4 FILLER_26_307 ();
 FILLCELL_X2 FILLER_26_311 ();
 FILLCELL_X1 FILLER_26_313 ();
 FILLCELL_X4 FILLER_26_345 ();
 FILLCELL_X1 FILLER_26_349 ();
 FILLCELL_X2 FILLER_26_355 ();
 FILLCELL_X2 FILLER_26_360 ();
 FILLCELL_X16 FILLER_26_379 ();
 FILLCELL_X8 FILLER_26_395 ();
 FILLCELL_X4 FILLER_26_403 ();
 FILLCELL_X2 FILLER_26_407 ();
 FILLCELL_X1 FILLER_26_409 ();
 FILLCELL_X1 FILLER_26_427 ();
 FILLCELL_X2 FILLER_26_445 ();
 FILLCELL_X1 FILLER_26_447 ();
 FILLCELL_X4 FILLER_26_465 ();
 FILLCELL_X1 FILLER_26_469 ();
 FILLCELL_X1 FILLER_26_475 ();
 FILLCELL_X8 FILLER_26_500 ();
 FILLCELL_X2 FILLER_26_508 ();
 FILLCELL_X1 FILLER_26_510 ();
 FILLCELL_X2 FILLER_26_553 ();
 FILLCELL_X1 FILLER_26_555 ();
 FILLCELL_X8 FILLER_26_563 ();
 FILLCELL_X16 FILLER_26_575 ();
 FILLCELL_X8 FILLER_26_591 ();
 FILLCELL_X4 FILLER_26_599 ();
 FILLCELL_X1 FILLER_26_621 ();
 FILLCELL_X2 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X2 FILLER_26_632 ();
 FILLCELL_X1 FILLER_26_634 ();
 FILLCELL_X8 FILLER_26_645 ();
 FILLCELL_X1 FILLER_26_653 ();
 FILLCELL_X4 FILLER_26_658 ();
 FILLCELL_X2 FILLER_26_662 ();
 FILLCELL_X8 FILLER_26_666 ();
 FILLCELL_X8 FILLER_26_694 ();
 FILLCELL_X4 FILLER_26_702 ();
 FILLCELL_X1 FILLER_26_706 ();
 FILLCELL_X2 FILLER_26_718 ();
 FILLCELL_X16 FILLER_26_734 ();
 FILLCELL_X2 FILLER_26_750 ();
 FILLCELL_X1 FILLER_26_752 ();
 FILLCELL_X2 FILLER_26_761 ();
 FILLCELL_X2 FILLER_26_768 ();
 FILLCELL_X1 FILLER_26_770 ();
 FILLCELL_X2 FILLER_26_778 ();
 FILLCELL_X1 FILLER_26_780 ();
 FILLCELL_X2 FILLER_26_786 ();
 FILLCELL_X1 FILLER_26_788 ();
 FILLCELL_X8 FILLER_26_811 ();
 FILLCELL_X8 FILLER_26_841 ();
 FILLCELL_X2 FILLER_26_849 ();
 FILLCELL_X1 FILLER_26_851 ();
 FILLCELL_X4 FILLER_26_893 ();
 FILLCELL_X1 FILLER_26_897 ();
 FILLCELL_X8 FILLER_26_938 ();
 FILLCELL_X4 FILLER_26_962 ();
 FILLCELL_X2 FILLER_26_966 ();
 FILLCELL_X2 FILLER_26_974 ();
 FILLCELL_X1 FILLER_26_976 ();
 FILLCELL_X2 FILLER_26_984 ();
 FILLCELL_X4 FILLER_26_990 ();
 FILLCELL_X2 FILLER_26_1008 ();
 FILLCELL_X2 FILLER_26_1030 ();
 FILLCELL_X8 FILLER_26_1039 ();
 FILLCELL_X2 FILLER_26_1061 ();
 FILLCELL_X1 FILLER_26_1063 ();
 FILLCELL_X2 FILLER_26_1091 ();
 FILLCELL_X1 FILLER_26_1093 ();
 FILLCELL_X16 FILLER_26_1116 ();
 FILLCELL_X8 FILLER_26_1134 ();
 FILLCELL_X4 FILLER_26_1142 ();
 FILLCELL_X2 FILLER_26_1146 ();
 FILLCELL_X1 FILLER_26_1168 ();
 FILLCELL_X8 FILLER_26_1195 ();
 FILLCELL_X1 FILLER_26_1203 ();
 FILLCELL_X8 FILLER_26_1211 ();
 FILLCELL_X1 FILLER_26_1219 ();
 FILLCELL_X8 FILLER_26_1247 ();
 FILLCELL_X4 FILLER_26_1255 ();
 FILLCELL_X1 FILLER_26_1259 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X8 FILLER_27_193 ();
 FILLCELL_X4 FILLER_27_201 ();
 FILLCELL_X1 FILLER_27_205 ();
 FILLCELL_X8 FILLER_27_230 ();
 FILLCELL_X1 FILLER_27_238 ();
 FILLCELL_X2 FILLER_27_268 ();
 FILLCELL_X8 FILLER_27_277 ();
 FILLCELL_X4 FILLER_27_285 ();
 FILLCELL_X8 FILLER_27_296 ();
 FILLCELL_X4 FILLER_27_314 ();
 FILLCELL_X2 FILLER_27_318 ();
 FILLCELL_X1 FILLER_27_320 ();
 FILLCELL_X4 FILLER_27_328 ();
 FILLCELL_X4 FILLER_27_346 ();
 FILLCELL_X2 FILLER_27_350 ();
 FILLCELL_X8 FILLER_27_371 ();
 FILLCELL_X16 FILLER_27_398 ();
 FILLCELL_X4 FILLER_27_414 ();
 FILLCELL_X2 FILLER_27_425 ();
 FILLCELL_X4 FILLER_27_434 ();
 FILLCELL_X1 FILLER_27_438 ();
 FILLCELL_X4 FILLER_27_446 ();
 FILLCELL_X1 FILLER_27_450 ();
 FILLCELL_X2 FILLER_27_458 ();
 FILLCELL_X1 FILLER_27_460 ();
 FILLCELL_X4 FILLER_27_468 ();
 FILLCELL_X16 FILLER_27_506 ();
 FILLCELL_X4 FILLER_27_522 ();
 FILLCELL_X2 FILLER_27_550 ();
 FILLCELL_X1 FILLER_27_552 ();
 FILLCELL_X4 FILLER_27_573 ();
 FILLCELL_X4 FILLER_27_599 ();
 FILLCELL_X1 FILLER_27_614 ();
 FILLCELL_X16 FILLER_27_643 ();
 FILLCELL_X2 FILLER_27_673 ();
 FILLCELL_X1 FILLER_27_675 ();
 FILLCELL_X4 FILLER_27_680 ();
 FILLCELL_X1 FILLER_27_684 ();
 FILLCELL_X2 FILLER_27_690 ();
 FILLCELL_X1 FILLER_27_696 ();
 FILLCELL_X2 FILLER_27_700 ();
 FILLCELL_X2 FILLER_27_704 ();
 FILLCELL_X2 FILLER_27_709 ();
 FILLCELL_X4 FILLER_27_724 ();
 FILLCELL_X1 FILLER_27_728 ();
 FILLCELL_X2 FILLER_27_735 ();
 FILLCELL_X4 FILLER_27_741 ();
 FILLCELL_X1 FILLER_27_745 ();
 FILLCELL_X2 FILLER_27_772 ();
 FILLCELL_X4 FILLER_27_788 ();
 FILLCELL_X16 FILLER_27_799 ();
 FILLCELL_X8 FILLER_27_815 ();
 FILLCELL_X2 FILLER_27_823 ();
 FILLCELL_X2 FILLER_27_855 ();
 FILLCELL_X1 FILLER_27_857 ();
 FILLCELL_X8 FILLER_27_861 ();
 FILLCELL_X4 FILLER_27_869 ();
 FILLCELL_X1 FILLER_27_873 ();
 FILLCELL_X16 FILLER_27_879 ();
 FILLCELL_X8 FILLER_27_895 ();
 FILLCELL_X4 FILLER_27_903 ();
 FILLCELL_X8 FILLER_27_914 ();
 FILLCELL_X1 FILLER_27_922 ();
 FILLCELL_X1 FILLER_27_925 ();
 FILLCELL_X1 FILLER_27_932 ();
 FILLCELL_X1 FILLER_27_953 ();
 FILLCELL_X1 FILLER_27_957 ();
 FILLCELL_X1 FILLER_27_1030 ();
 FILLCELL_X1 FILLER_27_1036 ();
 FILLCELL_X8 FILLER_27_1044 ();
 FILLCELL_X2 FILLER_27_1052 ();
 FILLCELL_X1 FILLER_27_1057 ();
 FILLCELL_X1 FILLER_27_1064 ();
 FILLCELL_X2 FILLER_27_1076 ();
 FILLCELL_X2 FILLER_27_1084 ();
 FILLCELL_X1 FILLER_27_1086 ();
 FILLCELL_X2 FILLER_27_1089 ();
 FILLCELL_X1 FILLER_27_1091 ();
 FILLCELL_X16 FILLER_27_1095 ();
 FILLCELL_X4 FILLER_27_1116 ();
 FILLCELL_X2 FILLER_27_1120 ();
 FILLCELL_X2 FILLER_27_1147 ();
 FILLCELL_X1 FILLER_27_1157 ();
 FILLCELL_X1 FILLER_27_1167 ();
 FILLCELL_X1 FILLER_27_1174 ();
 FILLCELL_X1 FILLER_27_1177 ();
 FILLCELL_X8 FILLER_27_1181 ();
 FILLCELL_X2 FILLER_27_1189 ();
 FILLCELL_X2 FILLER_27_1196 ();
 FILLCELL_X2 FILLER_27_1202 ();
 FILLCELL_X1 FILLER_27_1204 ();
 FILLCELL_X4 FILLER_27_1217 ();
 FILLCELL_X2 FILLER_27_1221 ();
 FILLCELL_X1 FILLER_27_1223 ();
 FILLCELL_X4 FILLER_27_1253 ();
 FILLCELL_X2 FILLER_27_1257 ();
 FILLCELL_X1 FILLER_27_1259 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X16 FILLER_28_193 ();
 FILLCELL_X2 FILLER_28_209 ();
 FILLCELL_X16 FILLER_28_235 ();
 FILLCELL_X2 FILLER_28_251 ();
 FILLCELL_X4 FILLER_28_267 ();
 FILLCELL_X1 FILLER_28_271 ();
 FILLCELL_X8 FILLER_28_279 ();
 FILLCELL_X1 FILLER_28_287 ();
 FILLCELL_X1 FILLER_28_325 ();
 FILLCELL_X2 FILLER_28_384 ();
 FILLCELL_X4 FILLER_28_393 ();
 FILLCELL_X1 FILLER_28_397 ();
 FILLCELL_X8 FILLER_28_405 ();
 FILLCELL_X1 FILLER_28_413 ();
 FILLCELL_X4 FILLER_28_447 ();
 FILLCELL_X1 FILLER_28_451 ();
 FILLCELL_X16 FILLER_28_515 ();
 FILLCELL_X8 FILLER_28_531 ();
 FILLCELL_X4 FILLER_28_539 ();
 FILLCELL_X2 FILLER_28_543 ();
 FILLCELL_X4 FILLER_28_569 ();
 FILLCELL_X1 FILLER_28_573 ();
 FILLCELL_X1 FILLER_28_594 ();
 FILLCELL_X2 FILLER_28_599 ();
 FILLCELL_X1 FILLER_28_601 ();
 FILLCELL_X1 FILLER_28_610 ();
 FILLCELL_X1 FILLER_28_614 ();
 FILLCELL_X2 FILLER_28_620 ();
 FILLCELL_X2 FILLER_28_678 ();
 FILLCELL_X1 FILLER_28_680 ();
 FILLCELL_X2 FILLER_28_683 ();
 FILLCELL_X1 FILLER_28_685 ();
 FILLCELL_X4 FILLER_28_689 ();
 FILLCELL_X1 FILLER_28_693 ();
 FILLCELL_X1 FILLER_28_704 ();
 FILLCELL_X2 FILLER_28_709 ();
 FILLCELL_X1 FILLER_28_711 ();
 FILLCELL_X2 FILLER_28_744 ();
 FILLCELL_X1 FILLER_28_757 ();
 FILLCELL_X2 FILLER_28_762 ();
 FILLCELL_X32 FILLER_28_773 ();
 FILLCELL_X4 FILLER_28_805 ();
 FILLCELL_X2 FILLER_28_809 ();
 FILLCELL_X1 FILLER_28_811 ();
 FILLCELL_X8 FILLER_28_832 ();
 FILLCELL_X1 FILLER_28_840 ();
 FILLCELL_X1 FILLER_28_878 ();
 FILLCELL_X2 FILLER_28_900 ();
 FILLCELL_X1 FILLER_28_902 ();
 FILLCELL_X4 FILLER_28_906 ();
 FILLCELL_X2 FILLER_28_910 ();
 FILLCELL_X16 FILLER_28_915 ();
 FILLCELL_X1 FILLER_28_931 ();
 FILLCELL_X4 FILLER_28_939 ();
 FILLCELL_X1 FILLER_28_943 ();
 FILLCELL_X1 FILLER_28_951 ();
 FILLCELL_X4 FILLER_28_965 ();
 FILLCELL_X1 FILLER_28_969 ();
 FILLCELL_X4 FILLER_28_978 ();
 FILLCELL_X8 FILLER_28_987 ();
 FILLCELL_X4 FILLER_28_995 ();
 FILLCELL_X8 FILLER_28_1006 ();
 FILLCELL_X16 FILLER_28_1023 ();
 FILLCELL_X2 FILLER_28_1039 ();
 FILLCELL_X1 FILLER_28_1041 ();
 FILLCELL_X1 FILLER_28_1046 ();
 FILLCELL_X1 FILLER_28_1052 ();
 FILLCELL_X4 FILLER_28_1081 ();
 FILLCELL_X1 FILLER_28_1085 ();
 FILLCELL_X2 FILLER_28_1124 ();
 FILLCELL_X2 FILLER_28_1146 ();
 FILLCELL_X1 FILLER_28_1148 ();
 FILLCELL_X1 FILLER_28_1152 ();
 FILLCELL_X1 FILLER_28_1160 ();
 FILLCELL_X1 FILLER_28_1168 ();
 FILLCELL_X2 FILLER_28_1172 ();
 FILLCELL_X2 FILLER_28_1182 ();
 FILLCELL_X1 FILLER_28_1184 ();
 FILLCELL_X2 FILLER_28_1199 ();
 FILLCELL_X2 FILLER_28_1228 ();
 FILLCELL_X16 FILLER_28_1235 ();
 FILLCELL_X8 FILLER_28_1251 ();
 FILLCELL_X1 FILLER_28_1259 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X16 FILLER_29_193 ();
 FILLCELL_X8 FILLER_29_209 ();
 FILLCELL_X4 FILLER_29_217 ();
 FILLCELL_X2 FILLER_29_252 ();
 FILLCELL_X4 FILLER_29_261 ();
 FILLCELL_X16 FILLER_29_282 ();
 FILLCELL_X2 FILLER_29_298 ();
 FILLCELL_X1 FILLER_29_300 ();
 FILLCELL_X4 FILLER_29_308 ();
 FILLCELL_X1 FILLER_29_334 ();
 FILLCELL_X1 FILLER_29_349 ();
 FILLCELL_X1 FILLER_29_357 ();
 FILLCELL_X1 FILLER_29_365 ();
 FILLCELL_X2 FILLER_29_373 ();
 FILLCELL_X16 FILLER_29_382 ();
 FILLCELL_X2 FILLER_29_402 ();
 FILLCELL_X2 FILLER_29_435 ();
 FILLCELL_X4 FILLER_29_454 ();
 FILLCELL_X2 FILLER_29_458 ();
 FILLCELL_X2 FILLER_29_467 ();
 FILLCELL_X8 FILLER_29_488 ();
 FILLCELL_X4 FILLER_29_496 ();
 FILLCELL_X2 FILLER_29_500 ();
 FILLCELL_X1 FILLER_29_502 ();
 FILLCELL_X16 FILLER_29_539 ();
 FILLCELL_X8 FILLER_29_575 ();
 FILLCELL_X4 FILLER_29_586 ();
 FILLCELL_X2 FILLER_29_590 ();
 FILLCELL_X1 FILLER_29_592 ();
 FILLCELL_X1 FILLER_29_611 ();
 FILLCELL_X1 FILLER_29_617 ();
 FILLCELL_X8 FILLER_29_640 ();
 FILLCELL_X2 FILLER_29_648 ();
 FILLCELL_X2 FILLER_29_652 ();
 FILLCELL_X4 FILLER_29_658 ();
 FILLCELL_X4 FILLER_29_666 ();
 FILLCELL_X1 FILLER_29_678 ();
 FILLCELL_X2 FILLER_29_713 ();
 FILLCELL_X2 FILLER_29_719 ();
 FILLCELL_X1 FILLER_29_721 ();
 FILLCELL_X2 FILLER_29_739 ();
 FILLCELL_X2 FILLER_29_746 ();
 FILLCELL_X1 FILLER_29_748 ();
 FILLCELL_X4 FILLER_29_752 ();
 FILLCELL_X8 FILLER_29_780 ();
 FILLCELL_X1 FILLER_29_788 ();
 FILLCELL_X4 FILLER_29_796 ();
 FILLCELL_X2 FILLER_29_800 ();
 FILLCELL_X1 FILLER_29_829 ();
 FILLCELL_X2 FILLER_29_837 ();
 FILLCELL_X1 FILLER_29_853 ();
 FILLCELL_X2 FILLER_29_862 ();
 FILLCELL_X4 FILLER_29_886 ();
 FILLCELL_X2 FILLER_29_890 ();
 FILLCELL_X8 FILLER_29_958 ();
 FILLCELL_X2 FILLER_29_966 ();
 FILLCELL_X1 FILLER_29_968 ();
 FILLCELL_X2 FILLER_29_976 ();
 FILLCELL_X1 FILLER_29_978 ();
 FILLCELL_X8 FILLER_29_1009 ();
 FILLCELL_X4 FILLER_29_1017 ();
 FILLCELL_X2 FILLER_29_1021 ();
 FILLCELL_X1 FILLER_29_1023 ();
 FILLCELL_X8 FILLER_29_1046 ();
 FILLCELL_X1 FILLER_29_1054 ();
 FILLCELL_X4 FILLER_29_1058 ();
 FILLCELL_X8 FILLER_29_1064 ();
 FILLCELL_X4 FILLER_29_1072 ();
 FILLCELL_X2 FILLER_29_1076 ();
 FILLCELL_X1 FILLER_29_1078 ();
 FILLCELL_X8 FILLER_29_1112 ();
 FILLCELL_X4 FILLER_29_1120 ();
 FILLCELL_X2 FILLER_29_1144 ();
 FILLCELL_X2 FILLER_29_1163 ();
 FILLCELL_X4 FILLER_29_1176 ();
 FILLCELL_X2 FILLER_29_1180 ();
 FILLCELL_X2 FILLER_29_1186 ();
 FILLCELL_X8 FILLER_29_1246 ();
 FILLCELL_X4 FILLER_29_1254 ();
 FILLCELL_X2 FILLER_29_1258 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X16 FILLER_30_193 ();
 FILLCELL_X4 FILLER_30_230 ();
 FILLCELL_X1 FILLER_30_234 ();
 FILLCELL_X4 FILLER_30_242 ();
 FILLCELL_X2 FILLER_30_263 ();
 FILLCELL_X2 FILLER_30_286 ();
 FILLCELL_X1 FILLER_30_288 ();
 FILLCELL_X2 FILLER_30_303 ();
 FILLCELL_X2 FILLER_30_314 ();
 FILLCELL_X2 FILLER_30_326 ();
 FILLCELL_X2 FILLER_30_347 ();
 FILLCELL_X4 FILLER_30_358 ();
 FILLCELL_X2 FILLER_30_379 ();
 FILLCELL_X2 FILLER_30_428 ();
 FILLCELL_X8 FILLER_30_437 ();
 FILLCELL_X2 FILLER_30_445 ();
 FILLCELL_X4 FILLER_30_461 ();
 FILLCELL_X2 FILLER_30_472 ();
 FILLCELL_X8 FILLER_30_480 ();
 FILLCELL_X2 FILLER_30_488 ();
 FILLCELL_X1 FILLER_30_490 ();
 FILLCELL_X4 FILLER_30_505 ();
 FILLCELL_X2 FILLER_30_509 ();
 FILLCELL_X1 FILLER_30_511 ();
 FILLCELL_X8 FILLER_30_514 ();
 FILLCELL_X4 FILLER_30_522 ();
 FILLCELL_X1 FILLER_30_526 ();
 FILLCELL_X2 FILLER_30_554 ();
 FILLCELL_X1 FILLER_30_611 ();
 FILLCELL_X2 FILLER_30_625 ();
 FILLCELL_X1 FILLER_30_627 ();
 FILLCELL_X4 FILLER_30_642 ();
 FILLCELL_X1 FILLER_30_651 ();
 FILLCELL_X2 FILLER_30_663 ();
 FILLCELL_X4 FILLER_30_670 ();
 FILLCELL_X1 FILLER_30_674 ();
 FILLCELL_X1 FILLER_30_694 ();
 FILLCELL_X4 FILLER_30_699 ();
 FILLCELL_X1 FILLER_30_703 ();
 FILLCELL_X1 FILLER_30_709 ();
 FILLCELL_X8 FILLER_30_713 ();
 FILLCELL_X4 FILLER_30_721 ();
 FILLCELL_X2 FILLER_30_740 ();
 FILLCELL_X4 FILLER_30_766 ();
 FILLCELL_X2 FILLER_30_770 ();
 FILLCELL_X1 FILLER_30_772 ();
 FILLCELL_X1 FILLER_30_785 ();
 FILLCELL_X1 FILLER_30_859 ();
 FILLCELL_X8 FILLER_30_863 ();
 FILLCELL_X2 FILLER_30_883 ();
 FILLCELL_X1 FILLER_30_885 ();
 FILLCELL_X2 FILLER_30_893 ();
 FILLCELL_X4 FILLER_30_921 ();
 FILLCELL_X2 FILLER_30_925 ();
 FILLCELL_X2 FILLER_30_935 ();
 FILLCELL_X1 FILLER_30_937 ();
 FILLCELL_X1 FILLER_30_984 ();
 FILLCELL_X2 FILLER_30_989 ();
 FILLCELL_X1 FILLER_30_991 ();
 FILLCELL_X1 FILLER_30_995 ();
 FILLCELL_X8 FILLER_30_1037 ();
 FILLCELL_X4 FILLER_30_1059 ();
 FILLCELL_X1 FILLER_30_1063 ();
 FILLCELL_X4 FILLER_30_1084 ();
 FILLCELL_X2 FILLER_30_1088 ();
 FILLCELL_X1 FILLER_30_1090 ();
 FILLCELL_X8 FILLER_30_1099 ();
 FILLCELL_X4 FILLER_30_1107 ();
 FILLCELL_X2 FILLER_30_1111 ();
 FILLCELL_X1 FILLER_30_1118 ();
 FILLCELL_X4 FILLER_30_1137 ();
 FILLCELL_X1 FILLER_30_1168 ();
 FILLCELL_X8 FILLER_30_1171 ();
 FILLCELL_X4 FILLER_30_1179 ();
 FILLCELL_X2 FILLER_30_1183 ();
 FILLCELL_X1 FILLER_30_1185 ();
 FILLCELL_X4 FILLER_30_1190 ();
 FILLCELL_X1 FILLER_30_1194 ();
 FILLCELL_X1 FILLER_30_1202 ();
 FILLCELL_X32 FILLER_30_1225 ();
 FILLCELL_X2 FILLER_30_1257 ();
 FILLCELL_X1 FILLER_30_1259 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X8 FILLER_31_193 ();
 FILLCELL_X4 FILLER_31_218 ();
 FILLCELL_X1 FILLER_31_222 ();
 FILLCELL_X16 FILLER_31_247 ();
 FILLCELL_X1 FILLER_31_263 ();
 FILLCELL_X4 FILLER_31_281 ();
 FILLCELL_X2 FILLER_31_285 ();
 FILLCELL_X2 FILLER_31_311 ();
 FILLCELL_X16 FILLER_31_357 ();
 FILLCELL_X2 FILLER_31_373 ();
 FILLCELL_X4 FILLER_31_392 ();
 FILLCELL_X2 FILLER_31_396 ();
 FILLCELL_X4 FILLER_31_419 ();
 FILLCELL_X8 FILLER_31_434 ();
 FILLCELL_X8 FILLER_31_466 ();
 FILLCELL_X2 FILLER_31_474 ();
 FILLCELL_X8 FILLER_31_487 ();
 FILLCELL_X2 FILLER_31_515 ();
 FILLCELL_X32 FILLER_31_522 ();
 FILLCELL_X8 FILLER_31_554 ();
 FILLCELL_X4 FILLER_31_562 ();
 FILLCELL_X2 FILLER_31_566 ();
 FILLCELL_X8 FILLER_31_576 ();
 FILLCELL_X4 FILLER_31_584 ();
 FILLCELL_X2 FILLER_31_588 ();
 FILLCELL_X1 FILLER_31_590 ();
 FILLCELL_X2 FILLER_31_595 ();
 FILLCELL_X8 FILLER_31_612 ();
 FILLCELL_X4 FILLER_31_620 ();
 FILLCELL_X2 FILLER_31_624 ();
 FILLCELL_X4 FILLER_31_635 ();
 FILLCELL_X2 FILLER_31_639 ();
 FILLCELL_X1 FILLER_31_641 ();
 FILLCELL_X2 FILLER_31_652 ();
 FILLCELL_X1 FILLER_31_663 ();
 FILLCELL_X1 FILLER_31_677 ();
 FILLCELL_X2 FILLER_31_703 ();
 FILLCELL_X8 FILLER_31_716 ();
 FILLCELL_X1 FILLER_31_724 ();
 FILLCELL_X2 FILLER_31_744 ();
 FILLCELL_X4 FILLER_31_768 ();
 FILLCELL_X2 FILLER_31_772 ();
 FILLCELL_X16 FILLER_31_787 ();
 FILLCELL_X8 FILLER_31_803 ();
 FILLCELL_X2 FILLER_31_811 ();
 FILLCELL_X4 FILLER_31_818 ();
 FILLCELL_X2 FILLER_31_827 ();
 FILLCELL_X8 FILLER_31_842 ();
 FILLCELL_X2 FILLER_31_850 ();
 FILLCELL_X2 FILLER_31_883 ();
 FILLCELL_X4 FILLER_31_901 ();
 FILLCELL_X2 FILLER_31_905 ();
 FILLCELL_X2 FILLER_31_916 ();
 FILLCELL_X1 FILLER_31_918 ();
 FILLCELL_X2 FILLER_31_924 ();
 FILLCELL_X2 FILLER_31_950 ();
 FILLCELL_X4 FILLER_31_963 ();
 FILLCELL_X2 FILLER_31_967 ();
 FILLCELL_X8 FILLER_31_973 ();
 FILLCELL_X4 FILLER_31_981 ();
 FILLCELL_X2 FILLER_31_995 ();
 FILLCELL_X1 FILLER_31_997 ();
 FILLCELL_X4 FILLER_31_1009 ();
 FILLCELL_X2 FILLER_31_1017 ();
 FILLCELL_X1 FILLER_31_1067 ();
 FILLCELL_X8 FILLER_31_1075 ();
 FILLCELL_X4 FILLER_31_1083 ();
 FILLCELL_X1 FILLER_31_1087 ();
 FILLCELL_X4 FILLER_31_1122 ();
 FILLCELL_X2 FILLER_31_1126 ();
 FILLCELL_X1 FILLER_31_1128 ();
 FILLCELL_X1 FILLER_31_1161 ();
 FILLCELL_X1 FILLER_31_1168 ();
 FILLCELL_X1 FILLER_31_1172 ();
 FILLCELL_X4 FILLER_31_1180 ();
 FILLCELL_X2 FILLER_31_1184 ();
 FILLCELL_X1 FILLER_31_1186 ();
 FILLCELL_X8 FILLER_31_1199 ();
 FILLCELL_X4 FILLER_31_1207 ();
 FILLCELL_X2 FILLER_31_1211 ();
 FILLCELL_X8 FILLER_31_1245 ();
 FILLCELL_X1 FILLER_31_1253 ();
 FILLCELL_X2 FILLER_31_1258 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X4 FILLER_32_193 ();
 FILLCELL_X1 FILLER_32_197 ();
 FILLCELL_X4 FILLER_32_215 ();
 FILLCELL_X2 FILLER_32_219 ();
 FILLCELL_X4 FILLER_32_267 ();
 FILLCELL_X16 FILLER_32_278 ();
 FILLCELL_X4 FILLER_32_294 ();
 FILLCELL_X1 FILLER_32_307 ();
 FILLCELL_X8 FILLER_32_325 ();
 FILLCELL_X4 FILLER_32_340 ();
 FILLCELL_X4 FILLER_32_360 ();
 FILLCELL_X2 FILLER_32_364 ();
 FILLCELL_X1 FILLER_32_399 ();
 FILLCELL_X2 FILLER_32_407 ();
 FILLCELL_X1 FILLER_32_409 ();
 FILLCELL_X4 FILLER_32_417 ();
 FILLCELL_X1 FILLER_32_421 ();
 FILLCELL_X2 FILLER_32_433 ();
 FILLCELL_X2 FILLER_32_444 ();
 FILLCELL_X1 FILLER_32_446 ();
 FILLCELL_X1 FILLER_32_451 ();
 FILLCELL_X2 FILLER_32_459 ();
 FILLCELL_X1 FILLER_32_461 ();
 FILLCELL_X2 FILLER_32_475 ();
 FILLCELL_X1 FILLER_32_489 ();
 FILLCELL_X2 FILLER_32_508 ();
 FILLCELL_X1 FILLER_32_510 ();
 FILLCELL_X1 FILLER_32_515 ();
 FILLCELL_X2 FILLER_32_523 ();
 FILLCELL_X1 FILLER_32_530 ();
 FILLCELL_X1 FILLER_32_535 ();
 FILLCELL_X1 FILLER_32_538 ();
 FILLCELL_X8 FILLER_32_543 ();
 FILLCELL_X4 FILLER_32_551 ();
 FILLCELL_X8 FILLER_32_562 ();
 FILLCELL_X2 FILLER_32_570 ();
 FILLCELL_X2 FILLER_32_594 ();
 FILLCELL_X2 FILLER_32_620 ();
 FILLCELL_X1 FILLER_32_622 ();
 FILLCELL_X1 FILLER_32_630 ();
 FILLCELL_X8 FILLER_32_632 ();
 FILLCELL_X2 FILLER_32_640 ();
 FILLCELL_X1 FILLER_32_642 ();
 FILLCELL_X8 FILLER_32_650 ();
 FILLCELL_X8 FILLER_32_671 ();
 FILLCELL_X2 FILLER_32_679 ();
 FILLCELL_X1 FILLER_32_681 ();
 FILLCELL_X16 FILLER_32_686 ();
 FILLCELL_X2 FILLER_32_702 ();
 FILLCELL_X4 FILLER_32_714 ();
 FILLCELL_X8 FILLER_32_732 ();
 FILLCELL_X4 FILLER_32_740 ();
 FILLCELL_X1 FILLER_32_744 ();
 FILLCELL_X8 FILLER_32_752 ();
 FILLCELL_X8 FILLER_32_767 ();
 FILLCELL_X1 FILLER_32_775 ();
 FILLCELL_X4 FILLER_32_792 ();
 FILLCELL_X2 FILLER_32_796 ();
 FILLCELL_X1 FILLER_32_798 ();
 FILLCELL_X1 FILLER_32_802 ();
 FILLCELL_X32 FILLER_32_851 ();
 FILLCELL_X2 FILLER_32_883 ();
 FILLCELL_X1 FILLER_32_885 ();
 FILLCELL_X16 FILLER_32_893 ();
 FILLCELL_X8 FILLER_32_909 ();
 FILLCELL_X2 FILLER_32_917 ();
 FILLCELL_X1 FILLER_32_919 ();
 FILLCELL_X4 FILLER_32_924 ();
 FILLCELL_X2 FILLER_32_928 ();
 FILLCELL_X1 FILLER_32_930 ();
 FILLCELL_X4 FILLER_32_974 ();
 FILLCELL_X8 FILLER_32_1002 ();
 FILLCELL_X4 FILLER_32_1010 ();
 FILLCELL_X2 FILLER_32_1014 ();
 FILLCELL_X1 FILLER_32_1046 ();
 FILLCELL_X1 FILLER_32_1069 ();
 FILLCELL_X8 FILLER_32_1094 ();
 FILLCELL_X2 FILLER_32_1102 ();
 FILLCELL_X1 FILLER_32_1104 ();
 FILLCELL_X2 FILLER_32_1132 ();
 FILLCELL_X1 FILLER_32_1156 ();
 FILLCELL_X4 FILLER_32_1168 ();
 FILLCELL_X2 FILLER_32_1172 ();
 FILLCELL_X1 FILLER_32_1196 ();
 FILLCELL_X1 FILLER_32_1217 ();
 FILLCELL_X4 FILLER_32_1221 ();
 FILLCELL_X2 FILLER_32_1225 ();
 FILLCELL_X1 FILLER_32_1227 ();
 FILLCELL_X16 FILLER_32_1235 ();
 FILLCELL_X4 FILLER_32_1251 ();
 FILLCELL_X2 FILLER_32_1255 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X8 FILLER_33_193 ();
 FILLCELL_X4 FILLER_33_201 ();
 FILLCELL_X2 FILLER_33_205 ();
 FILLCELL_X2 FILLER_33_224 ();
 FILLCELL_X1 FILLER_33_226 ();
 FILLCELL_X8 FILLER_33_241 ();
 FILLCELL_X2 FILLER_33_249 ();
 FILLCELL_X2 FILLER_33_272 ();
 FILLCELL_X1 FILLER_33_274 ();
 FILLCELL_X8 FILLER_33_299 ();
 FILLCELL_X16 FILLER_33_333 ();
 FILLCELL_X1 FILLER_33_349 ();
 FILLCELL_X8 FILLER_33_374 ();
 FILLCELL_X2 FILLER_33_389 ();
 FILLCELL_X1 FILLER_33_391 ();
 FILLCELL_X8 FILLER_33_399 ();
 FILLCELL_X1 FILLER_33_407 ();
 FILLCELL_X2 FILLER_33_412 ();
 FILLCELL_X1 FILLER_33_414 ();
 FILLCELL_X4 FILLER_33_424 ();
 FILLCELL_X2 FILLER_33_428 ();
 FILLCELL_X2 FILLER_33_443 ();
 FILLCELL_X1 FILLER_33_445 ();
 FILLCELL_X4 FILLER_33_453 ();
 FILLCELL_X2 FILLER_33_457 ();
 FILLCELL_X2 FILLER_33_479 ();
 FILLCELL_X1 FILLER_33_481 ();
 FILLCELL_X1 FILLER_33_487 ();
 FILLCELL_X2 FILLER_33_499 ();
 FILLCELL_X2 FILLER_33_505 ();
 FILLCELL_X1 FILLER_33_507 ();
 FILLCELL_X1 FILLER_33_511 ();
 FILLCELL_X1 FILLER_33_519 ();
 FILLCELL_X1 FILLER_33_527 ();
 FILLCELL_X2 FILLER_33_532 ();
 FILLCELL_X2 FILLER_33_541 ();
 FILLCELL_X1 FILLER_33_543 ();
 FILLCELL_X4 FILLER_33_564 ();
 FILLCELL_X1 FILLER_33_568 ();
 FILLCELL_X2 FILLER_33_589 ();
 FILLCELL_X4 FILLER_33_595 ();
 FILLCELL_X1 FILLER_33_599 ();
 FILLCELL_X16 FILLER_33_603 ();
 FILLCELL_X2 FILLER_33_619 ();
 FILLCELL_X1 FILLER_33_621 ();
 FILLCELL_X4 FILLER_33_636 ();
 FILLCELL_X2 FILLER_33_640 ();
 FILLCELL_X8 FILLER_33_656 ();
 FILLCELL_X8 FILLER_33_684 ();
 FILLCELL_X4 FILLER_33_716 ();
 FILLCELL_X2 FILLER_33_720 ();
 FILLCELL_X8 FILLER_33_744 ();
 FILLCELL_X8 FILLER_33_759 ();
 FILLCELL_X1 FILLER_33_767 ();
 FILLCELL_X1 FILLER_33_775 ();
 FILLCELL_X1 FILLER_33_786 ();
 FILLCELL_X1 FILLER_33_791 ();
 FILLCELL_X2 FILLER_33_799 ();
 FILLCELL_X8 FILLER_33_808 ();
 FILLCELL_X1 FILLER_33_824 ();
 FILLCELL_X2 FILLER_33_829 ();
 FILLCELL_X2 FILLER_33_837 ();
 FILLCELL_X4 FILLER_33_843 ();
 FILLCELL_X1 FILLER_33_847 ();
 FILLCELL_X2 FILLER_33_852 ();
 FILLCELL_X1 FILLER_33_854 ();
 FILLCELL_X4 FILLER_33_869 ();
 FILLCELL_X2 FILLER_33_873 ();
 FILLCELL_X1 FILLER_33_875 ();
 FILLCELL_X2 FILLER_33_879 ();
 FILLCELL_X1 FILLER_33_881 ();
 FILLCELL_X4 FILLER_33_889 ();
 FILLCELL_X2 FILLER_33_917 ();
 FILLCELL_X4 FILLER_33_953 ();
 FILLCELL_X4 FILLER_33_972 ();
 FILLCELL_X2 FILLER_33_976 ();
 FILLCELL_X4 FILLER_33_984 ();
 FILLCELL_X1 FILLER_33_988 ();
 FILLCELL_X8 FILLER_33_991 ();
 FILLCELL_X4 FILLER_33_999 ();
 FILLCELL_X2 FILLER_33_1003 ();
 FILLCELL_X2 FILLER_33_1078 ();
 FILLCELL_X4 FILLER_33_1085 ();
 FILLCELL_X1 FILLER_33_1089 ();
 FILLCELL_X2 FILLER_33_1101 ();
 FILLCELL_X16 FILLER_33_1119 ();
 FILLCELL_X1 FILLER_33_1135 ();
 FILLCELL_X4 FILLER_33_1141 ();
 FILLCELL_X1 FILLER_33_1145 ();
 FILLCELL_X4 FILLER_33_1154 ();
 FILLCELL_X4 FILLER_33_1169 ();
 FILLCELL_X4 FILLER_33_1182 ();
 FILLCELL_X2 FILLER_33_1186 ();
 FILLCELL_X4 FILLER_33_1197 ();
 FILLCELL_X2 FILLER_33_1201 ();
 FILLCELL_X2 FILLER_33_1210 ();
 FILLCELL_X1 FILLER_33_1234 ();
 FILLCELL_X4 FILLER_33_1255 ();
 FILLCELL_X1 FILLER_33_1259 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X16 FILLER_34_193 ();
 FILLCELL_X2 FILLER_34_209 ();
 FILLCELL_X1 FILLER_34_211 ();
 FILLCELL_X4 FILLER_34_226 ();
 FILLCELL_X2 FILLER_34_230 ();
 FILLCELL_X1 FILLER_34_232 ();
 FILLCELL_X1 FILLER_34_250 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X8 FILLER_34_321 ();
 FILLCELL_X4 FILLER_34_329 ();
 FILLCELL_X16 FILLER_34_357 ();
 FILLCELL_X4 FILLER_34_373 ();
 FILLCELL_X8 FILLER_34_394 ();
 FILLCELL_X1 FILLER_34_409 ();
 FILLCELL_X16 FILLER_34_423 ();
 FILLCELL_X8 FILLER_34_439 ();
 FILLCELL_X4 FILLER_34_447 ();
 FILLCELL_X2 FILLER_34_451 ();
 FILLCELL_X1 FILLER_34_453 ();
 FILLCELL_X4 FILLER_34_461 ();
 FILLCELL_X2 FILLER_34_465 ();
 FILLCELL_X1 FILLER_34_467 ();
 FILLCELL_X32 FILLER_34_486 ();
 FILLCELL_X4 FILLER_34_518 ();
 FILLCELL_X2 FILLER_34_522 ();
 FILLCELL_X4 FILLER_34_550 ();
 FILLCELL_X8 FILLER_34_557 ();
 FILLCELL_X4 FILLER_34_565 ();
 FILLCELL_X2 FILLER_34_589 ();
 FILLCELL_X8 FILLER_34_595 ();
 FILLCELL_X8 FILLER_34_607 ();
 FILLCELL_X2 FILLER_34_626 ();
 FILLCELL_X2 FILLER_34_632 ();
 FILLCELL_X8 FILLER_34_638 ();
 FILLCELL_X4 FILLER_34_646 ();
 FILLCELL_X1 FILLER_34_650 ();
 FILLCELL_X4 FILLER_34_656 ();
 FILLCELL_X2 FILLER_34_660 ();
 FILLCELL_X1 FILLER_34_662 ();
 FILLCELL_X8 FILLER_34_670 ();
 FILLCELL_X2 FILLER_34_678 ();
 FILLCELL_X1 FILLER_34_680 ();
 FILLCELL_X16 FILLER_34_691 ();
 FILLCELL_X1 FILLER_34_707 ();
 FILLCELL_X4 FILLER_34_726 ();
 FILLCELL_X1 FILLER_34_730 ();
 FILLCELL_X16 FILLER_34_740 ();
 FILLCELL_X2 FILLER_34_756 ();
 FILLCELL_X1 FILLER_34_758 ();
 FILLCELL_X4 FILLER_34_761 ();
 FILLCELL_X2 FILLER_34_765 ();
 FILLCELL_X1 FILLER_34_767 ();
 FILLCELL_X2 FILLER_34_782 ();
 FILLCELL_X1 FILLER_34_811 ();
 FILLCELL_X1 FILLER_34_815 ();
 FILLCELL_X1 FILLER_34_822 ();
 FILLCELL_X1 FILLER_34_830 ();
 FILLCELL_X8 FILLER_34_836 ();
 FILLCELL_X1 FILLER_34_844 ();
 FILLCELL_X1 FILLER_34_852 ();
 FILLCELL_X2 FILLER_34_862 ();
 FILLCELL_X1 FILLER_34_864 ();
 FILLCELL_X2 FILLER_34_889 ();
 FILLCELL_X8 FILLER_34_910 ();
 FILLCELL_X4 FILLER_34_918 ();
 FILLCELL_X1 FILLER_34_922 ();
 FILLCELL_X2 FILLER_34_930 ();
 FILLCELL_X8 FILLER_34_946 ();
 FILLCELL_X2 FILLER_34_954 ();
 FILLCELL_X1 FILLER_34_956 ();
 FILLCELL_X1 FILLER_34_964 ();
 FILLCELL_X4 FILLER_34_993 ();
 FILLCELL_X1 FILLER_34_997 ();
 FILLCELL_X8 FILLER_34_1003 ();
 FILLCELL_X4 FILLER_34_1011 ();
 FILLCELL_X2 FILLER_34_1015 ();
 FILLCELL_X1 FILLER_34_1017 ();
 FILLCELL_X1 FILLER_34_1029 ();
 FILLCELL_X2 FILLER_34_1042 ();
 FILLCELL_X1 FILLER_34_1044 ();
 FILLCELL_X8 FILLER_34_1048 ();
 FILLCELL_X2 FILLER_34_1056 ();
 FILLCELL_X4 FILLER_34_1116 ();
 FILLCELL_X1 FILLER_34_1120 ();
 FILLCELL_X2 FILLER_34_1124 ();
 FILLCELL_X1 FILLER_34_1126 ();
 FILLCELL_X4 FILLER_34_1161 ();
 FILLCELL_X2 FILLER_34_1165 ();
 FILLCELL_X8 FILLER_34_1173 ();
 FILLCELL_X1 FILLER_34_1181 ();
 FILLCELL_X2 FILLER_34_1233 ();
 FILLCELL_X1 FILLER_34_1235 ();
 FILLCELL_X4 FILLER_34_1239 ();
 FILLCELL_X1 FILLER_34_1243 ();
 FILLCELL_X8 FILLER_34_1249 ();
 FILLCELL_X2 FILLER_34_1257 ();
 FILLCELL_X1 FILLER_34_1259 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X4 FILLER_35_193 ();
 FILLCELL_X2 FILLER_35_197 ();
 FILLCELL_X4 FILLER_35_220 ();
 FILLCELL_X2 FILLER_35_224 ();
 FILLCELL_X1 FILLER_35_226 ();
 FILLCELL_X2 FILLER_35_234 ();
 FILLCELL_X1 FILLER_35_236 ();
 FILLCELL_X4 FILLER_35_244 ();
 FILLCELL_X2 FILLER_35_248 ();
 FILLCELL_X1 FILLER_35_260 ();
 FILLCELL_X4 FILLER_35_270 ();
 FILLCELL_X1 FILLER_35_274 ();
 FILLCELL_X4 FILLER_35_282 ();
 FILLCELL_X2 FILLER_35_286 ();
 FILLCELL_X1 FILLER_35_288 ();
 FILLCELL_X16 FILLER_35_313 ();
 FILLCELL_X2 FILLER_35_329 ();
 FILLCELL_X2 FILLER_35_344 ();
 FILLCELL_X1 FILLER_35_346 ();
 FILLCELL_X1 FILLER_35_371 ();
 FILLCELL_X2 FILLER_35_386 ();
 FILLCELL_X1 FILLER_35_391 ();
 FILLCELL_X4 FILLER_35_399 ();
 FILLCELL_X2 FILLER_35_403 ();
 FILLCELL_X8 FILLER_35_410 ();
 FILLCELL_X4 FILLER_35_418 ();
 FILLCELL_X2 FILLER_35_422 ();
 FILLCELL_X4 FILLER_35_445 ();
 FILLCELL_X2 FILLER_35_449 ();
 FILLCELL_X1 FILLER_35_456 ();
 FILLCELL_X2 FILLER_35_462 ();
 FILLCELL_X1 FILLER_35_468 ();
 FILLCELL_X1 FILLER_35_473 ();
 FILLCELL_X2 FILLER_35_490 ();
 FILLCELL_X1 FILLER_35_492 ();
 FILLCELL_X8 FILLER_35_509 ();
 FILLCELL_X2 FILLER_35_517 ();
 FILLCELL_X16 FILLER_35_537 ();
 FILLCELL_X8 FILLER_35_553 ();
 FILLCELL_X1 FILLER_35_561 ();
 FILLCELL_X16 FILLER_35_569 ();
 FILLCELL_X8 FILLER_35_605 ();
 FILLCELL_X2 FILLER_35_613 ();
 FILLCELL_X1 FILLER_35_615 ();
 FILLCELL_X8 FILLER_35_636 ();
 FILLCELL_X32 FILLER_35_648 ();
 FILLCELL_X2 FILLER_35_680 ();
 FILLCELL_X2 FILLER_35_687 ();
 FILLCELL_X1 FILLER_35_689 ();
 FILLCELL_X1 FILLER_35_721 ();
 FILLCELL_X2 FILLER_35_727 ();
 FILLCELL_X1 FILLER_35_729 ();
 FILLCELL_X2 FILLER_35_748 ();
 FILLCELL_X1 FILLER_35_750 ();
 FILLCELL_X2 FILLER_35_760 ();
 FILLCELL_X1 FILLER_35_762 ();
 FILLCELL_X2 FILLER_35_776 ();
 FILLCELL_X1 FILLER_35_778 ();
 FILLCELL_X8 FILLER_35_793 ();
 FILLCELL_X1 FILLER_35_801 ();
 FILLCELL_X8 FILLER_35_807 ();
 FILLCELL_X1 FILLER_35_861 ();
 FILLCELL_X4 FILLER_35_871 ();
 FILLCELL_X2 FILLER_35_875 ();
 FILLCELL_X1 FILLER_35_877 ();
 FILLCELL_X4 FILLER_35_882 ();
 FILLCELL_X2 FILLER_35_886 ();
 FILLCELL_X1 FILLER_35_888 ();
 FILLCELL_X2 FILLER_35_896 ();
 FILLCELL_X1 FILLER_35_898 ();
 FILLCELL_X1 FILLER_35_916 ();
 FILLCELL_X2 FILLER_35_977 ();
 FILLCELL_X8 FILLER_35_985 ();
 FILLCELL_X1 FILLER_35_993 ();
 FILLCELL_X8 FILLER_35_1025 ();
 FILLCELL_X4 FILLER_35_1033 ();
 FILLCELL_X2 FILLER_35_1037 ();
 FILLCELL_X1 FILLER_35_1039 ();
 FILLCELL_X2 FILLER_35_1088 ();
 FILLCELL_X1 FILLER_35_1090 ();
 FILLCELL_X4 FILLER_35_1094 ();
 FILLCELL_X1 FILLER_35_1098 ();
 FILLCELL_X4 FILLER_35_1118 ();
 FILLCELL_X2 FILLER_35_1127 ();
 FILLCELL_X8 FILLER_35_1149 ();
 FILLCELL_X4 FILLER_35_1157 ();
 FILLCELL_X2 FILLER_35_1161 ();
 FILLCELL_X1 FILLER_35_1163 ();
 FILLCELL_X1 FILLER_35_1188 ();
 FILLCELL_X2 FILLER_35_1198 ();
 FILLCELL_X4 FILLER_35_1207 ();
 FILLCELL_X2 FILLER_35_1211 ();
 FILLCELL_X16 FILLER_35_1240 ();
 FILLCELL_X4 FILLER_35_1256 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X1 FILLER_36_193 ();
 FILLCELL_X2 FILLER_36_211 ();
 FILLCELL_X1 FILLER_36_213 ();
 FILLCELL_X2 FILLER_36_231 ();
 FILLCELL_X1 FILLER_36_233 ();
 FILLCELL_X1 FILLER_36_256 ();
 FILLCELL_X4 FILLER_36_266 ();
 FILLCELL_X2 FILLER_36_270 ();
 FILLCELL_X4 FILLER_36_289 ();
 FILLCELL_X1 FILLER_36_293 ();
 FILLCELL_X4 FILLER_36_308 ();
 FILLCELL_X2 FILLER_36_312 ();
 FILLCELL_X1 FILLER_36_314 ();
 FILLCELL_X1 FILLER_36_322 ();
 FILLCELL_X1 FILLER_36_326 ();
 FILLCELL_X1 FILLER_36_347 ();
 FILLCELL_X8 FILLER_36_362 ();
 FILLCELL_X2 FILLER_36_370 ();
 FILLCELL_X1 FILLER_36_372 ();
 FILLCELL_X1 FILLER_36_395 ();
 FILLCELL_X1 FILLER_36_403 ();
 FILLCELL_X16 FILLER_36_411 ();
 FILLCELL_X4 FILLER_36_429 ();
 FILLCELL_X2 FILLER_36_441 ();
 FILLCELL_X1 FILLER_36_452 ();
 FILLCELL_X1 FILLER_36_457 ();
 FILLCELL_X4 FILLER_36_491 ();
 FILLCELL_X4 FILLER_36_550 ();
 FILLCELL_X1 FILLER_36_554 ();
 FILLCELL_X4 FILLER_36_558 ();
 FILLCELL_X2 FILLER_36_562 ();
 FILLCELL_X1 FILLER_36_564 ();
 FILLCELL_X8 FILLER_36_592 ();
 FILLCELL_X4 FILLER_36_600 ();
 FILLCELL_X2 FILLER_36_604 ();
 FILLCELL_X8 FILLER_36_632 ();
 FILLCELL_X4 FILLER_36_640 ();
 FILLCELL_X2 FILLER_36_644 ();
 FILLCELL_X1 FILLER_36_660 ();
 FILLCELL_X2 FILLER_36_665 ();
 FILLCELL_X8 FILLER_36_670 ();
 FILLCELL_X1 FILLER_36_678 ();
 FILLCELL_X8 FILLER_36_683 ();
 FILLCELL_X4 FILLER_36_691 ();
 FILLCELL_X2 FILLER_36_695 ();
 FILLCELL_X1 FILLER_36_697 ();
 FILLCELL_X16 FILLER_36_701 ();
 FILLCELL_X1 FILLER_36_717 ();
 FILLCELL_X2 FILLER_36_740 ();
 FILLCELL_X1 FILLER_36_742 ();
 FILLCELL_X8 FILLER_36_756 ();
 FILLCELL_X4 FILLER_36_764 ();
 FILLCELL_X2 FILLER_36_776 ();
 FILLCELL_X1 FILLER_36_778 ();
 FILLCELL_X4 FILLER_36_781 ();
 FILLCELL_X1 FILLER_36_785 ();
 FILLCELL_X2 FILLER_36_791 ();
 FILLCELL_X8 FILLER_36_807 ();
 FILLCELL_X16 FILLER_36_820 ();
 FILLCELL_X2 FILLER_36_836 ();
 FILLCELL_X1 FILLER_36_852 ();
 FILLCELL_X4 FILLER_36_889 ();
 FILLCELL_X1 FILLER_36_893 ();
 FILLCELL_X4 FILLER_36_899 ();
 FILLCELL_X2 FILLER_36_903 ();
 FILLCELL_X1 FILLER_36_909 ();
 FILLCELL_X8 FILLER_36_929 ();
 FILLCELL_X4 FILLER_36_968 ();
 FILLCELL_X4 FILLER_36_994 ();
 FILLCELL_X4 FILLER_36_1004 ();
 FILLCELL_X2 FILLER_36_1008 ();
 FILLCELL_X2 FILLER_36_1039 ();
 FILLCELL_X1 FILLER_36_1041 ();
 FILLCELL_X4 FILLER_36_1047 ();
 FILLCELL_X1 FILLER_36_1051 ();
 FILLCELL_X16 FILLER_36_1060 ();
 FILLCELL_X2 FILLER_36_1076 ();
 FILLCELL_X8 FILLER_36_1111 ();
 FILLCELL_X4 FILLER_36_1119 ();
 FILLCELL_X2 FILLER_36_1123 ();
 FILLCELL_X8 FILLER_36_1139 ();
 FILLCELL_X2 FILLER_36_1147 ();
 FILLCELL_X1 FILLER_36_1149 ();
 FILLCELL_X2 FILLER_36_1165 ();
 FILLCELL_X1 FILLER_36_1167 ();
 FILLCELL_X4 FILLER_36_1171 ();
 FILLCELL_X2 FILLER_36_1175 ();
 FILLCELL_X1 FILLER_36_1177 ();
 FILLCELL_X1 FILLER_36_1183 ();
 FILLCELL_X32 FILLER_36_1227 ();
 FILLCELL_X1 FILLER_36_1259 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X8 FILLER_37_193 ();
 FILLCELL_X4 FILLER_37_201 ();
 FILLCELL_X32 FILLER_37_212 ();
 FILLCELL_X4 FILLER_37_244 ();
 FILLCELL_X1 FILLER_37_255 ();
 FILLCELL_X1 FILLER_37_263 ();
 FILLCELL_X1 FILLER_37_271 ();
 FILLCELL_X8 FILLER_37_289 ();
 FILLCELL_X2 FILLER_37_297 ();
 FILLCELL_X2 FILLER_37_315 ();
 FILLCELL_X1 FILLER_37_317 ();
 FILLCELL_X8 FILLER_37_325 ();
 FILLCELL_X4 FILLER_37_333 ();
 FILLCELL_X1 FILLER_37_344 ();
 FILLCELL_X8 FILLER_37_359 ();
 FILLCELL_X2 FILLER_37_367 ();
 FILLCELL_X8 FILLER_37_388 ();
 FILLCELL_X1 FILLER_37_396 ();
 FILLCELL_X1 FILLER_37_414 ();
 FILLCELL_X4 FILLER_37_447 ();
 FILLCELL_X1 FILLER_37_451 ();
 FILLCELL_X4 FILLER_37_457 ();
 FILLCELL_X1 FILLER_37_461 ();
 FILLCELL_X1 FILLER_37_466 ();
 FILLCELL_X1 FILLER_37_472 ();
 FILLCELL_X1 FILLER_37_477 ();
 FILLCELL_X4 FILLER_37_503 ();
 FILLCELL_X2 FILLER_37_511 ();
 FILLCELL_X1 FILLER_37_513 ();
 FILLCELL_X2 FILLER_37_521 ();
 FILLCELL_X1 FILLER_37_523 ();
 FILLCELL_X1 FILLER_37_528 ();
 FILLCELL_X1 FILLER_37_541 ();
 FILLCELL_X16 FILLER_37_547 ();
 FILLCELL_X1 FILLER_37_563 ();
 FILLCELL_X8 FILLER_37_606 ();
 FILLCELL_X2 FILLER_37_614 ();
 FILLCELL_X1 FILLER_37_621 ();
 FILLCELL_X1 FILLER_37_625 ();
 FILLCELL_X8 FILLER_37_630 ();
 FILLCELL_X2 FILLER_37_638 ();
 FILLCELL_X4 FILLER_37_645 ();
 FILLCELL_X2 FILLER_37_649 ();
 FILLCELL_X1 FILLER_37_651 ();
 FILLCELL_X1 FILLER_37_664 ();
 FILLCELL_X2 FILLER_37_670 ();
 FILLCELL_X1 FILLER_37_672 ();
 FILLCELL_X8 FILLER_37_687 ();
 FILLCELL_X2 FILLER_37_695 ();
 FILLCELL_X1 FILLER_37_697 ();
 FILLCELL_X2 FILLER_37_701 ();
 FILLCELL_X1 FILLER_37_703 ();
 FILLCELL_X4 FILLER_37_706 ();
 FILLCELL_X1 FILLER_37_710 ();
 FILLCELL_X8 FILLER_37_715 ();
 FILLCELL_X4 FILLER_37_723 ();
 FILLCELL_X2 FILLER_37_727 ();
 FILLCELL_X4 FILLER_37_747 ();
 FILLCELL_X1 FILLER_37_751 ();
 FILLCELL_X16 FILLER_37_754 ();
 FILLCELL_X8 FILLER_37_770 ();
 FILLCELL_X4 FILLER_37_778 ();
 FILLCELL_X1 FILLER_37_782 ();
 FILLCELL_X1 FILLER_37_797 ();
 FILLCELL_X2 FILLER_37_839 ();
 FILLCELL_X1 FILLER_37_841 ();
 FILLCELL_X8 FILLER_37_871 ();
 FILLCELL_X4 FILLER_37_879 ();
 FILLCELL_X2 FILLER_37_883 ();
 FILLCELL_X1 FILLER_37_885 ();
 FILLCELL_X4 FILLER_37_906 ();
 FILLCELL_X2 FILLER_37_910 ();
 FILLCELL_X4 FILLER_37_919 ();
 FILLCELL_X2 FILLER_37_923 ();
 FILLCELL_X2 FILLER_37_930 ();
 FILLCELL_X1 FILLER_37_932 ();
 FILLCELL_X4 FILLER_37_935 ();
 FILLCELL_X2 FILLER_37_939 ();
 FILLCELL_X4 FILLER_37_946 ();
 FILLCELL_X1 FILLER_37_950 ();
 FILLCELL_X8 FILLER_37_963 ();
 FILLCELL_X2 FILLER_37_971 ();
 FILLCELL_X4 FILLER_37_984 ();
 FILLCELL_X1 FILLER_37_988 ();
 FILLCELL_X4 FILLER_37_1036 ();
 FILLCELL_X2 FILLER_37_1047 ();
 FILLCELL_X1 FILLER_37_1062 ();
 FILLCELL_X4 FILLER_37_1092 ();
 FILLCELL_X2 FILLER_37_1096 ();
 FILLCELL_X1 FILLER_37_1098 ();
 FILLCELL_X16 FILLER_37_1103 ();
 FILLCELL_X8 FILLER_37_1119 ();
 FILLCELL_X1 FILLER_37_1127 ();
 FILLCELL_X1 FILLER_37_1146 ();
 FILLCELL_X2 FILLER_37_1163 ();
 FILLCELL_X1 FILLER_37_1165 ();
 FILLCELL_X2 FILLER_37_1214 ();
 FILLCELL_X16 FILLER_37_1236 ();
 FILLCELL_X8 FILLER_37_1252 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X1 FILLER_38_193 ();
 FILLCELL_X4 FILLER_38_225 ();
 FILLCELL_X2 FILLER_38_229 ();
 FILLCELL_X2 FILLER_38_245 ();
 FILLCELL_X1 FILLER_38_247 ();
 FILLCELL_X8 FILLER_38_262 ();
 FILLCELL_X2 FILLER_38_270 ();
 FILLCELL_X8 FILLER_38_310 ();
 FILLCELL_X1 FILLER_38_318 ();
 FILLCELL_X4 FILLER_38_326 ();
 FILLCELL_X2 FILLER_38_330 ();
 FILLCELL_X1 FILLER_38_332 ();
 FILLCELL_X2 FILLER_38_364 ();
 FILLCELL_X1 FILLER_38_403 ();
 FILLCELL_X1 FILLER_38_409 ();
 FILLCELL_X1 FILLER_38_419 ();
 FILLCELL_X2 FILLER_38_427 ();
 FILLCELL_X4 FILLER_38_458 ();
 FILLCELL_X1 FILLER_38_462 ();
 FILLCELL_X8 FILLER_38_468 ();
 FILLCELL_X4 FILLER_38_476 ();
 FILLCELL_X2 FILLER_38_480 ();
 FILLCELL_X1 FILLER_38_482 ();
 FILLCELL_X4 FILLER_38_489 ();
 FILLCELL_X2 FILLER_38_507 ();
 FILLCELL_X1 FILLER_38_509 ();
 FILLCELL_X4 FILLER_38_515 ();
 FILLCELL_X8 FILLER_38_546 ();
 FILLCELL_X2 FILLER_38_554 ();
 FILLCELL_X1 FILLER_38_556 ();
 FILLCELL_X8 FILLER_38_593 ();
 FILLCELL_X8 FILLER_38_605 ();
 FILLCELL_X4 FILLER_38_613 ();
 FILLCELL_X8 FILLER_38_620 ();
 FILLCELL_X2 FILLER_38_628 ();
 FILLCELL_X1 FILLER_38_630 ();
 FILLCELL_X8 FILLER_38_632 ();
 FILLCELL_X2 FILLER_38_640 ();
 FILLCELL_X1 FILLER_38_642 ();
 FILLCELL_X1 FILLER_38_668 ();
 FILLCELL_X4 FILLER_38_674 ();
 FILLCELL_X1 FILLER_38_678 ();
 FILLCELL_X4 FILLER_38_682 ();
 FILLCELL_X1 FILLER_38_686 ();
 FILLCELL_X8 FILLER_38_691 ();
 FILLCELL_X8 FILLER_38_714 ();
 FILLCELL_X1 FILLER_38_722 ();
 FILLCELL_X2 FILLER_38_727 ();
 FILLCELL_X1 FILLER_38_729 ();
 FILLCELL_X8 FILLER_38_744 ();
 FILLCELL_X2 FILLER_38_752 ();
 FILLCELL_X1 FILLER_38_754 ();
 FILLCELL_X16 FILLER_38_770 ();
 FILLCELL_X2 FILLER_38_786 ();
 FILLCELL_X1 FILLER_38_788 ();
 FILLCELL_X8 FILLER_38_803 ();
 FILLCELL_X4 FILLER_38_820 ();
 FILLCELL_X16 FILLER_38_833 ();
 FILLCELL_X8 FILLER_38_849 ();
 FILLCELL_X4 FILLER_38_857 ();
 FILLCELL_X2 FILLER_38_861 ();
 FILLCELL_X8 FILLER_38_896 ();
 FILLCELL_X4 FILLER_38_909 ();
 FILLCELL_X8 FILLER_38_976 ();
 FILLCELL_X8 FILLER_38_1004 ();
 FILLCELL_X4 FILLER_38_1012 ();
 FILLCELL_X2 FILLER_38_1016 ();
 FILLCELL_X1 FILLER_38_1018 ();
 FILLCELL_X4 FILLER_38_1055 ();
 FILLCELL_X4 FILLER_38_1155 ();
 FILLCELL_X1 FILLER_38_1173 ();
 FILLCELL_X8 FILLER_38_1176 ();
 FILLCELL_X2 FILLER_38_1184 ();
 FILLCELL_X1 FILLER_38_1186 ();
 FILLCELL_X8 FILLER_38_1199 ();
 FILLCELL_X1 FILLER_38_1207 ();
 FILLCELL_X4 FILLER_38_1215 ();
 FILLCELL_X2 FILLER_38_1219 ();
 FILLCELL_X1 FILLER_38_1221 ();
 FILLCELL_X8 FILLER_38_1252 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X16 FILLER_39_193 ();
 FILLCELL_X4 FILLER_39_209 ();
 FILLCELL_X2 FILLER_39_213 ();
 FILLCELL_X1 FILLER_39_215 ();
 FILLCELL_X4 FILLER_39_259 ();
 FILLCELL_X16 FILLER_39_270 ();
 FILLCELL_X8 FILLER_39_286 ();
 FILLCELL_X2 FILLER_39_294 ();
 FILLCELL_X1 FILLER_39_296 ();
 FILLCELL_X8 FILLER_39_314 ();
 FILLCELL_X4 FILLER_39_322 ();
 FILLCELL_X2 FILLER_39_326 ();
 FILLCELL_X4 FILLER_39_342 ();
 FILLCELL_X8 FILLER_39_363 ();
 FILLCELL_X2 FILLER_39_371 ();
 FILLCELL_X1 FILLER_39_373 ();
 FILLCELL_X1 FILLER_39_394 ();
 FILLCELL_X1 FILLER_39_407 ();
 FILLCELL_X2 FILLER_39_415 ();
 FILLCELL_X4 FILLER_39_426 ();
 FILLCELL_X2 FILLER_39_430 ();
 FILLCELL_X1 FILLER_39_432 ();
 FILLCELL_X2 FILLER_39_468 ();
 FILLCELL_X4 FILLER_39_479 ();
 FILLCELL_X1 FILLER_39_483 ();
 FILLCELL_X2 FILLER_39_493 ();
 FILLCELL_X1 FILLER_39_504 ();
 FILLCELL_X2 FILLER_39_510 ();
 FILLCELL_X8 FILLER_39_519 ();
 FILLCELL_X4 FILLER_39_527 ();
 FILLCELL_X1 FILLER_39_531 ();
 FILLCELL_X8 FILLER_39_554 ();
 FILLCELL_X4 FILLER_39_562 ();
 FILLCELL_X2 FILLER_39_566 ();
 FILLCELL_X1 FILLER_39_568 ();
 FILLCELL_X2 FILLER_39_593 ();
 FILLCELL_X32 FILLER_39_615 ();
 FILLCELL_X1 FILLER_39_647 ();
 FILLCELL_X16 FILLER_39_664 ();
 FILLCELL_X8 FILLER_39_680 ();
 FILLCELL_X1 FILLER_39_693 ();
 FILLCELL_X1 FILLER_39_725 ();
 FILLCELL_X4 FILLER_39_731 ();
 FILLCELL_X1 FILLER_39_748 ();
 FILLCELL_X2 FILLER_39_781 ();
 FILLCELL_X1 FILLER_39_783 ();
 FILLCELL_X4 FILLER_39_793 ();
 FILLCELL_X1 FILLER_39_797 ();
 FILLCELL_X2 FILLER_39_802 ();
 FILLCELL_X4 FILLER_39_811 ();
 FILLCELL_X2 FILLER_39_815 ();
 FILLCELL_X1 FILLER_39_817 ();
 FILLCELL_X8 FILLER_39_844 ();
 FILLCELL_X2 FILLER_39_852 ();
 FILLCELL_X1 FILLER_39_854 ();
 FILLCELL_X1 FILLER_39_864 ();
 FILLCELL_X8 FILLER_39_876 ();
 FILLCELL_X2 FILLER_39_884 ();
 FILLCELL_X1 FILLER_39_886 ();
 FILLCELL_X8 FILLER_39_896 ();
 FILLCELL_X1 FILLER_39_904 ();
 FILLCELL_X1 FILLER_39_909 ();
 FILLCELL_X2 FILLER_39_919 ();
 FILLCELL_X1 FILLER_39_921 ();
 FILLCELL_X8 FILLER_39_935 ();
 FILLCELL_X2 FILLER_39_943 ();
 FILLCELL_X1 FILLER_39_945 ();
 FILLCELL_X4 FILLER_39_960 ();
 FILLCELL_X2 FILLER_39_964 ();
 FILLCELL_X1 FILLER_39_966 ();
 FILLCELL_X4 FILLER_39_974 ();
 FILLCELL_X4 FILLER_39_981 ();
 FILLCELL_X2 FILLER_39_985 ();
 FILLCELL_X1 FILLER_39_987 ();
 FILLCELL_X8 FILLER_39_1009 ();
 FILLCELL_X1 FILLER_39_1017 ();
 FILLCELL_X8 FILLER_39_1025 ();
 FILLCELL_X4 FILLER_39_1033 ();
 FILLCELL_X2 FILLER_39_1037 ();
 FILLCELL_X1 FILLER_39_1039 ();
 FILLCELL_X16 FILLER_39_1044 ();
 FILLCELL_X8 FILLER_39_1060 ();
 FILLCELL_X4 FILLER_39_1068 ();
 FILLCELL_X1 FILLER_39_1088 ();
 FILLCELL_X2 FILLER_39_1110 ();
 FILLCELL_X2 FILLER_39_1117 ();
 FILLCELL_X32 FILLER_39_1124 ();
 FILLCELL_X1 FILLER_39_1156 ();
 FILLCELL_X2 FILLER_39_1171 ();
 FILLCELL_X8 FILLER_39_1181 ();
 FILLCELL_X2 FILLER_39_1189 ();
 FILLCELL_X1 FILLER_39_1191 ();
 FILLCELL_X1 FILLER_39_1208 ();
 FILLCELL_X16 FILLER_39_1236 ();
 FILLCELL_X8 FILLER_39_1252 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X8 FILLER_40_193 ();
 FILLCELL_X2 FILLER_40_201 ();
 FILLCELL_X1 FILLER_40_203 ();
 FILLCELL_X1 FILLER_40_218 ();
 FILLCELL_X4 FILLER_40_224 ();
 FILLCELL_X2 FILLER_40_228 ();
 FILLCELL_X2 FILLER_40_244 ();
 FILLCELL_X8 FILLER_40_253 ();
 FILLCELL_X4 FILLER_40_261 ();
 FILLCELL_X8 FILLER_40_282 ();
 FILLCELL_X1 FILLER_40_290 ();
 FILLCELL_X8 FILLER_40_315 ();
 FILLCELL_X2 FILLER_40_323 ();
 FILLCELL_X4 FILLER_40_339 ();
 FILLCELL_X2 FILLER_40_343 ();
 FILLCELL_X4 FILLER_40_359 ();
 FILLCELL_X2 FILLER_40_363 ();
 FILLCELL_X16 FILLER_40_381 ();
 FILLCELL_X8 FILLER_40_397 ();
 FILLCELL_X2 FILLER_40_405 ();
 FILLCELL_X8 FILLER_40_410 ();
 FILLCELL_X4 FILLER_40_422 ();
 FILLCELL_X1 FILLER_40_426 ();
 FILLCELL_X1 FILLER_40_434 ();
 FILLCELL_X4 FILLER_40_440 ();
 FILLCELL_X1 FILLER_40_451 ();
 FILLCELL_X2 FILLER_40_455 ();
 FILLCELL_X1 FILLER_40_461 ();
 FILLCELL_X2 FILLER_40_469 ();
 FILLCELL_X2 FILLER_40_474 ();
 FILLCELL_X4 FILLER_40_481 ();
 FILLCELL_X2 FILLER_40_485 ();
 FILLCELL_X1 FILLER_40_487 ();
 FILLCELL_X4 FILLER_40_493 ();
 FILLCELL_X1 FILLER_40_497 ();
 FILLCELL_X8 FILLER_40_521 ();
 FILLCELL_X1 FILLER_40_529 ();
 FILLCELL_X2 FILLER_40_547 ();
 FILLCELL_X1 FILLER_40_549 ();
 FILLCELL_X4 FILLER_40_555 ();
 FILLCELL_X2 FILLER_40_559 ();
 FILLCELL_X2 FILLER_40_588 ();
 FILLCELL_X1 FILLER_40_590 ();
 FILLCELL_X2 FILLER_40_595 ();
 FILLCELL_X1 FILLER_40_597 ();
 FILLCELL_X16 FILLER_40_603 ();
 FILLCELL_X8 FILLER_40_619 ();
 FILLCELL_X1 FILLER_40_627 ();
 FILLCELL_X8 FILLER_40_632 ();
 FILLCELL_X2 FILLER_40_644 ();
 FILLCELL_X1 FILLER_40_646 ();
 FILLCELL_X1 FILLER_40_650 ();
 FILLCELL_X1 FILLER_40_655 ();
 FILLCELL_X4 FILLER_40_670 ();
 FILLCELL_X2 FILLER_40_674 ();
 FILLCELL_X1 FILLER_40_678 ();
 FILLCELL_X2 FILLER_40_682 ();
 FILLCELL_X2 FILLER_40_687 ();
 FILLCELL_X2 FILLER_40_698 ();
 FILLCELL_X4 FILLER_40_713 ();
 FILLCELL_X1 FILLER_40_717 ();
 FILLCELL_X1 FILLER_40_734 ();
 FILLCELL_X2 FILLER_40_753 ();
 FILLCELL_X1 FILLER_40_755 ();
 FILLCELL_X1 FILLER_40_766 ();
 FILLCELL_X1 FILLER_40_777 ();
 FILLCELL_X1 FILLER_40_784 ();
 FILLCELL_X2 FILLER_40_790 ();
 FILLCELL_X2 FILLER_40_799 ();
 FILLCELL_X1 FILLER_40_836 ();
 FILLCELL_X2 FILLER_40_851 ();
 FILLCELL_X4 FILLER_40_858 ();
 FILLCELL_X2 FILLER_40_873 ();
 FILLCELL_X4 FILLER_40_893 ();
 FILLCELL_X4 FILLER_40_916 ();
 FILLCELL_X4 FILLER_40_931 ();
 FILLCELL_X8 FILLER_40_939 ();
 FILLCELL_X2 FILLER_40_1071 ();
 FILLCELL_X8 FILLER_40_1100 ();
 FILLCELL_X4 FILLER_40_1108 ();
 FILLCELL_X2 FILLER_40_1112 ();
 FILLCELL_X1 FILLER_40_1114 ();
 FILLCELL_X8 FILLER_40_1120 ();
 FILLCELL_X2 FILLER_40_1128 ();
 FILLCELL_X2 FILLER_40_1154 ();
 FILLCELL_X1 FILLER_40_1156 ();
 FILLCELL_X2 FILLER_40_1164 ();
 FILLCELL_X8 FILLER_40_1188 ();
 FILLCELL_X1 FILLER_40_1196 ();
 FILLCELL_X2 FILLER_40_1201 ();
 FILLCELL_X8 FILLER_40_1252 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X16 FILLER_41_161 ();
 FILLCELL_X8 FILLER_41_177 ();
 FILLCELL_X4 FILLER_41_185 ();
 FILLCELL_X1 FILLER_41_189 ();
 FILLCELL_X1 FILLER_41_207 ();
 FILLCELL_X1 FILLER_41_225 ();
 FILLCELL_X1 FILLER_41_250 ();
 FILLCELL_X2 FILLER_41_258 ();
 FILLCELL_X4 FILLER_41_291 ();
 FILLCELL_X1 FILLER_41_302 ();
 FILLCELL_X1 FILLER_41_310 ();
 FILLCELL_X1 FILLER_41_335 ();
 FILLCELL_X8 FILLER_41_343 ();
 FILLCELL_X2 FILLER_41_351 ();
 FILLCELL_X1 FILLER_41_353 ();
 FILLCELL_X4 FILLER_41_361 ();
 FILLCELL_X2 FILLER_41_389 ();
 FILLCELL_X1 FILLER_41_391 ();
 FILLCELL_X4 FILLER_41_396 ();
 FILLCELL_X2 FILLER_41_404 ();
 FILLCELL_X1 FILLER_41_423 ();
 FILLCELL_X8 FILLER_41_450 ();
 FILLCELL_X4 FILLER_41_458 ();
 FILLCELL_X1 FILLER_41_462 ();
 FILLCELL_X4 FILLER_41_474 ();
 FILLCELL_X4 FILLER_41_488 ();
 FILLCELL_X2 FILLER_41_492 ();
 FILLCELL_X8 FILLER_41_508 ();
 FILLCELL_X4 FILLER_41_516 ();
 FILLCELL_X2 FILLER_41_520 ();
 FILLCELL_X1 FILLER_41_522 ();
 FILLCELL_X8 FILLER_41_527 ();
 FILLCELL_X2 FILLER_41_539 ();
 FILLCELL_X1 FILLER_41_541 ();
 FILLCELL_X16 FILLER_41_553 ();
 FILLCELL_X8 FILLER_41_569 ();
 FILLCELL_X1 FILLER_41_577 ();
 FILLCELL_X2 FILLER_41_584 ();
 FILLCELL_X8 FILLER_41_588 ();
 FILLCELL_X2 FILLER_41_596 ();
 FILLCELL_X2 FILLER_41_603 ();
 FILLCELL_X16 FILLER_41_609 ();
 FILLCELL_X4 FILLER_41_625 ();
 FILLCELL_X2 FILLER_41_629 ();
 FILLCELL_X1 FILLER_41_641 ();
 FILLCELL_X2 FILLER_41_656 ();
 FILLCELL_X1 FILLER_41_658 ();
 FILLCELL_X2 FILLER_41_667 ();
 FILLCELL_X8 FILLER_41_688 ();
 FILLCELL_X2 FILLER_41_696 ();
 FILLCELL_X1 FILLER_41_698 ();
 FILLCELL_X4 FILLER_41_706 ();
 FILLCELL_X8 FILLER_41_724 ();
 FILLCELL_X4 FILLER_41_732 ();
 FILLCELL_X2 FILLER_41_736 ();
 FILLCELL_X1 FILLER_41_738 ();
 FILLCELL_X8 FILLER_41_748 ();
 FILLCELL_X2 FILLER_41_756 ();
 FILLCELL_X2 FILLER_41_762 ();
 FILLCELL_X1 FILLER_41_769 ();
 FILLCELL_X1 FILLER_41_791 ();
 FILLCELL_X2 FILLER_41_801 ();
 FILLCELL_X1 FILLER_41_803 ();
 FILLCELL_X2 FILLER_41_823 ();
 FILLCELL_X16 FILLER_41_829 ();
 FILLCELL_X2 FILLER_41_845 ();
 FILLCELL_X1 FILLER_41_872 ();
 FILLCELL_X2 FILLER_41_902 ();
 FILLCELL_X1 FILLER_41_904 ();
 FILLCELL_X4 FILLER_41_925 ();
 FILLCELL_X2 FILLER_41_929 ();
 FILLCELL_X4 FILLER_41_951 ();
 FILLCELL_X1 FILLER_41_955 ();
 FILLCELL_X8 FILLER_41_961 ();
 FILLCELL_X2 FILLER_41_969 ();
 FILLCELL_X8 FILLER_41_976 ();
 FILLCELL_X2 FILLER_41_984 ();
 FILLCELL_X4 FILLER_41_990 ();
 FILLCELL_X2 FILLER_41_994 ();
 FILLCELL_X1 FILLER_41_996 ();
 FILLCELL_X2 FILLER_41_1033 ();
 FILLCELL_X1 FILLER_41_1038 ();
 FILLCELL_X2 FILLER_41_1044 ();
 FILLCELL_X2 FILLER_41_1053 ();
 FILLCELL_X2 FILLER_41_1075 ();
 FILLCELL_X1 FILLER_41_1077 ();
 FILLCELL_X1 FILLER_41_1085 ();
 FILLCELL_X16 FILLER_41_1097 ();
 FILLCELL_X8 FILLER_41_1113 ();
 FILLCELL_X4 FILLER_41_1121 ();
 FILLCELL_X1 FILLER_41_1125 ();
 FILLCELL_X8 FILLER_41_1135 ();
 FILLCELL_X2 FILLER_41_1143 ();
 FILLCELL_X2 FILLER_41_1176 ();
 FILLCELL_X1 FILLER_41_1178 ();
 FILLCELL_X4 FILLER_41_1183 ();
 FILLCELL_X2 FILLER_41_1187 ();
 FILLCELL_X1 FILLER_41_1196 ();
 FILLCELL_X32 FILLER_41_1211 ();
 FILLCELL_X16 FILLER_41_1243 ();
 FILLCELL_X1 FILLER_41_1259 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X8 FILLER_42_193 ();
 FILLCELL_X2 FILLER_42_201 ();
 FILLCELL_X2 FILLER_42_210 ();
 FILLCELL_X8 FILLER_42_219 ();
 FILLCELL_X2 FILLER_42_227 ();
 FILLCELL_X1 FILLER_42_229 ();
 FILLCELL_X4 FILLER_42_237 ();
 FILLCELL_X2 FILLER_42_241 ();
 FILLCELL_X1 FILLER_42_243 ();
 FILLCELL_X4 FILLER_42_260 ();
 FILLCELL_X2 FILLER_42_264 ();
 FILLCELL_X1 FILLER_42_266 ();
 FILLCELL_X8 FILLER_42_281 ();
 FILLCELL_X2 FILLER_42_289 ();
 FILLCELL_X1 FILLER_42_291 ();
 FILLCELL_X1 FILLER_42_299 ();
 FILLCELL_X2 FILLER_42_307 ();
 FILLCELL_X1 FILLER_42_309 ();
 FILLCELL_X2 FILLER_42_317 ();
 FILLCELL_X1 FILLER_42_319 ();
 FILLCELL_X2 FILLER_42_334 ();
 FILLCELL_X1 FILLER_42_336 ();
 FILLCELL_X1 FILLER_42_341 ();
 FILLCELL_X1 FILLER_42_351 ();
 FILLCELL_X1 FILLER_42_359 ();
 FILLCELL_X1 FILLER_42_367 ();
 FILLCELL_X16 FILLER_42_375 ();
 FILLCELL_X1 FILLER_42_394 ();
 FILLCELL_X1 FILLER_42_408 ();
 FILLCELL_X2 FILLER_42_417 ();
 FILLCELL_X1 FILLER_42_419 ();
 FILLCELL_X8 FILLER_42_427 ();
 FILLCELL_X4 FILLER_42_435 ();
 FILLCELL_X1 FILLER_42_439 ();
 FILLCELL_X1 FILLER_42_444 ();
 FILLCELL_X4 FILLER_42_449 ();
 FILLCELL_X1 FILLER_42_457 ();
 FILLCELL_X2 FILLER_42_461 ();
 FILLCELL_X4 FILLER_42_474 ();
 FILLCELL_X1 FILLER_42_478 ();
 FILLCELL_X4 FILLER_42_486 ();
 FILLCELL_X4 FILLER_42_494 ();
 FILLCELL_X2 FILLER_42_505 ();
 FILLCELL_X4 FILLER_42_509 ();
 FILLCELL_X1 FILLER_42_513 ();
 FILLCELL_X4 FILLER_42_549 ();
 FILLCELL_X1 FILLER_42_560 ();
 FILLCELL_X1 FILLER_42_565 ();
 FILLCELL_X2 FILLER_42_595 ();
 FILLCELL_X2 FILLER_42_603 ();
 FILLCELL_X1 FILLER_42_605 ();
 FILLCELL_X8 FILLER_42_615 ();
 FILLCELL_X4 FILLER_42_623 ();
 FILLCELL_X4 FILLER_42_642 ();
 FILLCELL_X1 FILLER_42_646 ();
 FILLCELL_X4 FILLER_42_656 ();
 FILLCELL_X2 FILLER_42_660 ();
 FILLCELL_X1 FILLER_42_662 ();
 FILLCELL_X8 FILLER_42_667 ();
 FILLCELL_X4 FILLER_42_675 ();
 FILLCELL_X16 FILLER_42_683 ();
 FILLCELL_X8 FILLER_42_699 ();
 FILLCELL_X4 FILLER_42_707 ();
 FILLCELL_X1 FILLER_42_718 ();
 FILLCELL_X4 FILLER_42_728 ();
 FILLCELL_X2 FILLER_42_732 ();
 FILLCELL_X2 FILLER_42_738 ();
 FILLCELL_X16 FILLER_42_756 ();
 FILLCELL_X2 FILLER_42_772 ();
 FILLCELL_X8 FILLER_42_792 ();
 FILLCELL_X4 FILLER_42_800 ();
 FILLCELL_X16 FILLER_42_847 ();
 FILLCELL_X4 FILLER_42_863 ();
 FILLCELL_X1 FILLER_42_879 ();
 FILLCELL_X1 FILLER_42_894 ();
 FILLCELL_X2 FILLER_42_908 ();
 FILLCELL_X2 FILLER_42_915 ();
 FILLCELL_X8 FILLER_42_924 ();
 FILLCELL_X4 FILLER_42_932 ();
 FILLCELL_X1 FILLER_42_936 ();
 FILLCELL_X4 FILLER_42_949 ();
 FILLCELL_X2 FILLER_42_953 ();
 FILLCELL_X1 FILLER_42_955 ();
 FILLCELL_X1 FILLER_42_963 ();
 FILLCELL_X4 FILLER_42_1009 ();
 FILLCELL_X2 FILLER_42_1013 ();
 FILLCELL_X1 FILLER_42_1015 ();
 FILLCELL_X16 FILLER_42_1055 ();
 FILLCELL_X2 FILLER_42_1071 ();
 FILLCELL_X1 FILLER_42_1073 ();
 FILLCELL_X1 FILLER_42_1083 ();
 FILLCELL_X4 FILLER_42_1113 ();
 FILLCELL_X16 FILLER_42_1121 ();
 FILLCELL_X2 FILLER_42_1137 ();
 FILLCELL_X1 FILLER_42_1163 ();
 FILLCELL_X16 FILLER_42_1168 ();
 FILLCELL_X4 FILLER_42_1184 ();
 FILLCELL_X1 FILLER_42_1188 ();
 FILLCELL_X16 FILLER_42_1231 ();
 FILLCELL_X8 FILLER_42_1247 ();
 FILLCELL_X4 FILLER_42_1255 ();
 FILLCELL_X1 FILLER_42_1259 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X4 FILLER_43_193 ();
 FILLCELL_X1 FILLER_43_197 ();
 FILLCELL_X1 FILLER_43_229 ();
 FILLCELL_X2 FILLER_43_237 ();
 FILLCELL_X1 FILLER_43_239 ();
 FILLCELL_X4 FILLER_43_247 ();
 FILLCELL_X2 FILLER_43_251 ();
 FILLCELL_X4 FILLER_43_286 ();
 FILLCELL_X1 FILLER_43_290 ();
 FILLCELL_X16 FILLER_43_298 ();
 FILLCELL_X2 FILLER_43_314 ();
 FILLCELL_X4 FILLER_43_337 ();
 FILLCELL_X2 FILLER_43_341 ();
 FILLCELL_X4 FILLER_43_363 ();
 FILLCELL_X2 FILLER_43_367 ();
 FILLCELL_X4 FILLER_43_386 ();
 FILLCELL_X2 FILLER_43_404 ();
 FILLCELL_X1 FILLER_43_406 ();
 FILLCELL_X8 FILLER_43_426 ();
 FILLCELL_X4 FILLER_43_434 ();
 FILLCELL_X2 FILLER_43_438 ();
 FILLCELL_X8 FILLER_43_451 ();
 FILLCELL_X2 FILLER_43_459 ();
 FILLCELL_X1 FILLER_43_461 ();
 FILLCELL_X16 FILLER_43_471 ();
 FILLCELL_X1 FILLER_43_487 ();
 FILLCELL_X8 FILLER_43_493 ();
 FILLCELL_X2 FILLER_43_501 ();
 FILLCELL_X4 FILLER_43_515 ();
 FILLCELL_X2 FILLER_43_519 ();
 FILLCELL_X8 FILLER_43_525 ();
 FILLCELL_X4 FILLER_43_535 ();
 FILLCELL_X2 FILLER_43_539 ();
 FILLCELL_X1 FILLER_43_541 ();
 FILLCELL_X2 FILLER_43_551 ();
 FILLCELL_X1 FILLER_43_553 ();
 FILLCELL_X32 FILLER_43_557 ();
 FILLCELL_X4 FILLER_43_589 ();
 FILLCELL_X2 FILLER_43_593 ();
 FILLCELL_X2 FILLER_43_617 ();
 FILLCELL_X1 FILLER_43_619 ();
 FILLCELL_X2 FILLER_43_656 ();
 FILLCELL_X1 FILLER_43_658 ();
 FILLCELL_X4 FILLER_43_670 ();
 FILLCELL_X1 FILLER_43_674 ();
 FILLCELL_X2 FILLER_43_678 ();
 FILLCELL_X1 FILLER_43_680 ();
 FILLCELL_X2 FILLER_43_685 ();
 FILLCELL_X8 FILLER_43_691 ();
 FILLCELL_X4 FILLER_43_699 ();
 FILLCELL_X1 FILLER_43_703 ();
 FILLCELL_X2 FILLER_43_711 ();
 FILLCELL_X1 FILLER_43_713 ();
 FILLCELL_X2 FILLER_43_721 ();
 FILLCELL_X1 FILLER_43_723 ();
 FILLCELL_X4 FILLER_43_731 ();
 FILLCELL_X2 FILLER_43_748 ();
 FILLCELL_X1 FILLER_43_750 ();
 FILLCELL_X4 FILLER_43_768 ();
 FILLCELL_X1 FILLER_43_772 ();
 FILLCELL_X16 FILLER_43_795 ();
 FILLCELL_X8 FILLER_43_811 ();
 FILLCELL_X4 FILLER_43_819 ();
 FILLCELL_X8 FILLER_43_826 ();
 FILLCELL_X1 FILLER_43_834 ();
 FILLCELL_X8 FILLER_43_838 ();
 FILLCELL_X2 FILLER_43_846 ();
 FILLCELL_X1 FILLER_43_848 ();
 FILLCELL_X4 FILLER_43_870 ();
 FILLCELL_X1 FILLER_43_874 ();
 FILLCELL_X4 FILLER_43_897 ();
 FILLCELL_X1 FILLER_43_901 ();
 FILLCELL_X2 FILLER_43_922 ();
 FILLCELL_X4 FILLER_43_944 ();
 FILLCELL_X2 FILLER_43_948 ();
 FILLCELL_X4 FILLER_43_970 ();
 FILLCELL_X2 FILLER_43_974 ();
 FILLCELL_X1 FILLER_43_976 ();
 FILLCELL_X4 FILLER_43_984 ();
 FILLCELL_X2 FILLER_43_988 ();
 FILLCELL_X1 FILLER_43_990 ();
 FILLCELL_X2 FILLER_43_994 ();
 FILLCELL_X1 FILLER_43_996 ();
 FILLCELL_X16 FILLER_43_1019 ();
 FILLCELL_X4 FILLER_43_1035 ();
 FILLCELL_X1 FILLER_43_1039 ();
 FILLCELL_X2 FILLER_43_1045 ();
 FILLCELL_X1 FILLER_43_1074 ();
 FILLCELL_X2 FILLER_43_1108 ();
 FILLCELL_X2 FILLER_43_1165 ();
 FILLCELL_X1 FILLER_43_1167 ();
 FILLCELL_X16 FILLER_43_1194 ();
 FILLCELL_X4 FILLER_43_1210 ();
 FILLCELL_X1 FILLER_43_1214 ();
 FILLCELL_X32 FILLER_43_1220 ();
 FILLCELL_X8 FILLER_43_1252 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X16 FILLER_44_193 ();
 FILLCELL_X8 FILLER_44_209 ();
 FILLCELL_X2 FILLER_44_234 ();
 FILLCELL_X1 FILLER_44_236 ();
 FILLCELL_X1 FILLER_44_280 ();
 FILLCELL_X8 FILLER_44_288 ();
 FILLCELL_X4 FILLER_44_296 ();
 FILLCELL_X1 FILLER_44_300 ();
 FILLCELL_X32 FILLER_44_359 ();
 FILLCELL_X1 FILLER_44_391 ();
 FILLCELL_X4 FILLER_44_416 ();
 FILLCELL_X2 FILLER_44_420 ();
 FILLCELL_X4 FILLER_44_426 ();
 FILLCELL_X4 FILLER_44_463 ();
 FILLCELL_X2 FILLER_44_467 ();
 FILLCELL_X1 FILLER_44_469 ();
 FILLCELL_X1 FILLER_44_477 ();
 FILLCELL_X4 FILLER_44_482 ();
 FILLCELL_X2 FILLER_44_490 ();
 FILLCELL_X1 FILLER_44_492 ();
 FILLCELL_X2 FILLER_44_497 ();
 FILLCELL_X4 FILLER_44_509 ();
 FILLCELL_X2 FILLER_44_513 ();
 FILLCELL_X4 FILLER_44_530 ();
 FILLCELL_X1 FILLER_44_542 ();
 FILLCELL_X32 FILLER_44_554 ();
 FILLCELL_X8 FILLER_44_586 ();
 FILLCELL_X2 FILLER_44_601 ();
 FILLCELL_X1 FILLER_44_603 ();
 FILLCELL_X8 FILLER_44_611 ();
 FILLCELL_X4 FILLER_44_619 ();
 FILLCELL_X2 FILLER_44_623 ();
 FILLCELL_X1 FILLER_44_625 ();
 FILLCELL_X1 FILLER_44_630 ();
 FILLCELL_X1 FILLER_44_632 ();
 FILLCELL_X4 FILLER_44_640 ();
 FILLCELL_X4 FILLER_44_650 ();
 FILLCELL_X4 FILLER_44_675 ();
 FILLCELL_X1 FILLER_44_685 ();
 FILLCELL_X1 FILLER_44_707 ();
 FILLCELL_X1 FILLER_44_722 ();
 FILLCELL_X2 FILLER_44_737 ();
 FILLCELL_X4 FILLER_44_744 ();
 FILLCELL_X1 FILLER_44_748 ();
 FILLCELL_X8 FILLER_44_756 ();
 FILLCELL_X1 FILLER_44_764 ();
 FILLCELL_X16 FILLER_44_770 ();
 FILLCELL_X8 FILLER_44_798 ();
 FILLCELL_X2 FILLER_44_806 ();
 FILLCELL_X8 FILLER_44_841 ();
 FILLCELL_X2 FILLER_44_874 ();
 FILLCELL_X4 FILLER_44_878 ();
 FILLCELL_X4 FILLER_44_889 ();
 FILLCELL_X1 FILLER_44_893 ();
 FILLCELL_X2 FILLER_44_898 ();
 FILLCELL_X1 FILLER_44_900 ();
 FILLCELL_X4 FILLER_44_913 ();
 FILLCELL_X2 FILLER_44_917 ();
 FILLCELL_X1 FILLER_44_919 ();
 FILLCELL_X4 FILLER_44_925 ();
 FILLCELL_X2 FILLER_44_941 ();
 FILLCELL_X1 FILLER_44_943 ();
 FILLCELL_X2 FILLER_44_966 ();
 FILLCELL_X2 FILLER_44_973 ();
 FILLCELL_X2 FILLER_44_988 ();
 FILLCELL_X1 FILLER_44_990 ();
 FILLCELL_X1 FILLER_44_995 ();
 FILLCELL_X8 FILLER_44_1005 ();
 FILLCELL_X1 FILLER_44_1013 ();
 FILLCELL_X2 FILLER_44_1056 ();
 FILLCELL_X16 FILLER_44_1065 ();
 FILLCELL_X8 FILLER_44_1081 ();
 FILLCELL_X2 FILLER_44_1089 ();
 FILLCELL_X1 FILLER_44_1116 ();
 FILLCELL_X1 FILLER_44_1123 ();
 FILLCELL_X2 FILLER_44_1128 ();
 FILLCELL_X8 FILLER_44_1138 ();
 FILLCELL_X2 FILLER_44_1146 ();
 FILLCELL_X1 FILLER_44_1153 ();
 FILLCELL_X4 FILLER_44_1160 ();
 FILLCELL_X2 FILLER_44_1164 ();
 FILLCELL_X4 FILLER_44_1170 ();
 FILLCELL_X2 FILLER_44_1180 ();
 FILLCELL_X1 FILLER_44_1182 ();
 FILLCELL_X4 FILLER_44_1216 ();
 FILLCELL_X1 FILLER_44_1220 ();
 FILLCELL_X16 FILLER_44_1226 ();
 FILLCELL_X1 FILLER_44_1242 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X16 FILLER_45_225 ();
 FILLCELL_X8 FILLER_45_241 ();
 FILLCELL_X1 FILLER_45_249 ();
 FILLCELL_X4 FILLER_45_272 ();
 FILLCELL_X1 FILLER_45_276 ();
 FILLCELL_X32 FILLER_45_297 ();
 FILLCELL_X8 FILLER_45_329 ();
 FILLCELL_X4 FILLER_45_337 ();
 FILLCELL_X2 FILLER_45_341 ();
 FILLCELL_X16 FILLER_45_370 ();
 FILLCELL_X8 FILLER_45_386 ();
 FILLCELL_X2 FILLER_45_394 ();
 FILLCELL_X4 FILLER_45_399 ();
 FILLCELL_X2 FILLER_45_403 ();
 FILLCELL_X2 FILLER_45_408 ();
 FILLCELL_X1 FILLER_45_410 ();
 FILLCELL_X4 FILLER_45_423 ();
 FILLCELL_X2 FILLER_45_427 ();
 FILLCELL_X1 FILLER_45_429 ();
 FILLCELL_X2 FILLER_45_438 ();
 FILLCELL_X1 FILLER_45_440 ();
 FILLCELL_X2 FILLER_45_446 ();
 FILLCELL_X2 FILLER_45_451 ();
 FILLCELL_X1 FILLER_45_453 ();
 FILLCELL_X4 FILLER_45_475 ();
 FILLCELL_X1 FILLER_45_479 ();
 FILLCELL_X4 FILLER_45_488 ();
 FILLCELL_X1 FILLER_45_492 ();
 FILLCELL_X2 FILLER_45_507 ();
 FILLCELL_X4 FILLER_45_516 ();
 FILLCELL_X2 FILLER_45_520 ();
 FILLCELL_X2 FILLER_45_526 ();
 FILLCELL_X2 FILLER_45_532 ();
 FILLCELL_X4 FILLER_45_545 ();
 FILLCELL_X1 FILLER_45_582 ();
 FILLCELL_X2 FILLER_45_607 ();
 FILLCELL_X2 FILLER_45_618 ();
 FILLCELL_X1 FILLER_45_631 ();
 FILLCELL_X8 FILLER_45_635 ();
 FILLCELL_X4 FILLER_45_643 ();
 FILLCELL_X1 FILLER_45_651 ();
 FILLCELL_X1 FILLER_45_656 ();
 FILLCELL_X8 FILLER_45_666 ();
 FILLCELL_X4 FILLER_45_674 ();
 FILLCELL_X1 FILLER_45_683 ();
 FILLCELL_X2 FILLER_45_691 ();
 FILLCELL_X1 FILLER_45_693 ();
 FILLCELL_X2 FILLER_45_697 ();
 FILLCELL_X1 FILLER_45_699 ();
 FILLCELL_X2 FILLER_45_714 ();
 FILLCELL_X1 FILLER_45_716 ();
 FILLCELL_X2 FILLER_45_741 ();
 FILLCELL_X1 FILLER_45_743 ();
 FILLCELL_X4 FILLER_45_747 ();
 FILLCELL_X1 FILLER_45_751 ();
 FILLCELL_X4 FILLER_45_765 ();
 FILLCELL_X16 FILLER_45_782 ();
 FILLCELL_X8 FILLER_45_798 ();
 FILLCELL_X2 FILLER_45_806 ();
 FILLCELL_X1 FILLER_45_808 ();
 FILLCELL_X2 FILLER_45_814 ();
 FILLCELL_X4 FILLER_45_825 ();
 FILLCELL_X4 FILLER_45_840 ();
 FILLCELL_X4 FILLER_45_849 ();
 FILLCELL_X2 FILLER_45_853 ();
 FILLCELL_X4 FILLER_45_865 ();
 FILLCELL_X2 FILLER_45_912 ();
 FILLCELL_X4 FILLER_45_921 ();
 FILLCELL_X2 FILLER_45_957 ();
 FILLCELL_X1 FILLER_45_959 ();
 FILLCELL_X2 FILLER_45_965 ();
 FILLCELL_X2 FILLER_45_974 ();
 FILLCELL_X1 FILLER_45_976 ();
 FILLCELL_X8 FILLER_45_1004 ();
 FILLCELL_X2 FILLER_45_1032 ();
 FILLCELL_X1 FILLER_45_1034 ();
 FILLCELL_X2 FILLER_45_1055 ();
 FILLCELL_X2 FILLER_45_1066 ();
 FILLCELL_X1 FILLER_45_1068 ();
 FILLCELL_X8 FILLER_45_1100 ();
 FILLCELL_X4 FILLER_45_1108 ();
 FILLCELL_X2 FILLER_45_1112 ();
 FILLCELL_X1 FILLER_45_1114 ();
 FILLCELL_X4 FILLER_45_1120 ();
 FILLCELL_X2 FILLER_45_1124 ();
 FILLCELL_X8 FILLER_45_1130 ();
 FILLCELL_X4 FILLER_45_1138 ();
 FILLCELL_X2 FILLER_45_1142 ();
 FILLCELL_X1 FILLER_45_1144 ();
 FILLCELL_X4 FILLER_45_1151 ();
 FILLCELL_X2 FILLER_45_1155 ();
 FILLCELL_X1 FILLER_45_1157 ();
 FILLCELL_X2 FILLER_45_1182 ();
 FILLCELL_X4 FILLER_45_1204 ();
 FILLCELL_X1 FILLER_45_1232 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X2 FILLER_45_1257 ();
 FILLCELL_X1 FILLER_45_1259 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X8 FILLER_46_225 ();
 FILLCELL_X1 FILLER_46_233 ();
 FILLCELL_X4 FILLER_46_254 ();
 FILLCELL_X1 FILLER_46_278 ();
 FILLCELL_X16 FILLER_46_286 ();
 FILLCELL_X2 FILLER_46_302 ();
 FILLCELL_X1 FILLER_46_304 ();
 FILLCELL_X8 FILLER_46_312 ();
 FILLCELL_X4 FILLER_46_320 ();
 FILLCELL_X4 FILLER_46_351 ();
 FILLCELL_X8 FILLER_46_382 ();
 FILLCELL_X1 FILLER_46_394 ();
 FILLCELL_X1 FILLER_46_399 ();
 FILLCELL_X2 FILLER_46_404 ();
 FILLCELL_X1 FILLER_46_410 ();
 FILLCELL_X1 FILLER_46_419 ();
 FILLCELL_X1 FILLER_46_425 ();
 FILLCELL_X1 FILLER_46_445 ();
 FILLCELL_X2 FILLER_46_450 ();
 FILLCELL_X1 FILLER_46_455 ();
 FILLCELL_X16 FILLER_46_467 ();
 FILLCELL_X8 FILLER_46_483 ();
 FILLCELL_X4 FILLER_46_491 ();
 FILLCELL_X1 FILLER_46_503 ();
 FILLCELL_X8 FILLER_46_515 ();
 FILLCELL_X4 FILLER_46_523 ();
 FILLCELL_X8 FILLER_46_533 ();
 FILLCELL_X4 FILLER_46_541 ();
 FILLCELL_X1 FILLER_46_545 ();
 FILLCELL_X1 FILLER_46_552 ();
 FILLCELL_X16 FILLER_46_563 ();
 FILLCELL_X8 FILLER_46_579 ();
 FILLCELL_X4 FILLER_46_587 ();
 FILLCELL_X2 FILLER_46_591 ();
 FILLCELL_X4 FILLER_46_596 ();
 FILLCELL_X8 FILLER_46_607 ();
 FILLCELL_X4 FILLER_46_615 ();
 FILLCELL_X8 FILLER_46_632 ();
 FILLCELL_X2 FILLER_46_640 ();
 FILLCELL_X2 FILLER_46_651 ();
 FILLCELL_X1 FILLER_46_653 ();
 FILLCELL_X8 FILLER_46_671 ();
 FILLCELL_X1 FILLER_46_679 ();
 FILLCELL_X8 FILLER_46_682 ();
 FILLCELL_X2 FILLER_46_690 ();
 FILLCELL_X1 FILLER_46_692 ();
 FILLCELL_X8 FILLER_46_700 ();
 FILLCELL_X2 FILLER_46_708 ();
 FILLCELL_X1 FILLER_46_710 ();
 FILLCELL_X16 FILLER_46_718 ();
 FILLCELL_X2 FILLER_46_734 ();
 FILLCELL_X1 FILLER_46_741 ();
 FILLCELL_X4 FILLER_46_747 ();
 FILLCELL_X2 FILLER_46_756 ();
 FILLCELL_X1 FILLER_46_758 ();
 FILLCELL_X8 FILLER_46_764 ();
 FILLCELL_X4 FILLER_46_772 ();
 FILLCELL_X4 FILLER_46_814 ();
 FILLCELL_X1 FILLER_46_839 ();
 FILLCELL_X4 FILLER_46_849 ();
 FILLCELL_X4 FILLER_46_879 ();
 FILLCELL_X2 FILLER_46_883 ();
 FILLCELL_X1 FILLER_46_885 ();
 FILLCELL_X8 FILLER_46_890 ();
 FILLCELL_X4 FILLER_46_898 ();
 FILLCELL_X2 FILLER_46_922 ();
 FILLCELL_X1 FILLER_46_924 ();
 FILLCELL_X16 FILLER_46_932 ();
 FILLCELL_X4 FILLER_46_948 ();
 FILLCELL_X1 FILLER_46_952 ();
 FILLCELL_X8 FILLER_46_962 ();
 FILLCELL_X4 FILLER_46_970 ();
 FILLCELL_X1 FILLER_46_974 ();
 FILLCELL_X2 FILLER_46_985 ();
 FILLCELL_X2 FILLER_46_1034 ();
 FILLCELL_X2 FILLER_46_1041 ();
 FILLCELL_X1 FILLER_46_1043 ();
 FILLCELL_X2 FILLER_46_1050 ();
 FILLCELL_X1 FILLER_46_1052 ();
 FILLCELL_X2 FILLER_46_1055 ();
 FILLCELL_X4 FILLER_46_1071 ();
 FILLCELL_X2 FILLER_46_1075 ();
 FILLCELL_X1 FILLER_46_1077 ();
 FILLCELL_X1 FILLER_46_1124 ();
 FILLCELL_X1 FILLER_46_1136 ();
 FILLCELL_X4 FILLER_46_1159 ();
 FILLCELL_X8 FILLER_46_1169 ();
 FILLCELL_X1 FILLER_46_1177 ();
 FILLCELL_X2 FILLER_46_1192 ();
 FILLCELL_X8 FILLER_46_1205 ();
 FILLCELL_X2 FILLER_46_1213 ();
 FILLCELL_X1 FILLER_46_1215 ();
 FILLCELL_X1 FILLER_46_1242 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X8 FILLER_47_193 ();
 FILLCELL_X2 FILLER_47_201 ();
 FILLCELL_X1 FILLER_47_203 ();
 FILLCELL_X32 FILLER_47_231 ();
 FILLCELL_X1 FILLER_47_263 ();
 FILLCELL_X8 FILLER_47_284 ();
 FILLCELL_X2 FILLER_47_292 ();
 FILLCELL_X16 FILLER_47_314 ();
 FILLCELL_X4 FILLER_47_330 ();
 FILLCELL_X2 FILLER_47_334 ();
 FILLCELL_X16 FILLER_47_343 ();
 FILLCELL_X2 FILLER_47_359 ();
 FILLCELL_X8 FILLER_47_388 ();
 FILLCELL_X4 FILLER_47_396 ();
 FILLCELL_X1 FILLER_47_412 ();
 FILLCELL_X2 FILLER_47_417 ();
 FILLCELL_X2 FILLER_47_423 ();
 FILLCELL_X1 FILLER_47_425 ();
 FILLCELL_X1 FILLER_47_434 ();
 FILLCELL_X4 FILLER_47_442 ();
 FILLCELL_X2 FILLER_47_460 ();
 FILLCELL_X8 FILLER_47_467 ();
 FILLCELL_X2 FILLER_47_475 ();
 FILLCELL_X2 FILLER_47_482 ();
 FILLCELL_X1 FILLER_47_484 ();
 FILLCELL_X1 FILLER_47_493 ();
 FILLCELL_X16 FILLER_47_498 ();
 FILLCELL_X2 FILLER_47_514 ();
 FILLCELL_X1 FILLER_47_516 ();
 FILLCELL_X8 FILLER_47_526 ();
 FILLCELL_X4 FILLER_47_558 ();
 FILLCELL_X2 FILLER_47_593 ();
 FILLCELL_X1 FILLER_47_595 ();
 FILLCELL_X2 FILLER_47_607 ();
 FILLCELL_X4 FILLER_47_631 ();
 FILLCELL_X2 FILLER_47_635 ();
 FILLCELL_X4 FILLER_47_641 ();
 FILLCELL_X4 FILLER_47_659 ();
 FILLCELL_X8 FILLER_47_670 ();
 FILLCELL_X2 FILLER_47_678 ();
 FILLCELL_X4 FILLER_47_685 ();
 FILLCELL_X2 FILLER_47_689 ();
 FILLCELL_X1 FILLER_47_691 ();
 FILLCELL_X8 FILLER_47_701 ();
 FILLCELL_X1 FILLER_47_709 ();
 FILLCELL_X4 FILLER_47_719 ();
 FILLCELL_X2 FILLER_47_727 ();
 FILLCELL_X1 FILLER_47_729 ();
 FILLCELL_X2 FILLER_47_740 ();
 FILLCELL_X1 FILLER_47_742 ();
 FILLCELL_X2 FILLER_47_748 ();
 FILLCELL_X2 FILLER_47_755 ();
 FILLCELL_X2 FILLER_47_779 ();
 FILLCELL_X1 FILLER_47_781 ();
 FILLCELL_X16 FILLER_47_784 ();
 FILLCELL_X8 FILLER_47_800 ();
 FILLCELL_X2 FILLER_47_808 ();
 FILLCELL_X2 FILLER_47_813 ();
 FILLCELL_X4 FILLER_47_818 ();
 FILLCELL_X1 FILLER_47_825 ();
 FILLCELL_X8 FILLER_47_849 ();
 FILLCELL_X2 FILLER_47_857 ();
 FILLCELL_X4 FILLER_47_864 ();
 FILLCELL_X1 FILLER_47_868 ();
 FILLCELL_X1 FILLER_47_880 ();
 FILLCELL_X16 FILLER_47_901 ();
 FILLCELL_X1 FILLER_47_917 ();
 FILLCELL_X2 FILLER_47_928 ();
 FILLCELL_X1 FILLER_47_930 ();
 FILLCELL_X4 FILLER_47_935 ();
 FILLCELL_X2 FILLER_47_939 ();
 FILLCELL_X8 FILLER_47_967 ();
 FILLCELL_X2 FILLER_47_975 ();
 FILLCELL_X1 FILLER_47_977 ();
 FILLCELL_X4 FILLER_47_981 ();
 FILLCELL_X32 FILLER_47_990 ();
 FILLCELL_X16 FILLER_47_1022 ();
 FILLCELL_X8 FILLER_47_1038 ();
 FILLCELL_X2 FILLER_47_1046 ();
 FILLCELL_X1 FILLER_47_1048 ();
 FILLCELL_X2 FILLER_47_1063 ();
 FILLCELL_X2 FILLER_47_1085 ();
 FILLCELL_X2 FILLER_47_1093 ();
 FILLCELL_X4 FILLER_47_1097 ();
 FILLCELL_X4 FILLER_47_1123 ();
 FILLCELL_X2 FILLER_47_1127 ();
 FILLCELL_X2 FILLER_47_1132 ();
 FILLCELL_X8 FILLER_47_1136 ();
 FILLCELL_X2 FILLER_47_1144 ();
 FILLCELL_X2 FILLER_47_1182 ();
 FILLCELL_X1 FILLER_47_1184 ();
 FILLCELL_X8 FILLER_47_1205 ();
 FILLCELL_X4 FILLER_47_1213 ();
 FILLCELL_X1 FILLER_47_1217 ();
 FILLCELL_X2 FILLER_47_1224 ();
 FILLCELL_X2 FILLER_47_1250 ();
 FILLCELL_X1 FILLER_47_1252 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X16 FILLER_48_193 ();
 FILLCELL_X4 FILLER_48_209 ();
 FILLCELL_X8 FILLER_48_267 ();
 FILLCELL_X8 FILLER_48_282 ();
 FILLCELL_X2 FILLER_48_290 ();
 FILLCELL_X1 FILLER_48_292 ();
 FILLCELL_X1 FILLER_48_327 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X16 FILLER_48_385 ();
 FILLCELL_X2 FILLER_48_401 ();
 FILLCELL_X1 FILLER_48_403 ();
 FILLCELL_X1 FILLER_48_408 ();
 FILLCELL_X2 FILLER_48_418 ();
 FILLCELL_X8 FILLER_48_423 ();
 FILLCELL_X2 FILLER_48_431 ();
 FILLCELL_X1 FILLER_48_433 ();
 FILLCELL_X8 FILLER_48_437 ();
 FILLCELL_X4 FILLER_48_445 ();
 FILLCELL_X4 FILLER_48_456 ();
 FILLCELL_X4 FILLER_48_480 ();
 FILLCELL_X1 FILLER_48_488 ();
 FILLCELL_X2 FILLER_48_492 ();
 FILLCELL_X1 FILLER_48_500 ();
 FILLCELL_X2 FILLER_48_507 ();
 FILLCELL_X2 FILLER_48_514 ();
 FILLCELL_X1 FILLER_48_527 ();
 FILLCELL_X1 FILLER_48_539 ();
 FILLCELL_X2 FILLER_48_545 ();
 FILLCELL_X1 FILLER_48_547 ();
 FILLCELL_X2 FILLER_48_552 ();
 FILLCELL_X1 FILLER_48_554 ();
 FILLCELL_X4 FILLER_48_579 ();
 FILLCELL_X2 FILLER_48_583 ();
 FILLCELL_X1 FILLER_48_585 ();
 FILLCELL_X4 FILLER_48_603 ();
 FILLCELL_X1 FILLER_48_607 ();
 FILLCELL_X4 FILLER_48_613 ();
 FILLCELL_X1 FILLER_48_617 ();
 FILLCELL_X1 FILLER_48_620 ();
 FILLCELL_X4 FILLER_48_632 ();
 FILLCELL_X1 FILLER_48_636 ();
 FILLCELL_X2 FILLER_48_651 ();
 FILLCELL_X1 FILLER_48_653 ();
 FILLCELL_X2 FILLER_48_659 ();
 FILLCELL_X1 FILLER_48_661 ();
 FILLCELL_X4 FILLER_48_669 ();
 FILLCELL_X1 FILLER_48_673 ();
 FILLCELL_X2 FILLER_48_690 ();
 FILLCELL_X4 FILLER_48_694 ();
 FILLCELL_X4 FILLER_48_705 ();
 FILLCELL_X2 FILLER_48_709 ();
 FILLCELL_X2 FILLER_48_713 ();
 FILLCELL_X1 FILLER_48_715 ();
 FILLCELL_X2 FILLER_48_733 ();
 FILLCELL_X1 FILLER_48_735 ();
 FILLCELL_X2 FILLER_48_743 ();
 FILLCELL_X1 FILLER_48_745 ();
 FILLCELL_X1 FILLER_48_751 ();
 FILLCELL_X8 FILLER_48_774 ();
 FILLCELL_X4 FILLER_48_782 ();
 FILLCELL_X1 FILLER_48_786 ();
 FILLCELL_X16 FILLER_48_827 ();
 FILLCELL_X2 FILLER_48_861 ();
 FILLCELL_X1 FILLER_48_868 ();
 FILLCELL_X2 FILLER_48_872 ();
 FILLCELL_X2 FILLER_48_878 ();
 FILLCELL_X2 FILLER_48_884 ();
 FILLCELL_X4 FILLER_48_893 ();
 FILLCELL_X1 FILLER_48_929 ();
 FILLCELL_X4 FILLER_48_950 ();
 FILLCELL_X1 FILLER_48_954 ();
 FILLCELL_X16 FILLER_48_965 ();
 FILLCELL_X2 FILLER_48_988 ();
 FILLCELL_X2 FILLER_48_1010 ();
 FILLCELL_X2 FILLER_48_1017 ();
 FILLCELL_X1 FILLER_48_1019 ();
 FILLCELL_X2 FILLER_48_1024 ();
 FILLCELL_X1 FILLER_48_1026 ();
 FILLCELL_X2 FILLER_48_1049 ();
 FILLCELL_X4 FILLER_48_1056 ();
 FILLCELL_X2 FILLER_48_1060 ();
 FILLCELL_X1 FILLER_48_1062 ();
 FILLCELL_X16 FILLER_48_1070 ();
 FILLCELL_X1 FILLER_48_1086 ();
 FILLCELL_X1 FILLER_48_1109 ();
 FILLCELL_X1 FILLER_48_1141 ();
 FILLCELL_X1 FILLER_48_1158 ();
 FILLCELL_X1 FILLER_48_1163 ();
 FILLCELL_X1 FILLER_48_1190 ();
 FILLCELL_X1 FILLER_48_1217 ();
 FILLCELL_X16 FILLER_48_1242 ();
 FILLCELL_X2 FILLER_48_1258 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X16 FILLER_49_161 ();
 FILLCELL_X8 FILLER_49_177 ();
 FILLCELL_X2 FILLER_49_193 ();
 FILLCELL_X1 FILLER_49_195 ();
 FILLCELL_X4 FILLER_49_223 ();
 FILLCELL_X16 FILLER_49_234 ();
 FILLCELL_X4 FILLER_49_250 ();
 FILLCELL_X1 FILLER_49_254 ();
 FILLCELL_X4 FILLER_49_262 ();
 FILLCELL_X2 FILLER_49_266 ();
 FILLCELL_X4 FILLER_49_302 ();
 FILLCELL_X2 FILLER_49_306 ();
 FILLCELL_X1 FILLER_49_308 ();
 FILLCELL_X4 FILLER_49_316 ();
 FILLCELL_X2 FILLER_49_320 ();
 FILLCELL_X8 FILLER_49_369 ();
 FILLCELL_X4 FILLER_49_377 ();
 FILLCELL_X8 FILLER_49_388 ();
 FILLCELL_X4 FILLER_49_396 ();
 FILLCELL_X2 FILLER_49_400 ();
 FILLCELL_X1 FILLER_49_402 ();
 FILLCELL_X2 FILLER_49_437 ();
 FILLCELL_X8 FILLER_49_448 ();
 FILLCELL_X2 FILLER_49_456 ();
 FILLCELL_X1 FILLER_49_458 ();
 FILLCELL_X2 FILLER_49_474 ();
 FILLCELL_X4 FILLER_49_481 ();
 FILLCELL_X2 FILLER_49_485 ();
 FILLCELL_X2 FILLER_49_491 ();
 FILLCELL_X1 FILLER_49_497 ();
 FILLCELL_X2 FILLER_49_507 ();
 FILLCELL_X1 FILLER_49_509 ();
 FILLCELL_X32 FILLER_49_525 ();
 FILLCELL_X1 FILLER_49_557 ();
 FILLCELL_X8 FILLER_49_565 ();
 FILLCELL_X1 FILLER_49_573 ();
 FILLCELL_X8 FILLER_49_605 ();
 FILLCELL_X4 FILLER_49_613 ();
 FILLCELL_X4 FILLER_49_632 ();
 FILLCELL_X8 FILLER_49_641 ();
 FILLCELL_X4 FILLER_49_649 ();
 FILLCELL_X1 FILLER_49_653 ();
 FILLCELL_X4 FILLER_49_659 ();
 FILLCELL_X8 FILLER_49_679 ();
 FILLCELL_X4 FILLER_49_687 ();
 FILLCELL_X8 FILLER_49_694 ();
 FILLCELL_X1 FILLER_49_702 ();
 FILLCELL_X2 FILLER_49_712 ();
 FILLCELL_X8 FILLER_49_730 ();
 FILLCELL_X4 FILLER_49_738 ();
 FILLCELL_X4 FILLER_49_771 ();
 FILLCELL_X2 FILLER_49_775 ();
 FILLCELL_X1 FILLER_49_777 ();
 FILLCELL_X16 FILLER_49_792 ();
 FILLCELL_X2 FILLER_49_817 ();
 FILLCELL_X1 FILLER_49_819 ();
 FILLCELL_X2 FILLER_49_829 ();
 FILLCELL_X4 FILLER_49_889 ();
 FILLCELL_X2 FILLER_49_893 ();
 FILLCELL_X1 FILLER_49_895 ();
 FILLCELL_X4 FILLER_49_905 ();
 FILLCELL_X2 FILLER_49_909 ();
 FILLCELL_X1 FILLER_49_911 ();
 FILLCELL_X1 FILLER_49_920 ();
 FILLCELL_X4 FILLER_49_928 ();
 FILLCELL_X8 FILLER_49_944 ();
 FILLCELL_X1 FILLER_49_952 ();
 FILLCELL_X1 FILLER_49_975 ();
 FILLCELL_X2 FILLER_49_981 ();
 FILLCELL_X2 FILLER_49_988 ();
 FILLCELL_X2 FILLER_49_997 ();
 FILLCELL_X1 FILLER_49_999 ();
 FILLCELL_X1 FILLER_49_1007 ();
 FILLCELL_X2 FILLER_49_1028 ();
 FILLCELL_X1 FILLER_49_1030 ();
 FILLCELL_X1 FILLER_49_1039 ();
 FILLCELL_X2 FILLER_49_1048 ();
 FILLCELL_X1 FILLER_49_1053 ();
 FILLCELL_X1 FILLER_49_1092 ();
 FILLCELL_X8 FILLER_49_1123 ();
 FILLCELL_X2 FILLER_49_1145 ();
 FILLCELL_X16 FILLER_49_1167 ();
 FILLCELL_X4 FILLER_49_1183 ();
 FILLCELL_X2 FILLER_49_1187 ();
 FILLCELL_X1 FILLER_49_1189 ();
 FILLCELL_X4 FILLER_49_1195 ();
 FILLCELL_X2 FILLER_49_1199 ();
 FILLCELL_X8 FILLER_49_1203 ();
 FILLCELL_X1 FILLER_49_1221 ();
 FILLCELL_X2 FILLER_49_1225 ();
 FILLCELL_X1 FILLER_49_1227 ();
 FILLCELL_X8 FILLER_49_1245 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X8 FILLER_50_161 ();
 FILLCELL_X4 FILLER_50_169 ();
 FILLCELL_X2 FILLER_50_200 ();
 FILLCELL_X4 FILLER_50_209 ();
 FILLCELL_X1 FILLER_50_213 ();
 FILLCELL_X8 FILLER_50_261 ();
 FILLCELL_X4 FILLER_50_269 ();
 FILLCELL_X1 FILLER_50_280 ();
 FILLCELL_X1 FILLER_50_288 ();
 FILLCELL_X2 FILLER_50_296 ();
 FILLCELL_X1 FILLER_50_305 ();
 FILLCELL_X8 FILLER_50_313 ();
 FILLCELL_X4 FILLER_50_321 ();
 FILLCELL_X2 FILLER_50_332 ();
 FILLCELL_X1 FILLER_50_334 ();
 FILLCELL_X2 FILLER_50_355 ();
 FILLCELL_X4 FILLER_50_364 ();
 FILLCELL_X2 FILLER_50_368 ();
 FILLCELL_X1 FILLER_50_370 ();
 FILLCELL_X4 FILLER_50_378 ();
 FILLCELL_X16 FILLER_50_402 ();
 FILLCELL_X4 FILLER_50_425 ();
 FILLCELL_X8 FILLER_50_431 ();
 FILLCELL_X2 FILLER_50_439 ();
 FILLCELL_X1 FILLER_50_441 ();
 FILLCELL_X1 FILLER_50_463 ();
 FILLCELL_X1 FILLER_50_471 ();
 FILLCELL_X4 FILLER_50_476 ();
 FILLCELL_X2 FILLER_50_480 ();
 FILLCELL_X1 FILLER_50_482 ();
 FILLCELL_X4 FILLER_50_494 ();
 FILLCELL_X2 FILLER_50_498 ();
 FILLCELL_X1 FILLER_50_503 ();
 FILLCELL_X4 FILLER_50_508 ();
 FILLCELL_X4 FILLER_50_523 ();
 FILLCELL_X1 FILLER_50_527 ();
 FILLCELL_X2 FILLER_50_532 ();
 FILLCELL_X4 FILLER_50_549 ();
 FILLCELL_X1 FILLER_50_553 ();
 FILLCELL_X4 FILLER_50_571 ();
 FILLCELL_X4 FILLER_50_592 ();
 FILLCELL_X1 FILLER_50_596 ();
 FILLCELL_X16 FILLER_50_614 ();
 FILLCELL_X1 FILLER_50_630 ();
 FILLCELL_X8 FILLER_50_632 ();
 FILLCELL_X1 FILLER_50_640 ();
 FILLCELL_X4 FILLER_50_652 ();
 FILLCELL_X1 FILLER_50_656 ();
 FILLCELL_X1 FILLER_50_664 ();
 FILLCELL_X2 FILLER_50_685 ();
 FILLCELL_X1 FILLER_50_700 ();
 FILLCELL_X4 FILLER_50_706 ();
 FILLCELL_X2 FILLER_50_710 ();
 FILLCELL_X1 FILLER_50_712 ();
 FILLCELL_X8 FILLER_50_768 ();
 FILLCELL_X2 FILLER_50_776 ();
 FILLCELL_X4 FILLER_50_784 ();
 FILLCELL_X2 FILLER_50_788 ();
 FILLCELL_X1 FILLER_50_790 ();
 FILLCELL_X16 FILLER_50_815 ();
 FILLCELL_X4 FILLER_50_831 ();
 FILLCELL_X1 FILLER_50_835 ();
 FILLCELL_X8 FILLER_50_860 ();
 FILLCELL_X4 FILLER_50_871 ();
 FILLCELL_X1 FILLER_50_875 ();
 FILLCELL_X8 FILLER_50_885 ();
 FILLCELL_X4 FILLER_50_893 ();
 FILLCELL_X2 FILLER_50_897 ();
 FILLCELL_X2 FILLER_50_914 ();
 FILLCELL_X1 FILLER_50_916 ();
 FILLCELL_X1 FILLER_50_931 ();
 FILLCELL_X4 FILLER_50_946 ();
 FILLCELL_X1 FILLER_50_950 ();
 FILLCELL_X1 FILLER_50_966 ();
 FILLCELL_X4 FILLER_50_972 ();
 FILLCELL_X2 FILLER_50_996 ();
 FILLCELL_X1 FILLER_50_998 ();
 FILLCELL_X8 FILLER_50_1004 ();
 FILLCELL_X4 FILLER_50_1012 ();
 FILLCELL_X2 FILLER_50_1016 ();
 FILLCELL_X8 FILLER_50_1030 ();
 FILLCELL_X4 FILLER_50_1044 ();
 FILLCELL_X2 FILLER_50_1048 ();
 FILLCELL_X8 FILLER_50_1059 ();
 FILLCELL_X1 FILLER_50_1074 ();
 FILLCELL_X8 FILLER_50_1104 ();
 FILLCELL_X4 FILLER_50_1112 ();
 FILLCELL_X1 FILLER_50_1120 ();
 FILLCELL_X2 FILLER_50_1127 ();
 FILLCELL_X4 FILLER_50_1131 ();
 FILLCELL_X8 FILLER_50_1174 ();
 FILLCELL_X2 FILLER_50_1182 ();
 FILLCELL_X1 FILLER_50_1184 ();
 FILLCELL_X1 FILLER_50_1204 ();
 FILLCELL_X8 FILLER_50_1222 ();
 FILLCELL_X1 FILLER_50_1234 ();
 FILLCELL_X2 FILLER_50_1241 ();
 FILLCELL_X8 FILLER_50_1250 ();
 FILLCELL_X2 FILLER_50_1258 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X16 FILLER_51_129 ();
 FILLCELL_X8 FILLER_51_145 ();
 FILLCELL_X1 FILLER_51_153 ();
 FILLCELL_X8 FILLER_51_161 ();
 FILLCELL_X2 FILLER_51_176 ();
 FILLCELL_X1 FILLER_51_178 ();
 FILLCELL_X4 FILLER_51_199 ();
 FILLCELL_X2 FILLER_51_203 ();
 FILLCELL_X4 FILLER_51_225 ();
 FILLCELL_X2 FILLER_51_229 ();
 FILLCELL_X4 FILLER_51_238 ();
 FILLCELL_X1 FILLER_51_242 ();
 FILLCELL_X1 FILLER_51_264 ();
 FILLCELL_X1 FILLER_51_272 ();
 FILLCELL_X1 FILLER_51_293 ();
 FILLCELL_X1 FILLER_51_301 ();
 FILLCELL_X4 FILLER_51_316 ();
 FILLCELL_X1 FILLER_51_320 ();
 FILLCELL_X4 FILLER_51_341 ();
 FILLCELL_X2 FILLER_51_345 ();
 FILLCELL_X2 FILLER_51_387 ();
 FILLCELL_X1 FILLER_51_393 ();
 FILLCELL_X2 FILLER_51_421 ();
 FILLCELL_X4 FILLER_51_427 ();
 FILLCELL_X1 FILLER_51_431 ();
 FILLCELL_X4 FILLER_51_437 ();
 FILLCELL_X1 FILLER_51_441 ();
 FILLCELL_X8 FILLER_51_446 ();
 FILLCELL_X1 FILLER_51_454 ();
 FILLCELL_X2 FILLER_51_459 ();
 FILLCELL_X8 FILLER_51_475 ();
 FILLCELL_X1 FILLER_51_486 ();
 FILLCELL_X4 FILLER_51_494 ();
 FILLCELL_X1 FILLER_51_498 ();
 FILLCELL_X2 FILLER_51_515 ();
 FILLCELL_X2 FILLER_51_525 ();
 FILLCELL_X1 FILLER_51_527 ();
 FILLCELL_X2 FILLER_51_532 ();
 FILLCELL_X1 FILLER_51_534 ();
 FILLCELL_X1 FILLER_51_538 ();
 FILLCELL_X8 FILLER_51_556 ();
 FILLCELL_X2 FILLER_51_564 ();
 FILLCELL_X1 FILLER_51_566 ();
 FILLCELL_X4 FILLER_51_574 ();
 FILLCELL_X2 FILLER_51_578 ();
 FILLCELL_X1 FILLER_51_580 ();
 FILLCELL_X2 FILLER_51_601 ();
 FILLCELL_X1 FILLER_51_603 ();
 FILLCELL_X2 FILLER_51_609 ();
 FILLCELL_X2 FILLER_51_622 ();
 FILLCELL_X8 FILLER_51_627 ();
 FILLCELL_X4 FILLER_51_642 ();
 FILLCELL_X8 FILLER_51_657 ();
 FILLCELL_X4 FILLER_51_665 ();
 FILLCELL_X8 FILLER_51_690 ();
 FILLCELL_X2 FILLER_51_741 ();
 FILLCELL_X16 FILLER_51_755 ();
 FILLCELL_X4 FILLER_51_771 ();
 FILLCELL_X8 FILLER_51_797 ();
 FILLCELL_X2 FILLER_51_805 ();
 FILLCELL_X1 FILLER_51_807 ();
 FILLCELL_X4 FILLER_51_819 ();
 FILLCELL_X1 FILLER_51_823 ();
 FILLCELL_X4 FILLER_51_828 ();
 FILLCELL_X1 FILLER_51_832 ();
 FILLCELL_X2 FILLER_51_835 ();
 FILLCELL_X4 FILLER_51_841 ();
 FILLCELL_X32 FILLER_51_875 ();
 FILLCELL_X2 FILLER_51_907 ();
 FILLCELL_X1 FILLER_51_909 ();
 FILLCELL_X4 FILLER_51_930 ();
 FILLCELL_X4 FILLER_51_980 ();
 FILLCELL_X2 FILLER_51_984 ();
 FILLCELL_X1 FILLER_51_991 ();
 FILLCELL_X1 FILLER_51_999 ();
 FILLCELL_X1 FILLER_51_1022 ();
 FILLCELL_X1 FILLER_51_1032 ();
 FILLCELL_X1 FILLER_51_1037 ();
 FILLCELL_X1 FILLER_51_1049 ();
 FILLCELL_X2 FILLER_51_1072 ();
 FILLCELL_X8 FILLER_51_1079 ();
 FILLCELL_X1 FILLER_51_1087 ();
 FILLCELL_X4 FILLER_51_1102 ();
 FILLCELL_X2 FILLER_51_1109 ();
 FILLCELL_X1 FILLER_51_1137 ();
 FILLCELL_X2 FILLER_51_1165 ();
 FILLCELL_X2 FILLER_51_1177 ();
 FILLCELL_X1 FILLER_51_1179 ();
 FILLCELL_X4 FILLER_51_1186 ();
 FILLCELL_X2 FILLER_51_1204 ();
 FILLCELL_X2 FILLER_51_1222 ();
 FILLCELL_X1 FILLER_51_1224 ();
 FILLCELL_X4 FILLER_51_1232 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X16 FILLER_52_129 ();
 FILLCELL_X2 FILLER_52_145 ();
 FILLCELL_X1 FILLER_52_147 ();
 FILLCELL_X2 FILLER_52_195 ();
 FILLCELL_X8 FILLER_52_204 ();
 FILLCELL_X4 FILLER_52_212 ();
 FILLCELL_X1 FILLER_52_216 ();
 FILLCELL_X1 FILLER_52_229 ();
 FILLCELL_X1 FILLER_52_250 ();
 FILLCELL_X2 FILLER_52_265 ();
 FILLCELL_X1 FILLER_52_267 ();
 FILLCELL_X8 FILLER_52_275 ();
 FILLCELL_X4 FILLER_52_283 ();
 FILLCELL_X2 FILLER_52_318 ();
 FILLCELL_X4 FILLER_52_327 ();
 FILLCELL_X2 FILLER_52_331 ();
 FILLCELL_X1 FILLER_52_333 ();
 FILLCELL_X2 FILLER_52_348 ();
 FILLCELL_X16 FILLER_52_357 ();
 FILLCELL_X4 FILLER_52_373 ();
 FILLCELL_X2 FILLER_52_377 ();
 FILLCELL_X16 FILLER_52_393 ();
 FILLCELL_X8 FILLER_52_409 ();
 FILLCELL_X4 FILLER_52_417 ();
 FILLCELL_X2 FILLER_52_421 ();
 FILLCELL_X2 FILLER_52_456 ();
 FILLCELL_X1 FILLER_52_458 ();
 FILLCELL_X1 FILLER_52_493 ();
 FILLCELL_X1 FILLER_52_498 ();
 FILLCELL_X1 FILLER_52_508 ();
 FILLCELL_X1 FILLER_52_518 ();
 FILLCELL_X1 FILLER_52_532 ();
 FILLCELL_X1 FILLER_52_539 ();
 FILLCELL_X2 FILLER_52_552 ();
 FILLCELL_X2 FILLER_52_585 ();
 FILLCELL_X1 FILLER_52_587 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X2 FILLER_52_650 ();
 FILLCELL_X8 FILLER_52_655 ();
 FILLCELL_X4 FILLER_52_663 ();
 FILLCELL_X4 FILLER_52_670 ();
 FILLCELL_X1 FILLER_52_674 ();
 FILLCELL_X2 FILLER_52_695 ();
 FILLCELL_X1 FILLER_52_697 ();
 FILLCELL_X8 FILLER_52_700 ();
 FILLCELL_X1 FILLER_52_708 ();
 FILLCELL_X4 FILLER_52_722 ();
 FILLCELL_X2 FILLER_52_726 ();
 FILLCELL_X1 FILLER_52_728 ();
 FILLCELL_X2 FILLER_52_750 ();
 FILLCELL_X1 FILLER_52_752 ();
 FILLCELL_X32 FILLER_52_755 ();
 FILLCELL_X8 FILLER_52_787 ();
 FILLCELL_X2 FILLER_52_795 ();
 FILLCELL_X1 FILLER_52_813 ();
 FILLCELL_X1 FILLER_52_818 ();
 FILLCELL_X4 FILLER_52_823 ();
 FILLCELL_X2 FILLER_52_827 ();
 FILLCELL_X1 FILLER_52_829 ();
 FILLCELL_X4 FILLER_52_859 ();
 FILLCELL_X4 FILLER_52_868 ();
 FILLCELL_X1 FILLER_52_872 ();
 FILLCELL_X4 FILLER_52_880 ();
 FILLCELL_X2 FILLER_52_895 ();
 FILLCELL_X1 FILLER_52_911 ();
 FILLCELL_X8 FILLER_52_924 ();
 FILLCELL_X4 FILLER_52_932 ();
 FILLCELL_X2 FILLER_52_936 ();
 FILLCELL_X1 FILLER_52_938 ();
 FILLCELL_X4 FILLER_52_944 ();
 FILLCELL_X2 FILLER_52_948 ();
 FILLCELL_X1 FILLER_52_950 ();
 FILLCELL_X2 FILLER_52_1014 ();
 FILLCELL_X1 FILLER_52_1023 ();
 FILLCELL_X16 FILLER_52_1027 ();
 FILLCELL_X4 FILLER_52_1043 ();
 FILLCELL_X2 FILLER_52_1047 ();
 FILLCELL_X2 FILLER_52_1052 ();
 FILLCELL_X1 FILLER_52_1054 ();
 FILLCELL_X4 FILLER_52_1060 ();
 FILLCELL_X2 FILLER_52_1064 ();
 FILLCELL_X16 FILLER_52_1073 ();
 FILLCELL_X16 FILLER_52_1092 ();
 FILLCELL_X4 FILLER_52_1125 ();
 FILLCELL_X4 FILLER_52_1139 ();
 FILLCELL_X4 FILLER_52_1149 ();
 FILLCELL_X2 FILLER_52_1153 ();
 FILLCELL_X16 FILLER_52_1169 ();
 FILLCELL_X4 FILLER_52_1185 ();
 FILLCELL_X4 FILLER_52_1209 ();
 FILLCELL_X2 FILLER_52_1250 ();
 FILLCELL_X1 FILLER_52_1252 ();
 FILLCELL_X1 FILLER_52_1256 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X16 FILLER_53_161 ();
 FILLCELL_X4 FILLER_53_177 ();
 FILLCELL_X2 FILLER_53_181 ();
 FILLCELL_X1 FILLER_53_183 ();
 FILLCELL_X4 FILLER_53_198 ();
 FILLCELL_X1 FILLER_53_202 ();
 FILLCELL_X1 FILLER_53_224 ();
 FILLCELL_X8 FILLER_53_266 ();
 FILLCELL_X2 FILLER_53_274 ();
 FILLCELL_X1 FILLER_53_276 ();
 FILLCELL_X2 FILLER_53_297 ();
 FILLCELL_X1 FILLER_53_306 ();
 FILLCELL_X4 FILLER_53_314 ();
 FILLCELL_X2 FILLER_53_338 ();
 FILLCELL_X4 FILLER_53_354 ();
 FILLCELL_X2 FILLER_53_358 ();
 FILLCELL_X1 FILLER_53_360 ();
 FILLCELL_X2 FILLER_53_379 ();
 FILLCELL_X1 FILLER_53_381 ();
 FILLCELL_X1 FILLER_53_396 ();
 FILLCELL_X2 FILLER_53_422 ();
 FILLCELL_X4 FILLER_53_431 ();
 FILLCELL_X1 FILLER_53_435 ();
 FILLCELL_X4 FILLER_53_470 ();
 FILLCELL_X4 FILLER_53_479 ();
 FILLCELL_X1 FILLER_53_483 ();
 FILLCELL_X1 FILLER_53_495 ();
 FILLCELL_X8 FILLER_53_517 ();
 FILLCELL_X2 FILLER_53_525 ();
 FILLCELL_X4 FILLER_53_534 ();
 FILLCELL_X1 FILLER_53_538 ();
 FILLCELL_X2 FILLER_53_545 ();
 FILLCELL_X1 FILLER_53_547 ();
 FILLCELL_X4 FILLER_53_550 ();
 FILLCELL_X1 FILLER_53_561 ();
 FILLCELL_X4 FILLER_53_579 ();
 FILLCELL_X4 FILLER_53_585 ();
 FILLCELL_X1 FILLER_53_589 ();
 FILLCELL_X4 FILLER_53_603 ();
 FILLCELL_X2 FILLER_53_607 ();
 FILLCELL_X1 FILLER_53_614 ();
 FILLCELL_X8 FILLER_53_622 ();
 FILLCELL_X4 FILLER_53_630 ();
 FILLCELL_X1 FILLER_53_634 ();
 FILLCELL_X4 FILLER_53_642 ();
 FILLCELL_X2 FILLER_53_646 ();
 FILLCELL_X1 FILLER_53_648 ();
 FILLCELL_X8 FILLER_53_653 ();
 FILLCELL_X4 FILLER_53_661 ();
 FILLCELL_X32 FILLER_53_672 ();
 FILLCELL_X2 FILLER_53_704 ();
 FILLCELL_X1 FILLER_53_716 ();
 FILLCELL_X16 FILLER_53_720 ();
 FILLCELL_X2 FILLER_53_736 ();
 FILLCELL_X8 FILLER_53_746 ();
 FILLCELL_X16 FILLER_53_772 ();
 FILLCELL_X2 FILLER_53_788 ();
 FILLCELL_X1 FILLER_53_790 ();
 FILLCELL_X4 FILLER_53_796 ();
 FILLCELL_X1 FILLER_53_800 ();
 FILLCELL_X1 FILLER_53_823 ();
 FILLCELL_X1 FILLER_53_837 ();
 FILLCELL_X2 FILLER_53_842 ();
 FILLCELL_X8 FILLER_53_849 ();
 FILLCELL_X4 FILLER_53_857 ();
 FILLCELL_X1 FILLER_53_861 ();
 FILLCELL_X16 FILLER_53_869 ();
 FILLCELL_X2 FILLER_53_885 ();
 FILLCELL_X2 FILLER_53_894 ();
 FILLCELL_X1 FILLER_53_896 ();
 FILLCELL_X4 FILLER_53_949 ();
 FILLCELL_X2 FILLER_53_953 ();
 FILLCELL_X1 FILLER_53_970 ();
 FILLCELL_X1 FILLER_53_991 ();
 FILLCELL_X8 FILLER_53_999 ();
 FILLCELL_X2 FILLER_53_1007 ();
 FILLCELL_X1 FILLER_53_1009 ();
 FILLCELL_X4 FILLER_53_1042 ();
 FILLCELL_X2 FILLER_53_1046 ();
 FILLCELL_X2 FILLER_53_1052 ();
 FILLCELL_X1 FILLER_53_1054 ();
 FILLCELL_X2 FILLER_53_1059 ();
 FILLCELL_X2 FILLER_53_1092 ();
 FILLCELL_X8 FILLER_53_1105 ();
 FILLCELL_X2 FILLER_53_1113 ();
 FILLCELL_X1 FILLER_53_1115 ();
 FILLCELL_X8 FILLER_53_1146 ();
 FILLCELL_X4 FILLER_53_1154 ();
 FILLCELL_X2 FILLER_53_1158 ();
 FILLCELL_X1 FILLER_53_1160 ();
 FILLCELL_X2 FILLER_53_1168 ();
 FILLCELL_X1 FILLER_53_1170 ();
 FILLCELL_X8 FILLER_53_1188 ();
 FILLCELL_X4 FILLER_53_1196 ();
 FILLCELL_X1 FILLER_53_1207 ();
 FILLCELL_X1 FILLER_53_1217 ();
 FILLCELL_X2 FILLER_53_1221 ();
 FILLCELL_X1 FILLER_53_1230 ();
 FILLCELL_X2 FILLER_53_1233 ();
 FILLCELL_X4 FILLER_53_1252 ();
 FILLCELL_X1 FILLER_53_1256 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X16 FILLER_54_129 ();
 FILLCELL_X8 FILLER_54_145 ();
 FILLCELL_X2 FILLER_54_153 ();
 FILLCELL_X4 FILLER_54_162 ();
 FILLCELL_X4 FILLER_54_186 ();
 FILLCELL_X1 FILLER_54_211 ();
 FILLCELL_X8 FILLER_54_226 ();
 FILLCELL_X2 FILLER_54_234 ();
 FILLCELL_X8 FILLER_54_243 ();
 FILLCELL_X4 FILLER_54_251 ();
 FILLCELL_X2 FILLER_54_255 ();
 FILLCELL_X8 FILLER_54_264 ();
 FILLCELL_X2 FILLER_54_272 ();
 FILLCELL_X4 FILLER_54_308 ();
 FILLCELL_X8 FILLER_54_321 ();
 FILLCELL_X2 FILLER_54_329 ();
 FILLCELL_X1 FILLER_54_331 ();
 FILLCELL_X4 FILLER_54_346 ();
 FILLCELL_X1 FILLER_54_357 ();
 FILLCELL_X4 FILLER_54_379 ();
 FILLCELL_X8 FILLER_54_397 ();
 FILLCELL_X32 FILLER_54_413 ();
 FILLCELL_X8 FILLER_54_445 ();
 FILLCELL_X4 FILLER_54_453 ();
 FILLCELL_X16 FILLER_54_474 ();
 FILLCELL_X1 FILLER_54_490 ();
 FILLCELL_X2 FILLER_54_495 ();
 FILLCELL_X8 FILLER_54_500 ();
 FILLCELL_X4 FILLER_54_525 ();
 FILLCELL_X2 FILLER_54_534 ();
 FILLCELL_X1 FILLER_54_536 ();
 FILLCELL_X2 FILLER_54_568 ();
 FILLCELL_X1 FILLER_54_570 ();
 FILLCELL_X8 FILLER_54_578 ();
 FILLCELL_X4 FILLER_54_586 ();
 FILLCELL_X1 FILLER_54_621 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X8 FILLER_54_632 ();
 FILLCELL_X4 FILLER_54_640 ();
 FILLCELL_X2 FILLER_54_644 ();
 FILLCELL_X1 FILLER_54_646 ();
 FILLCELL_X4 FILLER_54_673 ();
 FILLCELL_X4 FILLER_54_684 ();
 FILLCELL_X1 FILLER_54_688 ();
 FILLCELL_X8 FILLER_54_691 ();
 FILLCELL_X2 FILLER_54_715 ();
 FILLCELL_X16 FILLER_54_726 ();
 FILLCELL_X8 FILLER_54_742 ();
 FILLCELL_X2 FILLER_54_750 ();
 FILLCELL_X2 FILLER_54_758 ();
 FILLCELL_X1 FILLER_54_760 ();
 FILLCELL_X2 FILLER_54_785 ();
 FILLCELL_X4 FILLER_54_804 ();
 FILLCELL_X1 FILLER_54_808 ();
 FILLCELL_X2 FILLER_54_813 ();
 FILLCELL_X2 FILLER_54_822 ();
 FILLCELL_X2 FILLER_54_827 ();
 FILLCELL_X2 FILLER_54_834 ();
 FILLCELL_X1 FILLER_54_836 ();
 FILLCELL_X4 FILLER_54_840 ();
 FILLCELL_X1 FILLER_54_844 ();
 FILLCELL_X1 FILLER_54_857 ();
 FILLCELL_X2 FILLER_54_863 ();
 FILLCELL_X1 FILLER_54_865 ();
 FILLCELL_X1 FILLER_54_869 ();
 FILLCELL_X4 FILLER_54_873 ();
 FILLCELL_X2 FILLER_54_877 ();
 FILLCELL_X1 FILLER_54_879 ();
 FILLCELL_X1 FILLER_54_897 ();
 FILLCELL_X1 FILLER_54_901 ();
 FILLCELL_X4 FILLER_54_911 ();
 FILLCELL_X4 FILLER_54_927 ();
 FILLCELL_X1 FILLER_54_938 ();
 FILLCELL_X1 FILLER_54_942 ();
 FILLCELL_X2 FILLER_54_953 ();
 FILLCELL_X16 FILLER_54_980 ();
 FILLCELL_X2 FILLER_54_996 ();
 FILLCELL_X4 FILLER_54_1007 ();
 FILLCELL_X1 FILLER_54_1011 ();
 FILLCELL_X1 FILLER_54_1029 ();
 FILLCELL_X2 FILLER_54_1037 ();
 FILLCELL_X1 FILLER_54_1039 ();
 FILLCELL_X1 FILLER_54_1068 ();
 FILLCELL_X1 FILLER_54_1073 ();
 FILLCELL_X1 FILLER_54_1078 ();
 FILLCELL_X1 FILLER_54_1083 ();
 FILLCELL_X1 FILLER_54_1088 ();
 FILLCELL_X4 FILLER_54_1093 ();
 FILLCELL_X1 FILLER_54_1097 ();
 FILLCELL_X8 FILLER_54_1102 ();
 FILLCELL_X1 FILLER_54_1110 ();
 FILLCELL_X1 FILLER_54_1118 ();
 FILLCELL_X8 FILLER_54_1133 ();
 FILLCELL_X8 FILLER_54_1146 ();
 FILLCELL_X2 FILLER_54_1154 ();
 FILLCELL_X1 FILLER_54_1156 ();
 FILLCELL_X4 FILLER_54_1164 ();
 FILLCELL_X1 FILLER_54_1168 ();
 FILLCELL_X8 FILLER_54_1171 ();
 FILLCELL_X4 FILLER_54_1179 ();
 FILLCELL_X4 FILLER_54_1207 ();
 FILLCELL_X4 FILLER_54_1217 ();
 FILLCELL_X1 FILLER_54_1221 ();
 FILLCELL_X1 FILLER_54_1242 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X16 FILLER_55_129 ();
 FILLCELL_X4 FILLER_55_145 ();
 FILLCELL_X2 FILLER_55_149 ();
 FILLCELL_X1 FILLER_55_151 ();
 FILLCELL_X4 FILLER_55_172 ();
 FILLCELL_X2 FILLER_55_176 ();
 FILLCELL_X4 FILLER_55_185 ();
 FILLCELL_X2 FILLER_55_189 ();
 FILLCELL_X1 FILLER_55_191 ();
 FILLCELL_X16 FILLER_55_196 ();
 FILLCELL_X8 FILLER_55_212 ();
 FILLCELL_X1 FILLER_55_220 ();
 FILLCELL_X8 FILLER_55_230 ();
 FILLCELL_X1 FILLER_55_238 ();
 FILLCELL_X2 FILLER_55_259 ();
 FILLCELL_X1 FILLER_55_261 ();
 FILLCELL_X1 FILLER_55_276 ();
 FILLCELL_X2 FILLER_55_302 ();
 FILLCELL_X2 FILLER_55_312 ();
 FILLCELL_X1 FILLER_55_314 ();
 FILLCELL_X8 FILLER_55_324 ();
 FILLCELL_X2 FILLER_55_332 ();
 FILLCELL_X1 FILLER_55_334 ();
 FILLCELL_X1 FILLER_55_349 ();
 FILLCELL_X8 FILLER_55_357 ();
 FILLCELL_X4 FILLER_55_365 ();
 FILLCELL_X4 FILLER_55_380 ();
 FILLCELL_X1 FILLER_55_384 ();
 FILLCELL_X2 FILLER_55_392 ();
 FILLCELL_X2 FILLER_55_411 ();
 FILLCELL_X1 FILLER_55_413 ();
 FILLCELL_X16 FILLER_55_463 ();
 FILLCELL_X1 FILLER_55_479 ();
 FILLCELL_X2 FILLER_55_487 ();
 FILLCELL_X1 FILLER_55_489 ();
 FILLCELL_X2 FILLER_55_512 ();
 FILLCELL_X1 FILLER_55_514 ();
 FILLCELL_X2 FILLER_55_520 ();
 FILLCELL_X1 FILLER_55_522 ();
 FILLCELL_X16 FILLER_55_540 ();
 FILLCELL_X2 FILLER_55_556 ();
 FILLCELL_X4 FILLER_55_565 ();
 FILLCELL_X1 FILLER_55_586 ();
 FILLCELL_X1 FILLER_55_590 ();
 FILLCELL_X1 FILLER_55_598 ();
 FILLCELL_X1 FILLER_55_606 ();
 FILLCELL_X1 FILLER_55_624 ();
 FILLCELL_X16 FILLER_55_645 ();
 FILLCELL_X8 FILLER_55_661 ();
 FILLCELL_X2 FILLER_55_669 ();
 FILLCELL_X4 FILLER_55_683 ();
 FILLCELL_X1 FILLER_55_687 ();
 FILLCELL_X2 FILLER_55_710 ();
 FILLCELL_X1 FILLER_55_717 ();
 FILLCELL_X1 FILLER_55_720 ();
 FILLCELL_X1 FILLER_55_728 ();
 FILLCELL_X8 FILLER_55_733 ();
 FILLCELL_X2 FILLER_55_741 ();
 FILLCELL_X8 FILLER_55_752 ();
 FILLCELL_X2 FILLER_55_763 ();
 FILLCELL_X1 FILLER_55_765 ();
 FILLCELL_X2 FILLER_55_769 ();
 FILLCELL_X4 FILLER_55_785 ();
 FILLCELL_X1 FILLER_55_789 ();
 FILLCELL_X8 FILLER_55_821 ();
 FILLCELL_X2 FILLER_55_829 ();
 FILLCELL_X1 FILLER_55_831 ();
 FILLCELL_X2 FILLER_55_853 ();
 FILLCELL_X4 FILLER_55_859 ();
 FILLCELL_X2 FILLER_55_863 ();
 FILLCELL_X1 FILLER_55_874 ();
 FILLCELL_X4 FILLER_55_884 ();
 FILLCELL_X1 FILLER_55_888 ();
 FILLCELL_X2 FILLER_55_897 ();
 FILLCELL_X1 FILLER_55_903 ();
 FILLCELL_X2 FILLER_55_908 ();
 FILLCELL_X1 FILLER_55_929 ();
 FILLCELL_X4 FILLER_55_941 ();
 FILLCELL_X2 FILLER_55_945 ();
 FILLCELL_X1 FILLER_55_947 ();
 FILLCELL_X4 FILLER_55_956 ();
 FILLCELL_X1 FILLER_55_960 ();
 FILLCELL_X1 FILLER_55_966 ();
 FILLCELL_X16 FILLER_55_974 ();
 FILLCELL_X4 FILLER_55_990 ();
 FILLCELL_X8 FILLER_55_1018 ();
 FILLCELL_X1 FILLER_55_1026 ();
 FILLCELL_X8 FILLER_55_1034 ();
 FILLCELL_X1 FILLER_55_1042 ();
 FILLCELL_X2 FILLER_55_1060 ();
 FILLCELL_X1 FILLER_55_1062 ();
 FILLCELL_X1 FILLER_55_1066 ();
 FILLCELL_X4 FILLER_55_1098 ();
 FILLCELL_X4 FILLER_55_1109 ();
 FILLCELL_X2 FILLER_55_1113 ();
 FILLCELL_X1 FILLER_55_1115 ();
 FILLCELL_X2 FILLER_55_1137 ();
 FILLCELL_X1 FILLER_55_1144 ();
 FILLCELL_X4 FILLER_55_1156 ();
 FILLCELL_X2 FILLER_55_1160 ();
 FILLCELL_X1 FILLER_55_1175 ();
 FILLCELL_X2 FILLER_55_1186 ();
 FILLCELL_X1 FILLER_55_1230 ();
 FILLCELL_X1 FILLER_55_1247 ();
 FILLCELL_X4 FILLER_55_1251 ();
 FILLCELL_X2 FILLER_55_1255 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X16 FILLER_56_65 ();
 FILLCELL_X16 FILLER_56_147 ();
 FILLCELL_X8 FILLER_56_163 ();
 FILLCELL_X2 FILLER_56_171 ();
 FILLCELL_X4 FILLER_56_184 ();
 FILLCELL_X4 FILLER_56_249 ();
 FILLCELL_X2 FILLER_56_253 ();
 FILLCELL_X16 FILLER_56_289 ();
 FILLCELL_X16 FILLER_56_309 ();
 FILLCELL_X2 FILLER_56_325 ();
 FILLCELL_X1 FILLER_56_327 ();
 FILLCELL_X4 FILLER_56_355 ();
 FILLCELL_X2 FILLER_56_359 ();
 FILLCELL_X2 FILLER_56_388 ();
 FILLCELL_X1 FILLER_56_390 ();
 FILLCELL_X4 FILLER_56_411 ();
 FILLCELL_X2 FILLER_56_415 ();
 FILLCELL_X4 FILLER_56_424 ();
 FILLCELL_X2 FILLER_56_428 ();
 FILLCELL_X8 FILLER_56_450 ();
 FILLCELL_X4 FILLER_56_458 ();
 FILLCELL_X4 FILLER_56_499 ();
 FILLCELL_X8 FILLER_56_534 ();
 FILLCELL_X2 FILLER_56_542 ();
 FILLCELL_X1 FILLER_56_544 ();
 FILLCELL_X4 FILLER_56_552 ();
 FILLCELL_X2 FILLER_56_556 ();
 FILLCELL_X8 FILLER_56_565 ();
 FILLCELL_X2 FILLER_56_573 ();
 FILLCELL_X1 FILLER_56_575 ();
 FILLCELL_X4 FILLER_56_583 ();
 FILLCELL_X2 FILLER_56_587 ();
 FILLCELL_X2 FILLER_56_596 ();
 FILLCELL_X1 FILLER_56_605 ();
 FILLCELL_X1 FILLER_56_616 ();
 FILLCELL_X1 FILLER_56_632 ();
 FILLCELL_X8 FILLER_56_652 ();
 FILLCELL_X2 FILLER_56_660 ();
 FILLCELL_X1 FILLER_56_662 ();
 FILLCELL_X16 FILLER_56_681 ();
 FILLCELL_X4 FILLER_56_697 ();
 FILLCELL_X1 FILLER_56_701 ();
 FILLCELL_X8 FILLER_56_723 ();
 FILLCELL_X2 FILLER_56_740 ();
 FILLCELL_X1 FILLER_56_742 ();
 FILLCELL_X2 FILLER_56_749 ();
 FILLCELL_X16 FILLER_56_785 ();
 FILLCELL_X1 FILLER_56_801 ();
 FILLCELL_X2 FILLER_56_812 ();
 FILLCELL_X1 FILLER_56_837 ();
 FILLCELL_X2 FILLER_56_878 ();
 FILLCELL_X1 FILLER_56_880 ();
 FILLCELL_X8 FILLER_56_886 ();
 FILLCELL_X2 FILLER_56_894 ();
 FILLCELL_X1 FILLER_56_896 ();
 FILLCELL_X8 FILLER_56_901 ();
 FILLCELL_X1 FILLER_56_913 ();
 FILLCELL_X2 FILLER_56_926 ();
 FILLCELL_X2 FILLER_56_935 ();
 FILLCELL_X1 FILLER_56_937 ();
 FILLCELL_X2 FILLER_56_944 ();
 FILLCELL_X1 FILLER_56_970 ();
 FILLCELL_X4 FILLER_56_978 ();
 FILLCELL_X1 FILLER_56_982 ();
 FILLCELL_X4 FILLER_56_997 ();
 FILLCELL_X4 FILLER_56_1008 ();
 FILLCELL_X4 FILLER_56_1040 ();
 FILLCELL_X2 FILLER_56_1044 ();
 FILLCELL_X1 FILLER_56_1046 ();
 FILLCELL_X8 FILLER_56_1051 ();
 FILLCELL_X1 FILLER_56_1059 ();
 FILLCELL_X4 FILLER_56_1072 ();
 FILLCELL_X1 FILLER_56_1076 ();
 FILLCELL_X4 FILLER_56_1083 ();
 FILLCELL_X2 FILLER_56_1087 ();
 FILLCELL_X1 FILLER_56_1104 ();
 FILLCELL_X2 FILLER_56_1109 ();
 FILLCELL_X1 FILLER_56_1111 ();
 FILLCELL_X4 FILLER_56_1150 ();
 FILLCELL_X4 FILLER_56_1165 ();
 FILLCELL_X2 FILLER_56_1169 ();
 FILLCELL_X1 FILLER_56_1171 ();
 FILLCELL_X8 FILLER_56_1182 ();
 FILLCELL_X4 FILLER_56_1190 ();
 FILLCELL_X2 FILLER_56_1194 ();
 FILLCELL_X1 FILLER_56_1196 ();
 FILLCELL_X2 FILLER_56_1201 ();
 FILLCELL_X2 FILLER_56_1207 ();
 FILLCELL_X1 FILLER_56_1209 ();
 FILLCELL_X1 FILLER_56_1213 ();
 FILLCELL_X2 FILLER_56_1217 ();
 FILLCELL_X1 FILLER_56_1219 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X16 FILLER_57_65 ();
 FILLCELL_X8 FILLER_57_81 ();
 FILLCELL_X2 FILLER_57_89 ();
 FILLCELL_X1 FILLER_57_91 ();
 FILLCELL_X2 FILLER_57_119 ();
 FILLCELL_X1 FILLER_57_121 ();
 FILLCELL_X1 FILLER_57_182 ();
 FILLCELL_X4 FILLER_57_214 ();
 FILLCELL_X1 FILLER_57_218 ();
 FILLCELL_X16 FILLER_57_246 ();
 FILLCELL_X2 FILLER_57_262 ();
 FILLCELL_X1 FILLER_57_264 ();
 FILLCELL_X16 FILLER_57_302 ();
 FILLCELL_X2 FILLER_57_318 ();
 FILLCELL_X4 FILLER_57_354 ();
 FILLCELL_X8 FILLER_57_365 ();
 FILLCELL_X4 FILLER_57_373 ();
 FILLCELL_X1 FILLER_57_377 ();
 FILLCELL_X8 FILLER_57_422 ();
 FILLCELL_X4 FILLER_57_430 ();
 FILLCELL_X2 FILLER_57_434 ();
 FILLCELL_X8 FILLER_57_450 ();
 FILLCELL_X4 FILLER_57_458 ();
 FILLCELL_X1 FILLER_57_462 ();
 FILLCELL_X8 FILLER_57_490 ();
 FILLCELL_X4 FILLER_57_498 ();
 FILLCELL_X1 FILLER_57_526 ();
 FILLCELL_X4 FILLER_57_534 ();
 FILLCELL_X2 FILLER_57_538 ();
 FILLCELL_X1 FILLER_57_540 ();
 FILLCELL_X16 FILLER_57_558 ();
 FILLCELL_X4 FILLER_57_574 ();
 FILLCELL_X1 FILLER_57_578 ();
 FILLCELL_X2 FILLER_57_624 ();
 FILLCELL_X1 FILLER_57_626 ();
 FILLCELL_X4 FILLER_57_636 ();
 FILLCELL_X8 FILLER_57_653 ();
 FILLCELL_X4 FILLER_57_661 ();
 FILLCELL_X1 FILLER_57_665 ();
 FILLCELL_X2 FILLER_57_671 ();
 FILLCELL_X8 FILLER_57_691 ();
 FILLCELL_X8 FILLER_57_706 ();
 FILLCELL_X2 FILLER_57_714 ();
 FILLCELL_X8 FILLER_57_719 ();
 FILLCELL_X4 FILLER_57_727 ();
 FILLCELL_X4 FILLER_57_742 ();
 FILLCELL_X2 FILLER_57_746 ();
 FILLCELL_X16 FILLER_57_758 ();
 FILLCELL_X16 FILLER_57_788 ();
 FILLCELL_X2 FILLER_57_804 ();
 FILLCELL_X1 FILLER_57_806 ();
 FILLCELL_X8 FILLER_57_844 ();
 FILLCELL_X1 FILLER_57_852 ();
 FILLCELL_X4 FILLER_57_858 ();
 FILLCELL_X2 FILLER_57_869 ();
 FILLCELL_X4 FILLER_57_890 ();
 FILLCELL_X1 FILLER_57_894 ();
 FILLCELL_X16 FILLER_57_900 ();
 FILLCELL_X2 FILLER_57_916 ();
 FILLCELL_X2 FILLER_57_922 ();
 FILLCELL_X2 FILLER_57_945 ();
 FILLCELL_X1 FILLER_57_947 ();
 FILLCELL_X2 FILLER_57_952 ();
 FILLCELL_X4 FILLER_57_967 ();
 FILLCELL_X2 FILLER_57_971 ();
 FILLCELL_X8 FILLER_57_990 ();
 FILLCELL_X4 FILLER_57_998 ();
 FILLCELL_X1 FILLER_57_1002 ();
 FILLCELL_X4 FILLER_57_1036 ();
 FILLCELL_X1 FILLER_57_1059 ();
 FILLCELL_X4 FILLER_57_1066 ();
 FILLCELL_X2 FILLER_57_1097 ();
 FILLCELL_X8 FILLER_57_1109 ();
 FILLCELL_X2 FILLER_57_1117 ();
 FILLCELL_X2 FILLER_57_1129 ();
 FILLCELL_X4 FILLER_57_1145 ();
 FILLCELL_X1 FILLER_57_1149 ();
 FILLCELL_X8 FILLER_57_1155 ();
 FILLCELL_X2 FILLER_57_1174 ();
 FILLCELL_X2 FILLER_57_1198 ();
 FILLCELL_X1 FILLER_57_1200 ();
 FILLCELL_X1 FILLER_57_1205 ();
 FILLCELL_X4 FILLER_57_1216 ();
 FILLCELL_X4 FILLER_57_1226 ();
 FILLCELL_X2 FILLER_57_1230 ();
 FILLCELL_X2 FILLER_57_1246 ();
 FILLCELL_X2 FILLER_57_1255 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X4 FILLER_58_97 ();
 FILLCELL_X2 FILLER_58_101 ();
 FILLCELL_X8 FILLER_58_130 ();
 FILLCELL_X4 FILLER_58_138 ();
 FILLCELL_X1 FILLER_58_142 ();
 FILLCELL_X1 FILLER_58_150 ();
 FILLCELL_X2 FILLER_58_158 ();
 FILLCELL_X4 FILLER_58_167 ();
 FILLCELL_X8 FILLER_58_178 ();
 FILLCELL_X8 FILLER_58_193 ();
 FILLCELL_X1 FILLER_58_201 ();
 FILLCELL_X2 FILLER_58_209 ();
 FILLCELL_X4 FILLER_58_218 ();
 FILLCELL_X8 FILLER_58_229 ();
 FILLCELL_X1 FILLER_58_237 ();
 FILLCELL_X8 FILLER_58_258 ();
 FILLCELL_X4 FILLER_58_266 ();
 FILLCELL_X4 FILLER_58_277 ();
 FILLCELL_X2 FILLER_58_281 ();
 FILLCELL_X1 FILLER_58_283 ();
 FILLCELL_X2 FILLER_58_291 ();
 FILLCELL_X1 FILLER_58_300 ();
 FILLCELL_X2 FILLER_58_335 ();
 FILLCELL_X2 FILLER_58_344 ();
 FILLCELL_X1 FILLER_58_346 ();
 FILLCELL_X2 FILLER_58_374 ();
 FILLCELL_X1 FILLER_58_376 ();
 FILLCELL_X4 FILLER_58_405 ();
 FILLCELL_X2 FILLER_58_409 ();
 FILLCELL_X1 FILLER_58_411 ();
 FILLCELL_X4 FILLER_58_466 ();
 FILLCELL_X2 FILLER_58_470 ();
 FILLCELL_X1 FILLER_58_472 ();
 FILLCELL_X16 FILLER_58_486 ();
 FILLCELL_X4 FILLER_58_502 ();
 FILLCELL_X1 FILLER_58_523 ();
 FILLCELL_X8 FILLER_58_538 ();
 FILLCELL_X4 FILLER_58_546 ();
 FILLCELL_X1 FILLER_58_550 ();
 FILLCELL_X1 FILLER_58_558 ();
 FILLCELL_X4 FILLER_58_585 ();
 FILLCELL_X4 FILLER_58_608 ();
 FILLCELL_X2 FILLER_58_612 ();
 FILLCELL_X1 FILLER_58_614 ();
 FILLCELL_X2 FILLER_58_632 ();
 FILLCELL_X2 FILLER_58_643 ();
 FILLCELL_X1 FILLER_58_645 ();
 FILLCELL_X16 FILLER_58_660 ();
 FILLCELL_X4 FILLER_58_681 ();
 FILLCELL_X8 FILLER_58_692 ();
 FILLCELL_X2 FILLER_58_700 ();
 FILLCELL_X1 FILLER_58_720 ();
 FILLCELL_X2 FILLER_58_743 ();
 FILLCELL_X1 FILLER_58_745 ();
 FILLCELL_X8 FILLER_58_766 ();
 FILLCELL_X1 FILLER_58_774 ();
 FILLCELL_X16 FILLER_58_797 ();
 FILLCELL_X2 FILLER_58_813 ();
 FILLCELL_X1 FILLER_58_833 ();
 FILLCELL_X16 FILLER_58_840 ();
 FILLCELL_X8 FILLER_58_856 ();
 FILLCELL_X1 FILLER_58_881 ();
 FILLCELL_X4 FILLER_58_918 ();
 FILLCELL_X2 FILLER_58_922 ();
 FILLCELL_X1 FILLER_58_924 ();
 FILLCELL_X16 FILLER_58_928 ();
 FILLCELL_X8 FILLER_58_944 ();
 FILLCELL_X2 FILLER_58_952 ();
 FILLCELL_X1 FILLER_58_954 ();
 FILLCELL_X2 FILLER_58_958 ();
 FILLCELL_X1 FILLER_58_965 ();
 FILLCELL_X2 FILLER_58_971 ();
 FILLCELL_X2 FILLER_58_976 ();
 FILLCELL_X1 FILLER_58_981 ();
 FILLCELL_X2 FILLER_58_989 ();
 FILLCELL_X2 FILLER_58_997 ();
 FILLCELL_X8 FILLER_58_1023 ();
 FILLCELL_X8 FILLER_58_1038 ();
 FILLCELL_X2 FILLER_58_1046 ();
 FILLCELL_X1 FILLER_58_1048 ();
 FILLCELL_X4 FILLER_58_1056 ();
 FILLCELL_X2 FILLER_58_1060 ();
 FILLCELL_X1 FILLER_58_1062 ();
 FILLCELL_X4 FILLER_58_1067 ();
 FILLCELL_X2 FILLER_58_1071 ();
 FILLCELL_X1 FILLER_58_1073 ();
 FILLCELL_X4 FILLER_58_1081 ();
 FILLCELL_X1 FILLER_58_1085 ();
 FILLCELL_X1 FILLER_58_1112 ();
 FILLCELL_X4 FILLER_58_1117 ();
 FILLCELL_X8 FILLER_58_1128 ();
 FILLCELL_X1 FILLER_58_1144 ();
 FILLCELL_X1 FILLER_58_1150 ();
 FILLCELL_X1 FILLER_58_1156 ();
 FILLCELL_X2 FILLER_58_1164 ();
 FILLCELL_X4 FILLER_58_1183 ();
 FILLCELL_X4 FILLER_58_1193 ();
 FILLCELL_X1 FILLER_58_1197 ();
 FILLCELL_X1 FILLER_58_1223 ();
 FILLCELL_X1 FILLER_58_1231 ();
 FILLCELL_X1 FILLER_58_1259 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X16 FILLER_59_33 ();
 FILLCELL_X2 FILLER_59_49 ();
 FILLCELL_X2 FILLER_59_58 ();
 FILLCELL_X1 FILLER_59_60 ();
 FILLCELL_X16 FILLER_59_88 ();
 FILLCELL_X2 FILLER_59_104 ();
 FILLCELL_X1 FILLER_59_106 ();
 FILLCELL_X2 FILLER_59_115 ();
 FILLCELL_X1 FILLER_59_117 ();
 FILLCELL_X4 FILLER_59_145 ();
 FILLCELL_X2 FILLER_59_189 ();
 FILLCELL_X2 FILLER_59_198 ();
 FILLCELL_X4 FILLER_59_207 ();
 FILLCELL_X1 FILLER_59_211 ();
 FILLCELL_X1 FILLER_59_226 ();
 FILLCELL_X1 FILLER_59_255 ();
 FILLCELL_X8 FILLER_59_302 ();
 FILLCELL_X4 FILLER_59_310 ();
 FILLCELL_X2 FILLER_59_314 ();
 FILLCELL_X16 FILLER_59_323 ();
 FILLCELL_X1 FILLER_59_339 ();
 FILLCELL_X2 FILLER_59_360 ();
 FILLCELL_X1 FILLER_59_362 ();
 FILLCELL_X2 FILLER_59_397 ();
 FILLCELL_X16 FILLER_59_419 ();
 FILLCELL_X8 FILLER_59_469 ();
 FILLCELL_X2 FILLER_59_477 ();
 FILLCELL_X8 FILLER_59_513 ();
 FILLCELL_X2 FILLER_59_538 ();
 FILLCELL_X1 FILLER_59_540 ();
 FILLCELL_X8 FILLER_59_597 ();
 FILLCELL_X2 FILLER_59_605 ();
 FILLCELL_X1 FILLER_59_637 ();
 FILLCELL_X8 FILLER_59_647 ();
 FILLCELL_X1 FILLER_59_655 ();
 FILLCELL_X2 FILLER_59_672 ();
 FILLCELL_X1 FILLER_59_674 ();
 FILLCELL_X2 FILLER_59_691 ();
 FILLCELL_X1 FILLER_59_693 ();
 FILLCELL_X8 FILLER_59_715 ();
 FILLCELL_X2 FILLER_59_723 ();
 FILLCELL_X1 FILLER_59_725 ();
 FILLCELL_X32 FILLER_59_730 ();
 FILLCELL_X1 FILLER_59_762 ();
 FILLCELL_X4 FILLER_59_785 ();
 FILLCELL_X1 FILLER_59_789 ();
 FILLCELL_X8 FILLER_59_793 ();
 FILLCELL_X32 FILLER_59_819 ();
 FILLCELL_X8 FILLER_59_851 ();
 FILLCELL_X8 FILLER_59_892 ();
 FILLCELL_X2 FILLER_59_900 ();
 FILLCELL_X1 FILLER_59_902 ();
 FILLCELL_X4 FILLER_59_915 ();
 FILLCELL_X1 FILLER_59_919 ();
 FILLCELL_X4 FILLER_59_924 ();
 FILLCELL_X1 FILLER_59_974 ();
 FILLCELL_X1 FILLER_59_985 ();
 FILLCELL_X2 FILLER_59_991 ();
 FILLCELL_X1 FILLER_59_993 ();
 FILLCELL_X1 FILLER_59_1011 ();
 FILLCELL_X2 FILLER_59_1019 ();
 FILLCELL_X8 FILLER_59_1028 ();
 FILLCELL_X2 FILLER_59_1036 ();
 FILLCELL_X1 FILLER_59_1038 ();
 FILLCELL_X8 FILLER_59_1046 ();
 FILLCELL_X2 FILLER_59_1054 ();
 FILLCELL_X1 FILLER_59_1056 ();
 FILLCELL_X8 FILLER_59_1078 ();
 FILLCELL_X4 FILLER_59_1086 ();
 FILLCELL_X1 FILLER_59_1098 ();
 FILLCELL_X4 FILLER_59_1103 ();
 FILLCELL_X1 FILLER_59_1129 ();
 FILLCELL_X1 FILLER_59_1136 ();
 FILLCELL_X4 FILLER_59_1157 ();
 FILLCELL_X2 FILLER_59_1161 ();
 FILLCELL_X4 FILLER_59_1190 ();
 FILLCELL_X2 FILLER_59_1221 ();
 FILLCELL_X2 FILLER_59_1257 ();
 FILLCELL_X1 FILLER_59_1259 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X8 FILLER_60_33 ();
 FILLCELL_X4 FILLER_60_41 ();
 FILLCELL_X2 FILLER_60_45 ();
 FILLCELL_X1 FILLER_60_67 ();
 FILLCELL_X2 FILLER_60_88 ();
 FILLCELL_X4 FILLER_60_124 ();
 FILLCELL_X1 FILLER_60_128 ();
 FILLCELL_X32 FILLER_60_143 ();
 FILLCELL_X1 FILLER_60_175 ();
 FILLCELL_X4 FILLER_60_183 ();
 FILLCELL_X2 FILLER_60_187 ();
 FILLCELL_X8 FILLER_60_209 ();
 FILLCELL_X1 FILLER_60_231 ();
 FILLCELL_X16 FILLER_60_260 ();
 FILLCELL_X2 FILLER_60_276 ();
 FILLCELL_X8 FILLER_60_291 ();
 FILLCELL_X2 FILLER_60_299 ();
 FILLCELL_X2 FILLER_60_344 ();
 FILLCELL_X1 FILLER_60_346 ();
 FILLCELL_X1 FILLER_60_354 ();
 FILLCELL_X2 FILLER_60_382 ();
 FILLCELL_X1 FILLER_60_384 ();
 FILLCELL_X8 FILLER_60_399 ();
 FILLCELL_X2 FILLER_60_407 ();
 FILLCELL_X2 FILLER_60_456 ();
 FILLCELL_X1 FILLER_60_458 ();
 FILLCELL_X16 FILLER_60_485 ();
 FILLCELL_X4 FILLER_60_501 ();
 FILLCELL_X2 FILLER_60_505 ();
 FILLCELL_X4 FILLER_60_524 ();
 FILLCELL_X1 FILLER_60_528 ();
 FILLCELL_X16 FILLER_60_540 ();
 FILLCELL_X8 FILLER_60_592 ();
 FILLCELL_X4 FILLER_60_600 ();
 FILLCELL_X2 FILLER_60_604 ();
 FILLCELL_X4 FILLER_60_624 ();
 FILLCELL_X2 FILLER_60_628 ();
 FILLCELL_X1 FILLER_60_630 ();
 FILLCELL_X1 FILLER_60_632 ();
 FILLCELL_X4 FILLER_60_640 ();
 FILLCELL_X1 FILLER_60_644 ();
 FILLCELL_X2 FILLER_60_654 ();
 FILLCELL_X2 FILLER_60_669 ();
 FILLCELL_X4 FILLER_60_684 ();
 FILLCELL_X4 FILLER_60_706 ();
 FILLCELL_X2 FILLER_60_710 ();
 FILLCELL_X1 FILLER_60_712 ();
 FILLCELL_X2 FILLER_60_719 ();
 FILLCELL_X4 FILLER_60_725 ();
 FILLCELL_X8 FILLER_60_738 ();
 FILLCELL_X1 FILLER_60_746 ();
 FILLCELL_X4 FILLER_60_756 ();
 FILLCELL_X1 FILLER_60_778 ();
 FILLCELL_X4 FILLER_60_823 ();
 FILLCELL_X2 FILLER_60_844 ();
 FILLCELL_X4 FILLER_60_883 ();
 FILLCELL_X1 FILLER_60_887 ();
 FILLCELL_X1 FILLER_60_908 ();
 FILLCELL_X8 FILLER_60_927 ();
 FILLCELL_X1 FILLER_60_935 ();
 FILLCELL_X4 FILLER_60_947 ();
 FILLCELL_X2 FILLER_60_951 ();
 FILLCELL_X1 FILLER_60_980 ();
 FILLCELL_X1 FILLER_60_987 ();
 FILLCELL_X1 FILLER_60_991 ();
 FILLCELL_X1 FILLER_60_998 ();
 FILLCELL_X8 FILLER_60_1012 ();
 FILLCELL_X4 FILLER_60_1020 ();
 FILLCELL_X2 FILLER_60_1024 ();
 FILLCELL_X1 FILLER_60_1026 ();
 FILLCELL_X1 FILLER_60_1034 ();
 FILLCELL_X2 FILLER_60_1056 ();
 FILLCELL_X2 FILLER_60_1063 ();
 FILLCELL_X2 FILLER_60_1072 ();
 FILLCELL_X2 FILLER_60_1078 ();
 FILLCELL_X1 FILLER_60_1097 ();
 FILLCELL_X4 FILLER_60_1134 ();
 FILLCELL_X8 FILLER_60_1158 ();
 FILLCELL_X2 FILLER_60_1166 ();
 FILLCELL_X1 FILLER_60_1168 ();
 FILLCELL_X4 FILLER_60_1187 ();
 FILLCELL_X2 FILLER_60_1191 ();
 FILLCELL_X1 FILLER_60_1193 ();
 FILLCELL_X2 FILLER_60_1201 ();
 FILLCELL_X1 FILLER_60_1203 ();
 FILLCELL_X2 FILLER_60_1254 ();
 FILLCELL_X1 FILLER_60_1256 ();
 FILLCELL_X16 FILLER_61_1 ();
 FILLCELL_X8 FILLER_61_17 ();
 FILLCELL_X4 FILLER_61_25 ();
 FILLCELL_X16 FILLER_61_56 ();
 FILLCELL_X4 FILLER_61_72 ();
 FILLCELL_X8 FILLER_61_83 ();
 FILLCELL_X4 FILLER_61_91 ();
 FILLCELL_X2 FILLER_61_95 ();
 FILLCELL_X2 FILLER_61_104 ();
 FILLCELL_X1 FILLER_61_106 ();
 FILLCELL_X1 FILLER_61_121 ();
 FILLCELL_X8 FILLER_61_143 ();
 FILLCELL_X2 FILLER_61_151 ();
 FILLCELL_X2 FILLER_61_160 ();
 FILLCELL_X8 FILLER_61_189 ();
 FILLCELL_X2 FILLER_61_197 ();
 FILLCELL_X1 FILLER_61_199 ();
 FILLCELL_X8 FILLER_61_207 ();
 FILLCELL_X4 FILLER_61_215 ();
 FILLCELL_X2 FILLER_61_219 ();
 FILLCELL_X2 FILLER_61_241 ();
 FILLCELL_X2 FILLER_61_253 ();
 FILLCELL_X1 FILLER_61_255 ();
 FILLCELL_X8 FILLER_61_296 ();
 FILLCELL_X1 FILLER_61_304 ();
 FILLCELL_X2 FILLER_61_312 ();
 FILLCELL_X1 FILLER_61_334 ();
 FILLCELL_X1 FILLER_61_355 ();
 FILLCELL_X1 FILLER_61_380 ();
 FILLCELL_X8 FILLER_61_422 ();
 FILLCELL_X4 FILLER_61_430 ();
 FILLCELL_X2 FILLER_61_434 ();
 FILLCELL_X4 FILLER_61_443 ();
 FILLCELL_X2 FILLER_61_447 ();
 FILLCELL_X32 FILLER_61_488 ();
 FILLCELL_X8 FILLER_61_551 ();
 FILLCELL_X4 FILLER_61_559 ();
 FILLCELL_X1 FILLER_61_563 ();
 FILLCELL_X2 FILLER_61_583 ();
 FILLCELL_X8 FILLER_61_604 ();
 FILLCELL_X1 FILLER_61_612 ();
 FILLCELL_X1 FILLER_61_624 ();
 FILLCELL_X2 FILLER_61_661 ();
 FILLCELL_X1 FILLER_61_663 ();
 FILLCELL_X16 FILLER_61_668 ();
 FILLCELL_X2 FILLER_61_684 ();
 FILLCELL_X1 FILLER_61_719 ();
 FILLCELL_X16 FILLER_61_724 ();
 FILLCELL_X1 FILLER_61_740 ();
 FILLCELL_X8 FILLER_61_747 ();
 FILLCELL_X2 FILLER_61_755 ();
 FILLCELL_X16 FILLER_61_769 ();
 FILLCELL_X8 FILLER_61_792 ();
 FILLCELL_X1 FILLER_61_800 ();
 FILLCELL_X2 FILLER_61_808 ();
 FILLCELL_X1 FILLER_61_810 ();
 FILLCELL_X1 FILLER_61_828 ();
 FILLCELL_X8 FILLER_61_855 ();
 FILLCELL_X1 FILLER_61_863 ();
 FILLCELL_X8 FILLER_61_871 ();
 FILLCELL_X1 FILLER_61_879 ();
 FILLCELL_X2 FILLER_61_883 ();
 FILLCELL_X1 FILLER_61_892 ();
 FILLCELL_X1 FILLER_61_896 ();
 FILLCELL_X2 FILLER_61_904 ();
 FILLCELL_X1 FILLER_61_906 ();
 FILLCELL_X2 FILLER_61_934 ();
 FILLCELL_X4 FILLER_61_941 ();
 FILLCELL_X4 FILLER_61_952 ();
 FILLCELL_X4 FILLER_61_963 ();
 FILLCELL_X2 FILLER_61_972 ();
 FILLCELL_X1 FILLER_61_981 ();
 FILLCELL_X4 FILLER_61_993 ();
 FILLCELL_X1 FILLER_61_997 ();
 FILLCELL_X16 FILLER_61_1036 ();
 FILLCELL_X8 FILLER_61_1052 ();
 FILLCELL_X4 FILLER_61_1060 ();
 FILLCELL_X2 FILLER_61_1064 ();
 FILLCELL_X1 FILLER_61_1066 ();
 FILLCELL_X1 FILLER_61_1090 ();
 FILLCELL_X8 FILLER_61_1096 ();
 FILLCELL_X1 FILLER_61_1108 ();
 FILLCELL_X8 FILLER_61_1111 ();
 FILLCELL_X1 FILLER_61_1119 ();
 FILLCELL_X8 FILLER_61_1123 ();
 FILLCELL_X4 FILLER_61_1131 ();
 FILLCELL_X1 FILLER_61_1135 ();
 FILLCELL_X8 FILLER_61_1141 ();
 FILLCELL_X4 FILLER_61_1149 ();
 FILLCELL_X8 FILLER_61_1179 ();
 FILLCELL_X1 FILLER_61_1187 ();
 FILLCELL_X1 FILLER_61_1205 ();
 FILLCELL_X4 FILLER_61_1213 ();
 FILLCELL_X1 FILLER_61_1236 ();
 FILLCELL_X1 FILLER_61_1240 ();
 FILLCELL_X1 FILLER_61_1248 ();
 FILLCELL_X1 FILLER_61_1259 ();
 FILLCELL_X16 FILLER_62_1 ();
 FILLCELL_X8 FILLER_62_17 ();
 FILLCELL_X2 FILLER_62_25 ();
 FILLCELL_X1 FILLER_62_27 ();
 FILLCELL_X8 FILLER_62_69 ();
 FILLCELL_X1 FILLER_62_77 ();
 FILLCELL_X16 FILLER_62_99 ();
 FILLCELL_X1 FILLER_62_122 ();
 FILLCELL_X2 FILLER_62_130 ();
 FILLCELL_X4 FILLER_62_139 ();
 FILLCELL_X4 FILLER_62_150 ();
 FILLCELL_X2 FILLER_62_174 ();
 FILLCELL_X1 FILLER_62_176 ();
 FILLCELL_X4 FILLER_62_198 ();
 FILLCELL_X2 FILLER_62_202 ();
 FILLCELL_X1 FILLER_62_204 ();
 FILLCELL_X16 FILLER_62_225 ();
 FILLCELL_X8 FILLER_62_241 ();
 FILLCELL_X4 FILLER_62_249 ();
 FILLCELL_X1 FILLER_62_253 ();
 FILLCELL_X4 FILLER_62_281 ();
 FILLCELL_X2 FILLER_62_285 ();
 FILLCELL_X1 FILLER_62_287 ();
 FILLCELL_X2 FILLER_62_295 ();
 FILLCELL_X1 FILLER_62_297 ();
 FILLCELL_X16 FILLER_62_305 ();
 FILLCELL_X1 FILLER_62_321 ();
 FILLCELL_X1 FILLER_62_329 ();
 FILLCELL_X8 FILLER_62_335 ();
 FILLCELL_X1 FILLER_62_343 ();
 FILLCELL_X2 FILLER_62_351 ();
 FILLCELL_X1 FILLER_62_353 ();
 FILLCELL_X4 FILLER_62_358 ();
 FILLCELL_X1 FILLER_62_362 ();
 FILLCELL_X2 FILLER_62_385 ();
 FILLCELL_X4 FILLER_62_396 ();
 FILLCELL_X4 FILLER_62_405 ();
 FILLCELL_X1 FILLER_62_416 ();
 FILLCELL_X1 FILLER_62_444 ();
 FILLCELL_X2 FILLER_62_452 ();
 FILLCELL_X1 FILLER_62_461 ();
 FILLCELL_X2 FILLER_62_469 ();
 FILLCELL_X2 FILLER_62_478 ();
 FILLCELL_X1 FILLER_62_480 ();
 FILLCELL_X8 FILLER_62_508 ();
 FILLCELL_X4 FILLER_62_516 ();
 FILLCELL_X8 FILLER_62_525 ();
 FILLCELL_X2 FILLER_62_533 ();
 FILLCELL_X1 FILLER_62_535 ();
 FILLCELL_X2 FILLER_62_539 ();
 FILLCELL_X4 FILLER_62_545 ();
 FILLCELL_X2 FILLER_62_552 ();
 FILLCELL_X1 FILLER_62_554 ();
 FILLCELL_X2 FILLER_62_571 ();
 FILLCELL_X1 FILLER_62_624 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X2 FILLER_62_632 ();
 FILLCELL_X2 FILLER_62_637 ();
 FILLCELL_X1 FILLER_62_639 ();
 FILLCELL_X2 FILLER_62_653 ();
 FILLCELL_X1 FILLER_62_655 ();
 FILLCELL_X2 FILLER_62_663 ();
 FILLCELL_X8 FILLER_62_681 ();
 FILLCELL_X4 FILLER_62_689 ();
 FILLCELL_X1 FILLER_62_693 ();
 FILLCELL_X1 FILLER_62_700 ();
 FILLCELL_X8 FILLER_62_708 ();
 FILLCELL_X8 FILLER_62_721 ();
 FILLCELL_X2 FILLER_62_729 ();
 FILLCELL_X32 FILLER_62_738 ();
 FILLCELL_X2 FILLER_62_770 ();
 FILLCELL_X1 FILLER_62_772 ();
 FILLCELL_X16 FILLER_62_795 ();
 FILLCELL_X8 FILLER_62_825 ();
 FILLCELL_X4 FILLER_62_833 ();
 FILLCELL_X2 FILLER_62_869 ();
 FILLCELL_X1 FILLER_62_871 ();
 FILLCELL_X2 FILLER_62_879 ();
 FILLCELL_X1 FILLER_62_881 ();
 FILLCELL_X2 FILLER_62_885 ();
 FILLCELL_X1 FILLER_62_887 ();
 FILLCELL_X16 FILLER_62_908 ();
 FILLCELL_X2 FILLER_62_924 ();
 FILLCELL_X1 FILLER_62_926 ();
 FILLCELL_X1 FILLER_62_967 ();
 FILLCELL_X8 FILLER_62_975 ();
 FILLCELL_X2 FILLER_62_983 ();
 FILLCELL_X1 FILLER_62_985 ();
 FILLCELL_X4 FILLER_62_998 ();
 FILLCELL_X2 FILLER_62_1009 ();
 FILLCELL_X1 FILLER_62_1011 ();
 FILLCELL_X4 FILLER_62_1019 ();
 FILLCELL_X2 FILLER_62_1023 ();
 FILLCELL_X2 FILLER_62_1069 ();
 FILLCELL_X2 FILLER_62_1087 ();
 FILLCELL_X1 FILLER_62_1089 ();
 FILLCELL_X1 FILLER_62_1108 ();
 FILLCELL_X8 FILLER_62_1123 ();
 FILLCELL_X4 FILLER_62_1131 ();
 FILLCELL_X1 FILLER_62_1135 ();
 FILLCELL_X2 FILLER_62_1153 ();
 FILLCELL_X2 FILLER_62_1169 ();
 FILLCELL_X1 FILLER_62_1171 ();
 FILLCELL_X8 FILLER_62_1181 ();
 FILLCELL_X2 FILLER_62_1189 ();
 FILLCELL_X1 FILLER_62_1191 ();
 FILLCELL_X4 FILLER_62_1201 ();
 FILLCELL_X2 FILLER_62_1205 ();
 FILLCELL_X4 FILLER_62_1212 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X8 FILLER_63_33 ();
 FILLCELL_X4 FILLER_63_41 ();
 FILLCELL_X1 FILLER_63_45 ();
 FILLCELL_X1 FILLER_63_70 ();
 FILLCELL_X1 FILLER_63_78 ();
 FILLCELL_X1 FILLER_63_93 ();
 FILLCELL_X1 FILLER_63_101 ();
 FILLCELL_X2 FILLER_63_122 ();
 FILLCELL_X1 FILLER_63_124 ();
 FILLCELL_X2 FILLER_63_132 ();
 FILLCELL_X1 FILLER_63_134 ();
 FILLCELL_X4 FILLER_63_142 ();
 FILLCELL_X2 FILLER_63_146 ();
 FILLCELL_X1 FILLER_63_148 ();
 FILLCELL_X4 FILLER_63_202 ();
 FILLCELL_X1 FILLER_63_206 ();
 FILLCELL_X16 FILLER_63_214 ();
 FILLCELL_X4 FILLER_63_230 ();
 FILLCELL_X2 FILLER_63_234 ();
 FILLCELL_X4 FILLER_63_263 ();
 FILLCELL_X1 FILLER_63_267 ();
 FILLCELL_X2 FILLER_63_295 ();
 FILLCELL_X2 FILLER_63_304 ();
 FILLCELL_X1 FILLER_63_306 ();
 FILLCELL_X4 FILLER_63_327 ();
 FILLCELL_X2 FILLER_63_331 ();
 FILLCELL_X1 FILLER_63_333 ();
 FILLCELL_X4 FILLER_63_341 ();
 FILLCELL_X1 FILLER_63_345 ();
 FILLCELL_X1 FILLER_63_353 ();
 FILLCELL_X2 FILLER_63_358 ();
 FILLCELL_X1 FILLER_63_360 ();
 FILLCELL_X4 FILLER_63_368 ();
 FILLCELL_X1 FILLER_63_372 ();
 FILLCELL_X4 FILLER_63_411 ();
 FILLCELL_X8 FILLER_63_435 ();
 FILLCELL_X4 FILLER_63_443 ();
 FILLCELL_X2 FILLER_63_447 ();
 FILLCELL_X4 FILLER_63_463 ();
 FILLCELL_X1 FILLER_63_467 ();
 FILLCELL_X8 FILLER_63_488 ();
 FILLCELL_X2 FILLER_63_496 ();
 FILLCELL_X1 FILLER_63_498 ();
 FILLCELL_X1 FILLER_63_530 ();
 FILLCELL_X2 FILLER_63_553 ();
 FILLCELL_X1 FILLER_63_555 ();
 FILLCELL_X4 FILLER_63_586 ();
 FILLCELL_X4 FILLER_63_601 ();
 FILLCELL_X2 FILLER_63_605 ();
 FILLCELL_X1 FILLER_63_607 ();
 FILLCELL_X8 FILLER_63_613 ();
 FILLCELL_X1 FILLER_63_621 ();
 FILLCELL_X1 FILLER_63_625 ();
 FILLCELL_X1 FILLER_63_636 ();
 FILLCELL_X1 FILLER_63_644 ();
 FILLCELL_X1 FILLER_63_658 ();
 FILLCELL_X2 FILLER_63_668 ();
 FILLCELL_X8 FILLER_63_684 ();
 FILLCELL_X1 FILLER_63_701 ();
 FILLCELL_X1 FILLER_63_724 ();
 FILLCELL_X2 FILLER_63_730 ();
 FILLCELL_X1 FILLER_63_732 ();
 FILLCELL_X16 FILLER_63_747 ();
 FILLCELL_X8 FILLER_63_763 ();
 FILLCELL_X2 FILLER_63_771 ();
 FILLCELL_X1 FILLER_63_773 ();
 FILLCELL_X1 FILLER_63_779 ();
 FILLCELL_X8 FILLER_63_794 ();
 FILLCELL_X16 FILLER_63_923 ();
 FILLCELL_X8 FILLER_63_939 ();
 FILLCELL_X2 FILLER_63_947 ();
 FILLCELL_X1 FILLER_63_949 ();
 FILLCELL_X8 FILLER_63_955 ();
 FILLCELL_X4 FILLER_63_963 ();
 FILLCELL_X4 FILLER_63_987 ();
 FILLCELL_X2 FILLER_63_1008 ();
 FILLCELL_X1 FILLER_63_1010 ();
 FILLCELL_X2 FILLER_63_1028 ();
 FILLCELL_X2 FILLER_63_1037 ();
 FILLCELL_X16 FILLER_63_1046 ();
 FILLCELL_X2 FILLER_63_1069 ();
 FILLCELL_X1 FILLER_63_1108 ();
 FILLCELL_X1 FILLER_63_1180 ();
 FILLCELL_X2 FILLER_63_1211 ();
 FILLCELL_X1 FILLER_63_1219 ();
 FILLCELL_X2 FILLER_63_1258 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X2 FILLER_64_33 ();
 FILLCELL_X2 FILLER_64_55 ();
 FILLCELL_X1 FILLER_64_82 ();
 FILLCELL_X1 FILLER_64_90 ();
 FILLCELL_X4 FILLER_64_98 ();
 FILLCELL_X2 FILLER_64_102 ();
 FILLCELL_X4 FILLER_64_111 ();
 FILLCELL_X4 FILLER_64_129 ();
 FILLCELL_X2 FILLER_64_133 ();
 FILLCELL_X1 FILLER_64_135 ();
 FILLCELL_X4 FILLER_64_150 ();
 FILLCELL_X2 FILLER_64_154 ();
 FILLCELL_X8 FILLER_64_163 ();
 FILLCELL_X4 FILLER_64_171 ();
 FILLCELL_X2 FILLER_64_175 ();
 FILLCELL_X1 FILLER_64_177 ();
 FILLCELL_X1 FILLER_64_188 ();
 FILLCELL_X1 FILLER_64_196 ();
 FILLCELL_X4 FILLER_64_204 ();
 FILLCELL_X2 FILLER_64_208 ();
 FILLCELL_X1 FILLER_64_210 ();
 FILLCELL_X4 FILLER_64_259 ();
 FILLCELL_X1 FILLER_64_277 ();
 FILLCELL_X1 FILLER_64_288 ();
 FILLCELL_X2 FILLER_64_296 ();
 FILLCELL_X2 FILLER_64_305 ();
 FILLCELL_X2 FILLER_64_314 ();
 FILLCELL_X1 FILLER_64_316 ();
 FILLCELL_X8 FILLER_64_364 ();
 FILLCELL_X2 FILLER_64_372 ();
 FILLCELL_X1 FILLER_64_374 ();
 FILLCELL_X32 FILLER_64_382 ();
 FILLCELL_X2 FILLER_64_414 ();
 FILLCELL_X1 FILLER_64_416 ();
 FILLCELL_X4 FILLER_64_424 ();
 FILLCELL_X2 FILLER_64_428 ();
 FILLCELL_X1 FILLER_64_430 ();
 FILLCELL_X1 FILLER_64_438 ();
 FILLCELL_X1 FILLER_64_442 ();
 FILLCELL_X8 FILLER_64_463 ();
 FILLCELL_X1 FILLER_64_471 ();
 FILLCELL_X4 FILLER_64_479 ();
 FILLCELL_X16 FILLER_64_503 ();
 FILLCELL_X2 FILLER_64_519 ();
 FILLCELL_X16 FILLER_64_533 ();
 FILLCELL_X4 FILLER_64_549 ();
 FILLCELL_X1 FILLER_64_553 ();
 FILLCELL_X8 FILLER_64_561 ();
 FILLCELL_X4 FILLER_64_569 ();
 FILLCELL_X2 FILLER_64_573 ();
 FILLCELL_X1 FILLER_64_575 ();
 FILLCELL_X2 FILLER_64_594 ();
 FILLCELL_X2 FILLER_64_610 ();
 FILLCELL_X1 FILLER_64_612 ();
 FILLCELL_X8 FILLER_64_641 ();
 FILLCELL_X1 FILLER_64_649 ();
 FILLCELL_X2 FILLER_64_659 ();
 FILLCELL_X1 FILLER_64_661 ();
 FILLCELL_X16 FILLER_64_671 ();
 FILLCELL_X4 FILLER_64_687 ();
 FILLCELL_X2 FILLER_64_691 ();
 FILLCELL_X2 FILLER_64_695 ();
 FILLCELL_X16 FILLER_64_732 ();
 FILLCELL_X4 FILLER_64_748 ();
 FILLCELL_X2 FILLER_64_752 ();
 FILLCELL_X1 FILLER_64_754 ();
 FILLCELL_X2 FILLER_64_779 ();
 FILLCELL_X1 FILLER_64_781 ();
 FILLCELL_X2 FILLER_64_812 ();
 FILLCELL_X4 FILLER_64_827 ();
 FILLCELL_X1 FILLER_64_851 ();
 FILLCELL_X1 FILLER_64_880 ();
 FILLCELL_X1 FILLER_64_884 ();
 FILLCELL_X4 FILLER_64_920 ();
 FILLCELL_X1 FILLER_64_924 ();
 FILLCELL_X1 FILLER_64_928 ();
 FILLCELL_X1 FILLER_64_949 ();
 FILLCELL_X4 FILLER_64_957 ();
 FILLCELL_X2 FILLER_64_961 ();
 FILLCELL_X16 FILLER_64_966 ();
 FILLCELL_X2 FILLER_64_1006 ();
 FILLCELL_X1 FILLER_64_1016 ();
 FILLCELL_X2 FILLER_64_1056 ();
 FILLCELL_X1 FILLER_64_1058 ();
 FILLCELL_X2 FILLER_64_1078 ();
 FILLCELL_X16 FILLER_64_1087 ();
 FILLCELL_X4 FILLER_64_1103 ();
 FILLCELL_X2 FILLER_64_1107 ();
 FILLCELL_X4 FILLER_64_1114 ();
 FILLCELL_X1 FILLER_64_1118 ();
 FILLCELL_X8 FILLER_64_1123 ();
 FILLCELL_X4 FILLER_64_1131 ();
 FILLCELL_X2 FILLER_64_1150 ();
 FILLCELL_X2 FILLER_64_1159 ();
 FILLCELL_X1 FILLER_64_1165 ();
 FILLCELL_X8 FILLER_64_1186 ();
 FILLCELL_X4 FILLER_64_1194 ();
 FILLCELL_X1 FILLER_64_1198 ();
 FILLCELL_X4 FILLER_64_1213 ();
 FILLCELL_X2 FILLER_64_1217 ();
 FILLCELL_X1 FILLER_64_1219 ();
 FILLCELL_X2 FILLER_64_1225 ();
 FILLCELL_X2 FILLER_64_1234 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X8 FILLER_65_33 ();
 FILLCELL_X4 FILLER_65_41 ();
 FILLCELL_X2 FILLER_65_45 ();
 FILLCELL_X8 FILLER_65_54 ();
 FILLCELL_X8 FILLER_65_69 ();
 FILLCELL_X2 FILLER_65_77 ();
 FILLCELL_X1 FILLER_65_79 ();
 FILLCELL_X1 FILLER_65_100 ();
 FILLCELL_X2 FILLER_65_108 ();
 FILLCELL_X1 FILLER_65_110 ();
 FILLCELL_X4 FILLER_65_135 ();
 FILLCELL_X1 FILLER_65_139 ();
 FILLCELL_X4 FILLER_65_160 ();
 FILLCELL_X1 FILLER_65_164 ();
 FILLCELL_X4 FILLER_65_192 ();
 FILLCELL_X1 FILLER_65_196 ();
 FILLCELL_X2 FILLER_65_204 ();
 FILLCELL_X1 FILLER_65_233 ();
 FILLCELL_X2 FILLER_65_244 ();
 FILLCELL_X16 FILLER_65_255 ();
 FILLCELL_X2 FILLER_65_271 ();
 FILLCELL_X1 FILLER_65_273 ();
 FILLCELL_X8 FILLER_65_306 ();
 FILLCELL_X4 FILLER_65_314 ();
 FILLCELL_X4 FILLER_65_325 ();
 FILLCELL_X2 FILLER_65_329 ();
 FILLCELL_X8 FILLER_65_344 ();
 FILLCELL_X4 FILLER_65_352 ();
 FILLCELL_X2 FILLER_65_356 ();
 FILLCELL_X1 FILLER_65_358 ();
 FILLCELL_X8 FILLER_65_366 ();
 FILLCELL_X1 FILLER_65_374 ();
 FILLCELL_X1 FILLER_65_407 ();
 FILLCELL_X4 FILLER_65_422 ();
 FILLCELL_X1 FILLER_65_426 ();
 FILLCELL_X8 FILLER_65_453 ();
 FILLCELL_X4 FILLER_65_461 ();
 FILLCELL_X8 FILLER_65_478 ();
 FILLCELL_X8 FILLER_65_493 ();
 FILLCELL_X8 FILLER_65_515 ();
 FILLCELL_X2 FILLER_65_523 ();
 FILLCELL_X8 FILLER_65_556 ();
 FILLCELL_X2 FILLER_65_564 ();
 FILLCELL_X16 FILLER_65_569 ();
 FILLCELL_X4 FILLER_65_585 ();
 FILLCELL_X2 FILLER_65_589 ();
 FILLCELL_X1 FILLER_65_600 ();
 FILLCELL_X1 FILLER_65_628 ();
 FILLCELL_X1 FILLER_65_633 ();
 FILLCELL_X1 FILLER_65_646 ();
 FILLCELL_X1 FILLER_65_656 ();
 FILLCELL_X2 FILLER_65_664 ();
 FILLCELL_X8 FILLER_65_679 ();
 FILLCELL_X4 FILLER_65_687 ();
 FILLCELL_X1 FILLER_65_691 ();
 FILLCELL_X1 FILLER_65_695 ();
 FILLCELL_X8 FILLER_65_720 ();
 FILLCELL_X1 FILLER_65_728 ();
 FILLCELL_X1 FILLER_65_743 ();
 FILLCELL_X8 FILLER_65_761 ();
 FILLCELL_X1 FILLER_65_769 ();
 FILLCELL_X8 FILLER_65_777 ();
 FILLCELL_X2 FILLER_65_785 ();
 FILLCELL_X1 FILLER_65_787 ();
 FILLCELL_X16 FILLER_65_801 ();
 FILLCELL_X4 FILLER_65_817 ();
 FILLCELL_X2 FILLER_65_834 ();
 FILLCELL_X2 FILLER_65_843 ();
 FILLCELL_X1 FILLER_65_845 ();
 FILLCELL_X8 FILLER_65_859 ();
 FILLCELL_X1 FILLER_65_867 ();
 FILLCELL_X4 FILLER_65_880 ();
 FILLCELL_X2 FILLER_65_889 ();
 FILLCELL_X1 FILLER_65_891 ();
 FILLCELL_X8 FILLER_65_895 ();
 FILLCELL_X2 FILLER_65_920 ();
 FILLCELL_X4 FILLER_65_925 ();
 FILLCELL_X4 FILLER_65_981 ();
 FILLCELL_X1 FILLER_65_985 ();
 FILLCELL_X8 FILLER_65_1006 ();
 FILLCELL_X4 FILLER_65_1014 ();
 FILLCELL_X2 FILLER_65_1018 ();
 FILLCELL_X1 FILLER_65_1020 ();
 FILLCELL_X8 FILLER_65_1028 ();
 FILLCELL_X1 FILLER_65_1044 ();
 FILLCELL_X4 FILLER_65_1055 ();
 FILLCELL_X2 FILLER_65_1059 ();
 FILLCELL_X1 FILLER_65_1061 ();
 FILLCELL_X8 FILLER_65_1069 ();
 FILLCELL_X4 FILLER_65_1077 ();
 FILLCELL_X1 FILLER_65_1081 ();
 FILLCELL_X1 FILLER_65_1123 ();
 FILLCELL_X2 FILLER_65_1127 ();
 FILLCELL_X8 FILLER_65_1135 ();
 FILLCELL_X4 FILLER_65_1143 ();
 FILLCELL_X4 FILLER_65_1151 ();
 FILLCELL_X2 FILLER_65_1167 ();
 FILLCELL_X4 FILLER_65_1188 ();
 FILLCELL_X2 FILLER_65_1192 ();
 FILLCELL_X2 FILLER_65_1197 ();
 FILLCELL_X1 FILLER_65_1209 ();
 FILLCELL_X1 FILLER_65_1214 ();
 FILLCELL_X1 FILLER_65_1221 ();
 FILLCELL_X1 FILLER_65_1228 ();
 FILLCELL_X2 FILLER_65_1232 ();
 FILLCELL_X1 FILLER_65_1234 ();
 FILLCELL_X2 FILLER_65_1243 ();
 FILLCELL_X16 FILLER_66_1 ();
 FILLCELL_X2 FILLER_66_17 ();
 FILLCELL_X8 FILLER_66_46 ();
 FILLCELL_X4 FILLER_66_54 ();
 FILLCELL_X2 FILLER_66_58 ();
 FILLCELL_X1 FILLER_66_80 ();
 FILLCELL_X16 FILLER_66_88 ();
 FILLCELL_X4 FILLER_66_104 ();
 FILLCELL_X2 FILLER_66_108 ();
 FILLCELL_X1 FILLER_66_110 ();
 FILLCELL_X2 FILLER_66_118 ();
 FILLCELL_X8 FILLER_66_156 ();
 FILLCELL_X4 FILLER_66_164 ();
 FILLCELL_X2 FILLER_66_175 ();
 FILLCELL_X1 FILLER_66_177 ();
 FILLCELL_X4 FILLER_66_198 ();
 FILLCELL_X2 FILLER_66_202 ();
 FILLCELL_X2 FILLER_66_211 ();
 FILLCELL_X1 FILLER_66_213 ();
 FILLCELL_X4 FILLER_66_221 ();
 FILLCELL_X2 FILLER_66_225 ();
 FILLCELL_X2 FILLER_66_240 ();
 FILLCELL_X1 FILLER_66_242 ();
 FILLCELL_X2 FILLER_66_257 ();
 FILLCELL_X4 FILLER_66_286 ();
 FILLCELL_X1 FILLER_66_297 ();
 FILLCELL_X1 FILLER_66_325 ();
 FILLCELL_X16 FILLER_66_367 ();
 FILLCELL_X4 FILLER_66_383 ();
 FILLCELL_X1 FILLER_66_387 ();
 FILLCELL_X1 FILLER_66_415 ();
 FILLCELL_X8 FILLER_66_444 ();
 FILLCELL_X4 FILLER_66_452 ();
 FILLCELL_X2 FILLER_66_456 ();
 FILLCELL_X1 FILLER_66_485 ();
 FILLCELL_X2 FILLER_66_496 ();
 FILLCELL_X2 FILLER_66_505 ();
 FILLCELL_X4 FILLER_66_514 ();
 FILLCELL_X2 FILLER_66_518 ();
 FILLCELL_X1 FILLER_66_520 ();
 FILLCELL_X2 FILLER_66_571 ();
 FILLCELL_X2 FILLER_66_604 ();
 FILLCELL_X1 FILLER_66_606 ();
 FILLCELL_X8 FILLER_66_613 ();
 FILLCELL_X4 FILLER_66_624 ();
 FILLCELL_X4 FILLER_66_674 ();
 FILLCELL_X1 FILLER_66_678 ();
 FILLCELL_X1 FILLER_66_701 ();
 FILLCELL_X2 FILLER_66_725 ();
 FILLCELL_X1 FILLER_66_727 ();
 FILLCELL_X1 FILLER_66_733 ();
 FILLCELL_X4 FILLER_66_738 ();
 FILLCELL_X1 FILLER_66_753 ();
 FILLCELL_X8 FILLER_66_765 ();
 FILLCELL_X2 FILLER_66_773 ();
 FILLCELL_X4 FILLER_66_796 ();
 FILLCELL_X8 FILLER_66_827 ();
 FILLCELL_X4 FILLER_66_835 ();
 FILLCELL_X4 FILLER_66_846 ();
 FILLCELL_X4 FILLER_66_853 ();
 FILLCELL_X2 FILLER_66_857 ();
 FILLCELL_X1 FILLER_66_879 ();
 FILLCELL_X1 FILLER_66_891 ();
 FILLCELL_X2 FILLER_66_905 ();
 FILLCELL_X16 FILLER_66_932 ();
 FILLCELL_X2 FILLER_66_948 ();
 FILLCELL_X1 FILLER_66_960 ();
 FILLCELL_X2 FILLER_66_964 ();
 FILLCELL_X1 FILLER_66_966 ();
 FILLCELL_X1 FILLER_66_992 ();
 FILLCELL_X2 FILLER_66_999 ();
 FILLCELL_X1 FILLER_66_1001 ();
 FILLCELL_X4 FILLER_66_1009 ();
 FILLCELL_X2 FILLER_66_1013 ();
 FILLCELL_X1 FILLER_66_1015 ();
 FILLCELL_X4 FILLER_66_1023 ();
 FILLCELL_X2 FILLER_66_1027 ();
 FILLCELL_X1 FILLER_66_1029 ();
 FILLCELL_X8 FILLER_66_1055 ();
 FILLCELL_X1 FILLER_66_1063 ();
 FILLCELL_X8 FILLER_66_1085 ();
 FILLCELL_X4 FILLER_66_1093 ();
 FILLCELL_X2 FILLER_66_1097 ();
 FILLCELL_X1 FILLER_66_1108 ();
 FILLCELL_X1 FILLER_66_1113 ();
 FILLCELL_X1 FILLER_66_1120 ();
 FILLCELL_X8 FILLER_66_1136 ();
 FILLCELL_X4 FILLER_66_1144 ();
 FILLCELL_X2 FILLER_66_1148 ();
 FILLCELL_X1 FILLER_66_1150 ();
 FILLCELL_X8 FILLER_66_1170 ();
 FILLCELL_X4 FILLER_66_1178 ();
 FILLCELL_X2 FILLER_66_1182 ();
 FILLCELL_X1 FILLER_66_1184 ();
 FILLCELL_X1 FILLER_66_1208 ();
 FILLCELL_X2 FILLER_66_1223 ();
 FILLCELL_X2 FILLER_66_1258 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X4 FILLER_67_33 ();
 FILLCELL_X2 FILLER_67_37 ();
 FILLCELL_X4 FILLER_67_66 ();
 FILLCELL_X2 FILLER_67_70 ();
 FILLCELL_X1 FILLER_67_72 ();
 FILLCELL_X16 FILLER_67_80 ();
 FILLCELL_X4 FILLER_67_96 ();
 FILLCELL_X2 FILLER_67_100 ();
 FILLCELL_X2 FILLER_67_126 ();
 FILLCELL_X1 FILLER_67_128 ();
 FILLCELL_X4 FILLER_67_183 ();
 FILLCELL_X1 FILLER_67_187 ();
 FILLCELL_X4 FILLER_67_228 ();
 FILLCELL_X1 FILLER_67_232 ();
 FILLCELL_X2 FILLER_67_260 ();
 FILLCELL_X2 FILLER_67_269 ();
 FILLCELL_X32 FILLER_67_298 ();
 FILLCELL_X8 FILLER_67_330 ();
 FILLCELL_X2 FILLER_67_338 ();
 FILLCELL_X1 FILLER_67_340 ();
 FILLCELL_X8 FILLER_67_368 ();
 FILLCELL_X2 FILLER_67_376 ();
 FILLCELL_X4 FILLER_67_405 ();
 FILLCELL_X1 FILLER_67_409 ();
 FILLCELL_X2 FILLER_67_417 ();
 FILLCELL_X1 FILLER_67_426 ();
 FILLCELL_X4 FILLER_67_461 ();
 FILLCELL_X2 FILLER_67_469 ();
 FILLCELL_X1 FILLER_67_471 ();
 FILLCELL_X1 FILLER_67_476 ();
 FILLCELL_X1 FILLER_67_515 ();
 FILLCELL_X2 FILLER_67_523 ();
 FILLCELL_X1 FILLER_67_525 ();
 FILLCELL_X8 FILLER_67_533 ();
 FILLCELL_X2 FILLER_67_541 ();
 FILLCELL_X8 FILLER_67_567 ();
 FILLCELL_X8 FILLER_67_620 ();
 FILLCELL_X4 FILLER_67_628 ();
 FILLCELL_X1 FILLER_67_632 ();
 FILLCELL_X2 FILLER_67_641 ();
 FILLCELL_X1 FILLER_67_661 ();
 FILLCELL_X1 FILLER_67_665 ();
 FILLCELL_X2 FILLER_67_675 ();
 FILLCELL_X8 FILLER_67_727 ();
 FILLCELL_X1 FILLER_67_762 ();
 FILLCELL_X4 FILLER_67_772 ();
 FILLCELL_X1 FILLER_67_776 ();
 FILLCELL_X2 FILLER_67_801 ();
 FILLCELL_X1 FILLER_67_803 ();
 FILLCELL_X4 FILLER_67_825 ();
 FILLCELL_X1 FILLER_67_829 ();
 FILLCELL_X2 FILLER_67_854 ();
 FILLCELL_X2 FILLER_67_859 ();
 FILLCELL_X4 FILLER_67_865 ();
 FILLCELL_X8 FILLER_67_871 ();
 FILLCELL_X2 FILLER_67_879 ();
 FILLCELL_X2 FILLER_67_898 ();
 FILLCELL_X1 FILLER_67_903 ();
 FILLCELL_X1 FILLER_67_915 ();
 FILLCELL_X2 FILLER_67_934 ();
 FILLCELL_X1 FILLER_67_936 ();
 FILLCELL_X1 FILLER_67_942 ();
 FILLCELL_X8 FILLER_67_969 ();
 FILLCELL_X2 FILLER_67_977 ();
 FILLCELL_X2 FILLER_67_982 ();
 FILLCELL_X1 FILLER_67_984 ();
 FILLCELL_X1 FILLER_67_992 ();
 FILLCELL_X8 FILLER_67_997 ();
 FILLCELL_X4 FILLER_67_1005 ();
 FILLCELL_X1 FILLER_67_1009 ();
 FILLCELL_X4 FILLER_67_1035 ();
 FILLCELL_X2 FILLER_67_1039 ();
 FILLCELL_X1 FILLER_67_1045 ();
 FILLCELL_X8 FILLER_67_1057 ();
 FILLCELL_X2 FILLER_67_1065 ();
 FILLCELL_X8 FILLER_67_1074 ();
 FILLCELL_X2 FILLER_67_1082 ();
 FILLCELL_X1 FILLER_67_1084 ();
 FILLCELL_X2 FILLER_67_1109 ();
 FILLCELL_X1 FILLER_67_1125 ();
 FILLCELL_X4 FILLER_67_1146 ();
 FILLCELL_X16 FILLER_67_1167 ();
 FILLCELL_X8 FILLER_67_1183 ();
 FILLCELL_X4 FILLER_67_1191 ();
 FILLCELL_X1 FILLER_67_1195 ();
 FILLCELL_X2 FILLER_67_1203 ();
 FILLCELL_X4 FILLER_67_1212 ();
 FILLCELL_X2 FILLER_67_1219 ();
 FILLCELL_X4 FILLER_67_1228 ();
 FILLCELL_X4 FILLER_67_1239 ();
 FILLCELL_X8 FILLER_68_1 ();
 FILLCELL_X4 FILLER_68_9 ();
 FILLCELL_X2 FILLER_68_13 ();
 FILLCELL_X8 FILLER_68_42 ();
 FILLCELL_X1 FILLER_68_107 ();
 FILLCELL_X1 FILLER_68_112 ();
 FILLCELL_X4 FILLER_68_164 ();
 FILLCELL_X2 FILLER_68_168 ();
 FILLCELL_X1 FILLER_68_170 ();
 FILLCELL_X16 FILLER_68_178 ();
 FILLCELL_X2 FILLER_68_194 ();
 FILLCELL_X1 FILLER_68_196 ();
 FILLCELL_X1 FILLER_68_204 ();
 FILLCELL_X4 FILLER_68_207 ();
 FILLCELL_X1 FILLER_68_211 ();
 FILLCELL_X16 FILLER_68_219 ();
 FILLCELL_X8 FILLER_68_235 ();
 FILLCELL_X1 FILLER_68_243 ();
 FILLCELL_X8 FILLER_68_280 ();
 FILLCELL_X4 FILLER_68_288 ();
 FILLCELL_X8 FILLER_68_326 ();
 FILLCELL_X1 FILLER_68_334 ();
 FILLCELL_X4 FILLER_68_349 ();
 FILLCELL_X8 FILLER_68_369 ();
 FILLCELL_X1 FILLER_68_377 ();
 FILLCELL_X4 FILLER_68_405 ();
 FILLCELL_X8 FILLER_68_429 ();
 FILLCELL_X2 FILLER_68_437 ();
 FILLCELL_X8 FILLER_68_444 ();
 FILLCELL_X2 FILLER_68_452 ();
 FILLCELL_X1 FILLER_68_454 ();
 FILLCELL_X2 FILLER_68_463 ();
 FILLCELL_X1 FILLER_68_465 ();
 FILLCELL_X4 FILLER_68_473 ();
 FILLCELL_X2 FILLER_68_477 ();
 FILLCELL_X1 FILLER_68_489 ();
 FILLCELL_X4 FILLER_68_494 ();
 FILLCELL_X2 FILLER_68_498 ();
 FILLCELL_X8 FILLER_68_515 ();
 FILLCELL_X2 FILLER_68_523 ();
 FILLCELL_X1 FILLER_68_554 ();
 FILLCELL_X4 FILLER_68_562 ();
 FILLCELL_X1 FILLER_68_566 ();
 FILLCELL_X4 FILLER_68_574 ();
 FILLCELL_X8 FILLER_68_595 ();
 FILLCELL_X2 FILLER_68_603 ();
 FILLCELL_X1 FILLER_68_605 ();
 FILLCELL_X2 FILLER_68_610 ();
 FILLCELL_X1 FILLER_68_612 ();
 FILLCELL_X1 FILLER_68_643 ();
 FILLCELL_X16 FILLER_68_661 ();
 FILLCELL_X4 FILLER_68_677 ();
 FILLCELL_X1 FILLER_68_681 ();
 FILLCELL_X4 FILLER_68_715 ();
 FILLCELL_X2 FILLER_68_719 ();
 FILLCELL_X1 FILLER_68_728 ();
 FILLCELL_X8 FILLER_68_736 ();
 FILLCELL_X1 FILLER_68_744 ();
 FILLCELL_X8 FILLER_68_748 ();
 FILLCELL_X4 FILLER_68_756 ();
 FILLCELL_X8 FILLER_68_767 ();
 FILLCELL_X4 FILLER_68_775 ();
 FILLCELL_X1 FILLER_68_784 ();
 FILLCELL_X8 FILLER_68_805 ();
 FILLCELL_X2 FILLER_68_813 ();
 FILLCELL_X1 FILLER_68_815 ();
 FILLCELL_X8 FILLER_68_851 ();
 FILLCELL_X2 FILLER_68_873 ();
 FILLCELL_X1 FILLER_68_875 ();
 FILLCELL_X2 FILLER_68_881 ();
 FILLCELL_X1 FILLER_68_883 ();
 FILLCELL_X2 FILLER_68_895 ();
 FILLCELL_X4 FILLER_68_900 ();
 FILLCELL_X1 FILLER_68_904 ();
 FILLCELL_X2 FILLER_68_910 ();
 FILLCELL_X4 FILLER_68_915 ();
 FILLCELL_X4 FILLER_68_926 ();
 FILLCELL_X2 FILLER_68_930 ();
 FILLCELL_X1 FILLER_68_932 ();
 FILLCELL_X2 FILLER_68_954 ();
 FILLCELL_X2 FILLER_68_969 ();
 FILLCELL_X4 FILLER_68_977 ();
 FILLCELL_X4 FILLER_68_984 ();
 FILLCELL_X1 FILLER_68_994 ();
 FILLCELL_X1 FILLER_68_1002 ();
 FILLCELL_X2 FILLER_68_1008 ();
 FILLCELL_X4 FILLER_68_1017 ();
 FILLCELL_X1 FILLER_68_1021 ();
 FILLCELL_X8 FILLER_68_1028 ();
 FILLCELL_X4 FILLER_68_1036 ();
 FILLCELL_X2 FILLER_68_1040 ();
 FILLCELL_X1 FILLER_68_1050 ();
 FILLCELL_X4 FILLER_68_1058 ();
 FILLCELL_X2 FILLER_68_1062 ();
 FILLCELL_X4 FILLER_68_1071 ();
 FILLCELL_X1 FILLER_68_1075 ();
 FILLCELL_X8 FILLER_68_1083 ();
 FILLCELL_X2 FILLER_68_1091 ();
 FILLCELL_X1 FILLER_68_1093 ();
 FILLCELL_X2 FILLER_68_1101 ();
 FILLCELL_X1 FILLER_68_1103 ();
 FILLCELL_X1 FILLER_68_1108 ();
 FILLCELL_X4 FILLER_68_1130 ();
 FILLCELL_X2 FILLER_68_1134 ();
 FILLCELL_X1 FILLER_68_1157 ();
 FILLCELL_X1 FILLER_68_1175 ();
 FILLCELL_X2 FILLER_68_1190 ();
 FILLCELL_X8 FILLER_68_1220 ();
 FILLCELL_X1 FILLER_68_1228 ();
 FILLCELL_X1 FILLER_68_1253 ();
 FILLCELL_X2 FILLER_68_1257 ();
 FILLCELL_X1 FILLER_68_1259 ();
 FILLCELL_X8 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_9 ();
 FILLCELL_X1 FILLER_69_13 ();
 FILLCELL_X1 FILLER_69_96 ();
 FILLCELL_X16 FILLER_69_127 ();
 FILLCELL_X1 FILLER_69_143 ();
 FILLCELL_X2 FILLER_69_165 ();
 FILLCELL_X1 FILLER_69_207 ();
 FILLCELL_X1 FILLER_69_215 ();
 FILLCELL_X4 FILLER_69_230 ();
 FILLCELL_X2 FILLER_69_234 ();
 FILLCELL_X8 FILLER_69_261 ();
 FILLCELL_X4 FILLER_69_269 ();
 FILLCELL_X1 FILLER_69_273 ();
 FILLCELL_X4 FILLER_69_301 ();
 FILLCELL_X2 FILLER_69_305 ();
 FILLCELL_X16 FILLER_69_335 ();
 FILLCELL_X4 FILLER_69_351 ();
 FILLCELL_X2 FILLER_69_355 ();
 FILLCELL_X4 FILLER_69_364 ();
 FILLCELL_X2 FILLER_69_368 ();
 FILLCELL_X1 FILLER_69_370 ();
 FILLCELL_X1 FILLER_69_391 ();
 FILLCELL_X2 FILLER_69_398 ();
 FILLCELL_X2 FILLER_69_407 ();
 FILLCELL_X16 FILLER_69_416 ();
 FILLCELL_X4 FILLER_69_432 ();
 FILLCELL_X2 FILLER_69_436 ();
 FILLCELL_X1 FILLER_69_438 ();
 FILLCELL_X8 FILLER_69_480 ();
 FILLCELL_X8 FILLER_69_492 ();
 FILLCELL_X1 FILLER_69_500 ();
 FILLCELL_X32 FILLER_69_510 ();
 FILLCELL_X1 FILLER_69_542 ();
 FILLCELL_X8 FILLER_69_550 ();
 FILLCELL_X4 FILLER_69_558 ();
 FILLCELL_X1 FILLER_69_562 ();
 FILLCELL_X1 FILLER_69_567 ();
 FILLCELL_X16 FILLER_69_571 ();
 FILLCELL_X1 FILLER_69_587 ();
 FILLCELL_X2 FILLER_69_600 ();
 FILLCELL_X8 FILLER_69_619 ();
 FILLCELL_X4 FILLER_69_627 ();
 FILLCELL_X1 FILLER_69_631 ();
 FILLCELL_X4 FILLER_69_641 ();
 FILLCELL_X1 FILLER_69_645 ();
 FILLCELL_X16 FILLER_69_685 ();
 FILLCELL_X2 FILLER_69_701 ();
 FILLCELL_X8 FILLER_69_716 ();
 FILLCELL_X4 FILLER_69_724 ();
 FILLCELL_X2 FILLER_69_728 ();
 FILLCELL_X1 FILLER_69_730 ();
 FILLCELL_X4 FILLER_69_738 ();
 FILLCELL_X2 FILLER_69_742 ();
 FILLCELL_X1 FILLER_69_744 ();
 FILLCELL_X1 FILLER_69_762 ();
 FILLCELL_X2 FILLER_69_780 ();
 FILLCELL_X1 FILLER_69_782 ();
 FILLCELL_X2 FILLER_69_800 ();
 FILLCELL_X2 FILLER_69_822 ();
 FILLCELL_X1 FILLER_69_824 ();
 FILLCELL_X2 FILLER_69_852 ();
 FILLCELL_X1 FILLER_69_873 ();
 FILLCELL_X4 FILLER_69_892 ();
 FILLCELL_X4 FILLER_69_901 ();
 FILLCELL_X2 FILLER_69_921 ();
 FILLCELL_X1 FILLER_69_923 ();
 FILLCELL_X8 FILLER_69_950 ();
 FILLCELL_X2 FILLER_69_958 ();
 FILLCELL_X8 FILLER_69_967 ();
 FILLCELL_X4 FILLER_69_1002 ();
 FILLCELL_X2 FILLER_69_1006 ();
 FILLCELL_X2 FILLER_69_1034 ();
 FILLCELL_X1 FILLER_69_1036 ();
 FILLCELL_X1 FILLER_69_1070 ();
 FILLCELL_X4 FILLER_69_1092 ();
 FILLCELL_X1 FILLER_69_1096 ();
 FILLCELL_X16 FILLER_69_1100 ();
 FILLCELL_X1 FILLER_69_1123 ();
 FILLCELL_X4 FILLER_69_1129 ();
 FILLCELL_X4 FILLER_69_1137 ();
 FILLCELL_X2 FILLER_69_1141 ();
 FILLCELL_X4 FILLER_69_1178 ();
 FILLCELL_X2 FILLER_69_1182 ();
 FILLCELL_X1 FILLER_69_1184 ();
 FILLCELL_X4 FILLER_69_1238 ();
 FILLCELL_X2 FILLER_69_1249 ();
 FILLCELL_X4 FILLER_69_1254 ();
 FILLCELL_X2 FILLER_69_1258 ();
 FILLCELL_X4 FILLER_70_1 ();
 FILLCELL_X2 FILLER_70_5 ();
 FILLCELL_X1 FILLER_70_7 ();
 FILLCELL_X2 FILLER_70_22 ();
 FILLCELL_X2 FILLER_70_45 ();
 FILLCELL_X8 FILLER_70_54 ();
 FILLCELL_X4 FILLER_70_62 ();
 FILLCELL_X4 FILLER_70_79 ();
 FILLCELL_X8 FILLER_70_90 ();
 FILLCELL_X2 FILLER_70_102 ();
 FILLCELL_X1 FILLER_70_104 ();
 FILLCELL_X1 FILLER_70_112 ();
 FILLCELL_X2 FILLER_70_120 ();
 FILLCELL_X1 FILLER_70_122 ();
 FILLCELL_X1 FILLER_70_130 ();
 FILLCELL_X2 FILLER_70_138 ();
 FILLCELL_X1 FILLER_70_147 ();
 FILLCELL_X2 FILLER_70_155 ();
 FILLCELL_X8 FILLER_70_164 ();
 FILLCELL_X2 FILLER_70_175 ();
 FILLCELL_X1 FILLER_70_177 ();
 FILLCELL_X4 FILLER_70_181 ();
 FILLCELL_X2 FILLER_70_185 ();
 FILLCELL_X4 FILLER_70_227 ();
 FILLCELL_X1 FILLER_70_231 ();
 FILLCELL_X4 FILLER_70_252 ();
 FILLCELL_X2 FILLER_70_256 ();
 FILLCELL_X4 FILLER_70_300 ();
 FILLCELL_X4 FILLER_70_307 ();
 FILLCELL_X1 FILLER_70_311 ();
 FILLCELL_X1 FILLER_70_316 ();
 FILLCELL_X8 FILLER_70_322 ();
 FILLCELL_X4 FILLER_70_354 ();
 FILLCELL_X2 FILLER_70_371 ();
 FILLCELL_X2 FILLER_70_380 ();
 FILLCELL_X4 FILLER_70_402 ();
 FILLCELL_X1 FILLER_70_413 ();
 FILLCELL_X1 FILLER_70_445 ();
 FILLCELL_X2 FILLER_70_460 ();
 FILLCELL_X1 FILLER_70_462 ();
 FILLCELL_X2 FILLER_70_483 ();
 FILLCELL_X1 FILLER_70_485 ();
 FILLCELL_X1 FILLER_70_508 ();
 FILLCELL_X8 FILLER_70_524 ();
 FILLCELL_X2 FILLER_70_532 ();
 FILLCELL_X2 FILLER_70_584 ();
 FILLCELL_X1 FILLER_70_586 ();
 FILLCELL_X1 FILLER_70_600 ();
 FILLCELL_X8 FILLER_70_618 ();
 FILLCELL_X4 FILLER_70_626 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X4 FILLER_70_650 ();
 FILLCELL_X2 FILLER_70_654 ();
 FILLCELL_X1 FILLER_70_672 ();
 FILLCELL_X2 FILLER_70_680 ();
 FILLCELL_X8 FILLER_70_687 ();
 FILLCELL_X1 FILLER_70_695 ();
 FILLCELL_X8 FILLER_70_700 ();
 FILLCELL_X2 FILLER_70_708 ();
 FILLCELL_X8 FILLER_70_719 ();
 FILLCELL_X2 FILLER_70_727 ();
 FILLCELL_X8 FILLER_70_733 ();
 FILLCELL_X2 FILLER_70_741 ();
 FILLCELL_X1 FILLER_70_743 ();
 FILLCELL_X1 FILLER_70_751 ();
 FILLCELL_X8 FILLER_70_755 ();
 FILLCELL_X4 FILLER_70_763 ();
 FILLCELL_X1 FILLER_70_767 ();
 FILLCELL_X4 FILLER_70_779 ();
 FILLCELL_X2 FILLER_70_787 ();
 FILLCELL_X1 FILLER_70_789 ();
 FILLCELL_X8 FILLER_70_804 ();
 FILLCELL_X4 FILLER_70_812 ();
 FILLCELL_X2 FILLER_70_816 ();
 FILLCELL_X8 FILLER_70_835 ();
 FILLCELL_X2 FILLER_70_843 ();
 FILLCELL_X4 FILLER_70_848 ();
 FILLCELL_X2 FILLER_70_852 ();
 FILLCELL_X1 FILLER_70_854 ();
 FILLCELL_X4 FILLER_70_864 ();
 FILLCELL_X1 FILLER_70_868 ();
 FILLCELL_X2 FILLER_70_874 ();
 FILLCELL_X1 FILLER_70_887 ();
 FILLCELL_X16 FILLER_70_893 ();
 FILLCELL_X4 FILLER_70_916 ();
 FILLCELL_X8 FILLER_70_925 ();
 FILLCELL_X2 FILLER_70_933 ();
 FILLCELL_X1 FILLER_70_935 ();
 FILLCELL_X2 FILLER_70_991 ();
 FILLCELL_X1 FILLER_70_993 ();
 FILLCELL_X8 FILLER_70_997 ();
 FILLCELL_X2 FILLER_70_1005 ();
 FILLCELL_X2 FILLER_70_1018 ();
 FILLCELL_X8 FILLER_70_1031 ();
 FILLCELL_X1 FILLER_70_1039 ();
 FILLCELL_X2 FILLER_70_1047 ();
 FILLCELL_X2 FILLER_70_1059 ();
 FILLCELL_X4 FILLER_70_1063 ();
 FILLCELL_X1 FILLER_70_1067 ();
 FILLCELL_X8 FILLER_70_1071 ();
 FILLCELL_X2 FILLER_70_1079 ();
 FILLCELL_X8 FILLER_70_1114 ();
 FILLCELL_X1 FILLER_70_1122 ();
 FILLCELL_X16 FILLER_70_1164 ();
 FILLCELL_X8 FILLER_70_1180 ();
 FILLCELL_X4 FILLER_70_1191 ();
 FILLCELL_X1 FILLER_70_1195 ();
 FILLCELL_X1 FILLER_70_1199 ();
 FILLCELL_X4 FILLER_70_1250 ();
 FILLCELL_X2 FILLER_70_1254 ();
 FILLCELL_X1 FILLER_70_1256 ();
 FILLCELL_X8 FILLER_71_1 ();
 FILLCELL_X2 FILLER_71_9 ();
 FILLCELL_X16 FILLER_71_38 ();
 FILLCELL_X4 FILLER_71_54 ();
 FILLCELL_X2 FILLER_71_58 ();
 FILLCELL_X1 FILLER_71_60 ();
 FILLCELL_X2 FILLER_71_81 ();
 FILLCELL_X8 FILLER_71_90 ();
 FILLCELL_X4 FILLER_71_98 ();
 FILLCELL_X2 FILLER_71_122 ();
 FILLCELL_X8 FILLER_71_145 ();
 FILLCELL_X4 FILLER_71_153 ();
 FILLCELL_X2 FILLER_71_157 ();
 FILLCELL_X1 FILLER_71_159 ();
 FILLCELL_X2 FILLER_71_167 ();
 FILLCELL_X1 FILLER_71_203 ();
 FILLCELL_X2 FILLER_71_218 ();
 FILLCELL_X8 FILLER_71_227 ();
 FILLCELL_X2 FILLER_71_242 ();
 FILLCELL_X1 FILLER_71_244 ();
 FILLCELL_X16 FILLER_71_272 ();
 FILLCELL_X1 FILLER_71_288 ();
 FILLCELL_X8 FILLER_71_296 ();
 FILLCELL_X4 FILLER_71_304 ();
 FILLCELL_X2 FILLER_71_308 ();
 FILLCELL_X2 FILLER_71_334 ();
 FILLCELL_X8 FILLER_71_349 ();
 FILLCELL_X4 FILLER_71_357 ();
 FILLCELL_X1 FILLER_71_361 ();
 FILLCELL_X4 FILLER_71_373 ();
 FILLCELL_X1 FILLER_71_377 ();
 FILLCELL_X2 FILLER_71_398 ();
 FILLCELL_X1 FILLER_71_400 ();
 FILLCELL_X1 FILLER_71_415 ();
 FILLCELL_X1 FILLER_71_438 ();
 FILLCELL_X1 FILLER_71_459 ();
 FILLCELL_X4 FILLER_71_472 ();
 FILLCELL_X2 FILLER_71_476 ();
 FILLCELL_X4 FILLER_71_492 ();
 FILLCELL_X2 FILLER_71_496 ();
 FILLCELL_X2 FILLER_71_511 ();
 FILLCELL_X2 FILLER_71_545 ();
 FILLCELL_X1 FILLER_71_547 ();
 FILLCELL_X8 FILLER_71_555 ();
 FILLCELL_X2 FILLER_71_563 ();
 FILLCELL_X4 FILLER_71_567 ();
 FILLCELL_X2 FILLER_71_571 ();
 FILLCELL_X1 FILLER_71_573 ();
 FILLCELL_X4 FILLER_71_576 ();
 FILLCELL_X2 FILLER_71_580 ();
 FILLCELL_X1 FILLER_71_582 ();
 FILLCELL_X8 FILLER_71_586 ();
 FILLCELL_X4 FILLER_71_594 ();
 FILLCELL_X2 FILLER_71_598 ();
 FILLCELL_X1 FILLER_71_600 ();
 FILLCELL_X2 FILLER_71_627 ();
 FILLCELL_X1 FILLER_71_629 ();
 FILLCELL_X1 FILLER_71_633 ();
 FILLCELL_X2 FILLER_71_655 ();
 FILLCELL_X1 FILLER_71_670 ();
 FILLCELL_X2 FILLER_71_682 ();
 FILLCELL_X1 FILLER_71_684 ();
 FILLCELL_X4 FILLER_71_698 ();
 FILLCELL_X2 FILLER_71_707 ();
 FILLCELL_X1 FILLER_71_709 ();
 FILLCELL_X4 FILLER_71_714 ();
 FILLCELL_X2 FILLER_71_718 ();
 FILLCELL_X16 FILLER_71_734 ();
 FILLCELL_X8 FILLER_71_750 ();
 FILLCELL_X2 FILLER_71_758 ();
 FILLCELL_X8 FILLER_71_790 ();
 FILLCELL_X8 FILLER_71_801 ();
 FILLCELL_X4 FILLER_71_809 ();
 FILLCELL_X1 FILLER_71_813 ();
 FILLCELL_X2 FILLER_71_833 ();
 FILLCELL_X1 FILLER_71_835 ();
 FILLCELL_X1 FILLER_71_845 ();
 FILLCELL_X4 FILLER_71_873 ();
 FILLCELL_X2 FILLER_71_877 ();
 FILLCELL_X1 FILLER_71_893 ();
 FILLCELL_X2 FILLER_71_905 ();
 FILLCELL_X8 FILLER_71_910 ();
 FILLCELL_X4 FILLER_71_918 ();
 FILLCELL_X1 FILLER_71_946 ();
 FILLCELL_X1 FILLER_71_960 ();
 FILLCELL_X1 FILLER_71_968 ();
 FILLCELL_X1 FILLER_71_976 ();
 FILLCELL_X4 FILLER_71_991 ();
 FILLCELL_X1 FILLER_71_995 ();
 FILLCELL_X4 FILLER_71_999 ();
 FILLCELL_X2 FILLER_71_1003 ();
 FILLCELL_X1 FILLER_71_1005 ();
 FILLCELL_X4 FILLER_71_1087 ();
 FILLCELL_X1 FILLER_71_1109 ();
 FILLCELL_X4 FILLER_71_1123 ();
 FILLCELL_X4 FILLER_71_1137 ();
 FILLCELL_X1 FILLER_71_1148 ();
 FILLCELL_X8 FILLER_71_1159 ();
 FILLCELL_X1 FILLER_71_1167 ();
 FILLCELL_X1 FILLER_71_1192 ();
 FILLCELL_X1 FILLER_71_1199 ();
 FILLCELL_X1 FILLER_71_1203 ();
 FILLCELL_X4 FILLER_71_1232 ();
 FILLCELL_X4 FILLER_72_1 ();
 FILLCELL_X2 FILLER_72_5 ();
 FILLCELL_X1 FILLER_72_34 ();
 FILLCELL_X16 FILLER_72_104 ();
 FILLCELL_X8 FILLER_72_120 ();
 FILLCELL_X4 FILLER_72_128 ();
 FILLCELL_X1 FILLER_72_132 ();
 FILLCELL_X2 FILLER_72_138 ();
 FILLCELL_X1 FILLER_72_140 ();
 FILLCELL_X16 FILLER_72_168 ();
 FILLCELL_X2 FILLER_72_184 ();
 FILLCELL_X2 FILLER_72_213 ();
 FILLCELL_X4 FILLER_72_222 ();
 FILLCELL_X2 FILLER_72_226 ();
 FILLCELL_X8 FILLER_72_235 ();
 FILLCELL_X4 FILLER_72_243 ();
 FILLCELL_X2 FILLER_72_247 ();
 FILLCELL_X8 FILLER_72_304 ();
 FILLCELL_X1 FILLER_72_312 ();
 FILLCELL_X8 FILLER_72_321 ();
 FILLCELL_X8 FILLER_72_430 ();
 FILLCELL_X2 FILLER_72_438 ();
 FILLCELL_X1 FILLER_72_440 ();
 FILLCELL_X1 FILLER_72_448 ();
 FILLCELL_X2 FILLER_72_453 ();
 FILLCELL_X1 FILLER_72_462 ();
 FILLCELL_X2 FILLER_72_470 ();
 FILLCELL_X2 FILLER_72_479 ();
 FILLCELL_X2 FILLER_72_494 ();
 FILLCELL_X4 FILLER_72_509 ();
 FILLCELL_X2 FILLER_72_520 ();
 FILLCELL_X16 FILLER_72_552 ();
 FILLCELL_X1 FILLER_72_589 ();
 FILLCELL_X1 FILLER_72_607 ();
 FILLCELL_X4 FILLER_72_619 ();
 FILLCELL_X2 FILLER_72_623 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X2 FILLER_72_632 ();
 FILLCELL_X1 FILLER_72_634 ();
 FILLCELL_X2 FILLER_72_639 ();
 FILLCELL_X4 FILLER_72_672 ();
 FILLCELL_X2 FILLER_72_676 ();
 FILLCELL_X4 FILLER_72_704 ();
 FILLCELL_X1 FILLER_72_708 ();
 FILLCELL_X2 FILLER_72_727 ();
 FILLCELL_X16 FILLER_72_748 ();
 FILLCELL_X1 FILLER_72_764 ();
 FILLCELL_X4 FILLER_72_772 ();
 FILLCELL_X4 FILLER_72_789 ();
 FILLCELL_X1 FILLER_72_793 ();
 FILLCELL_X1 FILLER_72_807 ();
 FILLCELL_X2 FILLER_72_815 ();
 FILLCELL_X1 FILLER_72_817 ();
 FILLCELL_X4 FILLER_72_825 ();
 FILLCELL_X2 FILLER_72_846 ();
 FILLCELL_X1 FILLER_72_848 ();
 FILLCELL_X4 FILLER_72_863 ();
 FILLCELL_X1 FILLER_72_867 ();
 FILLCELL_X1 FILLER_72_875 ();
 FILLCELL_X1 FILLER_72_887 ();
 FILLCELL_X1 FILLER_72_891 ();
 FILLCELL_X2 FILLER_72_905 ();
 FILLCELL_X2 FILLER_72_918 ();
 FILLCELL_X1 FILLER_72_920 ();
 FILLCELL_X1 FILLER_72_950 ();
 FILLCELL_X1 FILLER_72_984 ();
 FILLCELL_X2 FILLER_72_988 ();
 FILLCELL_X1 FILLER_72_1010 ();
 FILLCELL_X2 FILLER_72_1022 ();
 FILLCELL_X4 FILLER_72_1033 ();
 FILLCELL_X1 FILLER_72_1043 ();
 FILLCELL_X1 FILLER_72_1049 ();
 FILLCELL_X1 FILLER_72_1063 ();
 FILLCELL_X2 FILLER_72_1081 ();
 FILLCELL_X4 FILLER_72_1110 ();
 FILLCELL_X1 FILLER_72_1114 ();
 FILLCELL_X2 FILLER_72_1137 ();
 FILLCELL_X1 FILLER_72_1144 ();
 FILLCELL_X1 FILLER_72_1149 ();
 FILLCELL_X1 FILLER_72_1154 ();
 FILLCELL_X1 FILLER_72_1172 ();
 FILLCELL_X8 FILLER_72_1176 ();
 FILLCELL_X4 FILLER_72_1184 ();
 FILLCELL_X2 FILLER_72_1188 ();
 FILLCELL_X1 FILLER_72_1190 ();
 FILLCELL_X1 FILLER_72_1205 ();
 FILLCELL_X4 FILLER_72_1217 ();
 FILLCELL_X1 FILLER_72_1228 ();
 FILLCELL_X4 FILLER_72_1235 ();
 FILLCELL_X1 FILLER_72_1239 ();
 FILLCELL_X4 FILLER_72_1253 ();
 FILLCELL_X2 FILLER_72_1257 ();
 FILLCELL_X1 FILLER_72_1259 ();
 FILLCELL_X16 FILLER_73_1 ();
 FILLCELL_X4 FILLER_73_17 ();
 FILLCELL_X2 FILLER_73_28 ();
 FILLCELL_X4 FILLER_73_37 ();
 FILLCELL_X2 FILLER_73_41 ();
 FILLCELL_X4 FILLER_73_50 ();
 FILLCELL_X2 FILLER_73_54 ();
 FILLCELL_X2 FILLER_73_71 ();
 FILLCELL_X1 FILLER_73_73 ();
 FILLCELL_X2 FILLER_73_101 ();
 FILLCELL_X1 FILLER_73_110 ();
 FILLCELL_X2 FILLER_73_138 ();
 FILLCELL_X1 FILLER_73_140 ();
 FILLCELL_X8 FILLER_73_148 ();
 FILLCELL_X4 FILLER_73_156 ();
 FILLCELL_X1 FILLER_73_160 ();
 FILLCELL_X8 FILLER_73_176 ();
 FILLCELL_X4 FILLER_73_184 ();
 FILLCELL_X2 FILLER_73_188 ();
 FILLCELL_X2 FILLER_73_203 ();
 FILLCELL_X4 FILLER_73_212 ();
 FILLCELL_X1 FILLER_73_225 ();
 FILLCELL_X16 FILLER_73_246 ();
 FILLCELL_X2 FILLER_73_269 ();
 FILLCELL_X4 FILLER_73_278 ();
 FILLCELL_X2 FILLER_73_282 ();
 FILLCELL_X4 FILLER_73_311 ();
 FILLCELL_X1 FILLER_73_315 ();
 FILLCELL_X2 FILLER_73_323 ();
 FILLCELL_X1 FILLER_73_325 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X2 FILLER_73_385 ();
 FILLCELL_X8 FILLER_73_394 ();
 FILLCELL_X4 FILLER_73_402 ();
 FILLCELL_X2 FILLER_73_406 ();
 FILLCELL_X1 FILLER_73_415 ();
 FILLCELL_X4 FILLER_73_418 ();
 FILLCELL_X1 FILLER_73_422 ();
 FILLCELL_X16 FILLER_73_499 ();
 FILLCELL_X8 FILLER_73_515 ();
 FILLCELL_X1 FILLER_73_523 ();
 FILLCELL_X4 FILLER_73_537 ();
 FILLCELL_X2 FILLER_73_541 ();
 FILLCELL_X1 FILLER_73_543 ();
 FILLCELL_X2 FILLER_73_548 ();
 FILLCELL_X8 FILLER_73_567 ();
 FILLCELL_X2 FILLER_73_575 ();
 FILLCELL_X4 FILLER_73_582 ();
 FILLCELL_X2 FILLER_73_586 ();
 FILLCELL_X1 FILLER_73_588 ();
 FILLCELL_X4 FILLER_73_606 ();
 FILLCELL_X1 FILLER_73_610 ();
 FILLCELL_X4 FILLER_73_624 ();
 FILLCELL_X1 FILLER_73_628 ();
 FILLCELL_X4 FILLER_73_634 ();
 FILLCELL_X8 FILLER_73_648 ();
 FILLCELL_X4 FILLER_73_674 ();
 FILLCELL_X4 FILLER_73_685 ();
 FILLCELL_X2 FILLER_73_689 ();
 FILLCELL_X4 FILLER_73_713 ();
 FILLCELL_X1 FILLER_73_717 ();
 FILLCELL_X16 FILLER_73_721 ();
 FILLCELL_X16 FILLER_73_774 ();
 FILLCELL_X8 FILLER_73_790 ();
 FILLCELL_X4 FILLER_73_801 ();
 FILLCELL_X16 FILLER_73_818 ();
 FILLCELL_X2 FILLER_73_834 ();
 FILLCELL_X1 FILLER_73_836 ();
 FILLCELL_X8 FILLER_73_842 ();
 FILLCELL_X1 FILLER_73_850 ();
 FILLCELL_X4 FILLER_73_864 ();
 FILLCELL_X16 FILLER_73_889 ();
 FILLCELL_X16 FILLER_73_912 ();
 FILLCELL_X1 FILLER_73_952 ();
 FILLCELL_X1 FILLER_73_956 ();
 FILLCELL_X1 FILLER_73_966 ();
 FILLCELL_X16 FILLER_73_987 ();
 FILLCELL_X8 FILLER_73_1003 ();
 FILLCELL_X2 FILLER_73_1011 ();
 FILLCELL_X1 FILLER_73_1016 ();
 FILLCELL_X16 FILLER_73_1020 ();
 FILLCELL_X2 FILLER_73_1055 ();
 FILLCELL_X8 FILLER_73_1078 ();
 FILLCELL_X8 FILLER_73_1100 ();
 FILLCELL_X2 FILLER_73_1108 ();
 FILLCELL_X1 FILLER_73_1110 ();
 FILLCELL_X2 FILLER_73_1122 ();
 FILLCELL_X1 FILLER_73_1128 ();
 FILLCELL_X2 FILLER_73_1141 ();
 FILLCELL_X1 FILLER_73_1143 ();
 FILLCELL_X2 FILLER_73_1147 ();
 FILLCELL_X1 FILLER_73_1149 ();
 FILLCELL_X2 FILLER_73_1154 ();
 FILLCELL_X1 FILLER_73_1156 ();
 FILLCELL_X2 FILLER_73_1165 ();
 FILLCELL_X1 FILLER_73_1167 ();
 FILLCELL_X2 FILLER_73_1200 ();
 FILLCELL_X2 FILLER_73_1213 ();
 FILLCELL_X1 FILLER_73_1224 ();
 FILLCELL_X4 FILLER_73_1230 ();
 FILLCELL_X1 FILLER_73_1234 ();
 FILLCELL_X2 FILLER_73_1242 ();
 FILLCELL_X2 FILLER_73_1251 ();
 FILLCELL_X1 FILLER_73_1253 ();
 FILLCELL_X8 FILLER_74_1 ();
 FILLCELL_X1 FILLER_74_9 ();
 FILLCELL_X4 FILLER_74_37 ();
 FILLCELL_X1 FILLER_74_88 ();
 FILLCELL_X2 FILLER_74_103 ();
 FILLCELL_X8 FILLER_74_126 ();
 FILLCELL_X1 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_180 ();
 FILLCELL_X1 FILLER_74_212 ();
 FILLCELL_X4 FILLER_74_227 ();
 FILLCELL_X1 FILLER_74_231 ();
 FILLCELL_X2 FILLER_74_259 ();
 FILLCELL_X8 FILLER_74_290 ();
 FILLCELL_X4 FILLER_74_298 ();
 FILLCELL_X1 FILLER_74_302 ();
 FILLCELL_X2 FILLER_74_316 ();
 FILLCELL_X1 FILLER_74_318 ();
 FILLCELL_X2 FILLER_74_339 ();
 FILLCELL_X1 FILLER_74_341 ();
 FILLCELL_X4 FILLER_74_346 ();
 FILLCELL_X1 FILLER_74_350 ();
 FILLCELL_X8 FILLER_74_394 ();
 FILLCELL_X8 FILLER_74_481 ();
 FILLCELL_X16 FILLER_74_525 ();
 FILLCELL_X1 FILLER_74_541 ();
 FILLCELL_X8 FILLER_74_563 ();
 FILLCELL_X2 FILLER_74_571 ();
 FILLCELL_X1 FILLER_74_573 ();
 FILLCELL_X4 FILLER_74_599 ();
 FILLCELL_X1 FILLER_74_603 ();
 FILLCELL_X4 FILLER_74_656 ();
 FILLCELL_X8 FILLER_74_664 ();
 FILLCELL_X2 FILLER_74_672 ();
 FILLCELL_X4 FILLER_74_687 ();
 FILLCELL_X1 FILLER_74_691 ();
 FILLCELL_X1 FILLER_74_699 ();
 FILLCELL_X4 FILLER_74_713 ();
 FILLCELL_X2 FILLER_74_717 ();
 FILLCELL_X4 FILLER_74_728 ();
 FILLCELL_X1 FILLER_74_732 ();
 FILLCELL_X1 FILLER_74_737 ();
 FILLCELL_X1 FILLER_74_743 ();
 FILLCELL_X2 FILLER_74_760 ();
 FILLCELL_X16 FILLER_74_785 ();
 FILLCELL_X8 FILLER_74_801 ();
 FILLCELL_X4 FILLER_74_809 ();
 FILLCELL_X2 FILLER_74_813 ();
 FILLCELL_X2 FILLER_74_818 ();
 FILLCELL_X2 FILLER_74_823 ();
 FILLCELL_X1 FILLER_74_825 ();
 FILLCELL_X2 FILLER_74_829 ();
 FILLCELL_X1 FILLER_74_831 ();
 FILLCELL_X4 FILLER_74_845 ();
 FILLCELL_X1 FILLER_74_849 ();
 FILLCELL_X8 FILLER_74_858 ();
 FILLCELL_X2 FILLER_74_866 ();
 FILLCELL_X1 FILLER_74_868 ();
 FILLCELL_X4 FILLER_74_929 ();
 FILLCELL_X1 FILLER_74_933 ();
 FILLCELL_X4 FILLER_74_942 ();
 FILLCELL_X1 FILLER_74_946 ();
 FILLCELL_X1 FILLER_74_952 ();
 FILLCELL_X8 FILLER_74_971 ();
 FILLCELL_X2 FILLER_74_979 ();
 FILLCELL_X1 FILLER_74_981 ();
 FILLCELL_X4 FILLER_74_1012 ();
 FILLCELL_X4 FILLER_74_1040 ();
 FILLCELL_X2 FILLER_74_1044 ();
 FILLCELL_X1 FILLER_74_1046 ();
 FILLCELL_X2 FILLER_74_1050 ();
 FILLCELL_X8 FILLER_74_1062 ();
 FILLCELL_X4 FILLER_74_1070 ();
 FILLCELL_X8 FILLER_74_1100 ();
 FILLCELL_X4 FILLER_74_1108 ();
 FILLCELL_X1 FILLER_74_1112 ();
 FILLCELL_X2 FILLER_74_1124 ();
 FILLCELL_X16 FILLER_74_1166 ();
 FILLCELL_X8 FILLER_74_1182 ();
 FILLCELL_X1 FILLER_74_1190 ();
 FILLCELL_X2 FILLER_74_1196 ();
 FILLCELL_X1 FILLER_74_1198 ();
 FILLCELL_X2 FILLER_74_1202 ();
 FILLCELL_X1 FILLER_74_1204 ();
 FILLCELL_X1 FILLER_74_1217 ();
 FILLCELL_X4 FILLER_74_1238 ();
 FILLCELL_X1 FILLER_74_1242 ();
 FILLCELL_X4 FILLER_75_21 ();
 FILLCELL_X2 FILLER_75_25 ();
 FILLCELL_X1 FILLER_75_54 ();
 FILLCELL_X1 FILLER_75_80 ();
 FILLCELL_X8 FILLER_75_108 ();
 FILLCELL_X2 FILLER_75_116 ();
 FILLCELL_X8 FILLER_75_145 ();
 FILLCELL_X8 FILLER_75_155 ();
 FILLCELL_X1 FILLER_75_163 ();
 FILLCELL_X2 FILLER_75_177 ();
 FILLCELL_X1 FILLER_75_179 ();
 FILLCELL_X1 FILLER_75_214 ();
 FILLCELL_X4 FILLER_75_229 ();
 FILLCELL_X1 FILLER_75_233 ();
 FILLCELL_X4 FILLER_75_241 ();
 FILLCELL_X2 FILLER_75_245 ();
 FILLCELL_X1 FILLER_75_249 ();
 FILLCELL_X16 FILLER_75_259 ();
 FILLCELL_X4 FILLER_75_275 ();
 FILLCELL_X2 FILLER_75_279 ();
 FILLCELL_X1 FILLER_75_281 ();
 FILLCELL_X2 FILLER_75_323 ();
 FILLCELL_X16 FILLER_75_361 ();
 FILLCELL_X2 FILLER_75_377 ();
 FILLCELL_X2 FILLER_75_406 ();
 FILLCELL_X2 FILLER_75_491 ();
 FILLCELL_X1 FILLER_75_493 ();
 FILLCELL_X16 FILLER_75_521 ();
 FILLCELL_X4 FILLER_75_572 ();
 FILLCELL_X2 FILLER_75_580 ();
 FILLCELL_X1 FILLER_75_582 ();
 FILLCELL_X2 FILLER_75_590 ();
 FILLCELL_X1 FILLER_75_592 ();
 FILLCELL_X2 FILLER_75_609 ();
 FILLCELL_X1 FILLER_75_647 ();
 FILLCELL_X2 FILLER_75_667 ();
 FILLCELL_X2 FILLER_75_682 ();
 FILLCELL_X2 FILLER_75_693 ();
 FILLCELL_X1 FILLER_75_695 ();
 FILLCELL_X2 FILLER_75_700 ();
 FILLCELL_X1 FILLER_75_702 ();
 FILLCELL_X2 FILLER_75_706 ();
 FILLCELL_X2 FILLER_75_715 ();
 FILLCELL_X8 FILLER_75_730 ();
 FILLCELL_X8 FILLER_75_745 ();
 FILLCELL_X4 FILLER_75_753 ();
 FILLCELL_X1 FILLER_75_757 ();
 FILLCELL_X4 FILLER_75_775 ();
 FILLCELL_X2 FILLER_75_779 ();
 FILLCELL_X4 FILLER_75_819 ();
 FILLCELL_X2 FILLER_75_823 ();
 FILLCELL_X2 FILLER_75_834 ();
 FILLCELL_X1 FILLER_75_839 ();
 FILLCELL_X1 FILLER_75_847 ();
 FILLCELL_X2 FILLER_75_853 ();
 FILLCELL_X4 FILLER_75_868 ();
 FILLCELL_X2 FILLER_75_872 ();
 FILLCELL_X8 FILLER_75_881 ();
 FILLCELL_X2 FILLER_75_889 ();
 FILLCELL_X16 FILLER_75_905 ();
 FILLCELL_X8 FILLER_75_921 ();
 FILLCELL_X2 FILLER_75_951 ();
 FILLCELL_X16 FILLER_75_960 ();
 FILLCELL_X2 FILLER_75_976 ();
 FILLCELL_X32 FILLER_75_991 ();
 FILLCELL_X8 FILLER_75_1023 ();
 FILLCELL_X2 FILLER_75_1031 ();
 FILLCELL_X2 FILLER_75_1043 ();
 FILLCELL_X1 FILLER_75_1045 ();
 FILLCELL_X1 FILLER_75_1049 ();
 FILLCELL_X32 FILLER_75_1055 ();
 FILLCELL_X4 FILLER_75_1087 ();
 FILLCELL_X1 FILLER_75_1128 ();
 FILLCELL_X4 FILLER_75_1136 ();
 FILLCELL_X2 FILLER_75_1140 ();
 FILLCELL_X2 FILLER_75_1150 ();
 FILLCELL_X4 FILLER_75_1161 ();
 FILLCELL_X1 FILLER_75_1172 ();
 FILLCELL_X1 FILLER_75_1181 ();
 FILLCELL_X1 FILLER_75_1187 ();
 FILLCELL_X1 FILLER_75_1191 ();
 FILLCELL_X2 FILLER_75_1211 ();
 FILLCELL_X16 FILLER_75_1243 ();
 FILLCELL_X1 FILLER_75_1259 ();
 FILLCELL_X8 FILLER_76_28 ();
 FILLCELL_X4 FILLER_76_36 ();
 FILLCELL_X4 FILLER_76_47 ();
 FILLCELL_X2 FILLER_76_51 ();
 FILLCELL_X1 FILLER_76_53 ();
 FILLCELL_X2 FILLER_76_68 ();
 FILLCELL_X2 FILLER_76_89 ();
 FILLCELL_X1 FILLER_76_91 ();
 FILLCELL_X1 FILLER_76_120 ();
 FILLCELL_X8 FILLER_76_123 ();
 FILLCELL_X2 FILLER_76_131 ();
 FILLCELL_X1 FILLER_76_133 ();
 FILLCELL_X1 FILLER_76_148 ();
 FILLCELL_X8 FILLER_76_158 ();
 FILLCELL_X4 FILLER_76_166 ();
 FILLCELL_X2 FILLER_76_170 ();
 FILLCELL_X1 FILLER_76_172 ();
 FILLCELL_X2 FILLER_76_192 ();
 FILLCELL_X1 FILLER_76_256 ();
 FILLCELL_X2 FILLER_76_277 ();
 FILLCELL_X2 FILLER_76_281 ();
 FILLCELL_X4 FILLER_76_302 ();
 FILLCELL_X2 FILLER_76_306 ();
 FILLCELL_X1 FILLER_76_308 ();
 FILLCELL_X2 FILLER_76_334 ();
 FILLCELL_X4 FILLER_76_339 ();
 FILLCELL_X8 FILLER_76_354 ();
 FILLCELL_X4 FILLER_76_362 ();
 FILLCELL_X2 FILLER_76_366 ();
 FILLCELL_X1 FILLER_76_368 ();
 FILLCELL_X2 FILLER_76_396 ();
 FILLCELL_X1 FILLER_76_398 ();
 FILLCELL_X8 FILLER_76_406 ();
 FILLCELL_X16 FILLER_76_448 ();
 FILLCELL_X4 FILLER_76_464 ();
 FILLCELL_X1 FILLER_76_468 ();
 FILLCELL_X1 FILLER_76_503 ();
 FILLCELL_X8 FILLER_76_531 ();
 FILLCELL_X4 FILLER_76_539 ();
 FILLCELL_X16 FILLER_76_552 ();
 FILLCELL_X8 FILLER_76_568 ();
 FILLCELL_X4 FILLER_76_576 ();
 FILLCELL_X2 FILLER_76_580 ();
 FILLCELL_X4 FILLER_76_594 ();
 FILLCELL_X8 FILLER_76_602 ();
 FILLCELL_X4 FILLER_76_610 ();
 FILLCELL_X2 FILLER_76_614 ();
 FILLCELL_X1 FILLER_76_616 ();
 FILLCELL_X1 FILLER_76_632 ();
 FILLCELL_X2 FILLER_76_640 ();
 FILLCELL_X2 FILLER_76_647 ();
 FILLCELL_X2 FILLER_76_662 ();
 FILLCELL_X1 FILLER_76_664 ();
 FILLCELL_X1 FILLER_76_681 ();
 FILLCELL_X1 FILLER_76_699 ();
 FILLCELL_X2 FILLER_76_713 ();
 FILLCELL_X2 FILLER_76_722 ();
 FILLCELL_X2 FILLER_76_733 ();
 FILLCELL_X1 FILLER_76_735 ();
 FILLCELL_X4 FILLER_76_743 ();
 FILLCELL_X1 FILLER_76_747 ();
 FILLCELL_X4 FILLER_76_756 ();
 FILLCELL_X2 FILLER_76_760 ();
 FILLCELL_X1 FILLER_76_762 ();
 FILLCELL_X4 FILLER_76_767 ();
 FILLCELL_X2 FILLER_76_771 ();
 FILLCELL_X1 FILLER_76_773 ();
 FILLCELL_X4 FILLER_76_781 ();
 FILLCELL_X2 FILLER_76_785 ();
 FILLCELL_X16 FILLER_76_815 ();
 FILLCELL_X4 FILLER_76_831 ();
 FILLCELL_X2 FILLER_76_835 ();
 FILLCELL_X1 FILLER_76_837 ();
 FILLCELL_X16 FILLER_76_848 ();
 FILLCELL_X16 FILLER_76_867 ();
 FILLCELL_X1 FILLER_76_883 ();
 FILLCELL_X4 FILLER_76_935 ();
 FILLCELL_X2 FILLER_76_939 ();
 FILLCELL_X1 FILLER_76_941 ();
 FILLCELL_X1 FILLER_76_949 ();
 FILLCELL_X1 FILLER_76_957 ();
 FILLCELL_X1 FILLER_76_978 ();
 FILLCELL_X8 FILLER_76_999 ();
 FILLCELL_X1 FILLER_76_1007 ();
 FILLCELL_X4 FILLER_76_1015 ();
 FILLCELL_X1 FILLER_76_1019 ();
 FILLCELL_X4 FILLER_76_1039 ();
 FILLCELL_X1 FILLER_76_1055 ();
 FILLCELL_X1 FILLER_76_1066 ();
 FILLCELL_X16 FILLER_76_1091 ();
 FILLCELL_X8 FILLER_76_1107 ();
 FILLCELL_X1 FILLER_76_1115 ();
 FILLCELL_X8 FILLER_76_1132 ();
 FILLCELL_X2 FILLER_76_1140 ();
 FILLCELL_X16 FILLER_76_1150 ();
 FILLCELL_X1 FILLER_76_1166 ();
 FILLCELL_X2 FILLER_76_1216 ();
 FILLCELL_X1 FILLER_76_1218 ();
 FILLCELL_X1 FILLER_76_1246 ();
 FILLCELL_X4 FILLER_76_1253 ();
 FILLCELL_X8 FILLER_77_1 ();
 FILLCELL_X2 FILLER_77_9 ();
 FILLCELL_X1 FILLER_77_11 ();
 FILLCELL_X2 FILLER_77_73 ();
 FILLCELL_X8 FILLER_77_89 ();
 FILLCELL_X1 FILLER_77_97 ();
 FILLCELL_X8 FILLER_77_119 ();
 FILLCELL_X4 FILLER_77_143 ();
 FILLCELL_X8 FILLER_77_149 ();
 FILLCELL_X4 FILLER_77_157 ();
 FILLCELL_X2 FILLER_77_161 ();
 FILLCELL_X8 FILLER_77_191 ();
 FILLCELL_X8 FILLER_77_231 ();
 FILLCELL_X4 FILLER_77_239 ();
 FILLCELL_X2 FILLER_77_243 ();
 FILLCELL_X1 FILLER_77_245 ();
 FILLCELL_X4 FILLER_77_249 ();
 FILLCELL_X2 FILLER_77_253 ();
 FILLCELL_X1 FILLER_77_262 ();
 FILLCELL_X2 FILLER_77_270 ();
 FILLCELL_X2 FILLER_77_286 ();
 FILLCELL_X1 FILLER_77_288 ();
 FILLCELL_X8 FILLER_77_296 ();
 FILLCELL_X2 FILLER_77_304 ();
 FILLCELL_X8 FILLER_77_342 ();
 FILLCELL_X1 FILLER_77_350 ();
 FILLCELL_X2 FILLER_77_378 ();
 FILLCELL_X1 FILLER_77_380 ();
 FILLCELL_X1 FILLER_77_388 ();
 FILLCELL_X1 FILLER_77_425 ();
 FILLCELL_X1 FILLER_77_436 ();
 FILLCELL_X4 FILLER_77_457 ();
 FILLCELL_X1 FILLER_77_461 ();
 FILLCELL_X8 FILLER_77_475 ();
 FILLCELL_X1 FILLER_77_483 ();
 FILLCELL_X2 FILLER_77_491 ();
 FILLCELL_X16 FILLER_77_527 ();
 FILLCELL_X1 FILLER_77_543 ();
 FILLCELL_X2 FILLER_77_556 ();
 FILLCELL_X4 FILLER_77_580 ();
 FILLCELL_X1 FILLER_77_584 ();
 FILLCELL_X2 FILLER_77_598 ();
 FILLCELL_X8 FILLER_77_619 ();
 FILLCELL_X1 FILLER_77_627 ();
 FILLCELL_X2 FILLER_77_641 ();
 FILLCELL_X1 FILLER_77_643 ();
 FILLCELL_X1 FILLER_77_656 ();
 FILLCELL_X2 FILLER_77_683 ();
 FILLCELL_X1 FILLER_77_685 ();
 FILLCELL_X1 FILLER_77_689 ();
 FILLCELL_X4 FILLER_77_705 ();
 FILLCELL_X1 FILLER_77_709 ();
 FILLCELL_X1 FILLER_77_715 ();
 FILLCELL_X2 FILLER_77_726 ();
 FILLCELL_X1 FILLER_77_728 ();
 FILLCELL_X4 FILLER_77_747 ();
 FILLCELL_X2 FILLER_77_754 ();
 FILLCELL_X1 FILLER_77_764 ();
 FILLCELL_X1 FILLER_77_780 ();
 FILLCELL_X1 FILLER_77_786 ();
 FILLCELL_X2 FILLER_77_790 ();
 FILLCELL_X2 FILLER_77_799 ();
 FILLCELL_X2 FILLER_77_805 ();
 FILLCELL_X2 FILLER_77_816 ();
 FILLCELL_X1 FILLER_77_818 ();
 FILLCELL_X8 FILLER_77_826 ();
 FILLCELL_X4 FILLER_77_834 ();
 FILLCELL_X2 FILLER_77_838 ();
 FILLCELL_X16 FILLER_77_842 ();
 FILLCELL_X4 FILLER_77_858 ();
 FILLCELL_X1 FILLER_77_862 ();
 FILLCELL_X1 FILLER_77_866 ();
 FILLCELL_X16 FILLER_77_869 ();
 FILLCELL_X4 FILLER_77_885 ();
 FILLCELL_X2 FILLER_77_889 ();
 FILLCELL_X1 FILLER_77_891 ();
 FILLCELL_X16 FILLER_77_895 ();
 FILLCELL_X4 FILLER_77_911 ();
 FILLCELL_X2 FILLER_77_924 ();
 FILLCELL_X4 FILLER_77_971 ();
 FILLCELL_X2 FILLER_77_975 ();
 FILLCELL_X8 FILLER_77_984 ();
 FILLCELL_X4 FILLER_77_992 ();
 FILLCELL_X1 FILLER_77_996 ();
 FILLCELL_X1 FILLER_77_1017 ();
 FILLCELL_X1 FILLER_77_1029 ();
 FILLCELL_X1 FILLER_77_1037 ();
 FILLCELL_X4 FILLER_77_1065 ();
 FILLCELL_X4 FILLER_77_1076 ();
 FILLCELL_X2 FILLER_77_1080 ();
 FILLCELL_X2 FILLER_77_1088 ();
 FILLCELL_X4 FILLER_77_1109 ();
 FILLCELL_X1 FILLER_77_1113 ();
 FILLCELL_X1 FILLER_77_1135 ();
 FILLCELL_X8 FILLER_77_1155 ();
 FILLCELL_X4 FILLER_77_1187 ();
 FILLCELL_X2 FILLER_77_1191 ();
 FILLCELL_X2 FILLER_77_1197 ();
 FILLCELL_X2 FILLER_77_1210 ();
 FILLCELL_X1 FILLER_77_1212 ();
 FILLCELL_X4 FILLER_77_1230 ();
 FILLCELL_X2 FILLER_77_1234 ();
 FILLCELL_X8 FILLER_78_1 ();
 FILLCELL_X4 FILLER_78_9 ();
 FILLCELL_X1 FILLER_78_13 ();
 FILLCELL_X8 FILLER_78_48 ();
 FILLCELL_X1 FILLER_78_56 ();
 FILLCELL_X1 FILLER_78_64 ();
 FILLCELL_X16 FILLER_78_67 ();
 FILLCELL_X4 FILLER_78_83 ();
 FILLCELL_X2 FILLER_78_87 ();
 FILLCELL_X1 FILLER_78_89 ();
 FILLCELL_X2 FILLER_78_97 ();
 FILLCELL_X2 FILLER_78_106 ();
 FILLCELL_X1 FILLER_78_108 ();
 FILLCELL_X4 FILLER_78_116 ();
 FILLCELL_X4 FILLER_78_178 ();
 FILLCELL_X8 FILLER_78_194 ();
 FILLCELL_X1 FILLER_78_202 ();
 FILLCELL_X1 FILLER_78_217 ();
 FILLCELL_X1 FILLER_78_240 ();
 FILLCELL_X1 FILLER_78_250 ();
 FILLCELL_X2 FILLER_78_262 ();
 FILLCELL_X1 FILLER_78_264 ();
 FILLCELL_X2 FILLER_78_285 ();
 FILLCELL_X1 FILLER_78_287 ();
 FILLCELL_X2 FILLER_78_302 ();
 FILLCELL_X4 FILLER_78_317 ();
 FILLCELL_X2 FILLER_78_328 ();
 FILLCELL_X1 FILLER_78_330 ();
 FILLCELL_X2 FILLER_78_334 ();
 FILLCELL_X1 FILLER_78_336 ();
 FILLCELL_X4 FILLER_78_342 ();
 FILLCELL_X2 FILLER_78_346 ();
 FILLCELL_X4 FILLER_78_357 ();
 FILLCELL_X2 FILLER_78_361 ();
 FILLCELL_X1 FILLER_78_363 ();
 FILLCELL_X8 FILLER_78_371 ();
 FILLCELL_X2 FILLER_78_379 ();
 FILLCELL_X1 FILLER_78_381 ();
 FILLCELL_X16 FILLER_78_408 ();
 FILLCELL_X1 FILLER_78_424 ();
 FILLCELL_X2 FILLER_78_487 ();
 FILLCELL_X4 FILLER_78_503 ();
 FILLCELL_X2 FILLER_78_507 ();
 FILLCELL_X1 FILLER_78_509 ();
 FILLCELL_X4 FILLER_78_531 ();
 FILLCELL_X2 FILLER_78_535 ();
 FILLCELL_X1 FILLER_78_537 ();
 FILLCELL_X1 FILLER_78_574 ();
 FILLCELL_X4 FILLER_78_579 ();
 FILLCELL_X2 FILLER_78_583 ();
 FILLCELL_X8 FILLER_78_619 ();
 FILLCELL_X4 FILLER_78_627 ();
 FILLCELL_X2 FILLER_78_632 ();
 FILLCELL_X1 FILLER_78_651 ();
 FILLCELL_X2 FILLER_78_659 ();
 FILLCELL_X4 FILLER_78_674 ();
 FILLCELL_X1 FILLER_78_678 ();
 FILLCELL_X1 FILLER_78_701 ();
 FILLCELL_X8 FILLER_78_706 ();
 FILLCELL_X2 FILLER_78_714 ();
 FILLCELL_X4 FILLER_78_728 ();
 FILLCELL_X2 FILLER_78_732 ();
 FILLCELL_X1 FILLER_78_734 ();
 FILLCELL_X4 FILLER_78_745 ();
 FILLCELL_X2 FILLER_78_749 ();
 FILLCELL_X1 FILLER_78_751 ();
 FILLCELL_X8 FILLER_78_761 ();
 FILLCELL_X1 FILLER_78_769 ();
 FILLCELL_X4 FILLER_78_779 ();
 FILLCELL_X1 FILLER_78_783 ();
 FILLCELL_X2 FILLER_78_796 ();
 FILLCELL_X16 FILLER_78_811 ();
 FILLCELL_X2 FILLER_78_827 ();
 FILLCELL_X4 FILLER_78_839 ();
 FILLCELL_X2 FILLER_78_843 ();
 FILLCELL_X16 FILLER_78_868 ();
 FILLCELL_X2 FILLER_78_884 ();
 FILLCELL_X1 FILLER_78_886 ();
 FILLCELL_X8 FILLER_78_901 ();
 FILLCELL_X1 FILLER_78_909 ();
 FILLCELL_X8 FILLER_78_944 ();
 FILLCELL_X2 FILLER_78_952 ();
 FILLCELL_X1 FILLER_78_954 ();
 FILLCELL_X16 FILLER_78_958 ();
 FILLCELL_X8 FILLER_78_974 ();
 FILLCELL_X4 FILLER_78_982 ();
 FILLCELL_X1 FILLER_78_998 ();
 FILLCELL_X2 FILLER_78_1011 ();
 FILLCELL_X1 FILLER_78_1017 ();
 FILLCELL_X1 FILLER_78_1027 ();
 FILLCELL_X1 FILLER_78_1036 ();
 FILLCELL_X2 FILLER_78_1045 ();
 FILLCELL_X1 FILLER_78_1047 ();
 FILLCELL_X1 FILLER_78_1060 ();
 FILLCELL_X4 FILLER_78_1068 ();
 FILLCELL_X4 FILLER_78_1076 ();
 FILLCELL_X2 FILLER_78_1080 ();
 FILLCELL_X1 FILLER_78_1082 ();
 FILLCELL_X16 FILLER_78_1107 ();
 FILLCELL_X4 FILLER_78_1127 ();
 FILLCELL_X2 FILLER_78_1131 ();
 FILLCELL_X8 FILLER_78_1147 ();
 FILLCELL_X2 FILLER_78_1155 ();
 FILLCELL_X2 FILLER_78_1160 ();
 FILLCELL_X16 FILLER_78_1169 ();
 FILLCELL_X4 FILLER_78_1191 ();
 FILLCELL_X1 FILLER_78_1195 ();
 FILLCELL_X1 FILLER_78_1199 ();
 FILLCELL_X8 FILLER_78_1231 ();
 FILLCELL_X2 FILLER_78_1239 ();
 FILLCELL_X1 FILLER_78_1241 ();
 FILLCELL_X8 FILLER_78_1252 ();
 FILLCELL_X8 FILLER_79_1 ();
 FILLCELL_X2 FILLER_79_9 ();
 FILLCELL_X1 FILLER_79_11 ();
 FILLCELL_X4 FILLER_79_39 ();
 FILLCELL_X2 FILLER_79_43 ();
 FILLCELL_X4 FILLER_79_52 ();
 FILLCELL_X2 FILLER_79_56 ();
 FILLCELL_X1 FILLER_79_58 ();
 FILLCELL_X1 FILLER_79_80 ();
 FILLCELL_X1 FILLER_79_88 ();
 FILLCELL_X32 FILLER_79_137 ();
 FILLCELL_X2 FILLER_79_169 ();
 FILLCELL_X2 FILLER_79_191 ();
 FILLCELL_X1 FILLER_79_193 ();
 FILLCELL_X2 FILLER_79_214 ();
 FILLCELL_X1 FILLER_79_216 ();
 FILLCELL_X1 FILLER_79_224 ();
 FILLCELL_X4 FILLER_79_279 ();
 FILLCELL_X2 FILLER_79_283 ();
 FILLCELL_X2 FILLER_79_299 ();
 FILLCELL_X1 FILLER_79_301 ();
 FILLCELL_X1 FILLER_79_327 ();
 FILLCELL_X1 FILLER_79_341 ();
 FILLCELL_X2 FILLER_79_348 ();
 FILLCELL_X16 FILLER_79_377 ();
 FILLCELL_X4 FILLER_79_393 ();
 FILLCELL_X1 FILLER_79_397 ();
 FILLCELL_X16 FILLER_79_439 ();
 FILLCELL_X8 FILLER_79_455 ();
 FILLCELL_X1 FILLER_79_463 ();
 FILLCELL_X1 FILLER_79_482 ();
 FILLCELL_X2 FILLER_79_518 ();
 FILLCELL_X4 FILLER_79_527 ();
 FILLCELL_X2 FILLER_79_531 ();
 FILLCELL_X4 FILLER_79_546 ();
 FILLCELL_X1 FILLER_79_550 ();
 FILLCELL_X1 FILLER_79_553 ();
 FILLCELL_X8 FILLER_79_558 ();
 FILLCELL_X1 FILLER_79_566 ();
 FILLCELL_X2 FILLER_79_581 ();
 FILLCELL_X1 FILLER_79_583 ();
 FILLCELL_X2 FILLER_79_613 ();
 FILLCELL_X1 FILLER_79_615 ();
 FILLCELL_X1 FILLER_79_620 ();
 FILLCELL_X2 FILLER_79_637 ();
 FILLCELL_X4 FILLER_79_648 ();
 FILLCELL_X4 FILLER_79_655 ();
 FILLCELL_X4 FILLER_79_664 ();
 FILLCELL_X1 FILLER_79_668 ();
 FILLCELL_X4 FILLER_79_683 ();
 FILLCELL_X2 FILLER_79_731 ();
 FILLCELL_X4 FILLER_79_740 ();
 FILLCELL_X2 FILLER_79_744 ();
 FILLCELL_X1 FILLER_79_746 ();
 FILLCELL_X4 FILLER_79_749 ();
 FILLCELL_X4 FILLER_79_778 ();
 FILLCELL_X2 FILLER_79_782 ();
 FILLCELL_X4 FILLER_79_814 ();
 FILLCELL_X1 FILLER_79_818 ();
 FILLCELL_X2 FILLER_79_832 ();
 FILLCELL_X2 FILLER_79_845 ();
 FILLCELL_X1 FILLER_79_847 ();
 FILLCELL_X8 FILLER_79_853 ();
 FILLCELL_X1 FILLER_79_861 ();
 FILLCELL_X8 FILLER_79_873 ();
 FILLCELL_X4 FILLER_79_881 ();
 FILLCELL_X2 FILLER_79_885 ();
 FILLCELL_X4 FILLER_79_903 ();
 FILLCELL_X2 FILLER_79_907 ();
 FILLCELL_X4 FILLER_79_924 ();
 FILLCELL_X2 FILLER_79_928 ();
 FILLCELL_X8 FILLER_79_932 ();
 FILLCELL_X16 FILLER_79_947 ();
 FILLCELL_X2 FILLER_79_963 ();
 FILLCELL_X1 FILLER_79_971 ();
 FILLCELL_X1 FILLER_79_981 ();
 FILLCELL_X4 FILLER_79_1041 ();
 FILLCELL_X2 FILLER_79_1045 ();
 FILLCELL_X1 FILLER_79_1047 ();
 FILLCELL_X2 FILLER_79_1063 ();
 FILLCELL_X1 FILLER_79_1065 ();
 FILLCELL_X1 FILLER_79_1073 ();
 FILLCELL_X2 FILLER_79_1077 ();
 FILLCELL_X1 FILLER_79_1079 ();
 FILLCELL_X4 FILLER_79_1083 ();
 FILLCELL_X2 FILLER_79_1087 ();
 FILLCELL_X2 FILLER_79_1094 ();
 FILLCELL_X8 FILLER_79_1109 ();
 FILLCELL_X4 FILLER_79_1117 ();
 FILLCELL_X2 FILLER_79_1130 ();
 FILLCELL_X1 FILLER_79_1132 ();
 FILLCELL_X2 FILLER_79_1136 ();
 FILLCELL_X1 FILLER_79_1138 ();
 FILLCELL_X1 FILLER_79_1165 ();
 FILLCELL_X4 FILLER_79_1190 ();
 FILLCELL_X2 FILLER_79_1207 ();
 FILLCELL_X2 FILLER_79_1214 ();
 FILLCELL_X4 FILLER_79_1222 ();
 FILLCELL_X1 FILLER_79_1226 ();
 FILLCELL_X2 FILLER_79_1234 ();
 FILLCELL_X16 FILLER_80_1 ();
 FILLCELL_X8 FILLER_80_17 ();
 FILLCELL_X1 FILLER_80_30 ();
 FILLCELL_X1 FILLER_80_51 ();
 FILLCELL_X1 FILLER_80_72 ();
 FILLCELL_X1 FILLER_80_80 ();
 FILLCELL_X16 FILLER_80_88 ();
 FILLCELL_X1 FILLER_80_104 ();
 FILLCELL_X32 FILLER_80_112 ();
 FILLCELL_X2 FILLER_80_144 ();
 FILLCELL_X1 FILLER_80_146 ();
 FILLCELL_X1 FILLER_80_170 ();
 FILLCELL_X2 FILLER_80_178 ();
 FILLCELL_X16 FILLER_80_188 ();
 FILLCELL_X1 FILLER_80_217 ();
 FILLCELL_X1 FILLER_80_252 ();
 FILLCELL_X2 FILLER_80_270 ();
 FILLCELL_X2 FILLER_80_292 ();
 FILLCELL_X4 FILLER_80_301 ();
 FILLCELL_X2 FILLER_80_305 ();
 FILLCELL_X1 FILLER_80_323 ();
 FILLCELL_X1 FILLER_80_362 ();
 FILLCELL_X2 FILLER_80_391 ();
 FILLCELL_X1 FILLER_80_400 ();
 FILLCELL_X1 FILLER_80_428 ();
 FILLCELL_X1 FILLER_80_438 ();
 FILLCELL_X4 FILLER_80_460 ();
 FILLCELL_X1 FILLER_80_464 ();
 FILLCELL_X8 FILLER_80_499 ();
 FILLCELL_X4 FILLER_80_523 ();
 FILLCELL_X2 FILLER_80_543 ();
 FILLCELL_X1 FILLER_80_545 ();
 FILLCELL_X1 FILLER_80_553 ();
 FILLCELL_X1 FILLER_80_558 ();
 FILLCELL_X1 FILLER_80_570 ();
 FILLCELL_X1 FILLER_80_577 ();
 FILLCELL_X2 FILLER_80_582 ();
 FILLCELL_X1 FILLER_80_603 ();
 FILLCELL_X2 FILLER_80_609 ();
 FILLCELL_X1 FILLER_80_611 ();
 FILLCELL_X1 FILLER_80_621 ();
 FILLCELL_X1 FILLER_80_642 ();
 FILLCELL_X2 FILLER_80_651 ();
 FILLCELL_X1 FILLER_80_653 ();
 FILLCELL_X2 FILLER_80_657 ();
 FILLCELL_X1 FILLER_80_678 ();
 FILLCELL_X8 FILLER_80_705 ();
 FILLCELL_X2 FILLER_80_713 ();
 FILLCELL_X1 FILLER_80_715 ();
 FILLCELL_X4 FILLER_80_720 ();
 FILLCELL_X2 FILLER_80_724 ();
 FILLCELL_X2 FILLER_80_742 ();
 FILLCELL_X2 FILLER_80_762 ();
 FILLCELL_X1 FILLER_80_764 ();
 FILLCELL_X8 FILLER_80_772 ();
 FILLCELL_X2 FILLER_80_780 ();
 FILLCELL_X1 FILLER_80_782 ();
 FILLCELL_X2 FILLER_80_794 ();
 FILLCELL_X1 FILLER_80_796 ();
 FILLCELL_X4 FILLER_80_804 ();
 FILLCELL_X8 FILLER_80_815 ();
 FILLCELL_X4 FILLER_80_833 ();
 FILLCELL_X16 FILLER_80_844 ();
 FILLCELL_X4 FILLER_80_860 ();
 FILLCELL_X2 FILLER_80_864 ();
 FILLCELL_X4 FILLER_80_883 ();
 FILLCELL_X2 FILLER_80_887 ();
 FILLCELL_X1 FILLER_80_889 ();
 FILLCELL_X1 FILLER_80_918 ();
 FILLCELL_X4 FILLER_80_922 ();
 FILLCELL_X2 FILLER_80_926 ();
 FILLCELL_X8 FILLER_80_931 ();
 FILLCELL_X4 FILLER_80_939 ();
 FILLCELL_X1 FILLER_80_943 ();
 FILLCELL_X8 FILLER_80_950 ();
 FILLCELL_X2 FILLER_80_958 ();
 FILLCELL_X1 FILLER_80_989 ();
 FILLCELL_X4 FILLER_80_1014 ();
 FILLCELL_X4 FILLER_80_1050 ();
 FILLCELL_X2 FILLER_80_1054 ();
 FILLCELL_X2 FILLER_80_1100 ();
 FILLCELL_X8 FILLER_80_1111 ();
 FILLCELL_X2 FILLER_80_1119 ();
 FILLCELL_X1 FILLER_80_1121 ();
 FILLCELL_X8 FILLER_80_1129 ();
 FILLCELL_X16 FILLER_80_1146 ();
 FILLCELL_X4 FILLER_80_1162 ();
 FILLCELL_X2 FILLER_80_1166 ();
 FILLCELL_X1 FILLER_80_1174 ();
 FILLCELL_X2 FILLER_80_1227 ();
 FILLCELL_X1 FILLER_80_1229 ();
 FILLCELL_X2 FILLER_80_1254 ();
 FILLCELL_X1 FILLER_80_1256 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X8 FILLER_81_33 ();
 FILLCELL_X4 FILLER_81_41 ();
 FILLCELL_X2 FILLER_81_45 ();
 FILLCELL_X8 FILLER_81_61 ();
 FILLCELL_X2 FILLER_81_69 ();
 FILLCELL_X1 FILLER_81_71 ();
 FILLCELL_X4 FILLER_81_79 ();
 FILLCELL_X4 FILLER_81_110 ();
 FILLCELL_X2 FILLER_81_114 ();
 FILLCELL_X1 FILLER_81_143 ();
 FILLCELL_X8 FILLER_81_151 ();
 FILLCELL_X2 FILLER_81_159 ();
 FILLCELL_X8 FILLER_81_163 ();
 FILLCELL_X1 FILLER_81_178 ();
 FILLCELL_X4 FILLER_81_185 ();
 FILLCELL_X2 FILLER_81_189 ();
 FILLCELL_X4 FILLER_81_208 ();
 FILLCELL_X2 FILLER_81_219 ();
 FILLCELL_X2 FILLER_81_235 ();
 FILLCELL_X2 FILLER_81_245 ();
 FILLCELL_X8 FILLER_81_274 ();
 FILLCELL_X2 FILLER_81_292 ();
 FILLCELL_X1 FILLER_81_294 ();
 FILLCELL_X4 FILLER_81_315 ();
 FILLCELL_X2 FILLER_81_319 ();
 FILLCELL_X8 FILLER_81_334 ();
 FILLCELL_X2 FILLER_81_342 ();
 FILLCELL_X1 FILLER_81_344 ();
 FILLCELL_X4 FILLER_81_364 ();
 FILLCELL_X2 FILLER_81_368 ();
 FILLCELL_X4 FILLER_81_384 ();
 FILLCELL_X1 FILLER_81_467 ();
 FILLCELL_X4 FILLER_81_502 ();
 FILLCELL_X4 FILLER_81_513 ();
 FILLCELL_X2 FILLER_81_517 ();
 FILLCELL_X1 FILLER_81_519 ();
 FILLCELL_X4 FILLER_81_527 ();
 FILLCELL_X2 FILLER_81_531 ();
 FILLCELL_X1 FILLER_81_533 ();
 FILLCELL_X2 FILLER_81_536 ();
 FILLCELL_X1 FILLER_81_538 ();
 FILLCELL_X8 FILLER_81_546 ();
 FILLCELL_X2 FILLER_81_554 ();
 FILLCELL_X1 FILLER_81_556 ();
 FILLCELL_X8 FILLER_81_568 ();
 FILLCELL_X4 FILLER_81_576 ();
 FILLCELL_X2 FILLER_81_590 ();
 FILLCELL_X1 FILLER_81_592 ();
 FILLCELL_X4 FILLER_81_596 ();
 FILLCELL_X1 FILLER_81_600 ();
 FILLCELL_X4 FILLER_81_606 ();
 FILLCELL_X1 FILLER_81_610 ();
 FILLCELL_X8 FILLER_81_620 ();
 FILLCELL_X2 FILLER_81_628 ();
 FILLCELL_X1 FILLER_81_630 ();
 FILLCELL_X4 FILLER_81_641 ();
 FILLCELL_X2 FILLER_81_654 ();
 FILLCELL_X1 FILLER_81_656 ();
 FILLCELL_X2 FILLER_81_679 ();
 FILLCELL_X1 FILLER_81_681 ();
 FILLCELL_X2 FILLER_81_684 ();
 FILLCELL_X1 FILLER_81_686 ();
 FILLCELL_X2 FILLER_81_691 ();
 FILLCELL_X16 FILLER_81_700 ();
 FILLCELL_X16 FILLER_81_741 ();
 FILLCELL_X4 FILLER_81_757 ();
 FILLCELL_X1 FILLER_81_761 ();
 FILLCELL_X1 FILLER_81_781 ();
 FILLCELL_X2 FILLER_81_795 ();
 FILLCELL_X1 FILLER_81_797 ();
 FILLCELL_X8 FILLER_81_813 ();
 FILLCELL_X4 FILLER_81_821 ();
 FILLCELL_X2 FILLER_81_825 ();
 FILLCELL_X1 FILLER_81_827 ();
 FILLCELL_X4 FILLER_81_841 ();
 FILLCELL_X2 FILLER_81_845 ();
 FILLCELL_X1 FILLER_81_847 ();
 FILLCELL_X8 FILLER_81_862 ();
 FILLCELL_X4 FILLER_81_891 ();
 FILLCELL_X1 FILLER_81_895 ();
 FILLCELL_X2 FILLER_81_911 ();
 FILLCELL_X1 FILLER_81_913 ();
 FILLCELL_X8 FILLER_81_925 ();
 FILLCELL_X2 FILLER_81_933 ();
 FILLCELL_X4 FILLER_81_947 ();
 FILLCELL_X8 FILLER_81_965 ();
 FILLCELL_X1 FILLER_81_973 ();
 FILLCELL_X1 FILLER_81_1074 ();
 FILLCELL_X4 FILLER_81_1099 ();
 FILLCELL_X2 FILLER_81_1103 ();
 FILLCELL_X1 FILLER_81_1105 ();
 FILLCELL_X4 FILLER_81_1128 ();
 FILLCELL_X2 FILLER_81_1132 ();
 FILLCELL_X1 FILLER_81_1142 ();
 FILLCELL_X4 FILLER_81_1155 ();
 FILLCELL_X1 FILLER_81_1159 ();
 FILLCELL_X1 FILLER_81_1178 ();
 FILLCELL_X4 FILLER_81_1188 ();
 FILLCELL_X2 FILLER_81_1207 ();
 FILLCELL_X1 FILLER_81_1209 ();
 FILLCELL_X1 FILLER_81_1256 ();
 FILLCELL_X16 FILLER_82_1 ();
 FILLCELL_X2 FILLER_82_17 ();
 FILLCELL_X1 FILLER_82_19 ();
 FILLCELL_X8 FILLER_82_54 ();
 FILLCELL_X2 FILLER_82_62 ();
 FILLCELL_X1 FILLER_82_78 ();
 FILLCELL_X8 FILLER_82_86 ();
 FILLCELL_X2 FILLER_82_94 ();
 FILLCELL_X1 FILLER_82_96 ();
 FILLCELL_X4 FILLER_82_152 ();
 FILLCELL_X1 FILLER_82_156 ();
 FILLCELL_X2 FILLER_82_166 ();
 FILLCELL_X8 FILLER_82_182 ();
 FILLCELL_X2 FILLER_82_190 ();
 FILLCELL_X1 FILLER_82_192 ();
 FILLCELL_X1 FILLER_82_233 ();
 FILLCELL_X4 FILLER_82_269 ();
 FILLCELL_X4 FILLER_82_277 ();
 FILLCELL_X2 FILLER_82_284 ();
 FILLCELL_X4 FILLER_82_293 ();
 FILLCELL_X8 FILLER_82_301 ();
 FILLCELL_X4 FILLER_82_309 ();
 FILLCELL_X2 FILLER_82_313 ();
 FILLCELL_X8 FILLER_82_322 ();
 FILLCELL_X4 FILLER_82_330 ();
 FILLCELL_X1 FILLER_82_334 ();
 FILLCELL_X2 FILLER_82_374 ();
 FILLCELL_X2 FILLER_82_403 ();
 FILLCELL_X1 FILLER_82_405 ();
 FILLCELL_X4 FILLER_82_420 ();
 FILLCELL_X2 FILLER_82_442 ();
 FILLCELL_X2 FILLER_82_451 ();
 FILLCELL_X1 FILLER_82_453 ();
 FILLCELL_X8 FILLER_82_467 ();
 FILLCELL_X2 FILLER_82_475 ();
 FILLCELL_X1 FILLER_82_477 ();
 FILLCELL_X8 FILLER_82_499 ();
 FILLCELL_X4 FILLER_82_507 ();
 FILLCELL_X2 FILLER_82_511 ();
 FILLCELL_X1 FILLER_82_513 ();
 FILLCELL_X1 FILLER_82_535 ();
 FILLCELL_X8 FILLER_82_543 ();
 FILLCELL_X4 FILLER_82_551 ();
 FILLCELL_X8 FILLER_82_623 ();
 FILLCELL_X8 FILLER_82_632 ();
 FILLCELL_X1 FILLER_82_640 ();
 FILLCELL_X1 FILLER_82_658 ();
 FILLCELL_X1 FILLER_82_662 ();
 FILLCELL_X2 FILLER_82_666 ();
 FILLCELL_X4 FILLER_82_683 ();
 FILLCELL_X2 FILLER_82_687 ();
 FILLCELL_X1 FILLER_82_689 ();
 FILLCELL_X4 FILLER_82_710 ();
 FILLCELL_X2 FILLER_82_714 ();
 FILLCELL_X1 FILLER_82_716 ();
 FILLCELL_X4 FILLER_82_720 ();
 FILLCELL_X1 FILLER_82_724 ();
 FILLCELL_X2 FILLER_82_732 ();
 FILLCELL_X4 FILLER_82_743 ();
 FILLCELL_X1 FILLER_82_747 ();
 FILLCELL_X16 FILLER_82_755 ();
 FILLCELL_X8 FILLER_82_771 ();
 FILLCELL_X1 FILLER_82_779 ();
 FILLCELL_X8 FILLER_82_787 ();
 FILLCELL_X1 FILLER_82_795 ();
 FILLCELL_X16 FILLER_82_810 ();
 FILLCELL_X8 FILLER_82_826 ();
 FILLCELL_X2 FILLER_82_834 ();
 FILLCELL_X8 FILLER_82_847 ();
 FILLCELL_X1 FILLER_82_860 ();
 FILLCELL_X4 FILLER_82_872 ();
 FILLCELL_X2 FILLER_82_876 ();
 FILLCELL_X1 FILLER_82_888 ();
 FILLCELL_X4 FILLER_82_892 ();
 FILLCELL_X4 FILLER_82_911 ();
 FILLCELL_X1 FILLER_82_915 ();
 FILLCELL_X8 FILLER_82_931 ();
 FILLCELL_X2 FILLER_82_951 ();
 FILLCELL_X1 FILLER_82_953 ();
 FILLCELL_X1 FILLER_82_968 ();
 FILLCELL_X4 FILLER_82_984 ();
 FILLCELL_X1 FILLER_82_988 ();
 FILLCELL_X8 FILLER_82_993 ();
 FILLCELL_X2 FILLER_82_1001 ();
 FILLCELL_X1 FILLER_82_1009 ();
 FILLCELL_X2 FILLER_82_1039 ();
 FILLCELL_X4 FILLER_82_1086 ();
 FILLCELL_X1 FILLER_82_1094 ();
 FILLCELL_X2 FILLER_82_1117 ();
 FILLCELL_X1 FILLER_82_1119 ();
 FILLCELL_X4 FILLER_82_1122 ();
 FILLCELL_X2 FILLER_82_1126 ();
 FILLCELL_X1 FILLER_82_1128 ();
 FILLCELL_X4 FILLER_82_1150 ();
 FILLCELL_X2 FILLER_82_1154 ();
 FILLCELL_X2 FILLER_82_1170 ();
 FILLCELL_X2 FILLER_82_1189 ();
 FILLCELL_X2 FILLER_82_1208 ();
 FILLCELL_X2 FILLER_82_1217 ();
 FILLCELL_X1 FILLER_82_1227 ();
 FILLCELL_X1 FILLER_82_1242 ();
 FILLCELL_X4 FILLER_83_4 ();
 FILLCELL_X1 FILLER_83_8 ();
 FILLCELL_X2 FILLER_83_49 ();
 FILLCELL_X8 FILLER_83_91 ();
 FILLCELL_X4 FILLER_83_99 ();
 FILLCELL_X8 FILLER_83_120 ();
 FILLCELL_X4 FILLER_83_165 ();
 FILLCELL_X1 FILLER_83_169 ();
 FILLCELL_X4 FILLER_83_174 ();
 FILLCELL_X2 FILLER_83_185 ();
 FILLCELL_X1 FILLER_83_187 ();
 FILLCELL_X2 FILLER_83_208 ();
 FILLCELL_X1 FILLER_83_210 ();
 FILLCELL_X2 FILLER_83_259 ();
 FILLCELL_X8 FILLER_83_295 ();
 FILLCELL_X1 FILLER_83_303 ();
 FILLCELL_X16 FILLER_83_306 ();
 FILLCELL_X2 FILLER_83_322 ();
 FILLCELL_X4 FILLER_83_337 ();
 FILLCELL_X2 FILLER_83_355 ();
 FILLCELL_X1 FILLER_83_357 ();
 FILLCELL_X16 FILLER_83_385 ();
 FILLCELL_X2 FILLER_83_415 ();
 FILLCELL_X1 FILLER_83_417 ();
 FILLCELL_X4 FILLER_83_434 ();
 FILLCELL_X2 FILLER_83_438 ();
 FILLCELL_X1 FILLER_83_447 ();
 FILLCELL_X4 FILLER_83_458 ();
 FILLCELL_X4 FILLER_83_489 ();
 FILLCELL_X1 FILLER_83_493 ();
 FILLCELL_X8 FILLER_83_521 ();
 FILLCELL_X1 FILLER_83_529 ();
 FILLCELL_X4 FILLER_83_550 ();
 FILLCELL_X2 FILLER_83_554 ();
 FILLCELL_X2 FILLER_83_565 ();
 FILLCELL_X1 FILLER_83_567 ();
 FILLCELL_X8 FILLER_83_573 ();
 FILLCELL_X4 FILLER_83_581 ();
 FILLCELL_X1 FILLER_83_606 ();
 FILLCELL_X8 FILLER_83_618 ();
 FILLCELL_X2 FILLER_83_626 ();
 FILLCELL_X1 FILLER_83_628 ();
 FILLCELL_X2 FILLER_83_643 ();
 FILLCELL_X1 FILLER_83_645 ();
 FILLCELL_X4 FILLER_83_670 ();
 FILLCELL_X1 FILLER_83_674 ();
 FILLCELL_X8 FILLER_83_695 ();
 FILLCELL_X4 FILLER_83_703 ();
 FILLCELL_X2 FILLER_83_707 ();
 FILLCELL_X4 FILLER_83_716 ();
 FILLCELL_X2 FILLER_83_720 ();
 FILLCELL_X8 FILLER_83_728 ();
 FILLCELL_X4 FILLER_83_736 ();
 FILLCELL_X2 FILLER_83_740 ();
 FILLCELL_X4 FILLER_83_752 ();
 FILLCELL_X2 FILLER_83_756 ();
 FILLCELL_X8 FILLER_83_765 ();
 FILLCELL_X8 FILLER_83_794 ();
 FILLCELL_X1 FILLER_83_802 ();
 FILLCELL_X1 FILLER_83_806 ();
 FILLCELL_X8 FILLER_83_818 ();
 FILLCELL_X4 FILLER_83_826 ();
 FILLCELL_X2 FILLER_83_830 ();
 FILLCELL_X8 FILLER_83_835 ();
 FILLCELL_X2 FILLER_83_843 ();
 FILLCELL_X4 FILLER_83_852 ();
 FILLCELL_X8 FILLER_83_866 ();
 FILLCELL_X2 FILLER_83_874 ();
 FILLCELL_X2 FILLER_83_878 ();
 FILLCELL_X8 FILLER_83_884 ();
 FILLCELL_X4 FILLER_83_892 ();
 FILLCELL_X2 FILLER_83_896 ();
 FILLCELL_X8 FILLER_83_933 ();
 FILLCELL_X4 FILLER_83_941 ();
 FILLCELL_X8 FILLER_83_958 ();
 FILLCELL_X4 FILLER_83_966 ();
 FILLCELL_X32 FILLER_83_981 ();
 FILLCELL_X2 FILLER_83_1048 ();
 FILLCELL_X1 FILLER_83_1088 ();
 FILLCELL_X1 FILLER_83_1102 ();
 FILLCELL_X1 FILLER_83_1121 ();
 FILLCELL_X2 FILLER_83_1129 ();
 FILLCELL_X1 FILLER_83_1131 ();
 FILLCELL_X2 FILLER_83_1144 ();
 FILLCELL_X4 FILLER_83_1148 ();
 FILLCELL_X1 FILLER_83_1152 ();
 FILLCELL_X2 FILLER_83_1158 ();
 FILLCELL_X1 FILLER_83_1160 ();
 FILLCELL_X16 FILLER_83_1175 ();
 FILLCELL_X1 FILLER_83_1191 ();
 FILLCELL_X8 FILLER_83_1199 ();
 FILLCELL_X4 FILLER_83_1207 ();
 FILLCELL_X1 FILLER_83_1211 ();
 FILLCELL_X8 FILLER_83_1219 ();
 FILLCELL_X4 FILLER_83_1227 ();
 FILLCELL_X2 FILLER_83_1231 ();
 FILLCELL_X2 FILLER_83_1257 ();
 FILLCELL_X1 FILLER_83_1259 ();
 FILLCELL_X2 FILLER_84_1 ();
 FILLCELL_X1 FILLER_84_3 ();
 FILLCELL_X2 FILLER_84_36 ();
 FILLCELL_X4 FILLER_84_59 ();
 FILLCELL_X1 FILLER_84_70 ();
 FILLCELL_X2 FILLER_84_78 ();
 FILLCELL_X1 FILLER_84_80 ();
 FILLCELL_X2 FILLER_84_102 ();
 FILLCELL_X8 FILLER_84_107 ();
 FILLCELL_X4 FILLER_84_115 ();
 FILLCELL_X2 FILLER_84_119 ();
 FILLCELL_X16 FILLER_84_138 ();
 FILLCELL_X2 FILLER_84_154 ();
 FILLCELL_X2 FILLER_84_176 ();
 FILLCELL_X1 FILLER_84_178 ();
 FILLCELL_X4 FILLER_84_190 ();
 FILLCELL_X2 FILLER_84_194 ();
 FILLCELL_X1 FILLER_84_196 ();
 FILLCELL_X8 FILLER_84_231 ();
 FILLCELL_X4 FILLER_84_239 ();
 FILLCELL_X16 FILLER_84_246 ();
 FILLCELL_X4 FILLER_84_262 ();
 FILLCELL_X1 FILLER_84_266 ();
 FILLCELL_X4 FILLER_84_274 ();
 FILLCELL_X1 FILLER_84_278 ();
 FILLCELL_X2 FILLER_84_287 ();
 FILLCELL_X1 FILLER_84_289 ();
 FILLCELL_X8 FILLER_84_297 ();
 FILLCELL_X1 FILLER_84_305 ();
 FILLCELL_X8 FILLER_84_327 ();
 FILLCELL_X4 FILLER_84_335 ();
 FILLCELL_X2 FILLER_84_339 ();
 FILLCELL_X4 FILLER_84_357 ();
 FILLCELL_X2 FILLER_84_361 ();
 FILLCELL_X1 FILLER_84_363 ();
 FILLCELL_X2 FILLER_84_373 ();
 FILLCELL_X1 FILLER_84_375 ();
 FILLCELL_X1 FILLER_84_383 ();
 FILLCELL_X16 FILLER_84_427 ();
 FILLCELL_X4 FILLER_84_443 ();
 FILLCELL_X4 FILLER_84_460 ();
 FILLCELL_X1 FILLER_84_464 ();
 FILLCELL_X1 FILLER_84_496 ();
 FILLCELL_X4 FILLER_84_532 ();
 FILLCELL_X2 FILLER_84_536 ();
 FILLCELL_X4 FILLER_84_545 ();
 FILLCELL_X1 FILLER_84_549 ();
 FILLCELL_X4 FILLER_84_552 ();
 FILLCELL_X2 FILLER_84_556 ();
 FILLCELL_X1 FILLER_84_558 ();
 FILLCELL_X2 FILLER_84_578 ();
 FILLCELL_X4 FILLER_84_590 ();
 FILLCELL_X1 FILLER_84_594 ();
 FILLCELL_X2 FILLER_84_602 ();
 FILLCELL_X1 FILLER_84_604 ();
 FILLCELL_X1 FILLER_84_608 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X4 FILLER_84_632 ();
 FILLCELL_X2 FILLER_84_636 ();
 FILLCELL_X4 FILLER_84_653 ();
 FILLCELL_X2 FILLER_84_657 ();
 FILLCELL_X1 FILLER_84_659 ();
 FILLCELL_X8 FILLER_84_673 ();
 FILLCELL_X4 FILLER_84_681 ();
 FILLCELL_X1 FILLER_84_685 ();
 FILLCELL_X8 FILLER_84_695 ();
 FILLCELL_X1 FILLER_84_703 ();
 FILLCELL_X4 FILLER_84_707 ();
 FILLCELL_X2 FILLER_84_711 ();
 FILLCELL_X1 FILLER_84_713 ();
 FILLCELL_X8 FILLER_84_717 ();
 FILLCELL_X1 FILLER_84_725 ();
 FILLCELL_X2 FILLER_84_733 ();
 FILLCELL_X1 FILLER_84_735 ();
 FILLCELL_X4 FILLER_84_753 ();
 FILLCELL_X2 FILLER_84_757 ();
 FILLCELL_X2 FILLER_84_766 ();
 FILLCELL_X1 FILLER_84_771 ();
 FILLCELL_X4 FILLER_84_779 ();
 FILLCELL_X8 FILLER_84_792 ();
 FILLCELL_X1 FILLER_84_800 ();
 FILLCELL_X8 FILLER_84_810 ();
 FILLCELL_X4 FILLER_84_818 ();
 FILLCELL_X1 FILLER_84_832 ();
 FILLCELL_X2 FILLER_84_836 ();
 FILLCELL_X2 FILLER_84_842 ();
 FILLCELL_X1 FILLER_84_844 ();
 FILLCELL_X8 FILLER_84_850 ();
 FILLCELL_X1 FILLER_84_858 ();
 FILLCELL_X4 FILLER_84_869 ();
 FILLCELL_X2 FILLER_84_898 ();
 FILLCELL_X1 FILLER_84_900 ();
 FILLCELL_X2 FILLER_84_903 ();
 FILLCELL_X4 FILLER_84_908 ();
 FILLCELL_X2 FILLER_84_916 ();
 FILLCELL_X2 FILLER_84_928 ();
 FILLCELL_X4 FILLER_84_932 ();
 FILLCELL_X1 FILLER_84_936 ();
 FILLCELL_X2 FILLER_84_950 ();
 FILLCELL_X1 FILLER_84_958 ();
 FILLCELL_X1 FILLER_84_966 ();
 FILLCELL_X8 FILLER_84_983 ();
 FILLCELL_X4 FILLER_84_991 ();
 FILLCELL_X2 FILLER_84_995 ();
 FILLCELL_X1 FILLER_84_997 ();
 FILLCELL_X4 FILLER_84_1015 ();
 FILLCELL_X1 FILLER_84_1019 ();
 FILLCELL_X2 FILLER_84_1032 ();
 FILLCELL_X1 FILLER_84_1034 ();
 FILLCELL_X2 FILLER_84_1045 ();
 FILLCELL_X1 FILLER_84_1054 ();
 FILLCELL_X1 FILLER_84_1059 ();
 FILLCELL_X1 FILLER_84_1092 ();
 FILLCELL_X1 FILLER_84_1107 ();
 FILLCELL_X8 FILLER_84_1118 ();
 FILLCELL_X2 FILLER_84_1134 ();
 FILLCELL_X2 FILLER_84_1144 ();
 FILLCELL_X2 FILLER_84_1151 ();
 FILLCELL_X1 FILLER_84_1153 ();
 FILLCELL_X4 FILLER_84_1157 ();
 FILLCELL_X1 FILLER_84_1161 ();
 FILLCELL_X1 FILLER_84_1175 ();
 FILLCELL_X4 FILLER_84_1200 ();
 FILLCELL_X1 FILLER_84_1204 ();
 FILLCELL_X4 FILLER_84_1222 ();
 FILLCELL_X2 FILLER_84_1226 ();
 FILLCELL_X16 FILLER_84_1235 ();
 FILLCELL_X8 FILLER_84_1251 ();
 FILLCELL_X1 FILLER_84_1259 ();
 FILLCELL_X1 FILLER_85_1 ();
 FILLCELL_X1 FILLER_85_22 ();
 FILLCELL_X1 FILLER_85_30 ();
 FILLCELL_X2 FILLER_85_38 ();
 FILLCELL_X16 FILLER_85_54 ();
 FILLCELL_X4 FILLER_85_91 ();
 FILLCELL_X2 FILLER_85_95 ();
 FILLCELL_X1 FILLER_85_97 ();
 FILLCELL_X8 FILLER_85_108 ();
 FILLCELL_X8 FILLER_85_129 ();
 FILLCELL_X16 FILLER_85_157 ();
 FILLCELL_X2 FILLER_85_173 ();
 FILLCELL_X8 FILLER_85_182 ();
 FILLCELL_X4 FILLER_85_197 ();
 FILLCELL_X2 FILLER_85_201 ();
 FILLCELL_X8 FILLER_85_229 ();
 FILLCELL_X4 FILLER_85_244 ();
 FILLCELL_X2 FILLER_85_248 ();
 FILLCELL_X1 FILLER_85_250 ();
 FILLCELL_X2 FILLER_85_259 ();
 FILLCELL_X1 FILLER_85_288 ();
 FILLCELL_X4 FILLER_85_309 ();
 FILLCELL_X1 FILLER_85_313 ();
 FILLCELL_X1 FILLER_85_336 ();
 FILLCELL_X1 FILLER_85_355 ();
 FILLCELL_X8 FILLER_85_363 ();
 FILLCELL_X4 FILLER_85_371 ();
 FILLCELL_X2 FILLER_85_375 ();
 FILLCELL_X1 FILLER_85_377 ();
 FILLCELL_X16 FILLER_85_398 ();
 FILLCELL_X1 FILLER_85_414 ();
 FILLCELL_X8 FILLER_85_436 ();
 FILLCELL_X2 FILLER_85_444 ();
 FILLCELL_X1 FILLER_85_446 ();
 FILLCELL_X4 FILLER_85_451 ();
 FILLCELL_X2 FILLER_85_455 ();
 FILLCELL_X16 FILLER_85_464 ();
 FILLCELL_X1 FILLER_85_480 ();
 FILLCELL_X1 FILLER_85_488 ();
 FILLCELL_X2 FILLER_85_492 ();
 FILLCELL_X16 FILLER_85_521 ();
 FILLCELL_X8 FILLER_85_537 ();
 FILLCELL_X4 FILLER_85_545 ();
 FILLCELL_X2 FILLER_85_549 ();
 FILLCELL_X8 FILLER_85_559 ();
 FILLCELL_X2 FILLER_85_583 ();
 FILLCELL_X1 FILLER_85_598 ();
 FILLCELL_X2 FILLER_85_613 ();
 FILLCELL_X1 FILLER_85_615 ();
 FILLCELL_X16 FILLER_85_624 ();
 FILLCELL_X8 FILLER_85_640 ();
 FILLCELL_X8 FILLER_85_665 ();
 FILLCELL_X1 FILLER_85_673 ();
 FILLCELL_X4 FILLER_85_679 ();
 FILLCELL_X2 FILLER_85_694 ();
 FILLCELL_X1 FILLER_85_714 ();
 FILLCELL_X8 FILLER_85_729 ();
 FILLCELL_X4 FILLER_85_737 ();
 FILLCELL_X4 FILLER_85_750 ();
 FILLCELL_X2 FILLER_85_754 ();
 FILLCELL_X2 FILLER_85_761 ();
 FILLCELL_X1 FILLER_85_767 ();
 FILLCELL_X2 FILLER_85_775 ();
 FILLCELL_X2 FILLER_85_784 ();
 FILLCELL_X4 FILLER_85_793 ();
 FILLCELL_X2 FILLER_85_804 ();
 FILLCELL_X4 FILLER_85_824 ();
 FILLCELL_X1 FILLER_85_849 ();
 FILLCELL_X2 FILLER_85_860 ();
 FILLCELL_X2 FILLER_85_872 ();
 FILLCELL_X1 FILLER_85_874 ();
 FILLCELL_X8 FILLER_85_880 ();
 FILLCELL_X2 FILLER_85_888 ();
 FILLCELL_X1 FILLER_85_901 ();
 FILLCELL_X8 FILLER_85_912 ();
 FILLCELL_X1 FILLER_85_966 ();
 FILLCELL_X2 FILLER_85_992 ();
 FILLCELL_X1 FILLER_85_994 ();
 FILLCELL_X1 FILLER_85_999 ();
 FILLCELL_X1 FILLER_85_1010 ();
 FILLCELL_X1 FILLER_85_1021 ();
 FILLCELL_X2 FILLER_85_1051 ();
 FILLCELL_X1 FILLER_85_1057 ();
 FILLCELL_X1 FILLER_85_1060 ();
 FILLCELL_X2 FILLER_85_1095 ();
 FILLCELL_X16 FILLER_85_1107 ();
 FILLCELL_X2 FILLER_85_1136 ();
 FILLCELL_X1 FILLER_85_1138 ();
 FILLCELL_X16 FILLER_85_1165 ();
 FILLCELL_X2 FILLER_85_1181 ();
 FILLCELL_X4 FILLER_85_1188 ();
 FILLCELL_X1 FILLER_85_1192 ();
 FILLCELL_X4 FILLER_85_1200 ();
 FILLCELL_X2 FILLER_85_1204 ();
 FILLCELL_X1 FILLER_85_1206 ();
 FILLCELL_X8 FILLER_85_1214 ();
 FILLCELL_X8 FILLER_85_1246 ();
 FILLCELL_X4 FILLER_85_1254 ();
 FILLCELL_X2 FILLER_85_1258 ();
 FILLCELL_X4 FILLER_86_1 ();
 FILLCELL_X1 FILLER_86_5 ();
 FILLCELL_X16 FILLER_86_36 ();
 FILLCELL_X1 FILLER_86_52 ();
 FILLCELL_X32 FILLER_86_80 ();
 FILLCELL_X1 FILLER_86_112 ();
 FILLCELL_X4 FILLER_86_120 ();
 FILLCELL_X2 FILLER_86_124 ();
 FILLCELL_X8 FILLER_86_183 ();
 FILLCELL_X1 FILLER_86_191 ();
 FILLCELL_X2 FILLER_86_213 ();
 FILLCELL_X4 FILLER_86_242 ();
 FILLCELL_X8 FILLER_86_273 ();
 FILLCELL_X4 FILLER_86_281 ();
 FILLCELL_X2 FILLER_86_287 ();
 FILLCELL_X1 FILLER_86_289 ();
 FILLCELL_X8 FILLER_86_297 ();
 FILLCELL_X4 FILLER_86_305 ();
 FILLCELL_X1 FILLER_86_309 ();
 FILLCELL_X8 FILLER_86_317 ();
 FILLCELL_X2 FILLER_86_325 ();
 FILLCELL_X4 FILLER_86_397 ();
 FILLCELL_X2 FILLER_86_401 ();
 FILLCELL_X1 FILLER_86_403 ();
 FILLCELL_X4 FILLER_86_407 ();
 FILLCELL_X2 FILLER_86_411 ();
 FILLCELL_X1 FILLER_86_413 ();
 FILLCELL_X8 FILLER_86_433 ();
 FILLCELL_X2 FILLER_86_441 ();
 FILLCELL_X2 FILLER_86_447 ();
 FILLCELL_X1 FILLER_86_449 ();
 FILLCELL_X2 FILLER_86_454 ();
 FILLCELL_X1 FILLER_86_460 ();
 FILLCELL_X2 FILLER_86_468 ();
 FILLCELL_X4 FILLER_86_477 ();
 FILLCELL_X2 FILLER_86_481 ();
 FILLCELL_X1 FILLER_86_488 ();
 FILLCELL_X1 FILLER_86_497 ();
 FILLCELL_X16 FILLER_86_516 ();
 FILLCELL_X4 FILLER_86_532 ();
 FILLCELL_X2 FILLER_86_536 ();
 FILLCELL_X1 FILLER_86_538 ();
 FILLCELL_X8 FILLER_86_573 ();
 FILLCELL_X2 FILLER_86_581 ();
 FILLCELL_X1 FILLER_86_590 ();
 FILLCELL_X2 FILLER_86_596 ();
 FILLCELL_X1 FILLER_86_601 ();
 FILLCELL_X1 FILLER_86_609 ();
 FILLCELL_X1 FILLER_86_613 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X2 FILLER_86_632 ();
 FILLCELL_X4 FILLER_86_641 ();
 FILLCELL_X2 FILLER_86_645 ();
 FILLCELL_X1 FILLER_86_647 ();
 FILLCELL_X4 FILLER_86_655 ();
 FILLCELL_X16 FILLER_86_671 ();
 FILLCELL_X4 FILLER_86_687 ();
 FILLCELL_X2 FILLER_86_691 ();
 FILLCELL_X1 FILLER_86_693 ();
 FILLCELL_X4 FILLER_86_707 ();
 FILLCELL_X8 FILLER_86_718 ();
 FILLCELL_X1 FILLER_86_726 ();
 FILLCELL_X16 FILLER_86_730 ();
 FILLCELL_X4 FILLER_86_760 ();
 FILLCELL_X2 FILLER_86_764 ();
 FILLCELL_X1 FILLER_86_766 ();
 FILLCELL_X8 FILLER_86_781 ();
 FILLCELL_X1 FILLER_86_789 ();
 FILLCELL_X8 FILLER_86_797 ();
 FILLCELL_X8 FILLER_86_812 ();
 FILLCELL_X1 FILLER_86_820 ();
 FILLCELL_X8 FILLER_86_828 ();
 FILLCELL_X2 FILLER_86_836 ();
 FILLCELL_X1 FILLER_86_838 ();
 FILLCELL_X8 FILLER_86_851 ();
 FILLCELL_X2 FILLER_86_859 ();
 FILLCELL_X1 FILLER_86_861 ();
 FILLCELL_X2 FILLER_86_866 ();
 FILLCELL_X1 FILLER_86_868 ();
 FILLCELL_X2 FILLER_86_876 ();
 FILLCELL_X2 FILLER_86_883 ();
 FILLCELL_X1 FILLER_86_885 ();
 FILLCELL_X8 FILLER_86_893 ();
 FILLCELL_X1 FILLER_86_901 ();
 FILLCELL_X4 FILLER_86_906 ();
 FILLCELL_X2 FILLER_86_915 ();
 FILLCELL_X8 FILLER_86_921 ();
 FILLCELL_X4 FILLER_86_933 ();
 FILLCELL_X8 FILLER_86_940 ();
 FILLCELL_X4 FILLER_86_948 ();
 FILLCELL_X2 FILLER_86_952 ();
 FILLCELL_X2 FILLER_86_961 ();
 FILLCELL_X2 FILLER_86_983 ();
 FILLCELL_X1 FILLER_86_985 ();
 FILLCELL_X2 FILLER_86_1008 ();
 FILLCELL_X4 FILLER_86_1014 ();
 FILLCELL_X2 FILLER_86_1018 ();
 FILLCELL_X1 FILLER_86_1020 ();
 FILLCELL_X2 FILLER_86_1038 ();
 FILLCELL_X4 FILLER_86_1054 ();
 FILLCELL_X8 FILLER_86_1068 ();
 FILLCELL_X4 FILLER_86_1076 ();
 FILLCELL_X1 FILLER_86_1080 ();
 FILLCELL_X16 FILLER_86_1091 ();
 FILLCELL_X1 FILLER_86_1130 ();
 FILLCELL_X2 FILLER_86_1140 ();
 FILLCELL_X2 FILLER_86_1149 ();
 FILLCELL_X1 FILLER_86_1164 ();
 FILLCELL_X1 FILLER_86_1205 ();
 FILLCELL_X16 FILLER_86_1237 ();
 FILLCELL_X4 FILLER_86_1253 ();
 FILLCELL_X2 FILLER_86_1257 ();
 FILLCELL_X1 FILLER_86_1259 ();
 FILLCELL_X4 FILLER_87_1 ();
 FILLCELL_X1 FILLER_87_5 ();
 FILLCELL_X8 FILLER_87_54 ();
 FILLCELL_X2 FILLER_87_89 ();
 FILLCELL_X2 FILLER_87_118 ();
 FILLCELL_X4 FILLER_87_134 ();
 FILLCELL_X4 FILLER_87_145 ();
 FILLCELL_X2 FILLER_87_149 ();
 FILLCELL_X8 FILLER_87_160 ();
 FILLCELL_X1 FILLER_87_178 ();
 FILLCELL_X2 FILLER_87_182 ();
 FILLCELL_X16 FILLER_87_198 ();
 FILLCELL_X2 FILLER_87_221 ();
 FILLCELL_X8 FILLER_87_230 ();
 FILLCELL_X1 FILLER_87_238 ();
 FILLCELL_X4 FILLER_87_253 ();
 FILLCELL_X2 FILLER_87_257 ();
 FILLCELL_X1 FILLER_87_259 ();
 FILLCELL_X2 FILLER_87_287 ();
 FILLCELL_X2 FILLER_87_320 ();
 FILLCELL_X1 FILLER_87_417 ();
 FILLCELL_X1 FILLER_87_425 ();
 FILLCELL_X2 FILLER_87_433 ();
 FILLCELL_X1 FILLER_87_435 ();
 FILLCELL_X1 FILLER_87_443 ();
 FILLCELL_X1 FILLER_87_474 ();
 FILLCELL_X1 FILLER_87_482 ();
 FILLCELL_X4 FILLER_87_529 ();
 FILLCELL_X2 FILLER_87_533 ();
 FILLCELL_X1 FILLER_87_535 ();
 FILLCELL_X2 FILLER_87_549 ();
 FILLCELL_X8 FILLER_87_565 ();
 FILLCELL_X2 FILLER_87_573 ();
 FILLCELL_X1 FILLER_87_613 ();
 FILLCELL_X32 FILLER_87_619 ();
 FILLCELL_X4 FILLER_87_651 ();
 FILLCELL_X8 FILLER_87_658 ();
 FILLCELL_X2 FILLER_87_666 ();
 FILLCELL_X4 FILLER_87_686 ();
 FILLCELL_X1 FILLER_87_690 ();
 FILLCELL_X1 FILLER_87_698 ();
 FILLCELL_X4 FILLER_87_735 ();
 FILLCELL_X2 FILLER_87_739 ();
 FILLCELL_X1 FILLER_87_741 ();
 FILLCELL_X4 FILLER_87_756 ();
 FILLCELL_X1 FILLER_87_760 ();
 FILLCELL_X16 FILLER_87_768 ();
 FILLCELL_X2 FILLER_87_784 ();
 FILLCELL_X1 FILLER_87_786 ();
 FILLCELL_X4 FILLER_87_815 ();
 FILLCELL_X2 FILLER_87_819 ();
 FILLCELL_X1 FILLER_87_821 ();
 FILLCELL_X4 FILLER_87_829 ();
 FILLCELL_X2 FILLER_87_833 ();
 FILLCELL_X1 FILLER_87_835 ();
 FILLCELL_X4 FILLER_87_840 ();
 FILLCELL_X2 FILLER_87_844 ();
 FILLCELL_X2 FILLER_87_849 ();
 FILLCELL_X1 FILLER_87_878 ();
 FILLCELL_X2 FILLER_87_904 ();
 FILLCELL_X4 FILLER_87_914 ();
 FILLCELL_X1 FILLER_87_918 ();
 FILLCELL_X4 FILLER_87_941 ();
 FILLCELL_X2 FILLER_87_957 ();
 FILLCELL_X8 FILLER_87_1015 ();
 FILLCELL_X2 FILLER_87_1023 ();
 FILLCELL_X1 FILLER_87_1025 ();
 FILLCELL_X1 FILLER_87_1033 ();
 FILLCELL_X4 FILLER_87_1043 ();
 FILLCELL_X4 FILLER_87_1056 ();
 FILLCELL_X8 FILLER_87_1082 ();
 FILLCELL_X4 FILLER_87_1090 ();
 FILLCELL_X4 FILLER_87_1097 ();
 FILLCELL_X1 FILLER_87_1101 ();
 FILLCELL_X2 FILLER_87_1142 ();
 FILLCELL_X1 FILLER_87_1144 ();
 FILLCELL_X16 FILLER_87_1185 ();
 FILLCELL_X4 FILLER_87_1201 ();
 FILLCELL_X1 FILLER_87_1205 ();
 FILLCELL_X32 FILLER_87_1223 ();
 FILLCELL_X4 FILLER_87_1255 ();
 FILLCELL_X1 FILLER_87_1259 ();
 FILLCELL_X16 FILLER_88_1 ();
 FILLCELL_X4 FILLER_88_17 ();
 FILLCELL_X2 FILLER_88_28 ();
 FILLCELL_X2 FILLER_88_80 ();
 FILLCELL_X1 FILLER_88_82 ();
 FILLCELL_X4 FILLER_88_95 ();
 FILLCELL_X1 FILLER_88_126 ();
 FILLCELL_X8 FILLER_88_187 ();
 FILLCELL_X2 FILLER_88_195 ();
 FILLCELL_X4 FILLER_88_237 ();
 FILLCELL_X2 FILLER_88_241 ();
 FILLCELL_X4 FILLER_88_268 ();
 FILLCELL_X16 FILLER_88_292 ();
 FILLCELL_X8 FILLER_88_308 ();
 FILLCELL_X2 FILLER_88_316 ();
 FILLCELL_X2 FILLER_88_332 ();
 FILLCELL_X1 FILLER_88_334 ();
 FILLCELL_X1 FILLER_88_344 ();
 FILLCELL_X2 FILLER_88_356 ();
 FILLCELL_X1 FILLER_88_358 ();
 FILLCELL_X2 FILLER_88_375 ();
 FILLCELL_X1 FILLER_88_377 ();
 FILLCELL_X1 FILLER_88_404 ();
 FILLCELL_X2 FILLER_88_437 ();
 FILLCELL_X1 FILLER_88_446 ();
 FILLCELL_X4 FILLER_88_460 ();
 FILLCELL_X2 FILLER_88_467 ();
 FILLCELL_X2 FILLER_88_507 ();
 FILLCELL_X1 FILLER_88_522 ();
 FILLCELL_X8 FILLER_88_536 ();
 FILLCELL_X1 FILLER_88_544 ();
 FILLCELL_X2 FILLER_88_557 ();
 FILLCELL_X8 FILLER_88_568 ();
 FILLCELL_X8 FILLER_88_581 ();
 FILLCELL_X2 FILLER_88_597 ();
 FILLCELL_X4 FILLER_88_616 ();
 FILLCELL_X2 FILLER_88_620 ();
 FILLCELL_X1 FILLER_88_622 ();
 FILLCELL_X1 FILLER_88_630 ();
 FILLCELL_X8 FILLER_88_632 ();
 FILLCELL_X16 FILLER_88_654 ();
 FILLCELL_X8 FILLER_88_670 ();
 FILLCELL_X2 FILLER_88_678 ();
 FILLCELL_X16 FILLER_88_706 ();
 FILLCELL_X16 FILLER_88_729 ();
 FILLCELL_X8 FILLER_88_756 ();
 FILLCELL_X2 FILLER_88_778 ();
 FILLCELL_X1 FILLER_88_787 ();
 FILLCELL_X2 FILLER_88_795 ();
 FILLCELL_X8 FILLER_88_804 ();
 FILLCELL_X4 FILLER_88_812 ();
 FILLCELL_X1 FILLER_88_816 ();
 FILLCELL_X2 FILLER_88_819 ();
 FILLCELL_X1 FILLER_88_821 ();
 FILLCELL_X2 FILLER_88_837 ();
 FILLCELL_X2 FILLER_88_846 ();
 FILLCELL_X1 FILLER_88_873 ();
 FILLCELL_X4 FILLER_88_877 ();
 FILLCELL_X2 FILLER_88_881 ();
 FILLCELL_X1 FILLER_88_883 ();
 FILLCELL_X2 FILLER_88_894 ();
 FILLCELL_X1 FILLER_88_896 ();
 FILLCELL_X1 FILLER_88_901 ();
 FILLCELL_X1 FILLER_88_905 ();
 FILLCELL_X1 FILLER_88_916 ();
 FILLCELL_X4 FILLER_88_922 ();
 FILLCELL_X1 FILLER_88_926 ();
 FILLCELL_X1 FILLER_88_932 ();
 FILLCELL_X2 FILLER_88_937 ();
 FILLCELL_X2 FILLER_88_945 ();
 FILLCELL_X1 FILLER_88_947 ();
 FILLCELL_X1 FILLER_88_955 ();
 FILLCELL_X2 FILLER_88_963 ();
 FILLCELL_X4 FILLER_88_977 ();
 FILLCELL_X4 FILLER_88_987 ();
 FILLCELL_X2 FILLER_88_991 ();
 FILLCELL_X1 FILLER_88_993 ();
 FILLCELL_X1 FILLER_88_1001 ();
 FILLCELL_X2 FILLER_88_1012 ();
 FILLCELL_X2 FILLER_88_1018 ();
 FILLCELL_X1 FILLER_88_1020 ();
 FILLCELL_X2 FILLER_88_1031 ();
 FILLCELL_X1 FILLER_88_1033 ();
 FILLCELL_X8 FILLER_88_1038 ();
 FILLCELL_X1 FILLER_88_1046 ();
 FILLCELL_X1 FILLER_88_1107 ();
 FILLCELL_X8 FILLER_88_1120 ();
 FILLCELL_X2 FILLER_88_1151 ();
 FILLCELL_X4 FILLER_88_1178 ();
 FILLCELL_X2 FILLER_88_1182 ();
 FILLCELL_X2 FILLER_88_1206 ();
 FILLCELL_X4 FILLER_88_1213 ();
 FILLCELL_X2 FILLER_88_1239 ();
 FILLCELL_X1 FILLER_88_1246 ();
 FILLCELL_X8 FILLER_88_1249 ();
 FILLCELL_X2 FILLER_88_1257 ();
 FILLCELL_X1 FILLER_88_1259 ();
 FILLCELL_X16 FILLER_89_1 ();
 FILLCELL_X2 FILLER_89_17 ();
 FILLCELL_X2 FILLER_89_39 ();
 FILLCELL_X1 FILLER_89_41 ();
 FILLCELL_X4 FILLER_89_47 ();
 FILLCELL_X4 FILLER_89_58 ();
 FILLCELL_X8 FILLER_89_69 ();
 FILLCELL_X4 FILLER_89_77 ();
 FILLCELL_X1 FILLER_89_81 ();
 FILLCELL_X16 FILLER_89_89 ();
 FILLCELL_X8 FILLER_89_105 ();
 FILLCELL_X1 FILLER_89_113 ();
 FILLCELL_X2 FILLER_89_135 ();
 FILLCELL_X1 FILLER_89_137 ();
 FILLCELL_X8 FILLER_89_140 ();
 FILLCELL_X4 FILLER_89_148 ();
 FILLCELL_X2 FILLER_89_152 ();
 FILLCELL_X2 FILLER_89_168 ();
 FILLCELL_X2 FILLER_89_176 ();
 FILLCELL_X1 FILLER_89_178 ();
 FILLCELL_X4 FILLER_89_193 ();
 FILLCELL_X1 FILLER_89_197 ();
 FILLCELL_X2 FILLER_89_205 ();
 FILLCELL_X8 FILLER_89_214 ();
 FILLCELL_X1 FILLER_89_222 ();
 FILLCELL_X8 FILLER_89_237 ();
 FILLCELL_X1 FILLER_89_248 ();
 FILLCELL_X1 FILLER_89_272 ();
 FILLCELL_X2 FILLER_89_280 ();
 FILLCELL_X1 FILLER_89_282 ();
 FILLCELL_X8 FILLER_89_290 ();
 FILLCELL_X2 FILLER_89_298 ();
 FILLCELL_X1 FILLER_89_300 ();
 FILLCELL_X8 FILLER_89_308 ();
 FILLCELL_X4 FILLER_89_316 ();
 FILLCELL_X2 FILLER_89_363 ();
 FILLCELL_X1 FILLER_89_365 ();
 FILLCELL_X1 FILLER_89_382 ();
 FILLCELL_X1 FILLER_89_394 ();
 FILLCELL_X1 FILLER_89_421 ();
 FILLCELL_X1 FILLER_89_450 ();
 FILLCELL_X2 FILLER_89_455 ();
 FILLCELL_X1 FILLER_89_457 ();
 FILLCELL_X2 FILLER_89_465 ();
 FILLCELL_X1 FILLER_89_467 ();
 FILLCELL_X1 FILLER_89_492 ();
 FILLCELL_X1 FILLER_89_513 ();
 FILLCELL_X1 FILLER_89_537 ();
 FILLCELL_X2 FILLER_89_551 ();
 FILLCELL_X16 FILLER_89_562 ();
 FILLCELL_X2 FILLER_89_578 ();
 FILLCELL_X1 FILLER_89_580 ();
 FILLCELL_X1 FILLER_89_595 ();
 FILLCELL_X8 FILLER_89_646 ();
 FILLCELL_X4 FILLER_89_654 ();
 FILLCELL_X8 FILLER_89_668 ();
 FILLCELL_X4 FILLER_89_676 ();
 FILLCELL_X2 FILLER_89_694 ();
 FILLCELL_X4 FILLER_89_724 ();
 FILLCELL_X2 FILLER_89_728 ();
 FILLCELL_X1 FILLER_89_741 ();
 FILLCELL_X8 FILLER_89_751 ();
 FILLCELL_X4 FILLER_89_759 ();
 FILLCELL_X4 FILLER_89_777 ();
 FILLCELL_X2 FILLER_89_781 ();
 FILLCELL_X1 FILLER_89_783 ();
 FILLCELL_X8 FILLER_89_791 ();
 FILLCELL_X4 FILLER_89_806 ();
 FILLCELL_X2 FILLER_89_810 ();
 FILLCELL_X1 FILLER_89_812 ();
 FILLCELL_X2 FILLER_89_827 ();
 FILLCELL_X8 FILLER_89_842 ();
 FILLCELL_X4 FILLER_89_850 ();
 FILLCELL_X1 FILLER_89_854 ();
 FILLCELL_X4 FILLER_89_857 ();
 FILLCELL_X2 FILLER_89_861 ();
 FILLCELL_X4 FILLER_89_874 ();
 FILLCELL_X8 FILLER_89_915 ();
 FILLCELL_X4 FILLER_89_923 ();
 FILLCELL_X2 FILLER_89_927 ();
 FILLCELL_X1 FILLER_89_933 ();
 FILLCELL_X2 FILLER_89_940 ();
 FILLCELL_X2 FILLER_89_948 ();
 FILLCELL_X2 FILLER_89_957 ();
 FILLCELL_X1 FILLER_89_959 ();
 FILLCELL_X16 FILLER_89_974 ();
 FILLCELL_X8 FILLER_89_990 ();
 FILLCELL_X2 FILLER_89_998 ();
 FILLCELL_X1 FILLER_89_1000 ();
 FILLCELL_X8 FILLER_89_1012 ();
 FILLCELL_X4 FILLER_89_1020 ();
 FILLCELL_X2 FILLER_89_1028 ();
 FILLCELL_X1 FILLER_89_1030 ();
 FILLCELL_X1 FILLER_89_1035 ();
 FILLCELL_X1 FILLER_89_1083 ();
 FILLCELL_X2 FILLER_89_1104 ();
 FILLCELL_X4 FILLER_89_1123 ();
 FILLCELL_X1 FILLER_89_1138 ();
 FILLCELL_X1 FILLER_89_1141 ();
 FILLCELL_X2 FILLER_89_1153 ();
 FILLCELL_X1 FILLER_89_1155 ();
 FILLCELL_X2 FILLER_89_1170 ();
 FILLCELL_X2 FILLER_89_1197 ();
 FILLCELL_X1 FILLER_89_1221 ();
 FILLCELL_X2 FILLER_89_1238 ();
 FILLCELL_X8 FILLER_90_28 ();
 FILLCELL_X4 FILLER_90_36 ();
 FILLCELL_X2 FILLER_90_40 ();
 FILLCELL_X2 FILLER_90_83 ();
 FILLCELL_X4 FILLER_90_153 ();
 FILLCELL_X2 FILLER_90_157 ();
 FILLCELL_X2 FILLER_90_169 ();
 FILLCELL_X2 FILLER_90_182 ();
 FILLCELL_X1 FILLER_90_184 ();
 FILLCELL_X8 FILLER_90_188 ();
 FILLCELL_X1 FILLER_90_221 ();
 FILLCELL_X2 FILLER_90_252 ();
 FILLCELL_X2 FILLER_90_265 ();
 FILLCELL_X2 FILLER_90_278 ();
 FILLCELL_X1 FILLER_90_280 ();
 FILLCELL_X4 FILLER_90_286 ();
 FILLCELL_X1 FILLER_90_290 ();
 FILLCELL_X8 FILLER_90_315 ();
 FILLCELL_X4 FILLER_90_323 ();
 FILLCELL_X1 FILLER_90_327 ();
 FILLCELL_X2 FILLER_90_342 ();
 FILLCELL_X1 FILLER_90_392 ();
 FILLCELL_X1 FILLER_90_400 ();
 FILLCELL_X1 FILLER_90_428 ();
 FILLCELL_X2 FILLER_90_461 ();
 FILLCELL_X2 FILLER_90_470 ();
 FILLCELL_X2 FILLER_90_479 ();
 FILLCELL_X1 FILLER_90_481 ();
 FILLCELL_X2 FILLER_90_512 ();
 FILLCELL_X1 FILLER_90_527 ();
 FILLCELL_X1 FILLER_90_531 ();
 FILLCELL_X2 FILLER_90_535 ();
 FILLCELL_X32 FILLER_90_562 ();
 FILLCELL_X8 FILLER_90_594 ();
 FILLCELL_X2 FILLER_90_602 ();
 FILLCELL_X8 FILLER_90_613 ();
 FILLCELL_X1 FILLER_90_621 ();
 FILLCELL_X1 FILLER_90_630 ();
 FILLCELL_X2 FILLER_90_632 ();
 FILLCELL_X8 FILLER_90_647 ();
 FILLCELL_X4 FILLER_90_655 ();
 FILLCELL_X1 FILLER_90_659 ();
 FILLCELL_X4 FILLER_90_670 ();
 FILLCELL_X2 FILLER_90_674 ();
 FILLCELL_X1 FILLER_90_676 ();
 FILLCELL_X4 FILLER_90_684 ();
 FILLCELL_X16 FILLER_90_709 ();
 FILLCELL_X1 FILLER_90_725 ();
 FILLCELL_X1 FILLER_90_733 ();
 FILLCELL_X4 FILLER_90_741 ();
 FILLCELL_X2 FILLER_90_745 ();
 FILLCELL_X8 FILLER_90_763 ();
 FILLCELL_X4 FILLER_90_771 ();
 FILLCELL_X1 FILLER_90_775 ();
 FILLCELL_X8 FILLER_90_783 ();
 FILLCELL_X4 FILLER_90_791 ();
 FILLCELL_X2 FILLER_90_795 ();
 FILLCELL_X1 FILLER_90_797 ();
 FILLCELL_X8 FILLER_90_805 ();
 FILLCELL_X4 FILLER_90_827 ();
 FILLCELL_X2 FILLER_90_831 ();
 FILLCELL_X1 FILLER_90_844 ();
 FILLCELL_X8 FILLER_90_867 ();
 FILLCELL_X2 FILLER_90_875 ();
 FILLCELL_X2 FILLER_90_897 ();
 FILLCELL_X1 FILLER_90_899 ();
 FILLCELL_X4 FILLER_90_917 ();
 FILLCELL_X2 FILLER_90_921 ();
 FILLCELL_X4 FILLER_90_927 ();
 FILLCELL_X2 FILLER_90_931 ();
 FILLCELL_X1 FILLER_90_933 ();
 FILLCELL_X2 FILLER_90_952 ();
 FILLCELL_X1 FILLER_90_954 ();
 FILLCELL_X4 FILLER_90_977 ();
 FILLCELL_X2 FILLER_90_981 ();
 FILLCELL_X1 FILLER_90_993 ();
 FILLCELL_X1 FILLER_90_999 ();
 FILLCELL_X8 FILLER_90_1013 ();
 FILLCELL_X4 FILLER_90_1021 ();
 FILLCELL_X1 FILLER_90_1100 ();
 FILLCELL_X1 FILLER_90_1122 ();
 FILLCELL_X2 FILLER_90_1132 ();
 FILLCELL_X1 FILLER_90_1134 ();
 FILLCELL_X1 FILLER_90_1148 ();
 FILLCELL_X4 FILLER_90_1182 ();
 FILLCELL_X1 FILLER_90_1188 ();
 FILLCELL_X1 FILLER_90_1196 ();
 FILLCELL_X8 FILLER_90_1204 ();
 FILLCELL_X2 FILLER_90_1212 ();
 FILLCELL_X8 FILLER_90_1221 ();
 FILLCELL_X2 FILLER_90_1236 ();
 FILLCELL_X1 FILLER_90_1238 ();
 FILLCELL_X8 FILLER_90_1248 ();
 FILLCELL_X4 FILLER_90_1256 ();
 FILLCELL_X8 FILLER_91_1 ();
 FILLCELL_X4 FILLER_91_9 ();
 FILLCELL_X2 FILLER_91_13 ();
 FILLCELL_X16 FILLER_91_49 ();
 FILLCELL_X2 FILLER_91_65 ();
 FILLCELL_X1 FILLER_91_67 ();
 FILLCELL_X4 FILLER_91_82 ();
 FILLCELL_X2 FILLER_91_86 ();
 FILLCELL_X1 FILLER_91_88 ();
 FILLCELL_X8 FILLER_91_93 ();
 FILLCELL_X1 FILLER_91_101 ();
 FILLCELL_X8 FILLER_91_109 ();
 FILLCELL_X1 FILLER_91_117 ();
 FILLCELL_X2 FILLER_91_125 ();
 FILLCELL_X1 FILLER_91_134 ();
 FILLCELL_X1 FILLER_91_142 ();
 FILLCELL_X4 FILLER_91_164 ();
 FILLCELL_X4 FILLER_91_175 ();
 FILLCELL_X1 FILLER_91_179 ();
 FILLCELL_X2 FILLER_91_193 ();
 FILLCELL_X1 FILLER_91_195 ();
 FILLCELL_X1 FILLER_91_203 ();
 FILLCELL_X16 FILLER_91_225 ();
 FILLCELL_X4 FILLER_91_241 ();
 FILLCELL_X1 FILLER_91_245 ();
 FILLCELL_X2 FILLER_91_256 ();
 FILLCELL_X2 FILLER_91_265 ();
 FILLCELL_X1 FILLER_91_267 ();
 FILLCELL_X2 FILLER_91_275 ();
 FILLCELL_X1 FILLER_91_277 ();
 FILLCELL_X4 FILLER_91_296 ();
 FILLCELL_X1 FILLER_91_300 ();
 FILLCELL_X4 FILLER_91_308 ();
 FILLCELL_X1 FILLER_91_312 ();
 FILLCELL_X4 FILLER_91_324 ();
 FILLCELL_X2 FILLER_91_328 ();
 FILLCELL_X8 FILLER_91_332 ();
 FILLCELL_X4 FILLER_91_340 ();
 FILLCELL_X2 FILLER_91_351 ();
 FILLCELL_X4 FILLER_91_358 ();
 FILLCELL_X4 FILLER_91_369 ();
 FILLCELL_X2 FILLER_91_377 ();
 FILLCELL_X1 FILLER_91_379 ();
 FILLCELL_X1 FILLER_91_387 ();
 FILLCELL_X4 FILLER_91_399 ();
 FILLCELL_X1 FILLER_91_403 ();
 FILLCELL_X8 FILLER_91_408 ();
 FILLCELL_X4 FILLER_91_416 ();
 FILLCELL_X1 FILLER_91_479 ();
 FILLCELL_X1 FILLER_91_500 ();
 FILLCELL_X4 FILLER_91_538 ();
 FILLCELL_X2 FILLER_91_542 ();
 FILLCELL_X4 FILLER_91_553 ();
 FILLCELL_X2 FILLER_91_557 ();
 FILLCELL_X1 FILLER_91_559 ();
 FILLCELL_X1 FILLER_91_574 ();
 FILLCELL_X4 FILLER_91_589 ();
 FILLCELL_X1 FILLER_91_593 ();
 FILLCELL_X16 FILLER_91_636 ();
 FILLCELL_X4 FILLER_91_652 ();
 FILLCELL_X1 FILLER_91_656 ();
 FILLCELL_X4 FILLER_91_664 ();
 FILLCELL_X1 FILLER_91_668 ();
 FILLCELL_X1 FILLER_91_676 ();
 FILLCELL_X1 FILLER_91_684 ();
 FILLCELL_X2 FILLER_91_692 ();
 FILLCELL_X1 FILLER_91_694 ();
 FILLCELL_X8 FILLER_91_719 ();
 FILLCELL_X4 FILLER_91_727 ();
 FILLCELL_X2 FILLER_91_731 ();
 FILLCELL_X8 FILLER_91_747 ();
 FILLCELL_X4 FILLER_91_755 ();
 FILLCELL_X2 FILLER_91_759 ();
 FILLCELL_X1 FILLER_91_761 ();
 FILLCELL_X4 FILLER_91_769 ();
 FILLCELL_X2 FILLER_91_773 ();
 FILLCELL_X1 FILLER_91_775 ();
 FILLCELL_X16 FILLER_91_783 ();
 FILLCELL_X4 FILLER_91_806 ();
 FILLCELL_X2 FILLER_91_810 ();
 FILLCELL_X1 FILLER_91_812 ();
 FILLCELL_X2 FILLER_91_827 ();
 FILLCELL_X4 FILLER_91_845 ();
 FILLCELL_X2 FILLER_91_849 ();
 FILLCELL_X16 FILLER_91_869 ();
 FILLCELL_X1 FILLER_91_885 ();
 FILLCELL_X4 FILLER_91_896 ();
 FILLCELL_X2 FILLER_91_900 ();
 FILLCELL_X1 FILLER_91_902 ();
 FILLCELL_X2 FILLER_91_920 ();
 FILLCELL_X4 FILLER_91_926 ();
 FILLCELL_X2 FILLER_91_930 ();
 FILLCELL_X1 FILLER_91_932 ();
 FILLCELL_X1 FILLER_91_937 ();
 FILLCELL_X2 FILLER_91_958 ();
 FILLCELL_X2 FILLER_91_967 ();
 FILLCELL_X2 FILLER_91_974 ();
 FILLCELL_X4 FILLER_91_981 ();
 FILLCELL_X2 FILLER_91_990 ();
 FILLCELL_X1 FILLER_91_992 ();
 FILLCELL_X4 FILLER_91_1036 ();
 FILLCELL_X1 FILLER_91_1040 ();
 FILLCELL_X4 FILLER_91_1045 ();
 FILLCELL_X1 FILLER_91_1080 ();
 FILLCELL_X4 FILLER_91_1144 ();
 FILLCELL_X1 FILLER_91_1148 ();
 FILLCELL_X2 FILLER_91_1171 ();
 FILLCELL_X2 FILLER_91_1178 ();
 FILLCELL_X4 FILLER_91_1182 ();
 FILLCELL_X2 FILLER_91_1186 ();
 FILLCELL_X1 FILLER_91_1188 ();
 FILLCELL_X1 FILLER_91_1196 ();
 FILLCELL_X2 FILLER_91_1199 ();
 FILLCELL_X1 FILLER_91_1201 ();
 FILLCELL_X4 FILLER_91_1224 ();
 FILLCELL_X1 FILLER_91_1228 ();
 FILLCELL_X2 FILLER_91_1258 ();
 FILLCELL_X16 FILLER_92_1 ();
 FILLCELL_X4 FILLER_92_24 ();
 FILLCELL_X2 FILLER_92_28 ();
 FILLCELL_X1 FILLER_92_30 ();
 FILLCELL_X4 FILLER_92_52 ();
 FILLCELL_X2 FILLER_92_56 ();
 FILLCELL_X1 FILLER_92_65 ();
 FILLCELL_X1 FILLER_92_73 ();
 FILLCELL_X1 FILLER_92_81 ();
 FILLCELL_X8 FILLER_92_89 ();
 FILLCELL_X4 FILLER_92_97 ();
 FILLCELL_X2 FILLER_92_101 ();
 FILLCELL_X1 FILLER_92_103 ();
 FILLCELL_X4 FILLER_92_115 ();
 FILLCELL_X2 FILLER_92_119 ();
 FILLCELL_X1 FILLER_92_121 ();
 FILLCELL_X32 FILLER_92_149 ();
 FILLCELL_X2 FILLER_92_181 ();
 FILLCELL_X1 FILLER_92_183 ();
 FILLCELL_X2 FILLER_92_204 ();
 FILLCELL_X4 FILLER_92_213 ();
 FILLCELL_X8 FILLER_92_238 ();
 FILLCELL_X2 FILLER_92_246 ();
 FILLCELL_X8 FILLER_92_255 ();
 FILLCELL_X2 FILLER_92_263 ();
 FILLCELL_X2 FILLER_92_268 ();
 FILLCELL_X4 FILLER_92_284 ();
 FILLCELL_X2 FILLER_92_295 ();
 FILLCELL_X1 FILLER_92_300 ();
 FILLCELL_X1 FILLER_92_311 ();
 FILLCELL_X4 FILLER_92_319 ();
 FILLCELL_X1 FILLER_92_323 ();
 FILLCELL_X2 FILLER_92_327 ();
 FILLCELL_X1 FILLER_92_329 ();
 FILLCELL_X8 FILLER_92_344 ();
 FILLCELL_X1 FILLER_92_393 ();
 FILLCELL_X2 FILLER_92_397 ();
 FILLCELL_X4 FILLER_92_406 ();
 FILLCELL_X2 FILLER_92_410 ();
 FILLCELL_X1 FILLER_92_416 ();
 FILLCELL_X1 FILLER_92_442 ();
 FILLCELL_X2 FILLER_92_456 ();
 FILLCELL_X2 FILLER_92_478 ();
 FILLCELL_X1 FILLER_92_540 ();
 FILLCELL_X4 FILLER_92_548 ();
 FILLCELL_X4 FILLER_92_575 ();
 FILLCELL_X32 FILLER_92_584 ();
 FILLCELL_X2 FILLER_92_628 ();
 FILLCELL_X1 FILLER_92_630 ();
 FILLCELL_X16 FILLER_92_642 ();
 FILLCELL_X4 FILLER_92_658 ();
 FILLCELL_X4 FILLER_92_667 ();
 FILLCELL_X1 FILLER_92_671 ();
 FILLCELL_X2 FILLER_92_676 ();
 FILLCELL_X4 FILLER_92_695 ();
 FILLCELL_X1 FILLER_92_706 ();
 FILLCELL_X4 FILLER_92_735 ();
 FILLCELL_X2 FILLER_92_739 ();
 FILLCELL_X2 FILLER_92_770 ();
 FILLCELL_X1 FILLER_92_784 ();
 FILLCELL_X1 FILLER_92_792 ();
 FILLCELL_X2 FILLER_92_806 ();
 FILLCELL_X4 FILLER_92_812 ();
 FILLCELL_X2 FILLER_92_816 ();
 FILLCELL_X4 FILLER_92_825 ();
 FILLCELL_X2 FILLER_92_835 ();
 FILLCELL_X16 FILLER_92_843 ();
 FILLCELL_X8 FILLER_92_859 ();
 FILLCELL_X8 FILLER_92_872 ();
 FILLCELL_X4 FILLER_92_880 ();
 FILLCELL_X2 FILLER_92_888 ();
 FILLCELL_X1 FILLER_92_890 ();
 FILLCELL_X1 FILLER_92_896 ();
 FILLCELL_X1 FILLER_92_924 ();
 FILLCELL_X8 FILLER_92_934 ();
 FILLCELL_X8 FILLER_92_949 ();
 FILLCELL_X1 FILLER_92_957 ();
 FILLCELL_X32 FILLER_92_971 ();
 FILLCELL_X8 FILLER_92_1003 ();
 FILLCELL_X4 FILLER_92_1011 ();
 FILLCELL_X2 FILLER_92_1015 ();
 FILLCELL_X1 FILLER_92_1017 ();
 FILLCELL_X2 FILLER_92_1022 ();
 FILLCELL_X1 FILLER_92_1034 ();
 FILLCELL_X1 FILLER_92_1045 ();
 FILLCELL_X1 FILLER_92_1053 ();
 FILLCELL_X1 FILLER_92_1071 ();
 FILLCELL_X8 FILLER_92_1077 ();
 FILLCELL_X4 FILLER_92_1085 ();
 FILLCELL_X1 FILLER_92_1089 ();
 FILLCELL_X2 FILLER_92_1116 ();
 FILLCELL_X2 FILLER_92_1131 ();
 FILLCELL_X2 FILLER_92_1140 ();
 FILLCELL_X1 FILLER_92_1155 ();
 FILLCELL_X2 FILLER_92_1164 ();
 FILLCELL_X4 FILLER_92_1247 ();
 FILLCELL_X1 FILLER_92_1251 ();
 FILLCELL_X4 FILLER_92_1254 ();
 FILLCELL_X2 FILLER_92_1258 ();
 FILLCELL_X8 FILLER_93_1 ();
 FILLCELL_X2 FILLER_93_9 ();
 FILLCELL_X1 FILLER_93_11 ();
 FILLCELL_X4 FILLER_93_19 ();
 FILLCELL_X1 FILLER_93_23 ();
 FILLCELL_X2 FILLER_93_31 ();
 FILLCELL_X2 FILLER_93_40 ();
 FILLCELL_X1 FILLER_93_42 ();
 FILLCELL_X1 FILLER_93_90 ();
 FILLCELL_X1 FILLER_93_95 ();
 FILLCELL_X8 FILLER_93_136 ();
 FILLCELL_X1 FILLER_93_144 ();
 FILLCELL_X8 FILLER_93_152 ();
 FILLCELL_X4 FILLER_93_160 ();
 FILLCELL_X2 FILLER_93_164 ();
 FILLCELL_X1 FILLER_93_166 ();
 FILLCELL_X4 FILLER_93_187 ();
 FILLCELL_X8 FILLER_93_226 ();
 FILLCELL_X4 FILLER_93_234 ();
 FILLCELL_X4 FILLER_93_245 ();
 FILLCELL_X2 FILLER_93_249 ();
 FILLCELL_X1 FILLER_93_258 ();
 FILLCELL_X8 FILLER_93_276 ();
 FILLCELL_X2 FILLER_93_305 ();
 FILLCELL_X4 FILLER_93_314 ();
 FILLCELL_X1 FILLER_93_318 ();
 FILLCELL_X16 FILLER_93_339 ();
 FILLCELL_X4 FILLER_93_355 ();
 FILLCELL_X1 FILLER_93_395 ();
 FILLCELL_X2 FILLER_93_454 ();
 FILLCELL_X1 FILLER_93_501 ();
 FILLCELL_X16 FILLER_93_543 ();
 FILLCELL_X8 FILLER_93_559 ();
 FILLCELL_X4 FILLER_93_567 ();
 FILLCELL_X1 FILLER_93_571 ();
 FILLCELL_X16 FILLER_93_586 ();
 FILLCELL_X1 FILLER_93_626 ();
 FILLCELL_X8 FILLER_93_650 ();
 FILLCELL_X4 FILLER_93_658 ();
 FILLCELL_X2 FILLER_93_662 ();
 FILLCELL_X4 FILLER_93_668 ();
 FILLCELL_X4 FILLER_93_676 ();
 FILLCELL_X2 FILLER_93_680 ();
 FILLCELL_X1 FILLER_93_682 ();
 FILLCELL_X2 FILLER_93_690 ();
 FILLCELL_X8 FILLER_93_702 ();
 FILLCELL_X1 FILLER_93_710 ();
 FILLCELL_X8 FILLER_93_717 ();
 FILLCELL_X1 FILLER_93_725 ();
 FILLCELL_X2 FILLER_93_737 ();
 FILLCELL_X1 FILLER_93_739 ();
 FILLCELL_X16 FILLER_93_747 ();
 FILLCELL_X8 FILLER_93_763 ();
 FILLCELL_X4 FILLER_93_771 ();
 FILLCELL_X2 FILLER_93_775 ();
 FILLCELL_X8 FILLER_93_791 ();
 FILLCELL_X2 FILLER_93_799 ();
 FILLCELL_X4 FILLER_93_808 ();
 FILLCELL_X1 FILLER_93_812 ();
 FILLCELL_X16 FILLER_93_816 ();
 FILLCELL_X1 FILLER_93_842 ();
 FILLCELL_X16 FILLER_93_847 ();
 FILLCELL_X2 FILLER_93_863 ();
 FILLCELL_X2 FILLER_93_874 ();
 FILLCELL_X4 FILLER_93_886 ();
 FILLCELL_X2 FILLER_93_890 ();
 FILLCELL_X2 FILLER_93_903 ();
 FILLCELL_X1 FILLER_93_905 ();
 FILLCELL_X1 FILLER_93_916 ();
 FILLCELL_X2 FILLER_93_921 ();
 FILLCELL_X1 FILLER_93_923 ();
 FILLCELL_X1 FILLER_93_949 ();
 FILLCELL_X4 FILLER_93_963 ();
 FILLCELL_X1 FILLER_93_967 ();
 FILLCELL_X2 FILLER_93_974 ();
 FILLCELL_X1 FILLER_93_976 ();
 FILLCELL_X4 FILLER_93_989 ();
 FILLCELL_X4 FILLER_93_998 ();
 FILLCELL_X4 FILLER_93_1017 ();
 FILLCELL_X2 FILLER_93_1021 ();
 FILLCELL_X8 FILLER_93_1035 ();
 FILLCELL_X4 FILLER_93_1043 ();
 FILLCELL_X2 FILLER_93_1047 ();
 FILLCELL_X2 FILLER_93_1053 ();
 FILLCELL_X2 FILLER_93_1059 ();
 FILLCELL_X1 FILLER_93_1061 ();
 FILLCELL_X2 FILLER_93_1078 ();
 FILLCELL_X1 FILLER_93_1080 ();
 FILLCELL_X4 FILLER_93_1091 ();
 FILLCELL_X2 FILLER_93_1095 ();
 FILLCELL_X2 FILLER_93_1149 ();
 FILLCELL_X8 FILLER_93_1161 ();
 FILLCELL_X4 FILLER_93_1169 ();
 FILLCELL_X4 FILLER_93_1178 ();
 FILLCELL_X2 FILLER_93_1184 ();
 FILLCELL_X4 FILLER_93_1188 ();
 FILLCELL_X1 FILLER_93_1192 ();
 FILLCELL_X16 FILLER_93_1200 ();
 FILLCELL_X2 FILLER_93_1216 ();
 FILLCELL_X1 FILLER_93_1218 ();
 FILLCELL_X8 FILLER_93_1221 ();
 FILLCELL_X2 FILLER_93_1229 ();
 FILLCELL_X2 FILLER_93_1238 ();
 FILLCELL_X8 FILLER_93_1247 ();
 FILLCELL_X4 FILLER_93_1255 ();
 FILLCELL_X1 FILLER_93_1259 ();
 FILLCELL_X2 FILLER_94_1 ();
 FILLCELL_X1 FILLER_94_3 ();
 FILLCELL_X16 FILLER_94_51 ();
 FILLCELL_X1 FILLER_94_67 ();
 FILLCELL_X4 FILLER_94_75 ();
 FILLCELL_X2 FILLER_94_79 ();
 FILLCELL_X1 FILLER_94_81 ();
 FILLCELL_X8 FILLER_94_89 ();
 FILLCELL_X1 FILLER_94_97 ();
 FILLCELL_X2 FILLER_94_112 ();
 FILLCELL_X1 FILLER_94_114 ();
 FILLCELL_X16 FILLER_94_122 ();
 FILLCELL_X8 FILLER_94_138 ();
 FILLCELL_X1 FILLER_94_146 ();
 FILLCELL_X8 FILLER_94_168 ();
 FILLCELL_X2 FILLER_94_210 ();
 FILLCELL_X1 FILLER_94_212 ();
 FILLCELL_X8 FILLER_94_234 ();
 FILLCELL_X4 FILLER_94_242 ();
 FILLCELL_X1 FILLER_94_246 ();
 FILLCELL_X1 FILLER_94_261 ();
 FILLCELL_X8 FILLER_94_296 ();
 FILLCELL_X4 FILLER_94_304 ();
 FILLCELL_X2 FILLER_94_308 ();
 FILLCELL_X4 FILLER_94_314 ();
 FILLCELL_X1 FILLER_94_318 ();
 FILLCELL_X2 FILLER_94_322 ();
 FILLCELL_X2 FILLER_94_338 ();
 FILLCELL_X2 FILLER_94_354 ();
 FILLCELL_X1 FILLER_94_356 ();
 FILLCELL_X4 FILLER_94_364 ();
 FILLCELL_X2 FILLER_94_368 ();
 FILLCELL_X1 FILLER_94_404 ();
 FILLCELL_X1 FILLER_94_527 ();
 FILLCELL_X2 FILLER_94_532 ();
 FILLCELL_X1 FILLER_94_534 ();
 FILLCELL_X4 FILLER_94_557 ();
 FILLCELL_X4 FILLER_94_589 ();
 FILLCELL_X1 FILLER_94_614 ();
 FILLCELL_X2 FILLER_94_628 ();
 FILLCELL_X1 FILLER_94_630 ();
 FILLCELL_X4 FILLER_94_632 ();
 FILLCELL_X16 FILLER_94_643 ();
 FILLCELL_X4 FILLER_94_659 ();
 FILLCELL_X1 FILLER_94_663 ();
 FILLCELL_X2 FILLER_94_669 ();
 FILLCELL_X1 FILLER_94_683 ();
 FILLCELL_X1 FILLER_94_721 ();
 FILLCELL_X4 FILLER_94_726 ();
 FILLCELL_X1 FILLER_94_730 ();
 FILLCELL_X4 FILLER_94_738 ();
 FILLCELL_X2 FILLER_94_742 ();
 FILLCELL_X8 FILLER_94_758 ();
 FILLCELL_X1 FILLER_94_766 ();
 FILLCELL_X8 FILLER_94_774 ();
 FILLCELL_X4 FILLER_94_782 ();
 FILLCELL_X1 FILLER_94_786 ();
 FILLCELL_X4 FILLER_94_794 ();
 FILLCELL_X2 FILLER_94_798 ();
 FILLCELL_X1 FILLER_94_800 ();
 FILLCELL_X4 FILLER_94_828 ();
 FILLCELL_X4 FILLER_94_840 ();
 FILLCELL_X2 FILLER_94_844 ();
 FILLCELL_X1 FILLER_94_850 ();
 FILLCELL_X1 FILLER_94_890 ();
 FILLCELL_X1 FILLER_94_903 ();
 FILLCELL_X2 FILLER_94_910 ();
 FILLCELL_X4 FILLER_94_922 ();
 FILLCELL_X1 FILLER_94_926 ();
 FILLCELL_X4 FILLER_94_941 ();
 FILLCELL_X2 FILLER_94_945 ();
 FILLCELL_X1 FILLER_94_947 ();
 FILLCELL_X8 FILLER_94_950 ();
 FILLCELL_X2 FILLER_94_958 ();
 FILLCELL_X1 FILLER_94_960 ();
 FILLCELL_X16 FILLER_94_968 ();
 FILLCELL_X1 FILLER_94_984 ();
 FILLCELL_X1 FILLER_94_990 ();
 FILLCELL_X4 FILLER_94_996 ();
 FILLCELL_X2 FILLER_94_1000 ();
 FILLCELL_X1 FILLER_94_1002 ();
 FILLCELL_X2 FILLER_94_1008 ();
 FILLCELL_X1 FILLER_94_1010 ();
 FILLCELL_X16 FILLER_94_1016 ();
 FILLCELL_X4 FILLER_94_1032 ();
 FILLCELL_X2 FILLER_94_1036 ();
 FILLCELL_X1 FILLER_94_1041 ();
 FILLCELL_X4 FILLER_94_1063 ();
 FILLCELL_X8 FILLER_94_1077 ();
 FILLCELL_X4 FILLER_94_1085 ();
 FILLCELL_X1 FILLER_94_1089 ();
 FILLCELL_X4 FILLER_94_1101 ();
 FILLCELL_X2 FILLER_94_1105 ();
 FILLCELL_X1 FILLER_94_1107 ();
 FILLCELL_X1 FILLER_94_1121 ();
 FILLCELL_X2 FILLER_94_1145 ();
 FILLCELL_X8 FILLER_94_1150 ();
 FILLCELL_X4 FILLER_94_1158 ();
 FILLCELL_X2 FILLER_94_1162 ();
 FILLCELL_X1 FILLER_94_1164 ();
 FILLCELL_X2 FILLER_94_1185 ();
 FILLCELL_X2 FILLER_94_1194 ();
 FILLCELL_X1 FILLER_94_1259 ();
 FILLCELL_X16 FILLER_95_1 ();
 FILLCELL_X2 FILLER_95_17 ();
 FILLCELL_X1 FILLER_95_19 ();
 FILLCELL_X2 FILLER_95_40 ();
 FILLCELL_X16 FILLER_95_47 ();
 FILLCELL_X2 FILLER_95_63 ();
 FILLCELL_X4 FILLER_95_92 ();
 FILLCELL_X4 FILLER_95_143 ();
 FILLCELL_X1 FILLER_95_147 ();
 FILLCELL_X8 FILLER_95_168 ();
 FILLCELL_X1 FILLER_95_176 ();
 FILLCELL_X4 FILLER_95_184 ();
 FILLCELL_X2 FILLER_95_188 ();
 FILLCELL_X1 FILLER_95_190 ();
 FILLCELL_X4 FILLER_95_198 ();
 FILLCELL_X2 FILLER_95_229 ();
 FILLCELL_X1 FILLER_95_231 ();
 FILLCELL_X8 FILLER_95_299 ();
 FILLCELL_X2 FILLER_95_307 ();
 FILLCELL_X1 FILLER_95_329 ();
 FILLCELL_X2 FILLER_95_337 ();
 FILLCELL_X1 FILLER_95_339 ();
 FILLCELL_X1 FILLER_95_385 ();
 FILLCELL_X1 FILLER_95_425 ();
 FILLCELL_X4 FILLER_95_540 ();
 FILLCELL_X2 FILLER_95_553 ();
 FILLCELL_X16 FILLER_95_573 ();
 FILLCELL_X8 FILLER_95_589 ();
 FILLCELL_X1 FILLER_95_602 ();
 FILLCELL_X8 FILLER_95_650 ();
 FILLCELL_X2 FILLER_95_658 ();
 FILLCELL_X1 FILLER_95_660 ();
 FILLCELL_X4 FILLER_95_682 ();
 FILLCELL_X2 FILLER_95_686 ();
 FILLCELL_X1 FILLER_95_691 ();
 FILLCELL_X1 FILLER_95_705 ();
 FILLCELL_X2 FILLER_95_709 ();
 FILLCELL_X4 FILLER_95_715 ();
 FILLCELL_X2 FILLER_95_719 ();
 FILLCELL_X1 FILLER_95_721 ();
 FILLCELL_X4 FILLER_95_729 ();
 FILLCELL_X1 FILLER_95_733 ();
 FILLCELL_X1 FILLER_95_741 ();
 FILLCELL_X8 FILLER_95_746 ();
 FILLCELL_X2 FILLER_95_754 ();
 FILLCELL_X4 FILLER_95_758 ();
 FILLCELL_X1 FILLER_95_762 ();
 FILLCELL_X8 FILLER_95_777 ();
 FILLCELL_X2 FILLER_95_785 ();
 FILLCELL_X4 FILLER_95_791 ();
 FILLCELL_X2 FILLER_95_815 ();
 FILLCELL_X1 FILLER_95_817 ();
 FILLCELL_X2 FILLER_95_822 ();
 FILLCELL_X1 FILLER_95_824 ();
 FILLCELL_X4 FILLER_95_828 ();
 FILLCELL_X2 FILLER_95_855 ();
 FILLCELL_X2 FILLER_95_885 ();
 FILLCELL_X1 FILLER_95_887 ();
 FILLCELL_X1 FILLER_95_892 ();
 FILLCELL_X1 FILLER_95_896 ();
 FILLCELL_X2 FILLER_95_921 ();
 FILLCELL_X2 FILLER_95_925 ();
 FILLCELL_X4 FILLER_95_935 ();
 FILLCELL_X2 FILLER_95_939 ();
 FILLCELL_X8 FILLER_95_970 ();
 FILLCELL_X4 FILLER_95_978 ();
 FILLCELL_X2 FILLER_95_987 ();
 FILLCELL_X2 FILLER_95_996 ();
 FILLCELL_X1 FILLER_95_998 ();
 FILLCELL_X1 FILLER_95_1008 ();
 FILLCELL_X1 FILLER_95_1013 ();
 FILLCELL_X2 FILLER_95_1039 ();
 FILLCELL_X4 FILLER_95_1046 ();
 FILLCELL_X2 FILLER_95_1050 ();
 FILLCELL_X4 FILLER_95_1057 ();
 FILLCELL_X1 FILLER_95_1061 ();
 FILLCELL_X4 FILLER_95_1066 ();
 FILLCELL_X2 FILLER_95_1070 ();
 FILLCELL_X8 FILLER_95_1077 ();
 FILLCELL_X8 FILLER_95_1095 ();
 FILLCELL_X4 FILLER_95_1103 ();
 FILLCELL_X1 FILLER_95_1107 ();
 FILLCELL_X4 FILLER_95_1113 ();
 FILLCELL_X2 FILLER_95_1121 ();
 FILLCELL_X4 FILLER_95_1143 ();
 FILLCELL_X8 FILLER_95_1167 ();
 FILLCELL_X4 FILLER_95_1192 ();
 FILLCELL_X8 FILLER_95_1205 ();
 FILLCELL_X4 FILLER_95_1213 ();
 FILLCELL_X1 FILLER_95_1236 ();
 FILLCELL_X1 FILLER_95_1244 ();
 FILLCELL_X2 FILLER_95_1252 ();
 FILLCELL_X16 FILLER_96_1 ();
 FILLCELL_X4 FILLER_96_17 ();
 FILLCELL_X2 FILLER_96_28 ();
 FILLCELL_X1 FILLER_96_52 ();
 FILLCELL_X2 FILLER_96_73 ();
 FILLCELL_X1 FILLER_96_75 ();
 FILLCELL_X4 FILLER_96_83 ();
 FILLCELL_X1 FILLER_96_87 ();
 FILLCELL_X2 FILLER_96_95 ();
 FILLCELL_X1 FILLER_96_97 ();
 FILLCELL_X4 FILLER_96_118 ();
 FILLCELL_X2 FILLER_96_122 ();
 FILLCELL_X4 FILLER_96_131 ();
 FILLCELL_X1 FILLER_96_169 ();
 FILLCELL_X2 FILLER_96_190 ();
 FILLCELL_X2 FILLER_96_196 ();
 FILLCELL_X1 FILLER_96_198 ();
 FILLCELL_X16 FILLER_96_219 ();
 FILLCELL_X4 FILLER_96_235 ();
 FILLCELL_X2 FILLER_96_239 ();
 FILLCELL_X1 FILLER_96_241 ();
 FILLCELL_X16 FILLER_96_249 ();
 FILLCELL_X1 FILLER_96_265 ();
 FILLCELL_X2 FILLER_96_273 ();
 FILLCELL_X1 FILLER_96_306 ();
 FILLCELL_X8 FILLER_96_341 ();
 FILLCELL_X4 FILLER_96_349 ();
 FILLCELL_X1 FILLER_96_353 ();
 FILLCELL_X2 FILLER_96_363 ();
 FILLCELL_X1 FILLER_96_404 ();
 FILLCELL_X1 FILLER_96_436 ();
 FILLCELL_X1 FILLER_96_524 ();
 FILLCELL_X2 FILLER_96_534 ();
 FILLCELL_X4 FILLER_96_546 ();
 FILLCELL_X1 FILLER_96_550 ();
 FILLCELL_X4 FILLER_96_560 ();
 FILLCELL_X8 FILLER_96_573 ();
 FILLCELL_X1 FILLER_96_619 ();
 FILLCELL_X1 FILLER_96_630 ();
 FILLCELL_X4 FILLER_96_632 ();
 FILLCELL_X1 FILLER_96_639 ();
 FILLCELL_X8 FILLER_96_653 ();
 FILLCELL_X2 FILLER_96_661 ();
 FILLCELL_X1 FILLER_96_663 ();
 FILLCELL_X2 FILLER_96_671 ();
 FILLCELL_X2 FILLER_96_680 ();
 FILLCELL_X1 FILLER_96_682 ();
 FILLCELL_X4 FILLER_96_690 ();
 FILLCELL_X1 FILLER_96_694 ();
 FILLCELL_X2 FILLER_96_716 ();
 FILLCELL_X1 FILLER_96_718 ();
 FILLCELL_X16 FILLER_96_733 ();
 FILLCELL_X4 FILLER_96_749 ();
 FILLCELL_X1 FILLER_96_753 ();
 FILLCELL_X1 FILLER_96_761 ();
 FILLCELL_X1 FILLER_96_765 ();
 FILLCELL_X4 FILLER_96_787 ();
 FILLCELL_X1 FILLER_96_791 ();
 FILLCELL_X1 FILLER_96_795 ();
 FILLCELL_X4 FILLER_96_807 ();
 FILLCELL_X4 FILLER_96_822 ();
 FILLCELL_X2 FILLER_96_826 ();
 FILLCELL_X4 FILLER_96_846 ();
 FILLCELL_X4 FILLER_96_866 ();
 FILLCELL_X1 FILLER_96_870 ();
 FILLCELL_X2 FILLER_96_888 ();
 FILLCELL_X1 FILLER_96_890 ();
 FILLCELL_X16 FILLER_96_904 ();
 FILLCELL_X8 FILLER_96_920 ();
 FILLCELL_X2 FILLER_96_941 ();
 FILLCELL_X16 FILLER_96_950 ();
 FILLCELL_X8 FILLER_96_966 ();
 FILLCELL_X4 FILLER_96_974 ();
 FILLCELL_X1 FILLER_96_992 ();
 FILLCELL_X1 FILLER_96_1006 ();
 FILLCELL_X2 FILLER_96_1020 ();
 FILLCELL_X1 FILLER_96_1022 ();
 FILLCELL_X1 FILLER_96_1032 ();
 FILLCELL_X2 FILLER_96_1038 ();
 FILLCELL_X1 FILLER_96_1040 ();
 FILLCELL_X2 FILLER_96_1046 ();
 FILLCELL_X1 FILLER_96_1063 ();
 FILLCELL_X8 FILLER_96_1069 ();
 FILLCELL_X4 FILLER_96_1077 ();
 FILLCELL_X4 FILLER_96_1099 ();
 FILLCELL_X2 FILLER_96_1103 ();
 FILLCELL_X1 FILLER_96_1105 ();
 FILLCELL_X2 FILLER_96_1135 ();
 FILLCELL_X1 FILLER_96_1137 ();
 FILLCELL_X2 FILLER_96_1142 ();
 FILLCELL_X8 FILLER_96_1151 ();
 FILLCELL_X4 FILLER_96_1159 ();
 FILLCELL_X1 FILLER_96_1176 ();
 FILLCELL_X2 FILLER_96_1207 ();
 FILLCELL_X1 FILLER_96_1209 ();
 FILLCELL_X2 FILLER_96_1237 ();
 FILLCELL_X1 FILLER_96_1239 ();
 FILLCELL_X8 FILLER_97_1 ();
 FILLCELL_X2 FILLER_97_9 ();
 FILLCELL_X4 FILLER_97_38 ();
 FILLCELL_X2 FILLER_97_42 ();
 FILLCELL_X8 FILLER_97_98 ();
 FILLCELL_X1 FILLER_97_106 ();
 FILLCELL_X4 FILLER_97_116 ();
 FILLCELL_X1 FILLER_97_120 ();
 FILLCELL_X1 FILLER_97_128 ();
 FILLCELL_X2 FILLER_97_136 ();
 FILLCELL_X1 FILLER_97_138 ();
 FILLCELL_X8 FILLER_97_155 ();
 FILLCELL_X2 FILLER_97_163 ();
 FILLCELL_X1 FILLER_97_165 ();
 FILLCELL_X4 FILLER_97_173 ();
 FILLCELL_X1 FILLER_97_197 ();
 FILLCELL_X2 FILLER_97_201 ();
 FILLCELL_X1 FILLER_97_210 ();
 FILLCELL_X2 FILLER_97_220 ();
 FILLCELL_X2 FILLER_97_269 ();
 FILLCELL_X8 FILLER_97_296 ();
 FILLCELL_X2 FILLER_97_304 ();
 FILLCELL_X1 FILLER_97_306 ();
 FILLCELL_X2 FILLER_97_319 ();
 FILLCELL_X8 FILLER_97_341 ();
 FILLCELL_X4 FILLER_97_349 ();
 FILLCELL_X2 FILLER_97_362 ();
 FILLCELL_X1 FILLER_97_364 ();
 FILLCELL_X2 FILLER_97_385 ();
 FILLCELL_X4 FILLER_97_413 ();
 FILLCELL_X1 FILLER_97_417 ();
 FILLCELL_X1 FILLER_97_532 ();
 FILLCELL_X1 FILLER_97_542 ();
 FILLCELL_X16 FILLER_97_574 ();
 FILLCELL_X8 FILLER_97_590 ();
 FILLCELL_X4 FILLER_97_598 ();
 FILLCELL_X2 FILLER_97_602 ();
 FILLCELL_X1 FILLER_97_604 ();
 FILLCELL_X2 FILLER_97_610 ();
 FILLCELL_X1 FILLER_97_612 ();
 FILLCELL_X8 FILLER_97_650 ();
 FILLCELL_X2 FILLER_97_658 ();
 FILLCELL_X1 FILLER_97_667 ();
 FILLCELL_X2 FILLER_97_675 ();
 FILLCELL_X2 FILLER_97_684 ();
 FILLCELL_X1 FILLER_97_686 ();
 FILLCELL_X8 FILLER_97_694 ();
 FILLCELL_X4 FILLER_97_702 ();
 FILLCELL_X2 FILLER_97_706 ();
 FILLCELL_X1 FILLER_97_708 ();
 FILLCELL_X2 FILLER_97_721 ();
 FILLCELL_X4 FILLER_97_730 ();
 FILLCELL_X2 FILLER_97_734 ();
 FILLCELL_X4 FILLER_97_747 ();
 FILLCELL_X1 FILLER_97_751 ();
 FILLCELL_X4 FILLER_97_757 ();
 FILLCELL_X1 FILLER_97_761 ();
 FILLCELL_X16 FILLER_97_766 ();
 FILLCELL_X2 FILLER_97_782 ();
 FILLCELL_X1 FILLER_97_784 ();
 FILLCELL_X2 FILLER_97_805 ();
 FILLCELL_X8 FILLER_97_810 ();
 FILLCELL_X1 FILLER_97_818 ();
 FILLCELL_X1 FILLER_97_826 ();
 FILLCELL_X2 FILLER_97_836 ();
 FILLCELL_X1 FILLER_97_838 ();
 FILLCELL_X2 FILLER_97_844 ();
 FILLCELL_X4 FILLER_97_850 ();
 FILLCELL_X2 FILLER_97_854 ();
 FILLCELL_X1 FILLER_97_861 ();
 FILLCELL_X1 FILLER_97_872 ();
 FILLCELL_X1 FILLER_97_877 ();
 FILLCELL_X1 FILLER_97_884 ();
 FILLCELL_X4 FILLER_97_899 ();
 FILLCELL_X1 FILLER_97_903 ();
 FILLCELL_X1 FILLER_97_908 ();
 FILLCELL_X1 FILLER_97_921 ();
 FILLCELL_X8 FILLER_97_926 ();
 FILLCELL_X2 FILLER_97_934 ();
 FILLCELL_X1 FILLER_97_936 ();
 FILLCELL_X2 FILLER_97_943 ();
 FILLCELL_X2 FILLER_97_952 ();
 FILLCELL_X1 FILLER_97_954 ();
 FILLCELL_X2 FILLER_97_967 ();
 FILLCELL_X16 FILLER_97_974 ();
 FILLCELL_X16 FILLER_97_997 ();
 FILLCELL_X2 FILLER_97_1013 ();
 FILLCELL_X2 FILLER_97_1019 ();
 FILLCELL_X4 FILLER_97_1051 ();
 FILLCELL_X4 FILLER_97_1062 ();
 FILLCELL_X1 FILLER_97_1066 ();
 FILLCELL_X1 FILLER_97_1069 ();
 FILLCELL_X4 FILLER_97_1077 ();
 FILLCELL_X4 FILLER_97_1102 ();
 FILLCELL_X2 FILLER_97_1120 ();
 FILLCELL_X16 FILLER_97_1138 ();
 FILLCELL_X2 FILLER_97_1154 ();
 FILLCELL_X8 FILLER_97_1203 ();
 FILLCELL_X4 FILLER_97_1211 ();
 FILLCELL_X1 FILLER_97_1215 ();
 FILLCELL_X4 FILLER_97_1248 ();
 FILLCELL_X1 FILLER_97_1252 ();
 FILLCELL_X4 FILLER_97_1255 ();
 FILLCELL_X1 FILLER_97_1259 ();
 FILLCELL_X2 FILLER_98_28 ();
 FILLCELL_X1 FILLER_98_30 ();
 FILLCELL_X1 FILLER_98_38 ();
 FILLCELL_X16 FILLER_98_46 ();
 FILLCELL_X4 FILLER_98_62 ();
 FILLCELL_X1 FILLER_98_66 ();
 FILLCELL_X2 FILLER_98_83 ();
 FILLCELL_X1 FILLER_98_85 ();
 FILLCELL_X4 FILLER_98_93 ();
 FILLCELL_X2 FILLER_98_97 ();
 FILLCELL_X2 FILLER_98_120 ();
 FILLCELL_X1 FILLER_98_122 ();
 FILLCELL_X16 FILLER_98_137 ();
 FILLCELL_X8 FILLER_98_153 ();
 FILLCELL_X4 FILLER_98_161 ();
 FILLCELL_X4 FILLER_98_186 ();
 FILLCELL_X1 FILLER_98_194 ();
 FILLCELL_X2 FILLER_98_202 ();
 FILLCELL_X1 FILLER_98_204 ();
 FILLCELL_X8 FILLER_98_235 ();
 FILLCELL_X2 FILLER_98_243 ();
 FILLCELL_X2 FILLER_98_252 ();
 FILLCELL_X1 FILLER_98_254 ();
 FILLCELL_X4 FILLER_98_302 ();
 FILLCELL_X2 FILLER_98_306 ();
 FILLCELL_X1 FILLER_98_315 ();
 FILLCELL_X2 FILLER_98_319 ();
 FILLCELL_X1 FILLER_98_325 ();
 FILLCELL_X2 FILLER_98_329 ();
 FILLCELL_X1 FILLER_98_331 ();
 FILLCELL_X4 FILLER_98_339 ();
 FILLCELL_X1 FILLER_98_343 ();
 FILLCELL_X4 FILLER_98_351 ();
 FILLCELL_X1 FILLER_98_364 ();
 FILLCELL_X2 FILLER_98_381 ();
 FILLCELL_X2 FILLER_98_395 ();
 FILLCELL_X1 FILLER_98_472 ();
 FILLCELL_X1 FILLER_98_490 ();
 FILLCELL_X8 FILLER_98_511 ();
 FILLCELL_X2 FILLER_98_519 ();
 FILLCELL_X1 FILLER_98_542 ();
 FILLCELL_X16 FILLER_98_552 ();
 FILLCELL_X2 FILLER_98_568 ();
 FILLCELL_X1 FILLER_98_570 ();
 FILLCELL_X8 FILLER_98_586 ();
 FILLCELL_X4 FILLER_98_594 ();
 FILLCELL_X2 FILLER_98_598 ();
 FILLCELL_X1 FILLER_98_600 ();
 FILLCELL_X2 FILLER_98_603 ();
 FILLCELL_X1 FILLER_98_605 ();
 FILLCELL_X1 FILLER_98_610 ();
 FILLCELL_X2 FILLER_98_628 ();
 FILLCELL_X1 FILLER_98_630 ();
 FILLCELL_X1 FILLER_98_632 ();
 FILLCELL_X16 FILLER_98_637 ();
 FILLCELL_X8 FILLER_98_653 ();
 FILLCELL_X4 FILLER_98_661 ();
 FILLCELL_X2 FILLER_98_674 ();
 FILLCELL_X1 FILLER_98_676 ();
 FILLCELL_X8 FILLER_98_687 ();
 FILLCELL_X2 FILLER_98_695 ();
 FILLCELL_X1 FILLER_98_704 ();
 FILLCELL_X2 FILLER_98_708 ();
 FILLCELL_X2 FILLER_98_714 ();
 FILLCELL_X1 FILLER_98_716 ();
 FILLCELL_X1 FILLER_98_724 ();
 FILLCELL_X2 FILLER_98_732 ();
 FILLCELL_X1 FILLER_98_734 ();
 FILLCELL_X8 FILLER_98_742 ();
 FILLCELL_X1 FILLER_98_750 ();
 FILLCELL_X16 FILLER_98_758 ();
 FILLCELL_X8 FILLER_98_774 ();
 FILLCELL_X2 FILLER_98_804 ();
 FILLCELL_X1 FILLER_98_806 ();
 FILLCELL_X2 FILLER_98_810 ();
 FILLCELL_X2 FILLER_98_823 ();
 FILLCELL_X2 FILLER_98_832 ();
 FILLCELL_X1 FILLER_98_834 ();
 FILLCELL_X2 FILLER_98_839 ();
 FILLCELL_X1 FILLER_98_841 ();
 FILLCELL_X2 FILLER_98_860 ();
 FILLCELL_X1 FILLER_98_862 ();
 FILLCELL_X4 FILLER_98_867 ();
 FILLCELL_X1 FILLER_98_871 ();
 FILLCELL_X1 FILLER_98_874 ();
 FILLCELL_X8 FILLER_98_896 ();
 FILLCELL_X1 FILLER_98_904 ();
 FILLCELL_X4 FILLER_98_919 ();
 FILLCELL_X2 FILLER_98_923 ();
 FILLCELL_X4 FILLER_98_931 ();
 FILLCELL_X2 FILLER_98_935 ();
 FILLCELL_X8 FILLER_98_944 ();
 FILLCELL_X1 FILLER_98_963 ();
 FILLCELL_X2 FILLER_98_967 ();
 FILLCELL_X1 FILLER_98_976 ();
 FILLCELL_X8 FILLER_98_980 ();
 FILLCELL_X1 FILLER_98_988 ();
 FILLCELL_X8 FILLER_98_996 ();
 FILLCELL_X4 FILLER_98_1004 ();
 FILLCELL_X2 FILLER_98_1008 ();
 FILLCELL_X1 FILLER_98_1010 ();
 FILLCELL_X1 FILLER_98_1014 ();
 FILLCELL_X4 FILLER_98_1062 ();
 FILLCELL_X1 FILLER_98_1066 ();
 FILLCELL_X4 FILLER_98_1078 ();
 FILLCELL_X1 FILLER_98_1106 ();
 FILLCELL_X1 FILLER_98_1114 ();
 FILLCELL_X1 FILLER_98_1119 ();
 FILLCELL_X1 FILLER_98_1127 ();
 FILLCELL_X2 FILLER_98_1132 ();
 FILLCELL_X16 FILLER_98_1140 ();
 FILLCELL_X2 FILLER_98_1156 ();
 FILLCELL_X4 FILLER_98_1165 ();
 FILLCELL_X1 FILLER_98_1174 ();
 FILLCELL_X4 FILLER_98_1177 ();
 FILLCELL_X1 FILLER_98_1181 ();
 FILLCELL_X1 FILLER_98_1193 ();
 FILLCELL_X8 FILLER_98_1196 ();
 FILLCELL_X2 FILLER_98_1204 ();
 FILLCELL_X1 FILLER_98_1206 ();
 FILLCELL_X8 FILLER_98_1212 ();
 FILLCELL_X2 FILLER_98_1220 ();
 FILLCELL_X4 FILLER_98_1236 ();
 FILLCELL_X4 FILLER_98_1242 ();
 FILLCELL_X2 FILLER_98_1246 ();
 FILLCELL_X8 FILLER_98_1252 ();
 FILLCELL_X8 FILLER_99_1 ();
 FILLCELL_X4 FILLER_99_9 ();
 FILLCELL_X1 FILLER_99_13 ();
 FILLCELL_X2 FILLER_99_41 ();
 FILLCELL_X1 FILLER_99_43 ();
 FILLCELL_X4 FILLER_99_51 ();
 FILLCELL_X2 FILLER_99_55 ();
 FILLCELL_X1 FILLER_99_82 ();
 FILLCELL_X16 FILLER_99_110 ();
 FILLCELL_X4 FILLER_99_126 ();
 FILLCELL_X2 FILLER_99_130 ();
 FILLCELL_X4 FILLER_99_179 ();
 FILLCELL_X2 FILLER_99_183 ();
 FILLCELL_X4 FILLER_99_199 ();
 FILLCELL_X2 FILLER_99_203 ();
 FILLCELL_X8 FILLER_99_212 ();
 FILLCELL_X32 FILLER_99_245 ();
 FILLCELL_X2 FILLER_99_277 ();
 FILLCELL_X4 FILLER_99_299 ();
 FILLCELL_X2 FILLER_99_307 ();
 FILLCELL_X4 FILLER_99_329 ();
 FILLCELL_X1 FILLER_99_333 ();
 FILLCELL_X8 FILLER_99_341 ();
 FILLCELL_X4 FILLER_99_363 ();
 FILLCELL_X1 FILLER_99_376 ();
 FILLCELL_X2 FILLER_99_380 ();
 FILLCELL_X2 FILLER_99_388 ();
 FILLCELL_X1 FILLER_99_402 ();
 FILLCELL_X1 FILLER_99_490 ();
 FILLCELL_X2 FILLER_99_504 ();
 FILLCELL_X1 FILLER_99_506 ();
 FILLCELL_X4 FILLER_99_519 ();
 FILLCELL_X2 FILLER_99_523 ();
 FILLCELL_X1 FILLER_99_550 ();
 FILLCELL_X16 FILLER_99_555 ();
 FILLCELL_X2 FILLER_99_571 ();
 FILLCELL_X1 FILLER_99_573 ();
 FILLCELL_X4 FILLER_99_581 ();
 FILLCELL_X1 FILLER_99_609 ();
 FILLCELL_X1 FILLER_99_614 ();
 FILLCELL_X1 FILLER_99_619 ();
 FILLCELL_X16 FILLER_99_636 ();
 FILLCELL_X8 FILLER_99_652 ();
 FILLCELL_X4 FILLER_99_660 ();
 FILLCELL_X2 FILLER_99_664 ();
 FILLCELL_X1 FILLER_99_666 ();
 FILLCELL_X2 FILLER_99_679 ();
 FILLCELL_X2 FILLER_99_695 ();
 FILLCELL_X1 FILLER_99_697 ();
 FILLCELL_X1 FILLER_99_714 ();
 FILLCELL_X2 FILLER_99_718 ();
 FILLCELL_X1 FILLER_99_720 ();
 FILLCELL_X1 FILLER_99_734 ();
 FILLCELL_X8 FILLER_99_742 ();
 FILLCELL_X1 FILLER_99_779 ();
 FILLCELL_X8 FILLER_99_783 ();
 FILLCELL_X2 FILLER_99_791 ();
 FILLCELL_X16 FILLER_99_796 ();
 FILLCELL_X4 FILLER_99_812 ();
 FILLCELL_X4 FILLER_99_827 ();
 FILLCELL_X4 FILLER_99_839 ();
 FILLCELL_X16 FILLER_99_854 ();
 FILLCELL_X8 FILLER_99_870 ();
 FILLCELL_X1 FILLER_99_878 ();
 FILLCELL_X4 FILLER_99_895 ();
 FILLCELL_X8 FILLER_99_911 ();
 FILLCELL_X1 FILLER_99_919 ();
 FILLCELL_X4 FILLER_99_950 ();
 FILLCELL_X4 FILLER_99_974 ();
 FILLCELL_X2 FILLER_99_978 ();
 FILLCELL_X1 FILLER_99_980 ();
 FILLCELL_X16 FILLER_99_1015 ();
 FILLCELL_X4 FILLER_99_1031 ();
 FILLCELL_X32 FILLER_99_1039 ();
 FILLCELL_X1 FILLER_99_1093 ();
 FILLCELL_X1 FILLER_99_1098 ();
 FILLCELL_X8 FILLER_99_1103 ();
 FILLCELL_X2 FILLER_99_1111 ();
 FILLCELL_X1 FILLER_99_1113 ();
 FILLCELL_X2 FILLER_99_1125 ();
 FILLCELL_X2 FILLER_99_1149 ();
 FILLCELL_X1 FILLER_99_1151 ();
 FILLCELL_X2 FILLER_99_1156 ();
 FILLCELL_X1 FILLER_99_1158 ();
 FILLCELL_X2 FILLER_99_1163 ();
 FILLCELL_X16 FILLER_99_1167 ();
 FILLCELL_X2 FILLER_99_1183 ();
 FILLCELL_X1 FILLER_99_1185 ();
 FILLCELL_X2 FILLER_99_1193 ();
 FILLCELL_X4 FILLER_99_1209 ();
 FILLCELL_X1 FILLER_99_1227 ();
 FILLCELL_X8 FILLER_99_1232 ();
 FILLCELL_X8 FILLER_100_1 ();
 FILLCELL_X1 FILLER_100_9 ();
 FILLCELL_X4 FILLER_100_18 ();
 FILLCELL_X2 FILLER_100_22 ();
 FILLCELL_X1 FILLER_100_24 ();
 FILLCELL_X1 FILLER_100_32 ();
 FILLCELL_X2 FILLER_100_47 ();
 FILLCELL_X4 FILLER_100_56 ();
 FILLCELL_X2 FILLER_100_60 ();
 FILLCELL_X1 FILLER_100_62 ();
 FILLCELL_X4 FILLER_100_70 ();
 FILLCELL_X4 FILLER_100_101 ();
 FILLCELL_X1 FILLER_100_119 ();
 FILLCELL_X1 FILLER_100_127 ();
 FILLCELL_X1 FILLER_100_135 ();
 FILLCELL_X1 FILLER_100_143 ();
 FILLCELL_X2 FILLER_100_159 ();
 FILLCELL_X4 FILLER_100_165 ();
 FILLCELL_X1 FILLER_100_169 ();
 FILLCELL_X8 FILLER_100_187 ();
 FILLCELL_X4 FILLER_100_228 ();
 FILLCELL_X2 FILLER_100_232 ();
 FILLCELL_X1 FILLER_100_234 ();
 FILLCELL_X8 FILLER_100_249 ();
 FILLCELL_X1 FILLER_100_257 ();
 FILLCELL_X4 FILLER_100_293 ();
 FILLCELL_X8 FILLER_100_345 ();
 FILLCELL_X2 FILLER_100_353 ();
 FILLCELL_X2 FILLER_100_364 ();
 FILLCELL_X1 FILLER_100_366 ();
 FILLCELL_X1 FILLER_100_371 ();
 FILLCELL_X2 FILLER_100_399 ();
 FILLCELL_X1 FILLER_100_401 ();
 FILLCELL_X2 FILLER_100_428 ();
 FILLCELL_X2 FILLER_100_439 ();
 FILLCELL_X4 FILLER_100_450 ();
 FILLCELL_X1 FILLER_100_477 ();
 FILLCELL_X1 FILLER_100_507 ();
 FILLCELL_X8 FILLER_100_529 ();
 FILLCELL_X4 FILLER_100_537 ();
 FILLCELL_X2 FILLER_100_541 ();
 FILLCELL_X1 FILLER_100_543 ();
 FILLCELL_X1 FILLER_100_565 ();
 FILLCELL_X4 FILLER_100_570 ();
 FILLCELL_X1 FILLER_100_574 ();
 FILLCELL_X8 FILLER_100_582 ();
 FILLCELL_X2 FILLER_100_597 ();
 FILLCELL_X1 FILLER_100_599 ();
 FILLCELL_X2 FILLER_100_604 ();
 FILLCELL_X2 FILLER_100_611 ();
 FILLCELL_X1 FILLER_100_617 ();
 FILLCELL_X2 FILLER_100_622 ();
 FILLCELL_X1 FILLER_100_624 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X16 FILLER_100_632 ();
 FILLCELL_X4 FILLER_100_648 ();
 FILLCELL_X1 FILLER_100_652 ();
 FILLCELL_X4 FILLER_100_656 ();
 FILLCELL_X2 FILLER_100_660 ();
 FILLCELL_X2 FILLER_100_679 ();
 FILLCELL_X1 FILLER_100_690 ();
 FILLCELL_X4 FILLER_100_695 ();
 FILLCELL_X1 FILLER_100_699 ();
 FILLCELL_X1 FILLER_100_722 ();
 FILLCELL_X8 FILLER_100_727 ();
 FILLCELL_X4 FILLER_100_735 ();
 FILLCELL_X8 FILLER_100_746 ();
 FILLCELL_X1 FILLER_100_754 ();
 FILLCELL_X8 FILLER_100_759 ();
 FILLCELL_X4 FILLER_100_767 ();
 FILLCELL_X1 FILLER_100_771 ();
 FILLCELL_X4 FILLER_100_783 ();
 FILLCELL_X1 FILLER_100_787 ();
 FILLCELL_X1 FILLER_100_799 ();
 FILLCELL_X1 FILLER_100_809 ();
 FILLCELL_X1 FILLER_100_824 ();
 FILLCELL_X2 FILLER_100_829 ();
 FILLCELL_X2 FILLER_100_836 ();
 FILLCELL_X2 FILLER_100_842 ();
 FILLCELL_X1 FILLER_100_848 ();
 FILLCELL_X8 FILLER_100_874 ();
 FILLCELL_X4 FILLER_100_882 ();
 FILLCELL_X2 FILLER_100_886 ();
 FILLCELL_X1 FILLER_100_888 ();
 FILLCELL_X4 FILLER_100_893 ();
 FILLCELL_X2 FILLER_100_897 ();
 FILLCELL_X1 FILLER_100_899 ();
 FILLCELL_X16 FILLER_100_903 ();
 FILLCELL_X4 FILLER_100_919 ();
 FILLCELL_X2 FILLER_100_923 ();
 FILLCELL_X1 FILLER_100_925 ();
 FILLCELL_X4 FILLER_100_933 ();
 FILLCELL_X1 FILLER_100_937 ();
 FILLCELL_X2 FILLER_100_942 ();
 FILLCELL_X1 FILLER_100_955 ();
 FILLCELL_X2 FILLER_100_962 ();
 FILLCELL_X2 FILLER_100_969 ();
 FILLCELL_X1 FILLER_100_971 ();
 FILLCELL_X1 FILLER_100_980 ();
 FILLCELL_X1 FILLER_100_988 ();
 FILLCELL_X2 FILLER_100_992 ();
 FILLCELL_X1 FILLER_100_994 ();
 FILLCELL_X2 FILLER_100_1002 ();
 FILLCELL_X1 FILLER_100_1006 ();
 FILLCELL_X1 FILLER_100_1010 ();
 FILLCELL_X1 FILLER_100_1018 ();
 FILLCELL_X1 FILLER_100_1035 ();
 FILLCELL_X2 FILLER_100_1039 ();
 FILLCELL_X2 FILLER_100_1061 ();
 FILLCELL_X1 FILLER_100_1063 ();
 FILLCELL_X2 FILLER_100_1086 ();
 FILLCELL_X1 FILLER_100_1088 ();
 FILLCELL_X1 FILLER_100_1093 ();
 FILLCELL_X1 FILLER_100_1098 ();
 FILLCELL_X4 FILLER_100_1103 ();
 FILLCELL_X1 FILLER_100_1107 ();
 FILLCELL_X2 FILLER_100_1125 ();
 FILLCELL_X8 FILLER_100_1131 ();
 FILLCELL_X4 FILLER_100_1148 ();
 FILLCELL_X8 FILLER_100_1183 ();
 FILLCELL_X2 FILLER_100_1191 ();
 FILLCELL_X8 FILLER_100_1230 ();
 FILLCELL_X4 FILLER_100_1252 ();
 FILLCELL_X1 FILLER_100_1256 ();
 FILLCELL_X1 FILLER_100_1259 ();
 FILLCELL_X1 FILLER_101_35 ();
 FILLCELL_X4 FILLER_101_50 ();
 FILLCELL_X1 FILLER_101_74 ();
 FILLCELL_X2 FILLER_101_82 ();
 FILLCELL_X4 FILLER_101_109 ();
 FILLCELL_X2 FILLER_101_127 ();
 FILLCELL_X8 FILLER_101_136 ();
 FILLCELL_X2 FILLER_101_144 ();
 FILLCELL_X1 FILLER_101_146 ();
 FILLCELL_X2 FILLER_101_161 ();
 FILLCELL_X2 FILLER_101_170 ();
 FILLCELL_X1 FILLER_101_172 ();
 FILLCELL_X2 FILLER_101_193 ();
 FILLCELL_X1 FILLER_101_195 ();
 FILLCELL_X1 FILLER_101_223 ();
 FILLCELL_X2 FILLER_101_244 ();
 FILLCELL_X1 FILLER_101_246 ();
 FILLCELL_X8 FILLER_101_254 ();
 FILLCELL_X1 FILLER_101_262 ();
 FILLCELL_X1 FILLER_101_283 ();
 FILLCELL_X2 FILLER_101_304 ();
 FILLCELL_X2 FILLER_101_310 ();
 FILLCELL_X2 FILLER_101_315 ();
 FILLCELL_X1 FILLER_101_320 ();
 FILLCELL_X1 FILLER_101_349 ();
 FILLCELL_X1 FILLER_101_360 ();
 FILLCELL_X1 FILLER_101_364 ();
 FILLCELL_X4 FILLER_101_374 ();
 FILLCELL_X1 FILLER_101_378 ();
 FILLCELL_X2 FILLER_101_386 ();
 FILLCELL_X1 FILLER_101_411 ();
 FILLCELL_X1 FILLER_101_416 ();
 FILLCELL_X8 FILLER_101_426 ();
 FILLCELL_X1 FILLER_101_434 ();
 FILLCELL_X8 FILLER_101_460 ();
 FILLCELL_X2 FILLER_101_468 ();
 FILLCELL_X1 FILLER_101_470 ();
 FILLCELL_X1 FILLER_101_478 ();
 FILLCELL_X2 FILLER_101_492 ();
 FILLCELL_X8 FILLER_101_497 ();
 FILLCELL_X2 FILLER_101_537 ();
 FILLCELL_X1 FILLER_101_539 ();
 FILLCELL_X4 FILLER_101_544 ();
 FILLCELL_X4 FILLER_101_578 ();
 FILLCELL_X4 FILLER_101_606 ();
 FILLCELL_X2 FILLER_101_610 ();
 FILLCELL_X1 FILLER_101_612 ();
 FILLCELL_X4 FILLER_101_640 ();
 FILLCELL_X2 FILLER_101_644 ();
 FILLCELL_X1 FILLER_101_646 ();
 FILLCELL_X16 FILLER_101_652 ();
 FILLCELL_X8 FILLER_101_668 ();
 FILLCELL_X2 FILLER_101_676 ();
 FILLCELL_X4 FILLER_101_685 ();
 FILLCELL_X2 FILLER_101_698 ();
 FILLCELL_X8 FILLER_101_707 ();
 FILLCELL_X4 FILLER_101_718 ();
 FILLCELL_X1 FILLER_101_722 ();
 FILLCELL_X8 FILLER_101_730 ();
 FILLCELL_X2 FILLER_101_738 ();
 FILLCELL_X8 FILLER_101_761 ();
 FILLCELL_X2 FILLER_101_769 ();
 FILLCELL_X16 FILLER_101_780 ();
 FILLCELL_X8 FILLER_101_796 ();
 FILLCELL_X4 FILLER_101_804 ();
 FILLCELL_X2 FILLER_101_812 ();
 FILLCELL_X1 FILLER_101_814 ();
 FILLCELL_X8 FILLER_101_826 ();
 FILLCELL_X2 FILLER_101_834 ();
 FILLCELL_X1 FILLER_101_836 ();
 FILLCELL_X1 FILLER_101_841 ();
 FILLCELL_X4 FILLER_101_853 ();
 FILLCELL_X2 FILLER_101_857 ();
 FILLCELL_X2 FILLER_101_862 ();
 FILLCELL_X8 FILLER_101_868 ();
 FILLCELL_X2 FILLER_101_876 ();
 FILLCELL_X1 FILLER_101_878 ();
 FILLCELL_X8 FILLER_101_883 ();
 FILLCELL_X4 FILLER_101_891 ();
 FILLCELL_X8 FILLER_101_917 ();
 FILLCELL_X2 FILLER_101_925 ();
 FILLCELL_X1 FILLER_101_931 ();
 FILLCELL_X4 FILLER_101_936 ();
 FILLCELL_X1 FILLER_101_950 ();
 FILLCELL_X4 FILLER_101_960 ();
 FILLCELL_X2 FILLER_101_964 ();
 FILLCELL_X1 FILLER_101_966 ();
 FILLCELL_X4 FILLER_101_971 ();
 FILLCELL_X1 FILLER_101_975 ();
 FILLCELL_X1 FILLER_101_982 ();
 FILLCELL_X4 FILLER_101_1058 ();
 FILLCELL_X2 FILLER_101_1062 ();
 FILLCELL_X1 FILLER_101_1064 ();
 FILLCELL_X4 FILLER_101_1069 ();
 FILLCELL_X1 FILLER_101_1073 ();
 FILLCELL_X2 FILLER_101_1081 ();
 FILLCELL_X1 FILLER_101_1083 ();
 FILLCELL_X2 FILLER_101_1088 ();
 FILLCELL_X2 FILLER_101_1113 ();
 FILLCELL_X1 FILLER_101_1118 ();
 FILLCELL_X4 FILLER_101_1123 ();
 FILLCELL_X1 FILLER_101_1136 ();
 FILLCELL_X8 FILLER_101_1166 ();
 FILLCELL_X4 FILLER_101_1174 ();
 FILLCELL_X2 FILLER_101_1178 ();
 FILLCELL_X1 FILLER_101_1180 ();
 FILLCELL_X8 FILLER_101_1185 ();
 FILLCELL_X8 FILLER_101_1211 ();
 FILLCELL_X4 FILLER_101_1256 ();
 FILLCELL_X8 FILLER_102_1 ();
 FILLCELL_X4 FILLER_102_9 ();
 FILLCELL_X2 FILLER_102_13 ();
 FILLCELL_X8 FILLER_102_42 ();
 FILLCELL_X1 FILLER_102_50 ();
 FILLCELL_X2 FILLER_102_78 ();
 FILLCELL_X1 FILLER_102_80 ();
 FILLCELL_X1 FILLER_102_120 ();
 FILLCELL_X1 FILLER_102_128 ();
 FILLCELL_X1 FILLER_102_132 ();
 FILLCELL_X1 FILLER_102_153 ();
 FILLCELL_X1 FILLER_102_174 ();
 FILLCELL_X32 FILLER_102_179 ();
 FILLCELL_X4 FILLER_102_211 ();
 FILLCELL_X1 FILLER_102_215 ();
 FILLCELL_X4 FILLER_102_223 ();
 FILLCELL_X2 FILLER_102_227 ();
 FILLCELL_X1 FILLER_102_229 ();
 FILLCELL_X8 FILLER_102_244 ();
 FILLCELL_X4 FILLER_102_252 ();
 FILLCELL_X1 FILLER_102_256 ();
 FILLCELL_X4 FILLER_102_275 ();
 FILLCELL_X1 FILLER_102_279 ();
 FILLCELL_X8 FILLER_102_287 ();
 FILLCELL_X4 FILLER_102_295 ();
 FILLCELL_X1 FILLER_102_303 ();
 FILLCELL_X1 FILLER_102_324 ();
 FILLCELL_X4 FILLER_102_332 ();
 FILLCELL_X2 FILLER_102_336 ();
 FILLCELL_X1 FILLER_102_338 ();
 FILLCELL_X16 FILLER_102_367 ();
 FILLCELL_X2 FILLER_102_383 ();
 FILLCELL_X1 FILLER_102_385 ();
 FILLCELL_X4 FILLER_102_411 ();
 FILLCELL_X8 FILLER_102_422 ();
 FILLCELL_X2 FILLER_102_430 ();
 FILLCELL_X8 FILLER_102_437 ();
 FILLCELL_X4 FILLER_102_452 ();
 FILLCELL_X2 FILLER_102_456 ();
 FILLCELL_X4 FILLER_102_478 ();
 FILLCELL_X4 FILLER_102_489 ();
 FILLCELL_X2 FILLER_102_493 ();
 FILLCELL_X1 FILLER_102_495 ();
 FILLCELL_X1 FILLER_102_553 ();
 FILLCELL_X4 FILLER_102_578 ();
 FILLCELL_X2 FILLER_102_582 ();
 FILLCELL_X8 FILLER_102_604 ();
 FILLCELL_X8 FILLER_102_619 ();
 FILLCELL_X4 FILLER_102_627 ();
 FILLCELL_X8 FILLER_102_639 ();
 FILLCELL_X1 FILLER_102_647 ();
 FILLCELL_X2 FILLER_102_661 ();
 FILLCELL_X1 FILLER_102_663 ();
 FILLCELL_X4 FILLER_102_684 ();
 FILLCELL_X4 FILLER_102_725 ();
 FILLCELL_X4 FILLER_102_745 ();
 FILLCELL_X1 FILLER_102_749 ();
 FILLCELL_X32 FILLER_102_755 ();
 FILLCELL_X2 FILLER_102_794 ();
 FILLCELL_X1 FILLER_102_796 ();
 FILLCELL_X4 FILLER_102_800 ();
 FILLCELL_X16 FILLER_102_807 ();
 FILLCELL_X8 FILLER_102_823 ();
 FILLCELL_X2 FILLER_102_831 ();
 FILLCELL_X1 FILLER_102_833 ();
 FILLCELL_X2 FILLER_102_838 ();
 FILLCELL_X2 FILLER_102_844 ();
 FILLCELL_X1 FILLER_102_846 ();
 FILLCELL_X2 FILLER_102_858 ();
 FILLCELL_X1 FILLER_102_860 ();
 FILLCELL_X8 FILLER_102_864 ();
 FILLCELL_X4 FILLER_102_872 ();
 FILLCELL_X2 FILLER_102_876 ();
 FILLCELL_X1 FILLER_102_878 ();
 FILLCELL_X4 FILLER_102_886 ();
 FILLCELL_X2 FILLER_102_890 ();
 FILLCELL_X1 FILLER_102_892 ();
 FILLCELL_X4 FILLER_102_897 ();
 FILLCELL_X2 FILLER_102_921 ();
 FILLCELL_X1 FILLER_102_939 ();
 FILLCELL_X2 FILLER_102_958 ();
 FILLCELL_X2 FILLER_102_971 ();
 FILLCELL_X1 FILLER_102_973 ();
 FILLCELL_X16 FILLER_102_977 ();
 FILLCELL_X4 FILLER_102_993 ();
 FILLCELL_X8 FILLER_102_1008 ();
 FILLCELL_X8 FILLER_102_1020 ();
 FILLCELL_X1 FILLER_102_1028 ();
 FILLCELL_X4 FILLER_102_1048 ();
 FILLCELL_X2 FILLER_102_1052 ();
 FILLCELL_X1 FILLER_102_1054 ();
 FILLCELL_X8 FILLER_102_1068 ();
 FILLCELL_X1 FILLER_102_1076 ();
 FILLCELL_X1 FILLER_102_1084 ();
 FILLCELL_X1 FILLER_102_1092 ();
 FILLCELL_X1 FILLER_102_1096 ();
 FILLCELL_X1 FILLER_102_1101 ();
 FILLCELL_X1 FILLER_102_1109 ();
 FILLCELL_X2 FILLER_102_1113 ();
 FILLCELL_X1 FILLER_102_1115 ();
 FILLCELL_X8 FILLER_102_1119 ();
 FILLCELL_X1 FILLER_102_1127 ();
 FILLCELL_X16 FILLER_102_1160 ();
 FILLCELL_X8 FILLER_102_1230 ();
 FILLCELL_X1 FILLER_102_1238 ();
 FILLCELL_X1 FILLER_102_1259 ();
 FILLCELL_X4 FILLER_103_21 ();
 FILLCELL_X2 FILLER_103_32 ();
 FILLCELL_X16 FILLER_103_48 ();
 FILLCELL_X8 FILLER_103_64 ();
 FILLCELL_X4 FILLER_103_72 ();
 FILLCELL_X1 FILLER_103_76 ();
 FILLCELL_X4 FILLER_103_104 ();
 FILLCELL_X2 FILLER_103_108 ();
 FILLCELL_X2 FILLER_103_131 ();
 FILLCELL_X2 FILLER_103_140 ();
 FILLCELL_X16 FILLER_103_155 ();
 FILLCELL_X1 FILLER_103_171 ();
 FILLCELL_X1 FILLER_103_181 ();
 FILLCELL_X1 FILLER_103_188 ();
 FILLCELL_X2 FILLER_103_193 ();
 FILLCELL_X1 FILLER_103_195 ();
 FILLCELL_X1 FILLER_103_198 ();
 FILLCELL_X8 FILLER_103_209 ();
 FILLCELL_X4 FILLER_103_217 ();
 FILLCELL_X4 FILLER_103_228 ();
 FILLCELL_X2 FILLER_103_232 ();
 FILLCELL_X1 FILLER_103_258 ();
 FILLCELL_X2 FILLER_103_266 ();
 FILLCELL_X1 FILLER_103_268 ();
 FILLCELL_X4 FILLER_103_276 ();
 FILLCELL_X2 FILLER_103_280 ();
 FILLCELL_X1 FILLER_103_282 ();
 FILLCELL_X8 FILLER_103_313 ();
 FILLCELL_X8 FILLER_103_342 ();
 FILLCELL_X1 FILLER_103_350 ();
 FILLCELL_X1 FILLER_103_362 ();
 FILLCELL_X1 FILLER_103_367 ();
 FILLCELL_X2 FILLER_103_387 ();
 FILLCELL_X2 FILLER_103_401 ();
 FILLCELL_X16 FILLER_103_406 ();
 FILLCELL_X4 FILLER_103_422 ();
 FILLCELL_X16 FILLER_103_446 ();
 FILLCELL_X16 FILLER_103_469 ();
 FILLCELL_X2 FILLER_103_485 ();
 FILLCELL_X2 FILLER_103_507 ();
 FILLCELL_X1 FILLER_103_509 ();
 FILLCELL_X1 FILLER_103_518 ();
 FILLCELL_X16 FILLER_103_526 ();
 FILLCELL_X8 FILLER_103_545 ();
 FILLCELL_X4 FILLER_103_553 ();
 FILLCELL_X2 FILLER_103_557 ();
 FILLCELL_X4 FILLER_103_563 ();
 FILLCELL_X1 FILLER_103_567 ();
 FILLCELL_X2 FILLER_103_578 ();
 FILLCELL_X4 FILLER_103_587 ();
 FILLCELL_X2 FILLER_103_591 ();
 FILLCELL_X1 FILLER_103_593 ();
 FILLCELL_X8 FILLER_103_619 ();
 FILLCELL_X1 FILLER_103_627 ();
 FILLCELL_X8 FILLER_103_650 ();
 FILLCELL_X1 FILLER_103_658 ();
 FILLCELL_X8 FILLER_103_664 ();
 FILLCELL_X8 FILLER_103_679 ();
 FILLCELL_X4 FILLER_103_687 ();
 FILLCELL_X1 FILLER_103_695 ();
 FILLCELL_X2 FILLER_103_703 ();
 FILLCELL_X1 FILLER_103_705 ();
 FILLCELL_X1 FILLER_103_710 ();
 FILLCELL_X8 FILLER_103_737 ();
 FILLCELL_X4 FILLER_103_745 ();
 FILLCELL_X2 FILLER_103_749 ();
 FILLCELL_X8 FILLER_103_770 ();
 FILLCELL_X2 FILLER_103_778 ();
 FILLCELL_X8 FILLER_103_797 ();
 FILLCELL_X4 FILLER_103_805 ();
 FILLCELL_X1 FILLER_103_809 ();
 FILLCELL_X2 FILLER_103_828 ();
 FILLCELL_X4 FILLER_103_837 ();
 FILLCELL_X1 FILLER_103_844 ();
 FILLCELL_X4 FILLER_103_859 ();
 FILLCELL_X2 FILLER_103_863 ();
 FILLCELL_X2 FILLER_103_885 ();
 FILLCELL_X1 FILLER_103_887 ();
 FILLCELL_X8 FILLER_103_901 ();
 FILLCELL_X4 FILLER_103_909 ();
 FILLCELL_X2 FILLER_103_913 ();
 FILLCELL_X2 FILLER_103_918 ();
 FILLCELL_X1 FILLER_103_920 ();
 FILLCELL_X1 FILLER_103_945 ();
 FILLCELL_X1 FILLER_103_960 ();
 FILLCELL_X2 FILLER_103_968 ();
 FILLCELL_X1 FILLER_103_984 ();
 FILLCELL_X8 FILLER_103_996 ();
 FILLCELL_X4 FILLER_103_1004 ();
 FILLCELL_X2 FILLER_103_1008 ();
 FILLCELL_X4 FILLER_103_1035 ();
 FILLCELL_X2 FILLER_103_1039 ();
 FILLCELL_X1 FILLER_103_1073 ();
 FILLCELL_X1 FILLER_103_1088 ();
 FILLCELL_X1 FILLER_103_1096 ();
 FILLCELL_X4 FILLER_103_1118 ();
 FILLCELL_X2 FILLER_103_1125 ();
 FILLCELL_X1 FILLER_103_1137 ();
 FILLCELL_X8 FILLER_103_1141 ();
 FILLCELL_X4 FILLER_103_1149 ();
 FILLCELL_X16 FILLER_103_1163 ();
 FILLCELL_X1 FILLER_103_1179 ();
 FILLCELL_X1 FILLER_103_1186 ();
 FILLCELL_X2 FILLER_103_1192 ();
 FILLCELL_X2 FILLER_103_1201 ();
 FILLCELL_X1 FILLER_103_1203 ();
 FILLCELL_X1 FILLER_103_1216 ();
 FILLCELL_X2 FILLER_103_1231 ();
 FILLCELL_X8 FILLER_103_1240 ();
 FILLCELL_X2 FILLER_103_1248 ();
 FILLCELL_X8 FILLER_104_1 ();
 FILLCELL_X2 FILLER_104_43 ();
 FILLCELL_X1 FILLER_104_45 ();
 FILLCELL_X16 FILLER_104_60 ();
 FILLCELL_X4 FILLER_104_76 ();
 FILLCELL_X1 FILLER_104_80 ();
 FILLCELL_X2 FILLER_104_93 ();
 FILLCELL_X16 FILLER_104_105 ();
 FILLCELL_X4 FILLER_104_121 ();
 FILLCELL_X2 FILLER_104_125 ();
 FILLCELL_X1 FILLER_104_127 ();
 FILLCELL_X1 FILLER_104_138 ();
 FILLCELL_X8 FILLER_104_150 ();
 FILLCELL_X8 FILLER_104_220 ();
 FILLCELL_X4 FILLER_104_228 ();
 FILLCELL_X2 FILLER_104_232 ();
 FILLCELL_X1 FILLER_104_234 ();
 FILLCELL_X16 FILLER_104_254 ();
 FILLCELL_X4 FILLER_104_270 ();
 FILLCELL_X2 FILLER_104_274 ();
 FILLCELL_X2 FILLER_104_297 ();
 FILLCELL_X4 FILLER_104_326 ();
 FILLCELL_X4 FILLER_104_337 ();
 FILLCELL_X2 FILLER_104_341 ();
 FILLCELL_X1 FILLER_104_343 ();
 FILLCELL_X2 FILLER_104_349 ();
 FILLCELL_X8 FILLER_104_374 ();
 FILLCELL_X2 FILLER_104_382 ();
 FILLCELL_X1 FILLER_104_384 ();
 FILLCELL_X1 FILLER_104_405 ();
 FILLCELL_X4 FILLER_104_413 ();
 FILLCELL_X2 FILLER_104_417 ();
 FILLCELL_X1 FILLER_104_419 ();
 FILLCELL_X2 FILLER_104_433 ();
 FILLCELL_X1 FILLER_104_496 ();
 FILLCELL_X2 FILLER_104_500 ();
 FILLCELL_X1 FILLER_104_502 ();
 FILLCELL_X4 FILLER_104_507 ();
 FILLCELL_X2 FILLER_104_511 ();
 FILLCELL_X1 FILLER_104_513 ();
 FILLCELL_X2 FILLER_104_516 ();
 FILLCELL_X8 FILLER_104_528 ();
 FILLCELL_X2 FILLER_104_536 ();
 FILLCELL_X1 FILLER_104_545 ();
 FILLCELL_X8 FILLER_104_578 ();
 FILLCELL_X1 FILLER_104_586 ();
 FILLCELL_X8 FILLER_104_594 ();
 FILLCELL_X4 FILLER_104_602 ();
 FILLCELL_X2 FILLER_104_606 ();
 FILLCELL_X1 FILLER_104_608 ();
 FILLCELL_X2 FILLER_104_616 ();
 FILLCELL_X1 FILLER_104_618 ();
 FILLCELL_X8 FILLER_104_622 ();
 FILLCELL_X1 FILLER_104_630 ();
 FILLCELL_X2 FILLER_104_632 ();
 FILLCELL_X16 FILLER_104_639 ();
 FILLCELL_X8 FILLER_104_655 ();
 FILLCELL_X4 FILLER_104_663 ();
 FILLCELL_X2 FILLER_104_667 ();
 FILLCELL_X1 FILLER_104_669 ();
 FILLCELL_X2 FILLER_104_682 ();
 FILLCELL_X8 FILLER_104_687 ();
 FILLCELL_X4 FILLER_104_695 ();
 FILLCELL_X2 FILLER_104_710 ();
 FILLCELL_X2 FILLER_104_715 ();
 FILLCELL_X1 FILLER_104_748 ();
 FILLCELL_X2 FILLER_104_756 ();
 FILLCELL_X1 FILLER_104_758 ();
 FILLCELL_X8 FILLER_104_762 ();
 FILLCELL_X2 FILLER_104_770 ();
 FILLCELL_X1 FILLER_104_772 ();
 FILLCELL_X8 FILLER_104_778 ();
 FILLCELL_X2 FILLER_104_786 ();
 FILLCELL_X1 FILLER_104_788 ();
 FILLCELL_X2 FILLER_104_794 ();
 FILLCELL_X8 FILLER_104_804 ();
 FILLCELL_X2 FILLER_104_812 ();
 FILLCELL_X1 FILLER_104_814 ();
 FILLCELL_X1 FILLER_104_821 ();
 FILLCELL_X4 FILLER_104_827 ();
 FILLCELL_X2 FILLER_104_831 ();
 FILLCELL_X1 FILLER_104_833 ();
 FILLCELL_X2 FILLER_104_845 ();
 FILLCELL_X4 FILLER_104_860 ();
 FILLCELL_X2 FILLER_104_864 ();
 FILLCELL_X1 FILLER_104_880 ();
 FILLCELL_X2 FILLER_104_885 ();
 FILLCELL_X1 FILLER_104_887 ();
 FILLCELL_X2 FILLER_104_895 ();
 FILLCELL_X1 FILLER_104_897 ();
 FILLCELL_X4 FILLER_104_901 ();
 FILLCELL_X1 FILLER_104_908 ();
 FILLCELL_X1 FILLER_104_916 ();
 FILLCELL_X2 FILLER_104_920 ();
 FILLCELL_X8 FILLER_104_926 ();
 FILLCELL_X2 FILLER_104_934 ();
 FILLCELL_X1 FILLER_104_936 ();
 FILLCELL_X4 FILLER_104_940 ();
 FILLCELL_X2 FILLER_104_944 ();
 FILLCELL_X2 FILLER_104_949 ();
 FILLCELL_X1 FILLER_104_951 ();
 FILLCELL_X1 FILLER_104_958 ();
 FILLCELL_X2 FILLER_104_969 ();
 FILLCELL_X1 FILLER_104_971 ();
 FILLCELL_X4 FILLER_104_976 ();
 FILLCELL_X1 FILLER_104_980 ();
 FILLCELL_X8 FILLER_104_992 ();
 FILLCELL_X2 FILLER_104_1000 ();
 FILLCELL_X1 FILLER_104_1002 ();
 FILLCELL_X1 FILLER_104_1015 ();
 FILLCELL_X1 FILLER_104_1021 ();
 FILLCELL_X2 FILLER_104_1026 ();
 FILLCELL_X2 FILLER_104_1041 ();
 FILLCELL_X1 FILLER_104_1043 ();
 FILLCELL_X4 FILLER_104_1050 ();
 FILLCELL_X8 FILLER_104_1064 ();
 FILLCELL_X2 FILLER_104_1072 ();
 FILLCELL_X2 FILLER_104_1130 ();
 FILLCELL_X1 FILLER_104_1139 ();
 FILLCELL_X2 FILLER_104_1200 ();
 FILLCELL_X1 FILLER_104_1205 ();
 FILLCELL_X4 FILLER_105_21 ();
 FILLCELL_X1 FILLER_105_25 ();
 FILLCELL_X4 FILLER_105_33 ();
 FILLCELL_X2 FILLER_105_37 ();
 FILLCELL_X1 FILLER_105_39 ();
 FILLCELL_X8 FILLER_105_67 ();
 FILLCELL_X4 FILLER_105_75 ();
 FILLCELL_X2 FILLER_105_79 ();
 FILLCELL_X1 FILLER_105_81 ();
 FILLCELL_X1 FILLER_105_109 ();
 FILLCELL_X2 FILLER_105_117 ();
 FILLCELL_X4 FILLER_105_133 ();
 FILLCELL_X2 FILLER_105_137 ();
 FILLCELL_X1 FILLER_105_139 ();
 FILLCELL_X8 FILLER_105_179 ();
 FILLCELL_X2 FILLER_105_187 ();
 FILLCELL_X8 FILLER_105_207 ();
 FILLCELL_X2 FILLER_105_215 ();
 FILLCELL_X4 FILLER_105_224 ();
 FILLCELL_X2 FILLER_105_228 ();
 FILLCELL_X1 FILLER_105_230 ();
 FILLCELL_X4 FILLER_105_245 ();
 FILLCELL_X2 FILLER_105_249 ();
 FILLCELL_X1 FILLER_105_251 ();
 FILLCELL_X8 FILLER_105_266 ();
 FILLCELL_X4 FILLER_105_274 ();
 FILLCELL_X4 FILLER_105_285 ();
 FILLCELL_X1 FILLER_105_289 ();
 FILLCELL_X16 FILLER_105_297 ();
 FILLCELL_X4 FILLER_105_313 ();
 FILLCELL_X8 FILLER_105_345 ();
 FILLCELL_X2 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_375 ();
 FILLCELL_X1 FILLER_105_407 ();
 FILLCELL_X8 FILLER_105_442 ();
 FILLCELL_X1 FILLER_105_450 ();
 FILLCELL_X1 FILLER_105_486 ();
 FILLCELL_X2 FILLER_105_494 ();
 FILLCELL_X2 FILLER_105_523 ();
 FILLCELL_X8 FILLER_105_555 ();
 FILLCELL_X1 FILLER_105_630 ();
 FILLCELL_X2 FILLER_105_644 ();
 FILLCELL_X1 FILLER_105_650 ();
 FILLCELL_X4 FILLER_105_664 ();
 FILLCELL_X2 FILLER_105_668 ();
 FILLCELL_X2 FILLER_105_673 ();
 FILLCELL_X1 FILLER_105_675 ();
 FILLCELL_X4 FILLER_105_683 ();
 FILLCELL_X8 FILLER_105_696 ();
 FILLCELL_X2 FILLER_105_711 ();
 FILLCELL_X2 FILLER_105_724 ();
 FILLCELL_X1 FILLER_105_726 ();
 FILLCELL_X4 FILLER_105_731 ();
 FILLCELL_X16 FILLER_105_740 ();
 FILLCELL_X1 FILLER_105_763 ();
 FILLCELL_X4 FILLER_105_771 ();
 FILLCELL_X8 FILLER_105_786 ();
 FILLCELL_X2 FILLER_105_794 ();
 FILLCELL_X1 FILLER_105_799 ();
 FILLCELL_X2 FILLER_105_808 ();
 FILLCELL_X4 FILLER_105_821 ();
 FILLCELL_X1 FILLER_105_825 ();
 FILLCELL_X4 FILLER_105_844 ();
 FILLCELL_X1 FILLER_105_848 ();
 FILLCELL_X4 FILLER_105_853 ();
 FILLCELL_X4 FILLER_105_870 ();
 FILLCELL_X8 FILLER_105_877 ();
 FILLCELL_X1 FILLER_105_888 ();
 FILLCELL_X1 FILLER_105_896 ();
 FILLCELL_X2 FILLER_105_910 ();
 FILLCELL_X2 FILLER_105_932 ();
 FILLCELL_X1 FILLER_105_934 ();
 FILLCELL_X2 FILLER_105_947 ();
 FILLCELL_X4 FILLER_105_957 ();
 FILLCELL_X2 FILLER_105_961 ();
 FILLCELL_X1 FILLER_105_963 ();
 FILLCELL_X8 FILLER_105_971 ();
 FILLCELL_X4 FILLER_105_988 ();
 FILLCELL_X1 FILLER_105_1033 ();
 FILLCELL_X8 FILLER_105_1064 ();
 FILLCELL_X2 FILLER_105_1072 ();
 FILLCELL_X2 FILLER_105_1099 ();
 FILLCELL_X2 FILLER_105_1104 ();
 FILLCELL_X16 FILLER_105_1113 ();
 FILLCELL_X4 FILLER_105_1133 ();
 FILLCELL_X1 FILLER_105_1137 ();
 FILLCELL_X2 FILLER_105_1145 ();
 FILLCELL_X4 FILLER_105_1154 ();
 FILLCELL_X1 FILLER_105_1158 ();
 FILLCELL_X1 FILLER_105_1166 ();
 FILLCELL_X8 FILLER_105_1172 ();
 FILLCELL_X4 FILLER_105_1180 ();
 FILLCELL_X4 FILLER_105_1189 ();
 FILLCELL_X1 FILLER_105_1193 ();
 FILLCELL_X1 FILLER_105_1210 ();
 FILLCELL_X2 FILLER_105_1214 ();
 FILLCELL_X2 FILLER_105_1221 ();
 FILLCELL_X4 FILLER_105_1230 ();
 FILLCELL_X2 FILLER_105_1234 ();
 FILLCELL_X4 FILLER_105_1243 ();
 FILLCELL_X2 FILLER_105_1254 ();
 FILLCELL_X1 FILLER_105_1259 ();
 FILLCELL_X4 FILLER_106_1 ();
 FILLCELL_X2 FILLER_106_5 ();
 FILLCELL_X16 FILLER_106_41 ();
 FILLCELL_X4 FILLER_106_84 ();
 FILLCELL_X2 FILLER_106_88 ();
 FILLCELL_X8 FILLER_106_118 ();
 FILLCELL_X2 FILLER_106_146 ();
 FILLCELL_X2 FILLER_106_155 ();
 FILLCELL_X4 FILLER_106_173 ();
 FILLCELL_X2 FILLER_106_177 ();
 FILLCELL_X1 FILLER_106_179 ();
 FILLCELL_X2 FILLER_106_207 ();
 FILLCELL_X8 FILLER_106_229 ();
 FILLCELL_X8 FILLER_106_244 ();
 FILLCELL_X2 FILLER_106_252 ();
 FILLCELL_X2 FILLER_106_281 ();
 FILLCELL_X1 FILLER_106_290 ();
 FILLCELL_X4 FILLER_106_358 ();
 FILLCELL_X1 FILLER_106_362 ();
 FILLCELL_X8 FILLER_106_370 ();
 FILLCELL_X4 FILLER_106_412 ();
 FILLCELL_X16 FILLER_106_463 ();
 FILLCELL_X2 FILLER_106_479 ();
 FILLCELL_X1 FILLER_106_481 ();
 FILLCELL_X16 FILLER_106_496 ();
 FILLCELL_X8 FILLER_106_519 ();
 FILLCELL_X2 FILLER_106_527 ();
 FILLCELL_X1 FILLER_106_529 ();
 FILLCELL_X2 FILLER_106_534 ();
 FILLCELL_X16 FILLER_106_574 ();
 FILLCELL_X2 FILLER_106_590 ();
 FILLCELL_X1 FILLER_106_592 ();
 FILLCELL_X16 FILLER_106_600 ();
 FILLCELL_X8 FILLER_106_616 ();
 FILLCELL_X4 FILLER_106_624 ();
 FILLCELL_X2 FILLER_106_628 ();
 FILLCELL_X1 FILLER_106_630 ();
 FILLCELL_X4 FILLER_106_632 ();
 FILLCELL_X1 FILLER_106_636 ();
 FILLCELL_X8 FILLER_106_687 ();
 FILLCELL_X4 FILLER_106_695 ();
 FILLCELL_X2 FILLER_106_699 ();
 FILLCELL_X1 FILLER_106_705 ();
 FILLCELL_X1 FILLER_106_714 ();
 FILLCELL_X4 FILLER_106_718 ();
 FILLCELL_X2 FILLER_106_722 ();
 FILLCELL_X2 FILLER_106_745 ();
 FILLCELL_X1 FILLER_106_747 ();
 FILLCELL_X4 FILLER_106_754 ();
 FILLCELL_X1 FILLER_106_758 ();
 FILLCELL_X4 FILLER_106_778 ();
 FILLCELL_X8 FILLER_106_786 ();
 FILLCELL_X4 FILLER_106_794 ();
 FILLCELL_X2 FILLER_106_798 ();
 FILLCELL_X16 FILLER_106_807 ();
 FILLCELL_X4 FILLER_106_823 ();
 FILLCELL_X1 FILLER_106_827 ();
 FILLCELL_X2 FILLER_106_831 ();
 FILLCELL_X4 FILLER_106_841 ();
 FILLCELL_X2 FILLER_106_849 ();
 FILLCELL_X1 FILLER_106_851 ();
 FILLCELL_X8 FILLER_106_857 ();
 FILLCELL_X4 FILLER_106_865 ();
 FILLCELL_X4 FILLER_106_878 ();
 FILLCELL_X2 FILLER_106_895 ();
 FILLCELL_X8 FILLER_106_931 ();
 FILLCELL_X2 FILLER_106_939 ();
 FILLCELL_X2 FILLER_106_948 ();
 FILLCELL_X2 FILLER_106_958 ();
 FILLCELL_X1 FILLER_106_960 ();
 FILLCELL_X1 FILLER_106_965 ();
 FILLCELL_X1 FILLER_106_981 ();
 FILLCELL_X16 FILLER_106_987 ();
 FILLCELL_X4 FILLER_106_1003 ();
 FILLCELL_X1 FILLER_106_1007 ();
 FILLCELL_X8 FILLER_106_1010 ();
 FILLCELL_X2 FILLER_106_1018 ();
 FILLCELL_X1 FILLER_106_1020 ();
 FILLCELL_X8 FILLER_106_1033 ();
 FILLCELL_X4 FILLER_106_1041 ();
 FILLCELL_X2 FILLER_106_1045 ();
 FILLCELL_X8 FILLER_106_1082 ();
 FILLCELL_X2 FILLER_106_1090 ();
 FILLCELL_X1 FILLER_106_1099 ();
 FILLCELL_X1 FILLER_106_1104 ();
 FILLCELL_X1 FILLER_106_1107 ();
 FILLCELL_X4 FILLER_106_1121 ();
 FILLCELL_X1 FILLER_106_1125 ();
 FILLCELL_X4 FILLER_106_1138 ();
 FILLCELL_X1 FILLER_106_1142 ();
 FILLCELL_X8 FILLER_106_1170 ();
 FILLCELL_X4 FILLER_106_1178 ();
 FILLCELL_X1 FILLER_106_1199 ();
 FILLCELL_X1 FILLER_106_1205 ();
 FILLCELL_X1 FILLER_106_1213 ();
 FILLCELL_X4 FILLER_106_1221 ();
 FILLCELL_X1 FILLER_106_1225 ();
 FILLCELL_X1 FILLER_106_1236 ();
 FILLCELL_X1 FILLER_106_1259 ();
 FILLCELL_X2 FILLER_107_1 ();
 FILLCELL_X1 FILLER_107_3 ();
 FILLCELL_X1 FILLER_107_45 ();
 FILLCELL_X1 FILLER_107_53 ();
 FILLCELL_X1 FILLER_107_81 ();
 FILLCELL_X32 FILLER_107_102 ();
 FILLCELL_X4 FILLER_107_141 ();
 FILLCELL_X1 FILLER_107_145 ();
 FILLCELL_X4 FILLER_107_153 ();
 FILLCELL_X4 FILLER_107_178 ();
 FILLCELL_X1 FILLER_107_182 ();
 FILLCELL_X16 FILLER_107_186 ();
 FILLCELL_X1 FILLER_107_202 ();
 FILLCELL_X2 FILLER_107_214 ();
 FILLCELL_X2 FILLER_107_219 ();
 FILLCELL_X1 FILLER_107_221 ();
 FILLCELL_X4 FILLER_107_229 ();
 FILLCELL_X2 FILLER_107_233 ();
 FILLCELL_X8 FILLER_107_262 ();
 FILLCELL_X2 FILLER_107_270 ();
 FILLCELL_X8 FILLER_107_306 ();
 FILLCELL_X8 FILLER_107_349 ();
 FILLCELL_X2 FILLER_107_396 ();
 FILLCELL_X8 FILLER_107_418 ();
 FILLCELL_X4 FILLER_107_426 ();
 FILLCELL_X2 FILLER_107_430 ();
 FILLCELL_X1 FILLER_107_432 ();
 FILLCELL_X1 FILLER_107_440 ();
 FILLCELL_X1 FILLER_107_448 ();
 FILLCELL_X1 FILLER_107_456 ();
 FILLCELL_X4 FILLER_107_477 ();
 FILLCELL_X2 FILLER_107_481 ();
 FILLCELL_X2 FILLER_107_490 ();
 FILLCELL_X4 FILLER_107_512 ();
 FILLCELL_X1 FILLER_107_546 ();
 FILLCELL_X1 FILLER_107_554 ();
 FILLCELL_X8 FILLER_107_558 ();
 FILLCELL_X4 FILLER_107_566 ();
 FILLCELL_X2 FILLER_107_570 ();
 FILLCELL_X8 FILLER_107_579 ();
 FILLCELL_X2 FILLER_107_587 ();
 FILLCELL_X32 FILLER_107_610 ();
 FILLCELL_X32 FILLER_107_642 ();
 FILLCELL_X8 FILLER_107_674 ();
 FILLCELL_X8 FILLER_107_691 ();
 FILLCELL_X2 FILLER_107_699 ();
 FILLCELL_X1 FILLER_107_704 ();
 FILLCELL_X4 FILLER_107_712 ();
 FILLCELL_X2 FILLER_107_716 ();
 FILLCELL_X16 FILLER_107_725 ();
 FILLCELL_X4 FILLER_107_741 ();
 FILLCELL_X1 FILLER_107_745 ();
 FILLCELL_X2 FILLER_107_753 ();
 FILLCELL_X16 FILLER_107_759 ();
 FILLCELL_X4 FILLER_107_775 ();
 FILLCELL_X1 FILLER_107_779 ();
 FILLCELL_X16 FILLER_107_789 ();
 FILLCELL_X4 FILLER_107_805 ();
 FILLCELL_X2 FILLER_107_827 ();
 FILLCELL_X1 FILLER_107_829 ();
 FILLCELL_X8 FILLER_107_835 ();
 FILLCELL_X1 FILLER_107_843 ();
 FILLCELL_X2 FILLER_107_848 ();
 FILLCELL_X1 FILLER_107_850 ();
 FILLCELL_X8 FILLER_107_867 ();
 FILLCELL_X1 FILLER_107_875 ();
 FILLCELL_X4 FILLER_107_930 ();
 FILLCELL_X1 FILLER_107_934 ();
 FILLCELL_X4 FILLER_107_949 ();
 FILLCELL_X1 FILLER_107_953 ();
 FILLCELL_X1 FILLER_107_958 ();
 FILLCELL_X1 FILLER_107_962 ();
 FILLCELL_X2 FILLER_107_997 ();
 FILLCELL_X1 FILLER_107_1002 ();
 FILLCELL_X1 FILLER_107_1028 ();
 FILLCELL_X4 FILLER_107_1051 ();
 FILLCELL_X1 FILLER_107_1055 ();
 FILLCELL_X4 FILLER_107_1060 ();
 FILLCELL_X2 FILLER_107_1064 ();
 FILLCELL_X1 FILLER_107_1098 ();
 FILLCELL_X2 FILLER_107_1104 ();
 FILLCELL_X1 FILLER_107_1106 ();
 FILLCELL_X2 FILLER_107_1125 ();
 FILLCELL_X4 FILLER_107_1134 ();
 FILLCELL_X2 FILLER_107_1138 ();
 FILLCELL_X8 FILLER_107_1145 ();
 FILLCELL_X4 FILLER_107_1153 ();
 FILLCELL_X1 FILLER_107_1157 ();
 FILLCELL_X1 FILLER_107_1195 ();
 FILLCELL_X1 FILLER_107_1201 ();
 FILLCELL_X1 FILLER_107_1212 ();
 FILLCELL_X4 FILLER_107_1235 ();
 FILLCELL_X2 FILLER_107_1244 ();
 FILLCELL_X2 FILLER_107_1253 ();
 FILLCELL_X8 FILLER_108_1 ();
 FILLCELL_X4 FILLER_108_9 ();
 FILLCELL_X1 FILLER_108_13 ();
 FILLCELL_X4 FILLER_108_28 ();
 FILLCELL_X1 FILLER_108_32 ();
 FILLCELL_X2 FILLER_108_40 ();
 FILLCELL_X1 FILLER_108_42 ();
 FILLCELL_X1 FILLER_108_50 ();
 FILLCELL_X8 FILLER_108_58 ();
 FILLCELL_X1 FILLER_108_66 ();
 FILLCELL_X8 FILLER_108_87 ();
 FILLCELL_X2 FILLER_108_95 ();
 FILLCELL_X2 FILLER_108_111 ();
 FILLCELL_X2 FILLER_108_134 ();
 FILLCELL_X1 FILLER_108_136 ();
 FILLCELL_X4 FILLER_108_144 ();
 FILLCELL_X1 FILLER_108_148 ();
 FILLCELL_X4 FILLER_108_169 ();
 FILLCELL_X1 FILLER_108_173 ();
 FILLCELL_X4 FILLER_108_177 ();
 FILLCELL_X2 FILLER_108_195 ();
 FILLCELL_X1 FILLER_108_215 ();
 FILLCELL_X16 FILLER_108_230 ();
 FILLCELL_X1 FILLER_108_246 ();
 FILLCELL_X4 FILLER_108_254 ();
 FILLCELL_X4 FILLER_108_285 ();
 FILLCELL_X2 FILLER_108_289 ();
 FILLCELL_X4 FILLER_108_319 ();
 FILLCELL_X1 FILLER_108_323 ();
 FILLCELL_X2 FILLER_108_331 ();
 FILLCELL_X1 FILLER_108_333 ();
 FILLCELL_X16 FILLER_108_381 ();
 FILLCELL_X4 FILLER_108_397 ();
 FILLCELL_X1 FILLER_108_401 ();
 FILLCELL_X1 FILLER_108_423 ();
 FILLCELL_X8 FILLER_108_450 ();
 FILLCELL_X4 FILLER_108_458 ();
 FILLCELL_X1 FILLER_108_462 ();
 FILLCELL_X1 FILLER_108_490 ();
 FILLCELL_X2 FILLER_108_498 ();
 FILLCELL_X8 FILLER_108_507 ();
 FILLCELL_X2 FILLER_108_515 ();
 FILLCELL_X1 FILLER_108_517 ();
 FILLCELL_X4 FILLER_108_538 ();
 FILLCELL_X1 FILLER_108_542 ();
 FILLCELL_X2 FILLER_108_568 ();
 FILLCELL_X2 FILLER_108_594 ();
 FILLCELL_X1 FILLER_108_603 ();
 FILLCELL_X8 FILLER_108_632 ();
 FILLCELL_X4 FILLER_108_640 ();
 FILLCELL_X2 FILLER_108_644 ();
 FILLCELL_X8 FILLER_108_656 ();
 FILLCELL_X1 FILLER_108_664 ();
 FILLCELL_X16 FILLER_108_676 ();
 FILLCELL_X8 FILLER_108_692 ();
 FILLCELL_X4 FILLER_108_705 ();
 FILLCELL_X1 FILLER_108_709 ();
 FILLCELL_X4 FILLER_108_731 ();
 FILLCELL_X1 FILLER_108_742 ();
 FILLCELL_X2 FILLER_108_746 ();
 FILLCELL_X4 FILLER_108_750 ();
 FILLCELL_X1 FILLER_108_754 ();
 FILLCELL_X2 FILLER_108_759 ();
 FILLCELL_X1 FILLER_108_761 ();
 FILLCELL_X2 FILLER_108_774 ();
 FILLCELL_X4 FILLER_108_781 ();
 FILLCELL_X2 FILLER_108_785 ();
 FILLCELL_X1 FILLER_108_787 ();
 FILLCELL_X1 FILLER_108_791 ();
 FILLCELL_X16 FILLER_108_801 ();
 FILLCELL_X4 FILLER_108_821 ();
 FILLCELL_X16 FILLER_108_829 ();
 FILLCELL_X4 FILLER_108_845 ();
 FILLCELL_X1 FILLER_108_849 ();
 FILLCELL_X8 FILLER_108_853 ();
 FILLCELL_X2 FILLER_108_861 ();
 FILLCELL_X4 FILLER_108_878 ();
 FILLCELL_X2 FILLER_108_882 ();
 FILLCELL_X1 FILLER_108_884 ();
 FILLCELL_X1 FILLER_108_913 ();
 FILLCELL_X2 FILLER_108_924 ();
 FILLCELL_X1 FILLER_108_926 ();
 FILLCELL_X8 FILLER_108_967 ();
 FILLCELL_X2 FILLER_108_995 ();
 FILLCELL_X8 FILLER_108_1008 ();
 FILLCELL_X2 FILLER_108_1016 ();
 FILLCELL_X2 FILLER_108_1062 ();
 FILLCELL_X1 FILLER_108_1064 ();
 FILLCELL_X8 FILLER_108_1069 ();
 FILLCELL_X4 FILLER_108_1077 ();
 FILLCELL_X1 FILLER_108_1102 ();
 FILLCELL_X2 FILLER_108_1114 ();
 FILLCELL_X4 FILLER_108_1139 ();
 FILLCELL_X16 FILLER_108_1161 ();
 FILLCELL_X2 FILLER_108_1177 ();
 FILLCELL_X1 FILLER_108_1179 ();
 FILLCELL_X8 FILLER_108_1187 ();
 FILLCELL_X2 FILLER_108_1195 ();
 FILLCELL_X4 FILLER_108_1204 ();
 FILLCELL_X1 FILLER_108_1208 ();
 FILLCELL_X4 FILLER_108_1216 ();
 FILLCELL_X4 FILLER_108_1223 ();
 FILLCELL_X2 FILLER_108_1227 ();
 FILLCELL_X2 FILLER_108_1239 ();
 FILLCELL_X8 FILLER_109_1 ();
 FILLCELL_X4 FILLER_109_9 ();
 FILLCELL_X1 FILLER_109_40 ();
 FILLCELL_X16 FILLER_109_48 ();
 FILLCELL_X4 FILLER_109_64 ();
 FILLCELL_X2 FILLER_109_102 ();
 FILLCELL_X4 FILLER_109_111 ();
 FILLCELL_X2 FILLER_109_129 ();
 FILLCELL_X1 FILLER_109_131 ();
 FILLCELL_X1 FILLER_109_135 ();
 FILLCELL_X4 FILLER_109_156 ();
 FILLCELL_X1 FILLER_109_160 ();
 FILLCELL_X1 FILLER_109_211 ();
 FILLCELL_X4 FILLER_109_216 ();
 FILLCELL_X1 FILLER_109_220 ();
 FILLCELL_X1 FILLER_109_228 ();
 FILLCELL_X2 FILLER_109_243 ();
 FILLCELL_X1 FILLER_109_245 ();
 FILLCELL_X4 FILLER_109_266 ();
 FILLCELL_X2 FILLER_109_270 ();
 FILLCELL_X1 FILLER_109_272 ();
 FILLCELL_X4 FILLER_109_300 ();
 FILLCELL_X2 FILLER_109_304 ();
 FILLCELL_X8 FILLER_109_320 ();
 FILLCELL_X1 FILLER_109_335 ();
 FILLCELL_X1 FILLER_109_343 ();
 FILLCELL_X1 FILLER_109_351 ();
 FILLCELL_X1 FILLER_109_359 ();
 FILLCELL_X2 FILLER_109_367 ();
 FILLCELL_X1 FILLER_109_369 ();
 FILLCELL_X16 FILLER_109_431 ();
 FILLCELL_X1 FILLER_109_447 ();
 FILLCELL_X16 FILLER_109_452 ();
 FILLCELL_X2 FILLER_109_468 ();
 FILLCELL_X8 FILLER_109_481 ();
 FILLCELL_X4 FILLER_109_489 ();
 FILLCELL_X1 FILLER_109_493 ();
 FILLCELL_X16 FILLER_109_521 ();
 FILLCELL_X4 FILLER_109_537 ();
 FILLCELL_X2 FILLER_109_541 ();
 FILLCELL_X1 FILLER_109_543 ();
 FILLCELL_X8 FILLER_109_578 ();
 FILLCELL_X4 FILLER_109_586 ();
 FILLCELL_X2 FILLER_109_590 ();
 FILLCELL_X4 FILLER_109_599 ();
 FILLCELL_X2 FILLER_109_603 ();
 FILLCELL_X8 FILLER_109_612 ();
 FILLCELL_X4 FILLER_109_620 ();
 FILLCELL_X8 FILLER_109_634 ();
 FILLCELL_X4 FILLER_109_642 ();
 FILLCELL_X2 FILLER_109_666 ();
 FILLCELL_X1 FILLER_109_688 ();
 FILLCELL_X16 FILLER_109_694 ();
 FILLCELL_X8 FILLER_109_710 ();
 FILLCELL_X4 FILLER_109_718 ();
 FILLCELL_X2 FILLER_109_722 ();
 FILLCELL_X1 FILLER_109_724 ();
 FILLCELL_X8 FILLER_109_734 ();
 FILLCELL_X2 FILLER_109_742 ();
 FILLCELL_X8 FILLER_109_753 ();
 FILLCELL_X4 FILLER_109_761 ();
 FILLCELL_X2 FILLER_109_765 ();
 FILLCELL_X2 FILLER_109_770 ();
 FILLCELL_X1 FILLER_109_772 ();
 FILLCELL_X2 FILLER_109_789 ();
 FILLCELL_X4 FILLER_109_813 ();
 FILLCELL_X1 FILLER_109_817 ();
 FILLCELL_X4 FILLER_109_822 ();
 FILLCELL_X1 FILLER_109_844 ();
 FILLCELL_X8 FILLER_109_852 ();
 FILLCELL_X4 FILLER_109_860 ();
 FILLCELL_X2 FILLER_109_864 ();
 FILLCELL_X1 FILLER_109_866 ();
 FILLCELL_X4 FILLER_109_876 ();
 FILLCELL_X1 FILLER_109_880 ();
 FILLCELL_X8 FILLER_109_895 ();
 FILLCELL_X4 FILLER_109_903 ();
 FILLCELL_X16 FILLER_109_914 ();
 FILLCELL_X8 FILLER_109_930 ();
 FILLCELL_X4 FILLER_109_938 ();
 FILLCELL_X2 FILLER_109_942 ();
 FILLCELL_X1 FILLER_109_944 ();
 FILLCELL_X4 FILLER_109_959 ();
 FILLCELL_X8 FILLER_109_977 ();
 FILLCELL_X2 FILLER_109_985 ();
 FILLCELL_X1 FILLER_109_987 ();
 FILLCELL_X8 FILLER_109_996 ();
 FILLCELL_X2 FILLER_109_1004 ();
 FILLCELL_X1 FILLER_109_1006 ();
 FILLCELL_X8 FILLER_109_1028 ();
 FILLCELL_X2 FILLER_109_1036 ();
 FILLCELL_X4 FILLER_109_1062 ();
 FILLCELL_X2 FILLER_109_1066 ();
 FILLCELL_X1 FILLER_109_1068 ();
 FILLCELL_X1 FILLER_109_1086 ();
 FILLCELL_X2 FILLER_109_1098 ();
 FILLCELL_X8 FILLER_109_1104 ();
 FILLCELL_X1 FILLER_109_1115 ();
 FILLCELL_X2 FILLER_109_1122 ();
 FILLCELL_X4 FILLER_109_1137 ();
 FILLCELL_X1 FILLER_109_1141 ();
 FILLCELL_X2 FILLER_109_1147 ();
 FILLCELL_X1 FILLER_109_1149 ();
 FILLCELL_X16 FILLER_109_1154 ();
 FILLCELL_X2 FILLER_109_1192 ();
 FILLCELL_X1 FILLER_109_1194 ();
 FILLCELL_X1 FILLER_109_1224 ();
 FILLCELL_X2 FILLER_109_1249 ();
 FILLCELL_X2 FILLER_109_1258 ();
 FILLCELL_X1 FILLER_110_1 ();
 FILLCELL_X1 FILLER_110_22 ();
 FILLCELL_X1 FILLER_110_30 ();
 FILLCELL_X1 FILLER_110_38 ();
 FILLCELL_X4 FILLER_110_53 ();
 FILLCELL_X8 FILLER_110_84 ();
 FILLCELL_X1 FILLER_110_92 ();
 FILLCELL_X8 FILLER_110_100 ();
 FILLCELL_X1 FILLER_110_108 ();
 FILLCELL_X4 FILLER_110_123 ();
 FILLCELL_X2 FILLER_110_127 ();
 FILLCELL_X4 FILLER_110_156 ();
 FILLCELL_X8 FILLER_110_167 ();
 FILLCELL_X2 FILLER_110_175 ();
 FILLCELL_X1 FILLER_110_177 ();
 FILLCELL_X1 FILLER_110_182 ();
 FILLCELL_X8 FILLER_110_190 ();
 FILLCELL_X8 FILLER_110_212 ();
 FILLCELL_X8 FILLER_110_222 ();
 FILLCELL_X2 FILLER_110_230 ();
 FILLCELL_X1 FILLER_110_232 ();
 FILLCELL_X4 FILLER_110_267 ();
 FILLCELL_X2 FILLER_110_271 ();
 FILLCELL_X1 FILLER_110_273 ();
 FILLCELL_X4 FILLER_110_308 ();
 FILLCELL_X2 FILLER_110_319 ();
 FILLCELL_X2 FILLER_110_324 ();
 FILLCELL_X1 FILLER_110_326 ();
 FILLCELL_X2 FILLER_110_347 ();
 FILLCELL_X4 FILLER_110_356 ();
 FILLCELL_X4 FILLER_110_367 ();
 FILLCELL_X2 FILLER_110_378 ();
 FILLCELL_X1 FILLER_110_380 ();
 FILLCELL_X1 FILLER_110_396 ();
 FILLCELL_X4 FILLER_110_404 ();
 FILLCELL_X4 FILLER_110_442 ();
 FILLCELL_X4 FILLER_110_453 ();
 FILLCELL_X1 FILLER_110_457 ();
 FILLCELL_X4 FILLER_110_501 ();
 FILLCELL_X2 FILLER_110_505 ();
 FILLCELL_X8 FILLER_110_555 ();
 FILLCELL_X4 FILLER_110_563 ();
 FILLCELL_X1 FILLER_110_598 ();
 FILLCELL_X2 FILLER_110_606 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X2 FILLER_110_637 ();
 FILLCELL_X2 FILLER_110_659 ();
 FILLCELL_X2 FILLER_110_668 ();
 FILLCELL_X16 FILLER_110_697 ();
 FILLCELL_X2 FILLER_110_713 ();
 FILLCELL_X1 FILLER_110_715 ();
 FILLCELL_X16 FILLER_110_723 ();
 FILLCELL_X4 FILLER_110_739 ();
 FILLCELL_X16 FILLER_110_750 ();
 FILLCELL_X4 FILLER_110_766 ();
 FILLCELL_X8 FILLER_110_774 ();
 FILLCELL_X4 FILLER_110_782 ();
 FILLCELL_X16 FILLER_110_793 ();
 FILLCELL_X4 FILLER_110_809 ();
 FILLCELL_X2 FILLER_110_813 ();
 FILLCELL_X1 FILLER_110_815 ();
 FILLCELL_X32 FILLER_110_839 ();
 FILLCELL_X2 FILLER_110_871 ();
 FILLCELL_X1 FILLER_110_879 ();
 FILLCELL_X8 FILLER_110_894 ();
 FILLCELL_X1 FILLER_110_902 ();
 FILLCELL_X8 FILLER_110_924 ();
 FILLCELL_X1 FILLER_110_932 ();
 FILLCELL_X8 FILLER_110_961 ();
 FILLCELL_X1 FILLER_110_1005 ();
 FILLCELL_X1 FILLER_110_1008 ();
 FILLCELL_X2 FILLER_110_1036 ();
 FILLCELL_X1 FILLER_110_1038 ();
 FILLCELL_X4 FILLER_110_1050 ();
 FILLCELL_X8 FILLER_110_1058 ();
 FILLCELL_X2 FILLER_110_1066 ();
 FILLCELL_X2 FILLER_110_1093 ();
 FILLCELL_X1 FILLER_110_1095 ();
 FILLCELL_X4 FILLER_110_1099 ();
 FILLCELL_X1 FILLER_110_1106 ();
 FILLCELL_X1 FILLER_110_1118 ();
 FILLCELL_X4 FILLER_110_1123 ();
 FILLCELL_X1 FILLER_110_1127 ();
 FILLCELL_X2 FILLER_110_1139 ();
 FILLCELL_X2 FILLER_110_1145 ();
 FILLCELL_X1 FILLER_110_1147 ();
 FILLCELL_X16 FILLER_110_1158 ();
 FILLCELL_X4 FILLER_110_1174 ();
 FILLCELL_X2 FILLER_110_1178 ();
 FILLCELL_X4 FILLER_110_1191 ();
 FILLCELL_X2 FILLER_110_1195 ();
 FILLCELL_X2 FILLER_110_1202 ();
 FILLCELL_X4 FILLER_110_1206 ();
 FILLCELL_X1 FILLER_110_1210 ();
 FILLCELL_X4 FILLER_110_1241 ();
 FILLCELL_X2 FILLER_110_1258 ();
 FILLCELL_X4 FILLER_111_1 ();
 FILLCELL_X2 FILLER_111_5 ();
 FILLCELL_X8 FILLER_111_48 ();
 FILLCELL_X4 FILLER_111_56 ();
 FILLCELL_X2 FILLER_111_60 ();
 FILLCELL_X2 FILLER_111_109 ();
 FILLCELL_X8 FILLER_111_132 ();
 FILLCELL_X4 FILLER_111_140 ();
 FILLCELL_X2 FILLER_111_144 ();
 FILLCELL_X4 FILLER_111_182 ();
 FILLCELL_X2 FILLER_111_197 ();
 FILLCELL_X2 FILLER_111_226 ();
 FILLCELL_X16 FILLER_111_276 ();
 FILLCELL_X1 FILLER_111_292 ();
 FILLCELL_X8 FILLER_111_312 ();
 FILLCELL_X1 FILLER_111_320 ();
 FILLCELL_X8 FILLER_111_335 ();
 FILLCELL_X2 FILLER_111_343 ();
 FILLCELL_X1 FILLER_111_345 ();
 FILLCELL_X1 FILLER_111_353 ();
 FILLCELL_X2 FILLER_111_361 ();
 FILLCELL_X1 FILLER_111_383 ();
 FILLCELL_X8 FILLER_111_404 ();
 FILLCELL_X1 FILLER_111_412 ();
 FILLCELL_X8 FILLER_111_420 ();
 FILLCELL_X4 FILLER_111_428 ();
 FILLCELL_X1 FILLER_111_432 ();
 FILLCELL_X8 FILLER_111_460 ();
 FILLCELL_X2 FILLER_111_475 ();
 FILLCELL_X1 FILLER_111_477 ();
 FILLCELL_X4 FILLER_111_540 ();
 FILLCELL_X2 FILLER_111_544 ();
 FILLCELL_X8 FILLER_111_553 ();
 FILLCELL_X4 FILLER_111_582 ();
 FILLCELL_X2 FILLER_111_586 ();
 FILLCELL_X1 FILLER_111_588 ();
 FILLCELL_X4 FILLER_111_618 ();
 FILLCELL_X16 FILLER_111_642 ();
 FILLCELL_X4 FILLER_111_665 ();
 FILLCELL_X2 FILLER_111_669 ();
 FILLCELL_X1 FILLER_111_671 ();
 FILLCELL_X4 FILLER_111_685 ();
 FILLCELL_X8 FILLER_111_700 ();
 FILLCELL_X4 FILLER_111_708 ();
 FILLCELL_X2 FILLER_111_712 ();
 FILLCELL_X2 FILLER_111_716 ();
 FILLCELL_X1 FILLER_111_718 ();
 FILLCELL_X8 FILLER_111_728 ();
 FILLCELL_X1 FILLER_111_736 ();
 FILLCELL_X8 FILLER_111_750 ();
 FILLCELL_X4 FILLER_111_762 ();
 FILLCELL_X1 FILLER_111_766 ();
 FILLCELL_X16 FILLER_111_774 ();
 FILLCELL_X2 FILLER_111_790 ();
 FILLCELL_X4 FILLER_111_807 ();
 FILLCELL_X1 FILLER_111_811 ();
 FILLCELL_X4 FILLER_111_816 ();
 FILLCELL_X2 FILLER_111_820 ();
 FILLCELL_X1 FILLER_111_838 ();
 FILLCELL_X8 FILLER_111_842 ();
 FILLCELL_X2 FILLER_111_850 ();
 FILLCELL_X1 FILLER_111_855 ();
 FILLCELL_X16 FILLER_111_865 ();
 FILLCELL_X4 FILLER_111_881 ();
 FILLCELL_X2 FILLER_111_885 ();
 FILLCELL_X1 FILLER_111_887 ();
 FILLCELL_X8 FILLER_111_908 ();
 FILLCELL_X2 FILLER_111_916 ();
 FILLCELL_X1 FILLER_111_918 ();
 FILLCELL_X8 FILLER_111_939 ();
 FILLCELL_X4 FILLER_111_947 ();
 FILLCELL_X1 FILLER_111_951 ();
 FILLCELL_X2 FILLER_111_957 ();
 FILLCELL_X4 FILLER_111_964 ();
 FILLCELL_X4 FILLER_111_975 ();
 FILLCELL_X2 FILLER_111_986 ();
 FILLCELL_X1 FILLER_111_988 ();
 FILLCELL_X4 FILLER_111_1005 ();
 FILLCELL_X1 FILLER_111_1009 ();
 FILLCELL_X4 FILLER_111_1016 ();
 FILLCELL_X1 FILLER_111_1020 ();
 FILLCELL_X16 FILLER_111_1025 ();
 FILLCELL_X2 FILLER_111_1041 ();
 FILLCELL_X1 FILLER_111_1056 ();
 FILLCELL_X4 FILLER_111_1069 ();
 FILLCELL_X2 FILLER_111_1073 ();
 FILLCELL_X1 FILLER_111_1075 ();
 FILLCELL_X1 FILLER_111_1086 ();
 FILLCELL_X1 FILLER_111_1094 ();
 FILLCELL_X1 FILLER_111_1102 ();
 FILLCELL_X1 FILLER_111_1110 ();
 FILLCELL_X1 FILLER_111_1122 ();
 FILLCELL_X1 FILLER_111_1134 ();
 FILLCELL_X2 FILLER_111_1146 ();
 FILLCELL_X16 FILLER_111_1162 ();
 FILLCELL_X2 FILLER_111_1178 ();
 FILLCELL_X1 FILLER_111_1180 ();
 FILLCELL_X1 FILLER_111_1186 ();
 FILLCELL_X1 FILLER_111_1191 ();
 FILLCELL_X4 FILLER_111_1212 ();
 FILLCELL_X1 FILLER_111_1216 ();
 FILLCELL_X1 FILLER_111_1222 ();
 FILLCELL_X2 FILLER_111_1225 ();
 FILLCELL_X2 FILLER_111_1229 ();
 FILLCELL_X2 FILLER_111_1249 ();
 FILLCELL_X1 FILLER_111_1251 ();
 FILLCELL_X1 FILLER_111_1255 ();
 FILLCELL_X16 FILLER_112_1 ();
 FILLCELL_X8 FILLER_112_17 ();
 FILLCELL_X4 FILLER_112_25 ();
 FILLCELL_X8 FILLER_112_56 ();
 FILLCELL_X8 FILLER_112_69 ();
 FILLCELL_X2 FILLER_112_77 ();
 FILLCELL_X4 FILLER_112_86 ();
 FILLCELL_X1 FILLER_112_110 ();
 FILLCELL_X4 FILLER_112_118 ();
 FILLCELL_X1 FILLER_112_122 ();
 FILLCELL_X16 FILLER_112_150 ();
 FILLCELL_X16 FILLER_112_203 ();
 FILLCELL_X8 FILLER_112_219 ();
 FILLCELL_X4 FILLER_112_227 ();
 FILLCELL_X1 FILLER_112_253 ();
 FILLCELL_X16 FILLER_112_275 ();
 FILLCELL_X8 FILLER_112_291 ();
 FILLCELL_X2 FILLER_112_299 ();
 FILLCELL_X4 FILLER_112_313 ();
 FILLCELL_X16 FILLER_112_351 ();
 FILLCELL_X4 FILLER_112_367 ();
 FILLCELL_X1 FILLER_112_371 ();
 FILLCELL_X4 FILLER_112_399 ();
 FILLCELL_X2 FILLER_112_403 ();
 FILLCELL_X1 FILLER_112_405 ();
 FILLCELL_X2 FILLER_112_413 ();
 FILLCELL_X1 FILLER_112_449 ();
 FILLCELL_X16 FILLER_112_457 ();
 FILLCELL_X1 FILLER_112_473 ();
 FILLCELL_X2 FILLER_112_479 ();
 FILLCELL_X8 FILLER_112_488 ();
 FILLCELL_X8 FILLER_112_503 ();
 FILLCELL_X1 FILLER_112_511 ();
 FILLCELL_X2 FILLER_112_539 ();
 FILLCELL_X1 FILLER_112_541 ();
 FILLCELL_X1 FILLER_112_569 ();
 FILLCELL_X4 FILLER_112_604 ();
 FILLCELL_X1 FILLER_112_608 ();
 FILLCELL_X1 FILLER_112_630 ();
 FILLCELL_X8 FILLER_112_634 ();
 FILLCELL_X1 FILLER_112_642 ();
 FILLCELL_X4 FILLER_112_663 ();
 FILLCELL_X8 FILLER_112_671 ();
 FILLCELL_X2 FILLER_112_679 ();
 FILLCELL_X1 FILLER_112_681 ();
 FILLCELL_X4 FILLER_112_687 ();
 FILLCELL_X1 FILLER_112_691 ();
 FILLCELL_X8 FILLER_112_699 ();
 FILLCELL_X8 FILLER_112_740 ();
 FILLCELL_X2 FILLER_112_768 ();
 FILLCELL_X1 FILLER_112_805 ();
 FILLCELL_X2 FILLER_112_831 ();
 FILLCELL_X1 FILLER_112_833 ();
 FILLCELL_X1 FILLER_112_837 ();
 FILLCELL_X4 FILLER_112_841 ();
 FILLCELL_X2 FILLER_112_845 ();
 FILLCELL_X16 FILLER_112_851 ();
 FILLCELL_X1 FILLER_112_867 ();
 FILLCELL_X4 FILLER_112_873 ();
 FILLCELL_X8 FILLER_112_880 ();
 FILLCELL_X4 FILLER_112_888 ();
 FILLCELL_X2 FILLER_112_892 ();
 FILLCELL_X8 FILLER_112_921 ();
 FILLCELL_X4 FILLER_112_929 ();
 FILLCELL_X1 FILLER_112_933 ();
 FILLCELL_X1 FILLER_112_948 ();
 FILLCELL_X8 FILLER_112_989 ();
 FILLCELL_X4 FILLER_112_997 ();
 FILLCELL_X2 FILLER_112_1001 ();
 FILLCELL_X1 FILLER_112_1010 ();
 FILLCELL_X4 FILLER_112_1019 ();
 FILLCELL_X2 FILLER_112_1023 ();
 FILLCELL_X1 FILLER_112_1025 ();
 FILLCELL_X32 FILLER_112_1030 ();
 FILLCELL_X2 FILLER_112_1073 ();
 FILLCELL_X1 FILLER_112_1090 ();
 FILLCELL_X4 FILLER_112_1098 ();
 FILLCELL_X1 FILLER_112_1102 ();
 FILLCELL_X4 FILLER_112_1113 ();
 FILLCELL_X4 FILLER_112_1125 ();
 FILLCELL_X2 FILLER_112_1129 ();
 FILLCELL_X4 FILLER_112_1137 ();
 FILLCELL_X1 FILLER_112_1141 ();
 FILLCELL_X2 FILLER_112_1145 ();
 FILLCELL_X1 FILLER_112_1147 ();
 FILLCELL_X4 FILLER_112_1203 ();
 FILLCELL_X1 FILLER_112_1217 ();
 FILLCELL_X1 FILLER_112_1223 ();
 FILLCELL_X16 FILLER_113_1 ();
 FILLCELL_X8 FILLER_113_17 ();
 FILLCELL_X4 FILLER_113_25 ();
 FILLCELL_X1 FILLER_113_29 ();
 FILLCELL_X16 FILLER_113_50 ();
 FILLCELL_X4 FILLER_113_66 ();
 FILLCELL_X1 FILLER_113_70 ();
 FILLCELL_X4 FILLER_113_98 ();
 FILLCELL_X2 FILLER_113_102 ();
 FILLCELL_X1 FILLER_113_104 ();
 FILLCELL_X2 FILLER_113_119 ();
 FILLCELL_X4 FILLER_113_148 ();
 FILLCELL_X2 FILLER_113_152 ();
 FILLCELL_X8 FILLER_113_174 ();
 FILLCELL_X8 FILLER_113_189 ();
 FILLCELL_X4 FILLER_113_204 ();
 FILLCELL_X2 FILLER_113_208 ();
 FILLCELL_X16 FILLER_113_217 ();
 FILLCELL_X1 FILLER_113_274 ();
 FILLCELL_X2 FILLER_113_282 ();
 FILLCELL_X4 FILLER_113_311 ();
 FILLCELL_X8 FILLER_113_322 ();
 FILLCELL_X4 FILLER_113_330 ();
 FILLCELL_X1 FILLER_113_334 ();
 FILLCELL_X8 FILLER_113_369 ();
 FILLCELL_X1 FILLER_113_377 ();
 FILLCELL_X8 FILLER_113_385 ();
 FILLCELL_X4 FILLER_113_393 ();
 FILLCELL_X2 FILLER_113_397 ();
 FILLCELL_X1 FILLER_113_406 ();
 FILLCELL_X8 FILLER_113_414 ();
 FILLCELL_X2 FILLER_113_422 ();
 FILLCELL_X1 FILLER_113_424 ();
 FILLCELL_X1 FILLER_113_427 ();
 FILLCELL_X2 FILLER_113_433 ();
 FILLCELL_X2 FILLER_113_442 ();
 FILLCELL_X2 FILLER_113_464 ();
 FILLCELL_X1 FILLER_113_466 ();
 FILLCELL_X4 FILLER_113_487 ();
 FILLCELL_X8 FILLER_113_518 ();
 FILLCELL_X1 FILLER_113_533 ();
 FILLCELL_X8 FILLER_113_541 ();
 FILLCELL_X2 FILLER_113_549 ();
 FILLCELL_X2 FILLER_113_558 ();
 FILLCELL_X1 FILLER_113_560 ();
 FILLCELL_X2 FILLER_113_588 ();
 FILLCELL_X16 FILLER_113_621 ();
 FILLCELL_X8 FILLER_113_637 ();
 FILLCELL_X1 FILLER_113_652 ();
 FILLCELL_X1 FILLER_113_672 ();
 FILLCELL_X1 FILLER_113_692 ();
 FILLCELL_X2 FILLER_113_709 ();
 FILLCELL_X8 FILLER_113_714 ();
 FILLCELL_X16 FILLER_113_742 ();
 FILLCELL_X1 FILLER_113_758 ();
 FILLCELL_X8 FILLER_113_776 ();
 FILLCELL_X2 FILLER_113_784 ();
 FILLCELL_X4 FILLER_113_799 ();
 FILLCELL_X2 FILLER_113_803 ();
 FILLCELL_X1 FILLER_113_805 ();
 FILLCELL_X8 FILLER_113_841 ();
 FILLCELL_X16 FILLER_113_880 ();
 FILLCELL_X4 FILLER_113_896 ();
 FILLCELL_X2 FILLER_113_900 ();
 FILLCELL_X1 FILLER_113_909 ();
 FILLCELL_X2 FILLER_113_917 ();
 FILLCELL_X16 FILLER_113_953 ();
 FILLCELL_X2 FILLER_113_969 ();
 FILLCELL_X4 FILLER_113_994 ();
 FILLCELL_X1 FILLER_113_998 ();
 FILLCELL_X4 FILLER_113_1059 ();
 FILLCELL_X1 FILLER_113_1083 ();
 FILLCELL_X4 FILLER_113_1096 ();
 FILLCELL_X2 FILLER_113_1100 ();
 FILLCELL_X1 FILLER_113_1102 ();
 FILLCELL_X1 FILLER_113_1111 ();
 FILLCELL_X1 FILLER_113_1115 ();
 FILLCELL_X1 FILLER_113_1130 ();
 FILLCELL_X1 FILLER_113_1142 ();
 FILLCELL_X1 FILLER_113_1147 ();
 FILLCELL_X8 FILLER_113_1179 ();
 FILLCELL_X2 FILLER_113_1187 ();
 FILLCELL_X1 FILLER_113_1189 ();
 FILLCELL_X2 FILLER_113_1207 ();
 FILLCELL_X1 FILLER_113_1209 ();
 FILLCELL_X4 FILLER_113_1232 ();
 FILLCELL_X1 FILLER_113_1256 ();
 FILLCELL_X8 FILLER_114_1 ();
 FILLCELL_X4 FILLER_114_9 ();
 FILLCELL_X2 FILLER_114_13 ();
 FILLCELL_X1 FILLER_114_15 ();
 FILLCELL_X1 FILLER_114_43 ();
 FILLCELL_X4 FILLER_114_51 ();
 FILLCELL_X1 FILLER_114_55 ();
 FILLCELL_X1 FILLER_114_103 ();
 FILLCELL_X4 FILLER_114_132 ();
 FILLCELL_X2 FILLER_114_136 ();
 FILLCELL_X8 FILLER_114_166 ();
 FILLCELL_X4 FILLER_114_174 ();
 FILLCELL_X1 FILLER_114_178 ();
 FILLCELL_X2 FILLER_114_222 ();
 FILLCELL_X8 FILLER_114_272 ();
 FILLCELL_X2 FILLER_114_280 ();
 FILLCELL_X16 FILLER_114_309 ();
 FILLCELL_X2 FILLER_114_325 ();
 FILLCELL_X1 FILLER_114_327 ();
 FILLCELL_X4 FILLER_114_335 ();
 FILLCELL_X2 FILLER_114_339 ();
 FILLCELL_X1 FILLER_114_341 ();
 FILLCELL_X2 FILLER_114_356 ();
 FILLCELL_X1 FILLER_114_358 ();
 FILLCELL_X2 FILLER_114_399 ();
 FILLCELL_X1 FILLER_114_401 ();
 FILLCELL_X4 FILLER_114_435 ();
 FILLCELL_X2 FILLER_114_446 ();
 FILLCELL_X1 FILLER_114_448 ();
 FILLCELL_X2 FILLER_114_462 ();
 FILLCELL_X2 FILLER_114_481 ();
 FILLCELL_X16 FILLER_114_510 ();
 FILLCELL_X4 FILLER_114_526 ();
 FILLCELL_X2 FILLER_114_530 ();
 FILLCELL_X4 FILLER_114_580 ();
 FILLCELL_X2 FILLER_114_584 ();
 FILLCELL_X4 FILLER_114_593 ();
 FILLCELL_X2 FILLER_114_597 ();
 FILLCELL_X1 FILLER_114_609 ();
 FILLCELL_X1 FILLER_114_630 ();
 FILLCELL_X1 FILLER_114_652 ();
 FILLCELL_X1 FILLER_114_660 ();
 FILLCELL_X2 FILLER_114_674 ();
 FILLCELL_X1 FILLER_114_676 ();
 FILLCELL_X2 FILLER_114_701 ();
 FILLCELL_X4 FILLER_114_710 ();
 FILLCELL_X1 FILLER_114_714 ();
 FILLCELL_X8 FILLER_114_729 ();
 FILLCELL_X1 FILLER_114_737 ();
 FILLCELL_X4 FILLER_114_751 ();
 FILLCELL_X16 FILLER_114_759 ();
 FILLCELL_X4 FILLER_114_775 ();
 FILLCELL_X2 FILLER_114_779 ();
 FILLCELL_X2 FILLER_114_796 ();
 FILLCELL_X1 FILLER_114_798 ();
 FILLCELL_X16 FILLER_114_823 ();
 FILLCELL_X8 FILLER_114_839 ();
 FILLCELL_X4 FILLER_114_847 ();
 FILLCELL_X2 FILLER_114_851 ();
 FILLCELL_X4 FILLER_114_856 ();
 FILLCELL_X2 FILLER_114_860 ();
 FILLCELL_X16 FILLER_114_866 ();
 FILLCELL_X2 FILLER_114_882 ();
 FILLCELL_X4 FILLER_114_947 ();
 FILLCELL_X2 FILLER_114_951 ();
 FILLCELL_X1 FILLER_114_953 ();
 FILLCELL_X2 FILLER_114_964 ();
 FILLCELL_X8 FILLER_114_973 ();
 FILLCELL_X1 FILLER_114_981 ();
 FILLCELL_X2 FILLER_114_987 ();
 FILLCELL_X16 FILLER_114_992 ();
 FILLCELL_X2 FILLER_114_1008 ();
 FILLCELL_X1 FILLER_114_1010 ();
 FILLCELL_X4 FILLER_114_1020 ();
 FILLCELL_X2 FILLER_114_1024 ();
 FILLCELL_X2 FILLER_114_1038 ();
 FILLCELL_X1 FILLER_114_1040 ();
 FILLCELL_X2 FILLER_114_1069 ();
 FILLCELL_X1 FILLER_114_1071 ();
 FILLCELL_X4 FILLER_114_1076 ();
 FILLCELL_X2 FILLER_114_1080 ();
 FILLCELL_X1 FILLER_114_1082 ();
 FILLCELL_X2 FILLER_114_1094 ();
 FILLCELL_X1 FILLER_114_1096 ();
 FILLCELL_X1 FILLER_114_1115 ();
 FILLCELL_X2 FILLER_114_1120 ();
 FILLCELL_X8 FILLER_114_1154 ();
 FILLCELL_X2 FILLER_114_1162 ();
 FILLCELL_X4 FILLER_114_1171 ();
 FILLCELL_X1 FILLER_114_1187 ();
 FILLCELL_X4 FILLER_114_1208 ();
 FILLCELL_X1 FILLER_114_1212 ();
 FILLCELL_X2 FILLER_114_1223 ();
 FILLCELL_X1 FILLER_114_1225 ();
 FILLCELL_X4 FILLER_114_1254 ();
 FILLCELL_X2 FILLER_114_1258 ();
 FILLCELL_X2 FILLER_115_28 ();
 FILLCELL_X1 FILLER_115_30 ();
 FILLCELL_X1 FILLER_115_38 ();
 FILLCELL_X2 FILLER_115_53 ();
 FILLCELL_X1 FILLER_115_55 ();
 FILLCELL_X2 FILLER_115_63 ();
 FILLCELL_X1 FILLER_115_65 ();
 FILLCELL_X2 FILLER_115_86 ();
 FILLCELL_X1 FILLER_115_88 ();
 FILLCELL_X8 FILLER_115_96 ();
 FILLCELL_X4 FILLER_115_111 ();
 FILLCELL_X2 FILLER_115_115 ();
 FILLCELL_X16 FILLER_115_161 ();
 FILLCELL_X8 FILLER_115_177 ();
 FILLCELL_X2 FILLER_115_185 ();
 FILLCELL_X4 FILLER_115_202 ();
 FILLCELL_X1 FILLER_115_206 ();
 FILLCELL_X4 FILLER_115_225 ();
 FILLCELL_X1 FILLER_115_229 ();
 FILLCELL_X4 FILLER_115_250 ();
 FILLCELL_X2 FILLER_115_254 ();
 FILLCELL_X8 FILLER_115_303 ();
 FILLCELL_X2 FILLER_115_311 ();
 FILLCELL_X1 FILLER_115_313 ();
 FILLCELL_X8 FILLER_115_327 ();
 FILLCELL_X2 FILLER_115_335 ();
 FILLCELL_X1 FILLER_115_337 ();
 FILLCELL_X2 FILLER_115_345 ();
 FILLCELL_X1 FILLER_115_347 ();
 FILLCELL_X8 FILLER_115_369 ();
 FILLCELL_X4 FILLER_115_384 ();
 FILLCELL_X8 FILLER_115_413 ();
 FILLCELL_X4 FILLER_115_421 ();
 FILLCELL_X2 FILLER_115_425 ();
 FILLCELL_X1 FILLER_115_427 ();
 FILLCELL_X4 FILLER_115_439 ();
 FILLCELL_X8 FILLER_115_457 ();
 FILLCELL_X2 FILLER_115_465 ();
 FILLCELL_X1 FILLER_115_467 ();
 FILLCELL_X1 FILLER_115_502 ();
 FILLCELL_X4 FILLER_115_537 ();
 FILLCELL_X4 FILLER_115_544 ();
 FILLCELL_X2 FILLER_115_548 ();
 FILLCELL_X1 FILLER_115_550 ();
 FILLCELL_X2 FILLER_115_623 ();
 FILLCELL_X8 FILLER_115_638 ();
 FILLCELL_X4 FILLER_115_646 ();
 FILLCELL_X2 FILLER_115_650 ();
 FILLCELL_X4 FILLER_115_686 ();
 FILLCELL_X2 FILLER_115_690 ();
 FILLCELL_X2 FILLER_115_696 ();
 FILLCELL_X1 FILLER_115_710 ();
 FILLCELL_X2 FILLER_115_724 ();
 FILLCELL_X1 FILLER_115_726 ();
 FILLCELL_X2 FILLER_115_731 ();
 FILLCELL_X8 FILLER_115_742 ();
 FILLCELL_X1 FILLER_115_750 ();
 FILLCELL_X1 FILLER_115_769 ();
 FILLCELL_X4 FILLER_115_778 ();
 FILLCELL_X1 FILLER_115_782 ();
 FILLCELL_X16 FILLER_115_787 ();
 FILLCELL_X4 FILLER_115_803 ();
 FILLCELL_X2 FILLER_115_807 ();
 FILLCELL_X2 FILLER_115_826 ();
 FILLCELL_X2 FILLER_115_860 ();
 FILLCELL_X4 FILLER_115_869 ();
 FILLCELL_X1 FILLER_115_873 ();
 FILLCELL_X2 FILLER_115_876 ();
 FILLCELL_X2 FILLER_115_898 ();
 FILLCELL_X16 FILLER_115_907 ();
 FILLCELL_X1 FILLER_115_930 ();
 FILLCELL_X1 FILLER_115_951 ();
 FILLCELL_X1 FILLER_115_974 ();
 FILLCELL_X1 FILLER_115_982 ();
 FILLCELL_X2 FILLER_115_987 ();
 FILLCELL_X1 FILLER_115_1007 ();
 FILLCELL_X2 FILLER_115_1013 ();
 FILLCELL_X16 FILLER_115_1019 ();
 FILLCELL_X4 FILLER_115_1035 ();
 FILLCELL_X2 FILLER_115_1039 ();
 FILLCELL_X1 FILLER_115_1041 ();
 FILLCELL_X1 FILLER_115_1070 ();
 FILLCELL_X4 FILLER_115_1078 ();
 FILLCELL_X4 FILLER_115_1100 ();
 FILLCELL_X1 FILLER_115_1115 ();
 FILLCELL_X2 FILLER_115_1140 ();
 FILLCELL_X16 FILLER_115_1145 ();
 FILLCELL_X1 FILLER_115_1161 ();
 FILLCELL_X1 FILLER_115_1169 ();
 FILLCELL_X8 FILLER_115_1190 ();
 FILLCELL_X4 FILLER_115_1198 ();
 FILLCELL_X4 FILLER_115_1209 ();
 FILLCELL_X1 FILLER_115_1213 ();
 FILLCELL_X4 FILLER_115_1234 ();
 FILLCELL_X2 FILLER_115_1249 ();
 FILLCELL_X2 FILLER_115_1254 ();
 FILLCELL_X1 FILLER_115_1256 ();
 FILLCELL_X8 FILLER_116_1 ();
 FILLCELL_X4 FILLER_116_9 ();
 FILLCELL_X1 FILLER_116_13 ();
 FILLCELL_X16 FILLER_116_48 ();
 FILLCELL_X32 FILLER_116_111 ();
 FILLCELL_X1 FILLER_116_150 ();
 FILLCELL_X1 FILLER_116_154 ();
 FILLCELL_X2 FILLER_116_163 ();
 FILLCELL_X8 FILLER_116_194 ();
 FILLCELL_X4 FILLER_116_212 ();
 FILLCELL_X8 FILLER_116_230 ();
 FILLCELL_X4 FILLER_116_238 ();
 FILLCELL_X1 FILLER_116_242 ();
 FILLCELL_X1 FILLER_116_270 ();
 FILLCELL_X4 FILLER_116_285 ();
 FILLCELL_X1 FILLER_116_289 ();
 FILLCELL_X4 FILLER_116_310 ();
 FILLCELL_X4 FILLER_116_344 ();
 FILLCELL_X1 FILLER_116_348 ();
 FILLCELL_X2 FILLER_116_356 ();
 FILLCELL_X8 FILLER_116_365 ();
 FILLCELL_X4 FILLER_116_373 ();
 FILLCELL_X2 FILLER_116_384 ();
 FILLCELL_X2 FILLER_116_392 ();
 FILLCELL_X1 FILLER_116_401 ();
 FILLCELL_X2 FILLER_116_405 ();
 FILLCELL_X4 FILLER_116_410 ();
 FILLCELL_X2 FILLER_116_421 ();
 FILLCELL_X4 FILLER_116_437 ();
 FILLCELL_X4 FILLER_116_458 ();
 FILLCELL_X1 FILLER_116_466 ();
 FILLCELL_X8 FILLER_116_470 ();
 FILLCELL_X1 FILLER_116_478 ();
 FILLCELL_X1 FILLER_116_518 ();
 FILLCELL_X1 FILLER_116_526 ();
 FILLCELL_X2 FILLER_116_534 ();
 FILLCELL_X2 FILLER_116_543 ();
 FILLCELL_X2 FILLER_116_558 ();
 FILLCELL_X1 FILLER_116_560 ();
 FILLCELL_X2 FILLER_116_581 ();
 FILLCELL_X4 FILLER_116_590 ();
 FILLCELL_X1 FILLER_116_594 ();
 FILLCELL_X4 FILLER_116_605 ();
 FILLCELL_X2 FILLER_116_609 ();
 FILLCELL_X1 FILLER_116_611 ();
 FILLCELL_X1 FILLER_116_619 ();
 FILLCELL_X8 FILLER_116_623 ();
 FILLCELL_X4 FILLER_116_673 ();
 FILLCELL_X1 FILLER_116_677 ();
 FILLCELL_X1 FILLER_116_689 ();
 FILLCELL_X2 FILLER_116_706 ();
 FILLCELL_X1 FILLER_116_708 ();
 FILLCELL_X8 FILLER_116_725 ();
 FILLCELL_X4 FILLER_116_733 ();
 FILLCELL_X16 FILLER_116_757 ();
 FILLCELL_X1 FILLER_116_773 ();
 FILLCELL_X32 FILLER_116_808 ();
 FILLCELL_X4 FILLER_116_840 ();
 FILLCELL_X2 FILLER_116_856 ();
 FILLCELL_X8 FILLER_116_868 ();
 FILLCELL_X2 FILLER_116_876 ();
 FILLCELL_X1 FILLER_116_878 ();
 FILLCELL_X1 FILLER_116_916 ();
 FILLCELL_X16 FILLER_116_929 ();
 FILLCELL_X2 FILLER_116_945 ();
 FILLCELL_X4 FILLER_116_961 ();
 FILLCELL_X1 FILLER_116_965 ();
 FILLCELL_X8 FILLER_116_973 ();
 FILLCELL_X2 FILLER_116_981 ();
 FILLCELL_X1 FILLER_116_983 ();
 FILLCELL_X1 FILLER_116_995 ();
 FILLCELL_X4 FILLER_116_1040 ();
 FILLCELL_X2 FILLER_116_1044 ();
 FILLCELL_X8 FILLER_116_1053 ();
 FILLCELL_X2 FILLER_116_1061 ();
 FILLCELL_X8 FILLER_116_1070 ();
 FILLCELL_X1 FILLER_116_1078 ();
 FILLCELL_X4 FILLER_116_1081 ();
 FILLCELL_X1 FILLER_116_1085 ();
 FILLCELL_X4 FILLER_116_1111 ();
 FILLCELL_X4 FILLER_116_1134 ();
 FILLCELL_X1 FILLER_116_1164 ();
 FILLCELL_X1 FILLER_116_1185 ();
 FILLCELL_X1 FILLER_116_1193 ();
 FILLCELL_X1 FILLER_116_1201 ();
 FILLCELL_X1 FILLER_116_1209 ();
 FILLCELL_X2 FILLER_116_1217 ();
 FILLCELL_X16 FILLER_116_1239 ();
 FILLCELL_X2 FILLER_116_1255 ();
 FILLCELL_X2 FILLER_117_21 ();
 FILLCELL_X1 FILLER_117_23 ();
 FILLCELL_X2 FILLER_117_36 ();
 FILLCELL_X2 FILLER_117_45 ();
 FILLCELL_X1 FILLER_117_47 ();
 FILLCELL_X4 FILLER_117_55 ();
 FILLCELL_X2 FILLER_117_59 ();
 FILLCELL_X2 FILLER_117_68 ();
 FILLCELL_X1 FILLER_117_70 ();
 FILLCELL_X4 FILLER_117_78 ();
 FILLCELL_X2 FILLER_117_82 ();
 FILLCELL_X1 FILLER_117_91 ();
 FILLCELL_X1 FILLER_117_120 ();
 FILLCELL_X1 FILLER_117_128 ();
 FILLCELL_X4 FILLER_117_139 ();
 FILLCELL_X2 FILLER_117_156 ();
 FILLCELL_X1 FILLER_117_158 ();
 FILLCELL_X2 FILLER_117_179 ();
 FILLCELL_X8 FILLER_117_188 ();
 FILLCELL_X4 FILLER_117_196 ();
 FILLCELL_X1 FILLER_117_200 ();
 FILLCELL_X8 FILLER_117_208 ();
 FILLCELL_X4 FILLER_117_216 ();
 FILLCELL_X1 FILLER_117_220 ();
 FILLCELL_X1 FILLER_117_251 ();
 FILLCELL_X2 FILLER_117_259 ();
 FILLCELL_X2 FILLER_117_268 ();
 FILLCELL_X1 FILLER_117_270 ();
 FILLCELL_X2 FILLER_117_298 ();
 FILLCELL_X8 FILLER_117_314 ();
 FILLCELL_X4 FILLER_117_322 ();
 FILLCELL_X2 FILLER_117_326 ();
 FILLCELL_X1 FILLER_117_328 ();
 FILLCELL_X1 FILLER_117_361 ();
 FILLCELL_X4 FILLER_117_369 ();
 FILLCELL_X2 FILLER_117_373 ();
 FILLCELL_X1 FILLER_117_375 ();
 FILLCELL_X4 FILLER_117_379 ();
 FILLCELL_X1 FILLER_117_390 ();
 FILLCELL_X2 FILLER_117_398 ();
 FILLCELL_X2 FILLER_117_403 ();
 FILLCELL_X2 FILLER_117_409 ();
 FILLCELL_X1 FILLER_117_411 ();
 FILLCELL_X2 FILLER_117_416 ();
 FILLCELL_X8 FILLER_117_449 ();
 FILLCELL_X2 FILLER_117_457 ();
 FILLCELL_X2 FILLER_117_466 ();
 FILLCELL_X1 FILLER_117_526 ();
 FILLCELL_X4 FILLER_117_547 ();
 FILLCELL_X2 FILLER_117_551 ();
 FILLCELL_X1 FILLER_117_553 ();
 FILLCELL_X8 FILLER_117_561 ();
 FILLCELL_X2 FILLER_117_569 ();
 FILLCELL_X1 FILLER_117_571 ();
 FILLCELL_X1 FILLER_117_579 ();
 FILLCELL_X4 FILLER_117_600 ();
 FILLCELL_X2 FILLER_117_604 ();
 FILLCELL_X1 FILLER_117_606 ();
 FILLCELL_X8 FILLER_117_627 ();
 FILLCELL_X4 FILLER_117_635 ();
 FILLCELL_X2 FILLER_117_646 ();
 FILLCELL_X1 FILLER_117_648 ();
 FILLCELL_X4 FILLER_117_663 ();
 FILLCELL_X1 FILLER_117_672 ();
 FILLCELL_X2 FILLER_117_681 ();
 FILLCELL_X1 FILLER_117_687 ();
 FILLCELL_X4 FILLER_117_697 ();
 FILLCELL_X1 FILLER_117_701 ();
 FILLCELL_X4 FILLER_117_705 ();
 FILLCELL_X2 FILLER_117_709 ();
 FILLCELL_X1 FILLER_117_711 ();
 FILLCELL_X8 FILLER_117_716 ();
 FILLCELL_X4 FILLER_117_724 ();
 FILLCELL_X1 FILLER_117_728 ();
 FILLCELL_X2 FILLER_117_733 ();
 FILLCELL_X4 FILLER_117_742 ();
 FILLCELL_X2 FILLER_117_753 ();
 FILLCELL_X1 FILLER_117_762 ();
 FILLCELL_X2 FILLER_117_770 ();
 FILLCELL_X1 FILLER_117_789 ();
 FILLCELL_X2 FILLER_117_804 ();
 FILLCELL_X8 FILLER_117_810 ();
 FILLCELL_X1 FILLER_117_818 ();
 FILLCELL_X8 FILLER_117_831 ();
 FILLCELL_X1 FILLER_117_839 ();
 FILLCELL_X4 FILLER_117_858 ();
 FILLCELL_X2 FILLER_117_862 ();
 FILLCELL_X16 FILLER_117_891 ();
 FILLCELL_X1 FILLER_117_917 ();
 FILLCELL_X8 FILLER_117_950 ();
 FILLCELL_X1 FILLER_117_958 ();
 FILLCELL_X4 FILLER_117_973 ();
 FILLCELL_X1 FILLER_117_977 ();
 FILLCELL_X2 FILLER_117_996 ();
 FILLCELL_X1 FILLER_117_998 ();
 FILLCELL_X4 FILLER_117_1004 ();
 FILLCELL_X1 FILLER_117_1008 ();
 FILLCELL_X4 FILLER_117_1014 ();
 FILLCELL_X2 FILLER_117_1018 ();
 FILLCELL_X16 FILLER_117_1025 ();
 FILLCELL_X2 FILLER_117_1041 ();
 FILLCELL_X1 FILLER_117_1048 ();
 FILLCELL_X2 FILLER_117_1057 ();
 FILLCELL_X1 FILLER_117_1068 ();
 FILLCELL_X1 FILLER_117_1074 ();
 FILLCELL_X4 FILLER_117_1082 ();
 FILLCELL_X1 FILLER_117_1093 ();
 FILLCELL_X2 FILLER_117_1097 ();
 FILLCELL_X8 FILLER_117_1108 ();
 FILLCELL_X1 FILLER_117_1116 ();
 FILLCELL_X32 FILLER_117_1124 ();
 FILLCELL_X8 FILLER_117_1156 ();
 FILLCELL_X1 FILLER_117_1164 ();
 FILLCELL_X8 FILLER_117_1172 ();
 FILLCELL_X4 FILLER_117_1180 ();
 FILLCELL_X1 FILLER_117_1184 ();
 FILLCELL_X8 FILLER_117_1192 ();
 FILLCELL_X2 FILLER_117_1207 ();
 FILLCELL_X1 FILLER_117_1209 ();
 FILLCELL_X1 FILLER_117_1224 ();
 FILLCELL_X8 FILLER_117_1237 ();
 FILLCELL_X4 FILLER_117_1245 ();
 FILLCELL_X2 FILLER_117_1249 ();
 FILLCELL_X1 FILLER_117_1251 ();
 FILLCELL_X4 FILLER_117_1255 ();
 FILLCELL_X1 FILLER_117_1259 ();
 FILLCELL_X4 FILLER_118_1 ();
 FILLCELL_X1 FILLER_118_5 ();
 FILLCELL_X1 FILLER_118_33 ();
 FILLCELL_X4 FILLER_118_48 ();
 FILLCELL_X2 FILLER_118_52 ();
 FILLCELL_X1 FILLER_118_54 ();
 FILLCELL_X1 FILLER_118_75 ();
 FILLCELL_X4 FILLER_118_96 ();
 FILLCELL_X2 FILLER_118_100 ();
 FILLCELL_X1 FILLER_118_109 ();
 FILLCELL_X8 FILLER_118_131 ();
 FILLCELL_X4 FILLER_118_139 ();
 FILLCELL_X2 FILLER_118_143 ();
 FILLCELL_X2 FILLER_118_167 ();
 FILLCELL_X1 FILLER_118_169 ();
 FILLCELL_X1 FILLER_118_181 ();
 FILLCELL_X2 FILLER_118_207 ();
 FILLCELL_X8 FILLER_118_229 ();
 FILLCELL_X2 FILLER_118_237 ();
 FILLCELL_X1 FILLER_118_239 ();
 FILLCELL_X16 FILLER_118_280 ();
 FILLCELL_X8 FILLER_118_316 ();
 FILLCELL_X2 FILLER_118_324 ();
 FILLCELL_X4 FILLER_118_333 ();
 FILLCELL_X1 FILLER_118_337 ();
 FILLCELL_X1 FILLER_118_342 ();
 FILLCELL_X1 FILLER_118_346 ();
 FILLCELL_X2 FILLER_118_354 ();
 FILLCELL_X1 FILLER_118_386 ();
 FILLCELL_X2 FILLER_118_391 ();
 FILLCELL_X2 FILLER_118_397 ();
 FILLCELL_X2 FILLER_118_421 ();
 FILLCELL_X1 FILLER_118_423 ();
 FILLCELL_X4 FILLER_118_455 ();
 FILLCELL_X1 FILLER_118_486 ();
 FILLCELL_X2 FILLER_118_549 ();
 FILLCELL_X1 FILLER_118_551 ();
 FILLCELL_X4 FILLER_118_572 ();
 FILLCELL_X4 FILLER_118_590 ();
 FILLCELL_X1 FILLER_118_594 ();
 FILLCELL_X8 FILLER_118_616 ();
 FILLCELL_X4 FILLER_118_624 ();
 FILLCELL_X2 FILLER_118_628 ();
 FILLCELL_X1 FILLER_118_630 ();
 FILLCELL_X1 FILLER_118_670 ();
 FILLCELL_X2 FILLER_118_681 ();
 FILLCELL_X8 FILLER_118_690 ();
 FILLCELL_X2 FILLER_118_707 ();
 FILLCELL_X1 FILLER_118_709 ();
 FILLCELL_X1 FILLER_118_715 ();
 FILLCELL_X2 FILLER_118_745 ();
 FILLCELL_X1 FILLER_118_747 ();
 FILLCELL_X1 FILLER_118_760 ();
 FILLCELL_X1 FILLER_118_775 ();
 FILLCELL_X1 FILLER_118_783 ();
 FILLCELL_X2 FILLER_118_820 ();
 FILLCELL_X4 FILLER_118_844 ();
 FILLCELL_X1 FILLER_118_848 ();
 FILLCELL_X16 FILLER_118_853 ();
 FILLCELL_X1 FILLER_118_869 ();
 FILLCELL_X1 FILLER_118_874 ();
 FILLCELL_X1 FILLER_118_882 ();
 FILLCELL_X1 FILLER_118_893 ();
 FILLCELL_X1 FILLER_118_927 ();
 FILLCELL_X8 FILLER_118_962 ();
 FILLCELL_X4 FILLER_118_970 ();
 FILLCELL_X4 FILLER_118_981 ();
 FILLCELL_X2 FILLER_118_985 ();
 FILLCELL_X1 FILLER_118_987 ();
 FILLCELL_X2 FILLER_118_995 ();
 FILLCELL_X8 FILLER_118_1010 ();
 FILLCELL_X2 FILLER_118_1022 ();
 FILLCELL_X1 FILLER_118_1024 ();
 FILLCELL_X8 FILLER_118_1029 ();
 FILLCELL_X4 FILLER_118_1037 ();
 FILLCELL_X2 FILLER_118_1041 ();
 FILLCELL_X1 FILLER_118_1043 ();
 FILLCELL_X1 FILLER_118_1080 ();
 FILLCELL_X2 FILLER_118_1085 ();
 FILLCELL_X1 FILLER_118_1087 ();
 FILLCELL_X2 FILLER_118_1092 ();
 FILLCELL_X2 FILLER_118_1098 ();
 FILLCELL_X16 FILLER_118_1111 ();
 FILLCELL_X8 FILLER_118_1127 ();
 FILLCELL_X4 FILLER_118_1135 ();
 FILLCELL_X2 FILLER_118_1139 ();
 FILLCELL_X16 FILLER_118_1173 ();
 FILLCELL_X8 FILLER_118_1189 ();
 FILLCELL_X2 FILLER_118_1197 ();
 FILLCELL_X1 FILLER_118_1199 ();
 FILLCELL_X8 FILLER_118_1220 ();
 FILLCELL_X4 FILLER_118_1228 ();
 FILLCELL_X2 FILLER_118_1235 ();
 FILLCELL_X1 FILLER_118_1240 ();
 FILLCELL_X8 FILLER_118_1247 ();
 FILLCELL_X4 FILLER_118_1255 ();
 FILLCELL_X1 FILLER_118_1259 ();
 FILLCELL_X8 FILLER_119_1 ();
 FILLCELL_X4 FILLER_119_9 ();
 FILLCELL_X8 FILLER_119_20 ();
 FILLCELL_X4 FILLER_119_28 ();
 FILLCELL_X1 FILLER_119_32 ();
 FILLCELL_X2 FILLER_119_40 ();
 FILLCELL_X16 FILLER_119_49 ();
 FILLCELL_X4 FILLER_119_65 ();
 FILLCELL_X2 FILLER_119_69 ();
 FILLCELL_X1 FILLER_119_112 ();
 FILLCELL_X2 FILLER_119_120 ();
 FILLCELL_X2 FILLER_119_129 ();
 FILLCELL_X8 FILLER_119_158 ();
 FILLCELL_X2 FILLER_119_166 ();
 FILLCELL_X1 FILLER_119_189 ();
 FILLCELL_X8 FILLER_119_207 ();
 FILLCELL_X4 FILLER_119_215 ();
 FILLCELL_X2 FILLER_119_219 ();
 FILLCELL_X1 FILLER_119_221 ();
 FILLCELL_X8 FILLER_119_259 ();
 FILLCELL_X4 FILLER_119_267 ();
 FILLCELL_X1 FILLER_119_271 ();
 FILLCELL_X2 FILLER_119_299 ();
 FILLCELL_X2 FILLER_119_308 ();
 FILLCELL_X2 FILLER_119_317 ();
 FILLCELL_X1 FILLER_119_319 ();
 FILLCELL_X2 FILLER_119_327 ();
 FILLCELL_X1 FILLER_119_329 ();
 FILLCELL_X2 FILLER_119_350 ();
 FILLCELL_X8 FILLER_119_366 ();
 FILLCELL_X2 FILLER_119_374 ();
 FILLCELL_X1 FILLER_119_393 ();
 FILLCELL_X4 FILLER_119_443 ();
 FILLCELL_X2 FILLER_119_501 ();
 FILLCELL_X2 FILLER_119_535 ();
 FILLCELL_X1 FILLER_119_537 ();
 FILLCELL_X1 FILLER_119_559 ();
 FILLCELL_X1 FILLER_119_570 ();
 FILLCELL_X1 FILLER_119_581 ();
 FILLCELL_X8 FILLER_119_589 ();
 FILLCELL_X1 FILLER_119_597 ();
 FILLCELL_X32 FILLER_119_611 ();
 FILLCELL_X8 FILLER_119_643 ();
 FILLCELL_X1 FILLER_119_651 ();
 FILLCELL_X4 FILLER_119_685 ();
 FILLCELL_X2 FILLER_119_689 ();
 FILLCELL_X1 FILLER_119_691 ();
 FILLCELL_X2 FILLER_119_699 ();
 FILLCELL_X1 FILLER_119_701 ();
 FILLCELL_X8 FILLER_119_707 ();
 FILLCELL_X2 FILLER_119_715 ();
 FILLCELL_X1 FILLER_119_717 ();
 FILLCELL_X1 FILLER_119_738 ();
 FILLCELL_X1 FILLER_119_745 ();
 FILLCELL_X4 FILLER_119_761 ();
 FILLCELL_X2 FILLER_119_772 ();
 FILLCELL_X2 FILLER_119_777 ();
 FILLCELL_X1 FILLER_119_779 ();
 FILLCELL_X1 FILLER_119_787 ();
 FILLCELL_X1 FILLER_119_801 ();
 FILLCELL_X2 FILLER_119_828 ();
 FILLCELL_X1 FILLER_119_830 ();
 FILLCELL_X4 FILLER_119_855 ();
 FILLCELL_X2 FILLER_119_859 ();
 FILLCELL_X1 FILLER_119_861 ();
 FILLCELL_X4 FILLER_119_939 ();
 FILLCELL_X1 FILLER_119_943 ();
 FILLCELL_X1 FILLER_119_958 ();
 FILLCELL_X1 FILLER_119_973 ();
 FILLCELL_X4 FILLER_119_977 ();
 FILLCELL_X2 FILLER_119_981 ();
 FILLCELL_X1 FILLER_119_983 ();
 FILLCELL_X8 FILLER_119_988 ();
 FILLCELL_X4 FILLER_119_996 ();
 FILLCELL_X2 FILLER_119_1000 ();
 FILLCELL_X1 FILLER_119_1002 ();
 FILLCELL_X1 FILLER_119_1016 ();
 FILLCELL_X16 FILLER_119_1025 ();
 FILLCELL_X2 FILLER_119_1041 ();
 FILLCELL_X1 FILLER_119_1043 ();
 FILLCELL_X4 FILLER_119_1049 ();
 FILLCELL_X1 FILLER_119_1053 ();
 FILLCELL_X4 FILLER_119_1070 ();
 FILLCELL_X2 FILLER_119_1074 ();
 FILLCELL_X16 FILLER_119_1083 ();
 FILLCELL_X16 FILLER_119_1106 ();
 FILLCELL_X8 FILLER_119_1122 ();
 FILLCELL_X2 FILLER_119_1130 ();
 FILLCELL_X2 FILLER_119_1159 ();
 FILLCELL_X1 FILLER_119_1161 ();
 FILLCELL_X2 FILLER_119_1176 ();
 FILLCELL_X4 FILLER_119_1198 ();
 FILLCELL_X2 FILLER_119_1202 ();
 FILLCELL_X1 FILLER_119_1204 ();
 FILLCELL_X8 FILLER_119_1245 ();
 FILLCELL_X4 FILLER_119_1253 ();
 FILLCELL_X2 FILLER_119_1257 ();
 FILLCELL_X1 FILLER_119_1259 ();
 FILLCELL_X1 FILLER_120_1 ();
 FILLCELL_X2 FILLER_120_22 ();
 FILLCELL_X2 FILLER_120_31 ();
 FILLCELL_X2 FILLER_120_40 ();
 FILLCELL_X4 FILLER_120_49 ();
 FILLCELL_X4 FILLER_120_73 ();
 FILLCELL_X4 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_115 ();
 FILLCELL_X2 FILLER_120_147 ();
 FILLCELL_X8 FILLER_120_203 ();
 FILLCELL_X2 FILLER_120_211 ();
 FILLCELL_X1 FILLER_120_213 ();
 FILLCELL_X1 FILLER_120_241 ();
 FILLCELL_X2 FILLER_120_256 ();
 FILLCELL_X1 FILLER_120_275 ();
 FILLCELL_X2 FILLER_120_280 ();
 FILLCELL_X8 FILLER_120_289 ();
 FILLCELL_X2 FILLER_120_297 ();
 FILLCELL_X1 FILLER_120_299 ();
 FILLCELL_X1 FILLER_120_307 ();
 FILLCELL_X1 FILLER_120_315 ();
 FILLCELL_X2 FILLER_120_323 ();
 FILLCELL_X2 FILLER_120_328 ();
 FILLCELL_X2 FILLER_120_335 ();
 FILLCELL_X1 FILLER_120_344 ();
 FILLCELL_X1 FILLER_120_352 ();
 FILLCELL_X4 FILLER_120_363 ();
 FILLCELL_X2 FILLER_120_367 ();
 FILLCELL_X8 FILLER_120_389 ();
 FILLCELL_X1 FILLER_120_397 ();
 FILLCELL_X8 FILLER_120_407 ();
 FILLCELL_X4 FILLER_120_415 ();
 FILLCELL_X2 FILLER_120_432 ();
 FILLCELL_X1 FILLER_120_506 ();
 FILLCELL_X8 FILLER_120_618 ();
 FILLCELL_X4 FILLER_120_632 ();
 FILLCELL_X2 FILLER_120_636 ();
 FILLCELL_X4 FILLER_120_641 ();
 FILLCELL_X4 FILLER_120_686 ();
 FILLCELL_X2 FILLER_120_690 ();
 FILLCELL_X1 FILLER_120_692 ();
 FILLCELL_X2 FILLER_120_709 ();
 FILLCELL_X4 FILLER_120_721 ();
 FILLCELL_X8 FILLER_120_730 ();
 FILLCELL_X4 FILLER_120_738 ();
 FILLCELL_X4 FILLER_120_746 ();
 FILLCELL_X2 FILLER_120_750 ();
 FILLCELL_X4 FILLER_120_759 ();
 FILLCELL_X1 FILLER_120_775 ();
 FILLCELL_X4 FILLER_120_793 ();
 FILLCELL_X4 FILLER_120_815 ();
 FILLCELL_X2 FILLER_120_819 ();
 FILLCELL_X1 FILLER_120_821 ();
 FILLCELL_X16 FILLER_120_839 ();
 FILLCELL_X2 FILLER_120_855 ();
 FILLCELL_X4 FILLER_120_921 ();
 FILLCELL_X2 FILLER_120_925 ();
 FILLCELL_X8 FILLER_120_934 ();
 FILLCELL_X2 FILLER_120_942 ();
 FILLCELL_X1 FILLER_120_944 ();
 FILLCELL_X8 FILLER_120_948 ();
 FILLCELL_X2 FILLER_120_956 ();
 FILLCELL_X1 FILLER_120_958 ();
 FILLCELL_X8 FILLER_120_973 ();
 FILLCELL_X2 FILLER_120_981 ();
 FILLCELL_X4 FILLER_120_997 ();
 FILLCELL_X1 FILLER_120_1001 ();
 FILLCELL_X4 FILLER_120_1016 ();
 FILLCELL_X1 FILLER_120_1020 ();
 FILLCELL_X8 FILLER_120_1025 ();
 FILLCELL_X4 FILLER_120_1033 ();
 FILLCELL_X8 FILLER_120_1042 ();
 FILLCELL_X2 FILLER_120_1050 ();
 FILLCELL_X1 FILLER_120_1052 ();
 FILLCELL_X8 FILLER_120_1061 ();
 FILLCELL_X2 FILLER_120_1069 ();
 FILLCELL_X1 FILLER_120_1071 ();
 FILLCELL_X2 FILLER_120_1086 ();
 FILLCELL_X4 FILLER_120_1101 ();
 FILLCELL_X2 FILLER_120_1105 ();
 FILLCELL_X1 FILLER_120_1107 ();
 FILLCELL_X8 FILLER_120_1123 ();
 FILLCELL_X4 FILLER_120_1131 ();
 FILLCELL_X1 FILLER_120_1135 ();
 FILLCELL_X1 FILLER_120_1163 ();
 FILLCELL_X2 FILLER_120_1200 ();
 FILLCELL_X1 FILLER_120_1202 ();
 FILLCELL_X4 FILLER_120_1210 ();
 FILLCELL_X1 FILLER_120_1214 ();
 FILLCELL_X8 FILLER_120_1222 ();
 FILLCELL_X1 FILLER_120_1230 ();
 FILLCELL_X4 FILLER_120_1238 ();
 FILLCELL_X1 FILLER_120_1242 ();
 FILLCELL_X1 FILLER_120_1246 ();
 FILLCELL_X2 FILLER_120_1250 ();
 FILLCELL_X1 FILLER_120_1252 ();
 FILLCELL_X4 FILLER_120_1256 ();
 FILLCELL_X4 FILLER_121_1 ();
 FILLCELL_X1 FILLER_121_5 ();
 FILLCELL_X8 FILLER_121_40 ();
 FILLCELL_X1 FILLER_121_48 ();
 FILLCELL_X2 FILLER_121_56 ();
 FILLCELL_X1 FILLER_121_58 ();
 FILLCELL_X8 FILLER_121_115 ();
 FILLCELL_X2 FILLER_121_123 ();
 FILLCELL_X2 FILLER_121_152 ();
 FILLCELL_X1 FILLER_121_154 ();
 FILLCELL_X2 FILLER_121_162 ();
 FILLCELL_X32 FILLER_121_180 ();
 FILLCELL_X8 FILLER_121_212 ();
 FILLCELL_X2 FILLER_121_220 ();
 FILLCELL_X1 FILLER_121_222 ();
 FILLCELL_X4 FILLER_121_235 ();
 FILLCELL_X1 FILLER_121_239 ();
 FILLCELL_X1 FILLER_121_247 ();
 FILLCELL_X2 FILLER_121_254 ();
 FILLCELL_X4 FILLER_121_279 ();
 FILLCELL_X8 FILLER_121_303 ();
 FILLCELL_X2 FILLER_121_311 ();
 FILLCELL_X1 FILLER_121_313 ();
 FILLCELL_X4 FILLER_121_321 ();
 FILLCELL_X1 FILLER_121_325 ();
 FILLCELL_X1 FILLER_121_349 ();
 FILLCELL_X2 FILLER_121_360 ();
 FILLCELL_X1 FILLER_121_362 ();
 FILLCELL_X2 FILLER_121_370 ();
 FILLCELL_X4 FILLER_121_379 ();
 FILLCELL_X4 FILLER_121_396 ();
 FILLCELL_X2 FILLER_121_400 ();
 FILLCELL_X1 FILLER_121_427 ();
 FILLCELL_X1 FILLER_121_434 ();
 FILLCELL_X2 FILLER_121_440 ();
 FILLCELL_X1 FILLER_121_442 ();
 FILLCELL_X2 FILLER_121_588 ();
 FILLCELL_X2 FILLER_121_597 ();
 FILLCELL_X8 FILLER_121_619 ();
 FILLCELL_X4 FILLER_121_629 ();
 FILLCELL_X1 FILLER_121_633 ();
 FILLCELL_X8 FILLER_121_661 ();
 FILLCELL_X2 FILLER_121_669 ();
 FILLCELL_X1 FILLER_121_685 ();
 FILLCELL_X4 FILLER_121_696 ();
 FILLCELL_X2 FILLER_121_700 ();
 FILLCELL_X1 FILLER_121_715 ();
 FILLCELL_X1 FILLER_121_720 ();
 FILLCELL_X2 FILLER_121_732 ();
 FILLCELL_X1 FILLER_121_734 ();
 FILLCELL_X1 FILLER_121_747 ();
 FILLCELL_X4 FILLER_121_753 ();
 FILLCELL_X1 FILLER_121_757 ();
 FILLCELL_X2 FILLER_121_791 ();
 FILLCELL_X1 FILLER_121_793 ();
 FILLCELL_X4 FILLER_121_797 ();
 FILLCELL_X1 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_809 ();
 FILLCELL_X4 FILLER_121_841 ();
 FILLCELL_X2 FILLER_121_845 ();
 FILLCELL_X4 FILLER_121_878 ();
 FILLCELL_X8 FILLER_121_886 ();
 FILLCELL_X1 FILLER_121_894 ();
 FILLCELL_X4 FILLER_121_902 ();
 FILLCELL_X2 FILLER_121_906 ();
 FILLCELL_X1 FILLER_121_908 ();
 FILLCELL_X4 FILLER_121_916 ();
 FILLCELL_X2 FILLER_121_920 ();
 FILLCELL_X1 FILLER_121_922 ();
 FILLCELL_X1 FILLER_121_930 ();
 FILLCELL_X2 FILLER_121_951 ();
 FILLCELL_X1 FILLER_121_953 ();
 FILLCELL_X16 FILLER_121_968 ();
 FILLCELL_X2 FILLER_121_984 ();
 FILLCELL_X1 FILLER_121_986 ();
 FILLCELL_X4 FILLER_121_992 ();
 FILLCELL_X2 FILLER_121_1000 ();
 FILLCELL_X1 FILLER_121_1002 ();
 FILLCELL_X1 FILLER_121_1041 ();
 FILLCELL_X2 FILLER_121_1046 ();
 FILLCELL_X1 FILLER_121_1048 ();
 FILLCELL_X2 FILLER_121_1051 ();
 FILLCELL_X8 FILLER_121_1064 ();
 FILLCELL_X1 FILLER_121_1072 ();
 FILLCELL_X8 FILLER_121_1077 ();
 FILLCELL_X1 FILLER_121_1085 ();
 FILLCELL_X1 FILLER_121_1093 ();
 FILLCELL_X1 FILLER_121_1096 ();
 FILLCELL_X2 FILLER_121_1101 ();
 FILLCELL_X2 FILLER_121_1127 ();
 FILLCELL_X2 FILLER_121_1156 ();
 FILLCELL_X4 FILLER_121_1165 ();
 FILLCELL_X2 FILLER_121_1210 ();
 FILLCELL_X1 FILLER_121_1212 ();
 FILLCELL_X2 FILLER_121_1240 ();
 FILLCELL_X4 FILLER_121_1245 ();
 FILLCELL_X2 FILLER_121_1249 ();
 FILLCELL_X2 FILLER_121_1257 ();
 FILLCELL_X1 FILLER_121_1259 ();
 FILLCELL_X4 FILLER_122_21 ();
 FILLCELL_X2 FILLER_122_25 ();
 FILLCELL_X8 FILLER_122_34 ();
 FILLCELL_X4 FILLER_122_42 ();
 FILLCELL_X2 FILLER_122_46 ();
 FILLCELL_X4 FILLER_122_55 ();
 FILLCELL_X1 FILLER_122_59 ();
 FILLCELL_X8 FILLER_122_87 ();
 FILLCELL_X1 FILLER_122_95 ();
 FILLCELL_X2 FILLER_122_103 ();
 FILLCELL_X1 FILLER_122_105 ();
 FILLCELL_X2 FILLER_122_133 ();
 FILLCELL_X1 FILLER_122_135 ();
 FILLCELL_X8 FILLER_122_194 ();
 FILLCELL_X4 FILLER_122_209 ();
 FILLCELL_X1 FILLER_122_240 ();
 FILLCELL_X2 FILLER_122_248 ();
 FILLCELL_X2 FILLER_122_254 ();
 FILLCELL_X2 FILLER_122_259 ();
 FILLCELL_X2 FILLER_122_268 ();
 FILLCELL_X2 FILLER_122_297 ();
 FILLCELL_X2 FILLER_122_306 ();
 FILLCELL_X1 FILLER_122_308 ();
 FILLCELL_X2 FILLER_122_316 ();
 FILLCELL_X1 FILLER_122_318 ();
 FILLCELL_X2 FILLER_122_333 ();
 FILLCELL_X1 FILLER_122_335 ();
 FILLCELL_X4 FILLER_122_356 ();
 FILLCELL_X2 FILLER_122_407 ();
 FILLCELL_X2 FILLER_122_426 ();
 FILLCELL_X8 FILLER_122_437 ();
 FILLCELL_X1 FILLER_122_489 ();
 FILLCELL_X1 FILLER_122_506 ();
 FILLCELL_X1 FILLER_122_630 ();
 FILLCELL_X4 FILLER_122_637 ();
 FILLCELL_X2 FILLER_122_641 ();
 FILLCELL_X1 FILLER_122_643 ();
 FILLCELL_X1 FILLER_122_651 ();
 FILLCELL_X2 FILLER_122_666 ();
 FILLCELL_X1 FILLER_122_681 ();
 FILLCELL_X4 FILLER_122_689 ();
 FILLCELL_X1 FILLER_122_693 ();
 FILLCELL_X2 FILLER_122_698 ();
 FILLCELL_X1 FILLER_122_700 ();
 FILLCELL_X2 FILLER_122_710 ();
 FILLCELL_X16 FILLER_122_717 ();
 FILLCELL_X1 FILLER_122_749 ();
 FILLCELL_X2 FILLER_122_757 ();
 FILLCELL_X1 FILLER_122_759 ();
 FILLCELL_X1 FILLER_122_773 ();
 FILLCELL_X8 FILLER_122_849 ();
 FILLCELL_X4 FILLER_122_857 ();
 FILLCELL_X2 FILLER_122_861 ();
 FILLCELL_X2 FILLER_122_866 ();
 FILLCELL_X2 FILLER_122_898 ();
 FILLCELL_X8 FILLER_122_907 ();
 FILLCELL_X4 FILLER_122_915 ();
 FILLCELL_X2 FILLER_122_919 ();
 FILLCELL_X2 FILLER_122_928 ();
 FILLCELL_X1 FILLER_122_930 ();
 FILLCELL_X4 FILLER_122_938 ();
 FILLCELL_X2 FILLER_122_942 ();
 FILLCELL_X2 FILLER_122_987 ();
 FILLCELL_X1 FILLER_122_993 ();
 FILLCELL_X8 FILLER_122_1003 ();
 FILLCELL_X4 FILLER_122_1011 ();
 FILLCELL_X1 FILLER_122_1020 ();
 FILLCELL_X8 FILLER_122_1036 ();
 FILLCELL_X1 FILLER_122_1058 ();
 FILLCELL_X4 FILLER_122_1070 ();
 FILLCELL_X2 FILLER_122_1074 ();
 FILLCELL_X2 FILLER_122_1079 ();
 FILLCELL_X2 FILLER_122_1094 ();
 FILLCELL_X1 FILLER_122_1096 ();
 FILLCELL_X4 FILLER_122_1102 ();
 FILLCELL_X1 FILLER_122_1106 ();
 FILLCELL_X1 FILLER_122_1114 ();
 FILLCELL_X16 FILLER_122_1122 ();
 FILLCELL_X8 FILLER_122_1138 ();
 FILLCELL_X4 FILLER_122_1146 ();
 FILLCELL_X1 FILLER_122_1150 ();
 FILLCELL_X16 FILLER_122_1156 ();
 FILLCELL_X8 FILLER_122_1172 ();
 FILLCELL_X2 FILLER_122_1180 ();
 FILLCELL_X4 FILLER_122_1189 ();
 FILLCELL_X2 FILLER_122_1200 ();
 FILLCELL_X1 FILLER_122_1202 ();
 FILLCELL_X32 FILLER_122_1210 ();
 FILLCELL_X8 FILLER_122_1242 ();
 FILLCELL_X4 FILLER_122_1250 ();
 FILLCELL_X4 FILLER_123_1 ();
 FILLCELL_X2 FILLER_123_5 ();
 FILLCELL_X1 FILLER_123_7 ();
 FILLCELL_X4 FILLER_123_35 ();
 FILLCELL_X2 FILLER_123_39 ();
 FILLCELL_X4 FILLER_123_68 ();
 FILLCELL_X2 FILLER_123_92 ();
 FILLCELL_X1 FILLER_123_101 ();
 FILLCELL_X2 FILLER_123_109 ();
 FILLCELL_X8 FILLER_123_118 ();
 FILLCELL_X4 FILLER_123_126 ();
 FILLCELL_X2 FILLER_123_130 ();
 FILLCELL_X1 FILLER_123_139 ();
 FILLCELL_X8 FILLER_123_147 ();
 FILLCELL_X1 FILLER_123_155 ();
 FILLCELL_X1 FILLER_123_170 ();
 FILLCELL_X2 FILLER_123_178 ();
 FILLCELL_X2 FILLER_123_200 ();
 FILLCELL_X8 FILLER_123_211 ();
 FILLCELL_X1 FILLER_123_219 ();
 FILLCELL_X1 FILLER_123_232 ();
 FILLCELL_X2 FILLER_123_240 ();
 FILLCELL_X4 FILLER_123_249 ();
 FILLCELL_X1 FILLER_123_253 ();
 FILLCELL_X16 FILLER_123_261 ();
 FILLCELL_X8 FILLER_123_277 ();
 FILLCELL_X1 FILLER_123_285 ();
 FILLCELL_X4 FILLER_123_293 ();
 FILLCELL_X2 FILLER_123_297 ();
 FILLCELL_X16 FILLER_123_313 ();
 FILLCELL_X4 FILLER_123_329 ();
 FILLCELL_X2 FILLER_123_333 ();
 FILLCELL_X1 FILLER_123_335 ();
 FILLCELL_X2 FILLER_123_339 ();
 FILLCELL_X4 FILLER_123_345 ();
 FILLCELL_X8 FILLER_123_357 ();
 FILLCELL_X4 FILLER_123_365 ();
 FILLCELL_X2 FILLER_123_369 ();
 FILLCELL_X1 FILLER_123_371 ();
 FILLCELL_X1 FILLER_123_401 ();
 FILLCELL_X1 FILLER_123_408 ();
 FILLCELL_X1 FILLER_123_433 ();
 FILLCELL_X1 FILLER_123_438 ();
 FILLCELL_X8 FILLER_123_442 ();
 FILLCELL_X2 FILLER_123_464 ();
 FILLCELL_X2 FILLER_123_495 ();
 FILLCELL_X1 FILLER_123_558 ();
 FILLCELL_X2 FILLER_123_615 ();
 FILLCELL_X8 FILLER_123_630 ();
 FILLCELL_X1 FILLER_123_638 ();
 FILLCELL_X2 FILLER_123_652 ();
 FILLCELL_X1 FILLER_123_654 ();
 FILLCELL_X1 FILLER_123_670 ();
 FILLCELL_X1 FILLER_123_708 ();
 FILLCELL_X4 FILLER_123_723 ();
 FILLCELL_X2 FILLER_123_727 ();
 FILLCELL_X2 FILLER_123_757 ();
 FILLCELL_X4 FILLER_123_766 ();
 FILLCELL_X2 FILLER_123_770 ();
 FILLCELL_X1 FILLER_123_779 ();
 FILLCELL_X8 FILLER_123_787 ();
 FILLCELL_X4 FILLER_123_795 ();
 FILLCELL_X1 FILLER_123_826 ();
 FILLCELL_X2 FILLER_123_837 ();
 FILLCELL_X2 FILLER_123_849 ();
 FILLCELL_X2 FILLER_123_886 ();
 FILLCELL_X2 FILLER_123_900 ();
 FILLCELL_X4 FILLER_123_922 ();
 FILLCELL_X2 FILLER_123_930 ();
 FILLCELL_X4 FILLER_123_952 ();
 FILLCELL_X2 FILLER_123_956 ();
 FILLCELL_X1 FILLER_123_958 ();
 FILLCELL_X2 FILLER_123_992 ();
 FILLCELL_X8 FILLER_123_1001 ();
 FILLCELL_X4 FILLER_123_1009 ();
 FILLCELL_X2 FILLER_123_1013 ();
 FILLCELL_X1 FILLER_123_1023 ();
 FILLCELL_X1 FILLER_123_1042 ();
 FILLCELL_X4 FILLER_123_1054 ();
 FILLCELL_X1 FILLER_123_1058 ();
 FILLCELL_X4 FILLER_123_1086 ();
 FILLCELL_X8 FILLER_123_1112 ();
 FILLCELL_X4 FILLER_123_1131 ();
 FILLCELL_X1 FILLER_123_1135 ();
 FILLCELL_X2 FILLER_123_1143 ();
 FILLCELL_X16 FILLER_123_1182 ();
 FILLCELL_X2 FILLER_123_1198 ();
 FILLCELL_X2 FILLER_123_1207 ();
 FILLCELL_X16 FILLER_123_1235 ();
 FILLCELL_X4 FILLER_123_1251 ();
 FILLCELL_X2 FILLER_123_1255 ();
 FILLCELL_X4 FILLER_124_1 ();
 FILLCELL_X2 FILLER_124_5 ();
 FILLCELL_X8 FILLER_124_12 ();
 FILLCELL_X4 FILLER_124_20 ();
 FILLCELL_X2 FILLER_124_24 ();
 FILLCELL_X4 FILLER_124_40 ();
 FILLCELL_X2 FILLER_124_44 ();
 FILLCELL_X1 FILLER_124_46 ();
 FILLCELL_X2 FILLER_124_74 ();
 FILLCELL_X1 FILLER_124_76 ();
 FILLCELL_X1 FILLER_124_103 ();
 FILLCELL_X8 FILLER_124_111 ();
 FILLCELL_X16 FILLER_124_147 ();
 FILLCELL_X4 FILLER_124_163 ();
 FILLCELL_X2 FILLER_124_174 ();
 FILLCELL_X4 FILLER_124_183 ();
 FILLCELL_X4 FILLER_124_198 ();
 FILLCELL_X2 FILLER_124_202 ();
 FILLCELL_X1 FILLER_124_204 ();
 FILLCELL_X2 FILLER_124_215 ();
 FILLCELL_X4 FILLER_124_230 ();
 FILLCELL_X2 FILLER_124_234 ();
 FILLCELL_X1 FILLER_124_236 ();
 FILLCELL_X4 FILLER_124_284 ();
 FILLCELL_X1 FILLER_124_288 ();
 FILLCELL_X1 FILLER_124_316 ();
 FILLCELL_X2 FILLER_124_321 ();
 FILLCELL_X1 FILLER_124_333 ();
 FILLCELL_X4 FILLER_124_359 ();
 FILLCELL_X8 FILLER_124_407 ();
 FILLCELL_X2 FILLER_124_415 ();
 FILLCELL_X4 FILLER_124_420 ();
 FILLCELL_X1 FILLER_124_424 ();
 FILLCELL_X4 FILLER_124_436 ();
 FILLCELL_X1 FILLER_124_529 ();
 FILLCELL_X2 FILLER_124_550 ();
 FILLCELL_X1 FILLER_124_556 ();
 FILLCELL_X1 FILLER_124_593 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X1 FILLER_124_692 ();
 FILLCELL_X2 FILLER_124_697 ();
 FILLCELL_X2 FILLER_124_703 ();
 FILLCELL_X2 FILLER_124_712 ();
 FILLCELL_X4 FILLER_124_721 ();
 FILLCELL_X2 FILLER_124_725 ();
 FILLCELL_X2 FILLER_124_751 ();
 FILLCELL_X1 FILLER_124_753 ();
 FILLCELL_X2 FILLER_124_768 ();
 FILLCELL_X32 FILLER_124_777 ();
 FILLCELL_X2 FILLER_124_809 ();
 FILLCELL_X1 FILLER_124_811 ();
 FILLCELL_X4 FILLER_124_821 ();
 FILLCELL_X1 FILLER_124_825 ();
 FILLCELL_X16 FILLER_124_842 ();
 FILLCELL_X8 FILLER_124_858 ();
 FILLCELL_X2 FILLER_124_866 ();
 FILLCELL_X2 FILLER_124_878 ();
 FILLCELL_X1 FILLER_124_880 ();
 FILLCELL_X1 FILLER_124_886 ();
 FILLCELL_X1 FILLER_124_915 ();
 FILLCELL_X8 FILLER_124_923 ();
 FILLCELL_X2 FILLER_124_931 ();
 FILLCELL_X1 FILLER_124_933 ();
 FILLCELL_X4 FILLER_124_942 ();
 FILLCELL_X8 FILLER_124_960 ();
 FILLCELL_X1 FILLER_124_968 ();
 FILLCELL_X1 FILLER_124_987 ();
 FILLCELL_X2 FILLER_124_995 ();
 FILLCELL_X1 FILLER_124_1004 ();
 FILLCELL_X2 FILLER_124_1015 ();
 FILLCELL_X1 FILLER_124_1017 ();
 FILLCELL_X8 FILLER_124_1025 ();
 FILLCELL_X2 FILLER_124_1033 ();
 FILLCELL_X1 FILLER_124_1035 ();
 FILLCELL_X4 FILLER_124_1041 ();
 FILLCELL_X4 FILLER_124_1053 ();
 FILLCELL_X2 FILLER_124_1057 ();
 FILLCELL_X16 FILLER_124_1074 ();
 FILLCELL_X4 FILLER_124_1090 ();
 FILLCELL_X1 FILLER_124_1094 ();
 FILLCELL_X2 FILLER_124_1105 ();
 FILLCELL_X4 FILLER_124_1125 ();
 FILLCELL_X1 FILLER_124_1129 ();
 FILLCELL_X1 FILLER_124_1172 ();
 FILLCELL_X1 FILLER_124_1200 ();
 FILLCELL_X16 FILLER_124_1233 ();
 FILLCELL_X8 FILLER_124_1249 ();
 FILLCELL_X2 FILLER_124_1257 ();
 FILLCELL_X1 FILLER_124_1259 ();
 FILLCELL_X4 FILLER_125_28 ();
 FILLCELL_X16 FILLER_125_46 ();
 FILLCELL_X4 FILLER_125_62 ();
 FILLCELL_X2 FILLER_125_66 ();
 FILLCELL_X2 FILLER_125_88 ();
 FILLCELL_X1 FILLER_125_131 ();
 FILLCELL_X8 FILLER_125_146 ();
 FILLCELL_X8 FILLER_125_181 ();
 FILLCELL_X2 FILLER_125_202 ();
 FILLCELL_X2 FILLER_125_230 ();
 FILLCELL_X1 FILLER_125_232 ();
 FILLCELL_X1 FILLER_125_259 ();
 FILLCELL_X8 FILLER_125_262 ();
 FILLCELL_X2 FILLER_125_270 ();
 FILLCELL_X1 FILLER_125_272 ();
 FILLCELL_X8 FILLER_125_293 ();
 FILLCELL_X2 FILLER_125_301 ();
 FILLCELL_X1 FILLER_125_310 ();
 FILLCELL_X2 FILLER_125_331 ();
 FILLCELL_X1 FILLER_125_333 ();
 FILLCELL_X8 FILLER_125_354 ();
 FILLCELL_X1 FILLER_125_378 ();
 FILLCELL_X8 FILLER_125_399 ();
 FILLCELL_X4 FILLER_125_407 ();
 FILLCELL_X8 FILLER_125_418 ();
 FILLCELL_X2 FILLER_125_426 ();
 FILLCELL_X1 FILLER_125_450 ();
 FILLCELL_X2 FILLER_125_492 ();
 FILLCELL_X1 FILLER_125_560 ();
 FILLCELL_X2 FILLER_125_609 ();
 FILLCELL_X1 FILLER_125_631 ();
 FILLCELL_X1 FILLER_125_672 ();
 FILLCELL_X2 FILLER_125_681 ();
 FILLCELL_X1 FILLER_125_683 ();
 FILLCELL_X1 FILLER_125_687 ();
 FILLCELL_X4 FILLER_125_695 ();
 FILLCELL_X1 FILLER_125_699 ();
 FILLCELL_X1 FILLER_125_703 ();
 FILLCELL_X2 FILLER_125_718 ();
 FILLCELL_X1 FILLER_125_720 ();
 FILLCELL_X4 FILLER_125_728 ();
 FILLCELL_X4 FILLER_125_750 ();
 FILLCELL_X16 FILLER_125_773 ();
 FILLCELL_X1 FILLER_125_789 ();
 FILLCELL_X2 FILLER_125_803 ();
 FILLCELL_X1 FILLER_125_808 ();
 FILLCELL_X1 FILLER_125_819 ();
 FILLCELL_X2 FILLER_125_843 ();
 FILLCELL_X1 FILLER_125_845 ();
 FILLCELL_X4 FILLER_125_859 ();
 FILLCELL_X2 FILLER_125_863 ();
 FILLCELL_X1 FILLER_125_865 ();
 FILLCELL_X2 FILLER_125_901 ();
 FILLCELL_X1 FILLER_125_910 ();
 FILLCELL_X8 FILLER_125_931 ();
 FILLCELL_X2 FILLER_125_939 ();
 FILLCELL_X16 FILLER_125_944 ();
 FILLCELL_X8 FILLER_125_960 ();
 FILLCELL_X4 FILLER_125_984 ();
 FILLCELL_X2 FILLER_125_988 ();
 FILLCELL_X1 FILLER_125_995 ();
 FILLCELL_X2 FILLER_125_1012 ();
 FILLCELL_X8 FILLER_125_1021 ();
 FILLCELL_X2 FILLER_125_1029 ();
 FILLCELL_X8 FILLER_125_1038 ();
 FILLCELL_X2 FILLER_125_1046 ();
 FILLCELL_X1 FILLER_125_1114 ();
 FILLCELL_X2 FILLER_125_1118 ();
 FILLCELL_X2 FILLER_125_1127 ();
 FILLCELL_X1 FILLER_125_1129 ();
 FILLCELL_X16 FILLER_125_1137 ();
 FILLCELL_X8 FILLER_125_1153 ();
 FILLCELL_X4 FILLER_125_1161 ();
 FILLCELL_X1 FILLER_125_1192 ();
 FILLCELL_X2 FILLER_125_1200 ();
 FILLCELL_X32 FILLER_125_1226 ();
 FILLCELL_X2 FILLER_125_1258 ();
 FILLCELL_X8 FILLER_126_1 ();
 FILLCELL_X4 FILLER_126_9 ();
 FILLCELL_X2 FILLER_126_13 ();
 FILLCELL_X4 FILLER_126_35 ();
 FILLCELL_X2 FILLER_126_39 ();
 FILLCELL_X4 FILLER_126_48 ();
 FILLCELL_X1 FILLER_126_79 ();
 FILLCELL_X1 FILLER_126_87 ();
 FILLCELL_X1 FILLER_126_95 ();
 FILLCELL_X1 FILLER_126_103 ();
 FILLCELL_X16 FILLER_126_112 ();
 FILLCELL_X8 FILLER_126_128 ();
 FILLCELL_X4 FILLER_126_136 ();
 FILLCELL_X2 FILLER_126_140 ();
 FILLCELL_X4 FILLER_126_155 ();
 FILLCELL_X2 FILLER_126_159 ();
 FILLCELL_X1 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_210 ();
 FILLCELL_X8 FILLER_126_258 ();
 FILLCELL_X2 FILLER_126_266 ();
 FILLCELL_X2 FILLER_126_275 ();
 FILLCELL_X1 FILLER_126_277 ();
 FILLCELL_X8 FILLER_126_285 ();
 FILLCELL_X4 FILLER_126_293 ();
 FILLCELL_X1 FILLER_126_297 ();
 FILLCELL_X1 FILLER_126_321 ();
 FILLCELL_X2 FILLER_126_329 ();
 FILLCELL_X4 FILLER_126_334 ();
 FILLCELL_X2 FILLER_126_338 ();
 FILLCELL_X1 FILLER_126_340 ();
 FILLCELL_X4 FILLER_126_387 ();
 FILLCELL_X1 FILLER_126_391 ();
 FILLCELL_X1 FILLER_126_396 ();
 FILLCELL_X4 FILLER_126_400 ();
 FILLCELL_X2 FILLER_126_404 ();
 FILLCELL_X2 FILLER_126_416 ();
 FILLCELL_X1 FILLER_126_418 ();
 FILLCELL_X1 FILLER_126_426 ();
 FILLCELL_X4 FILLER_126_434 ();
 FILLCELL_X1 FILLER_126_438 ();
 FILLCELL_X8 FILLER_126_462 ();
 FILLCELL_X2 FILLER_126_470 ();
 FILLCELL_X1 FILLER_126_510 ();
 FILLCELL_X2 FILLER_126_571 ();
 FILLCELL_X2 FILLER_126_636 ();
 FILLCELL_X1 FILLER_126_647 ();
 FILLCELL_X8 FILLER_126_660 ();
 FILLCELL_X8 FILLER_126_726 ();
 FILLCELL_X1 FILLER_126_734 ();
 FILLCELL_X1 FILLER_126_746 ();
 FILLCELL_X8 FILLER_126_781 ();
 FILLCELL_X2 FILLER_126_789 ();
 FILLCELL_X1 FILLER_126_791 ();
 FILLCELL_X2 FILLER_126_802 ();
 FILLCELL_X1 FILLER_126_804 ();
 FILLCELL_X4 FILLER_126_819 ();
 FILLCELL_X2 FILLER_126_823 ();
 FILLCELL_X1 FILLER_126_825 ();
 FILLCELL_X4 FILLER_126_829 ();
 FILLCELL_X2 FILLER_126_833 ();
 FILLCELL_X8 FILLER_126_838 ();
 FILLCELL_X4 FILLER_126_846 ();
 FILLCELL_X2 FILLER_126_850 ();
 FILLCELL_X8 FILLER_126_862 ();
 FILLCELL_X4 FILLER_126_892 ();
 FILLCELL_X2 FILLER_126_896 ();
 FILLCELL_X1 FILLER_126_898 ();
 FILLCELL_X8 FILLER_126_902 ();
 FILLCELL_X4 FILLER_126_910 ();
 FILLCELL_X2 FILLER_126_926 ();
 FILLCELL_X1 FILLER_126_928 ();
 FILLCELL_X2 FILLER_126_954 ();
 FILLCELL_X1 FILLER_126_956 ();
 FILLCELL_X4 FILLER_126_975 ();
 FILLCELL_X2 FILLER_126_979 ();
 FILLCELL_X1 FILLER_126_981 ();
 FILLCELL_X2 FILLER_126_1006 ();
 FILLCELL_X1 FILLER_126_1008 ();
 FILLCELL_X2 FILLER_126_1016 ();
 FILLCELL_X1 FILLER_126_1018 ();
 FILLCELL_X2 FILLER_126_1029 ();
 FILLCELL_X1 FILLER_126_1031 ();
 FILLCELL_X8 FILLER_126_1035 ();
 FILLCELL_X8 FILLER_126_1052 ();
 FILLCELL_X4 FILLER_126_1060 ();
 FILLCELL_X1 FILLER_126_1064 ();
 FILLCELL_X2 FILLER_126_1084 ();
 FILLCELL_X4 FILLER_126_1090 ();
 FILLCELL_X2 FILLER_126_1114 ();
 FILLCELL_X1 FILLER_126_1116 ();
 FILLCELL_X4 FILLER_126_1121 ();
 FILLCELL_X2 FILLER_126_1125 ();
 FILLCELL_X16 FILLER_126_1168 ();
 FILLCELL_X2 FILLER_126_1184 ();
 FILLCELL_X2 FILLER_126_1193 ();
 FILLCELL_X1 FILLER_126_1195 ();
 FILLCELL_X32 FILLER_126_1203 ();
 FILLCELL_X16 FILLER_126_1235 ();
 FILLCELL_X8 FILLER_126_1251 ();
 FILLCELL_X1 FILLER_126_1259 ();
 FILLCELL_X4 FILLER_127_21 ();
 FILLCELL_X2 FILLER_127_25 ();
 FILLCELL_X2 FILLER_127_41 ();
 FILLCELL_X1 FILLER_127_43 ();
 FILLCELL_X4 FILLER_127_56 ();
 FILLCELL_X1 FILLER_127_60 ();
 FILLCELL_X2 FILLER_127_68 ();
 FILLCELL_X1 FILLER_127_70 ();
 FILLCELL_X2 FILLER_127_98 ();
 FILLCELL_X1 FILLER_127_100 ();
 FILLCELL_X2 FILLER_127_143 ();
 FILLCELL_X2 FILLER_127_152 ();
 FILLCELL_X2 FILLER_127_174 ();
 FILLCELL_X1 FILLER_127_176 ();
 FILLCELL_X4 FILLER_127_195 ();
 FILLCELL_X2 FILLER_127_199 ();
 FILLCELL_X1 FILLER_127_201 ();
 FILLCELL_X1 FILLER_127_205 ();
 FILLCELL_X2 FILLER_127_215 ();
 FILLCELL_X4 FILLER_127_235 ();
 FILLCELL_X1 FILLER_127_239 ();
 FILLCELL_X4 FILLER_127_298 ();
 FILLCELL_X1 FILLER_127_302 ();
 FILLCELL_X2 FILLER_127_307 ();
 FILLCELL_X2 FILLER_127_312 ();
 FILLCELL_X1 FILLER_127_314 ();
 FILLCELL_X2 FILLER_127_319 ();
 FILLCELL_X1 FILLER_127_321 ();
 FILLCELL_X2 FILLER_127_329 ();
 FILLCELL_X1 FILLER_127_344 ();
 FILLCELL_X2 FILLER_127_356 ();
 FILLCELL_X1 FILLER_127_358 ();
 FILLCELL_X1 FILLER_127_376 ();
 FILLCELL_X2 FILLER_127_400 ();
 FILLCELL_X1 FILLER_127_402 ();
 FILLCELL_X1 FILLER_127_424 ();
 FILLCELL_X4 FILLER_127_435 ();
 FILLCELL_X2 FILLER_127_439 ();
 FILLCELL_X1 FILLER_127_441 ();
 FILLCELL_X2 FILLER_127_463 ();
 FILLCELL_X2 FILLER_127_470 ();
 FILLCELL_X2 FILLER_127_475 ();
 FILLCELL_X8 FILLER_127_606 ();
 FILLCELL_X2 FILLER_127_614 ();
 FILLCELL_X2 FILLER_127_644 ();
 FILLCELL_X4 FILLER_127_666 ();
 FILLCELL_X2 FILLER_127_670 ();
 FILLCELL_X1 FILLER_127_687 ();
 FILLCELL_X1 FILLER_127_695 ();
 FILLCELL_X2 FILLER_127_699 ();
 FILLCELL_X4 FILLER_127_706 ();
 FILLCELL_X8 FILLER_127_731 ();
 FILLCELL_X2 FILLER_127_739 ();
 FILLCELL_X16 FILLER_127_783 ();
 FILLCELL_X8 FILLER_127_799 ();
 FILLCELL_X2 FILLER_127_807 ();
 FILLCELL_X1 FILLER_127_834 ();
 FILLCELL_X4 FILLER_127_840 ();
 FILLCELL_X1 FILLER_127_844 ();
 FILLCELL_X2 FILLER_127_871 ();
 FILLCELL_X1 FILLER_127_873 ();
 FILLCELL_X2 FILLER_127_878 ();
 FILLCELL_X2 FILLER_127_900 ();
 FILLCELL_X1 FILLER_127_902 ();
 FILLCELL_X2 FILLER_127_912 ();
 FILLCELL_X1 FILLER_127_914 ();
 FILLCELL_X2 FILLER_127_918 ();
 FILLCELL_X1 FILLER_127_940 ();
 FILLCELL_X1 FILLER_127_958 ();
 FILLCELL_X8 FILLER_127_973 ();
 FILLCELL_X1 FILLER_127_981 ();
 FILLCELL_X2 FILLER_127_998 ();
 FILLCELL_X1 FILLER_127_1000 ();
 FILLCELL_X8 FILLER_127_1011 ();
 FILLCELL_X4 FILLER_127_1019 ();
 FILLCELL_X1 FILLER_127_1023 ();
 FILLCELL_X1 FILLER_127_1050 ();
 FILLCELL_X2 FILLER_127_1054 ();
 FILLCELL_X1 FILLER_127_1060 ();
 FILLCELL_X2 FILLER_127_1065 ();
 FILLCELL_X2 FILLER_127_1076 ();
 FILLCELL_X2 FILLER_127_1087 ();
 FILLCELL_X16 FILLER_127_1133 ();
 FILLCELL_X4 FILLER_127_1149 ();
 FILLCELL_X4 FILLER_127_1187 ();
 FILLCELL_X1 FILLER_127_1191 ();
 FILLCELL_X32 FILLER_127_1226 ();
 FILLCELL_X2 FILLER_127_1258 ();
 FILLCELL_X4 FILLER_128_1 ();
 FILLCELL_X2 FILLER_128_5 ();
 FILLCELL_X1 FILLER_128_7 ();
 FILLCELL_X16 FILLER_128_49 ();
 FILLCELL_X2 FILLER_128_65 ();
 FILLCELL_X4 FILLER_128_94 ();
 FILLCELL_X1 FILLER_128_98 ();
 FILLCELL_X1 FILLER_128_119 ();
 FILLCELL_X2 FILLER_128_165 ();
 FILLCELL_X2 FILLER_128_169 ();
 FILLCELL_X1 FILLER_128_171 ();
 FILLCELL_X2 FILLER_128_177 ();
 FILLCELL_X1 FILLER_128_179 ();
 FILLCELL_X2 FILLER_128_186 ();
 FILLCELL_X1 FILLER_128_188 ();
 FILLCELL_X1 FILLER_128_200 ();
 FILLCELL_X2 FILLER_128_204 ();
 FILLCELL_X2 FILLER_128_219 ();
 FILLCELL_X16 FILLER_128_250 ();
 FILLCELL_X4 FILLER_128_266 ();
 FILLCELL_X16 FILLER_128_277 ();
 FILLCELL_X1 FILLER_128_293 ();
 FILLCELL_X2 FILLER_128_335 ();
 FILLCELL_X4 FILLER_128_341 ();
 FILLCELL_X2 FILLER_128_345 ();
 FILLCELL_X1 FILLER_128_347 ();
 FILLCELL_X4 FILLER_128_355 ();
 FILLCELL_X2 FILLER_128_359 ();
 FILLCELL_X2 FILLER_128_371 ();
 FILLCELL_X2 FILLER_128_377 ();
 FILLCELL_X16 FILLER_128_384 ();
 FILLCELL_X4 FILLER_128_400 ();
 FILLCELL_X4 FILLER_128_456 ();
 FILLCELL_X1 FILLER_128_460 ();
 FILLCELL_X2 FILLER_128_481 ();
 FILLCELL_X4 FILLER_128_505 ();
 FILLCELL_X1 FILLER_128_533 ();
 FILLCELL_X2 FILLER_128_537 ();
 FILLCELL_X2 FILLER_128_560 ();
 FILLCELL_X1 FILLER_128_592 ();
 FILLCELL_X4 FILLER_128_613 ();
 FILLCELL_X2 FILLER_128_617 ();
 FILLCELL_X8 FILLER_128_622 ();
 FILLCELL_X1 FILLER_128_630 ();
 FILLCELL_X8 FILLER_128_632 ();
 FILLCELL_X2 FILLER_128_640 ();
 FILLCELL_X1 FILLER_128_642 ();
 FILLCELL_X16 FILLER_128_646 ();
 FILLCELL_X8 FILLER_128_662 ();
 FILLCELL_X2 FILLER_128_670 ();
 FILLCELL_X1 FILLER_128_672 ();
 FILLCELL_X1 FILLER_128_680 ();
 FILLCELL_X4 FILLER_128_701 ();
 FILLCELL_X2 FILLER_128_705 ();
 FILLCELL_X1 FILLER_128_707 ();
 FILLCELL_X2 FILLER_128_733 ();
 FILLCELL_X2 FILLER_128_751 ();
 FILLCELL_X2 FILLER_128_756 ();
 FILLCELL_X2 FILLER_128_782 ();
 FILLCELL_X4 FILLER_128_804 ();
 FILLCELL_X2 FILLER_128_822 ();
 FILLCELL_X4 FILLER_128_826 ();
 FILLCELL_X4 FILLER_128_844 ();
 FILLCELL_X2 FILLER_128_848 ();
 FILLCELL_X8 FILLER_128_855 ();
 FILLCELL_X1 FILLER_128_863 ();
 FILLCELL_X4 FILLER_128_869 ();
 FILLCELL_X2 FILLER_128_883 ();
 FILLCELL_X4 FILLER_128_888 ();
 FILLCELL_X1 FILLER_128_892 ();
 FILLCELL_X2 FILLER_128_901 ();
 FILLCELL_X1 FILLER_128_903 ();
 FILLCELL_X2 FILLER_128_911 ();
 FILLCELL_X1 FILLER_128_917 ();
 FILLCELL_X4 FILLER_128_932 ();
 FILLCELL_X1 FILLER_128_943 ();
 FILLCELL_X1 FILLER_128_958 ();
 FILLCELL_X1 FILLER_128_973 ();
 FILLCELL_X2 FILLER_128_981 ();
 FILLCELL_X4 FILLER_128_994 ();
 FILLCELL_X2 FILLER_128_998 ();
 FILLCELL_X1 FILLER_128_1000 ();
 FILLCELL_X2 FILLER_128_1022 ();
 FILLCELL_X1 FILLER_128_1032 ();
 FILLCELL_X1 FILLER_128_1046 ();
 FILLCELL_X1 FILLER_128_1051 ();
 FILLCELL_X1 FILLER_128_1056 ();
 FILLCELL_X8 FILLER_128_1078 ();
 FILLCELL_X4 FILLER_128_1086 ();
 FILLCELL_X2 FILLER_128_1117 ();
 FILLCELL_X2 FILLER_128_1138 ();
 FILLCELL_X1 FILLER_128_1140 ();
 FILLCELL_X4 FILLER_128_1148 ();
 FILLCELL_X2 FILLER_128_1152 ();
 FILLCELL_X1 FILLER_128_1154 ();
 FILLCELL_X1 FILLER_128_1175 ();
 FILLCELL_X2 FILLER_128_1203 ();
 FILLCELL_X1 FILLER_128_1205 ();
 FILLCELL_X32 FILLER_128_1226 ();
 FILLCELL_X2 FILLER_128_1258 ();
 FILLCELL_X4 FILLER_129_21 ();
 FILLCELL_X2 FILLER_129_25 ();
 FILLCELL_X2 FILLER_129_41 ();
 FILLCELL_X16 FILLER_129_50 ();
 FILLCELL_X8 FILLER_129_66 ();
 FILLCELL_X2 FILLER_129_74 ();
 FILLCELL_X2 FILLER_129_83 ();
 FILLCELL_X1 FILLER_129_85 ();
 FILLCELL_X8 FILLER_129_93 ();
 FILLCELL_X2 FILLER_129_101 ();
 FILLCELL_X4 FILLER_129_110 ();
 FILLCELL_X2 FILLER_129_114 ();
 FILLCELL_X1 FILLER_129_116 ();
 FILLCELL_X1 FILLER_129_131 ();
 FILLCELL_X1 FILLER_129_139 ();
 FILLCELL_X1 FILLER_129_151 ();
 FILLCELL_X4 FILLER_129_182 ();
 FILLCELL_X1 FILLER_129_186 ();
 FILLCELL_X32 FILLER_129_201 ();
 FILLCELL_X1 FILLER_129_236 ();
 FILLCELL_X2 FILLER_129_244 ();
 FILLCELL_X1 FILLER_129_246 ();
 FILLCELL_X4 FILLER_129_274 ();
 FILLCELL_X1 FILLER_129_278 ();
 FILLCELL_X2 FILLER_129_286 ();
 FILLCELL_X1 FILLER_129_288 ();
 FILLCELL_X8 FILLER_129_291 ();
 FILLCELL_X2 FILLER_129_299 ();
 FILLCELL_X1 FILLER_129_301 ();
 FILLCELL_X4 FILLER_129_329 ();
 FILLCELL_X2 FILLER_129_333 ();
 FILLCELL_X1 FILLER_129_335 ();
 FILLCELL_X2 FILLER_129_340 ();
 FILLCELL_X1 FILLER_129_345 ();
 FILLCELL_X1 FILLER_129_366 ();
 FILLCELL_X4 FILLER_129_407 ();
 FILLCELL_X8 FILLER_129_415 ();
 FILLCELL_X2 FILLER_129_423 ();
 FILLCELL_X2 FILLER_129_436 ();
 FILLCELL_X4 FILLER_129_440 ();
 FILLCELL_X2 FILLER_129_444 ();
 FILLCELL_X2 FILLER_129_453 ();
 FILLCELL_X1 FILLER_129_455 ();
 FILLCELL_X2 FILLER_129_460 ();
 FILLCELL_X8 FILLER_129_469 ();
 FILLCELL_X1 FILLER_129_477 ();
 FILLCELL_X2 FILLER_129_520 ();
 FILLCELL_X4 FILLER_129_565 ();
 FILLCELL_X8 FILLER_129_595 ();
 FILLCELL_X2 FILLER_129_603 ();
 FILLCELL_X2 FILLER_129_619 ();
 FILLCELL_X8 FILLER_129_628 ();
 FILLCELL_X1 FILLER_129_636 ();
 FILLCELL_X4 FILLER_129_644 ();
 FILLCELL_X4 FILLER_129_655 ();
 FILLCELL_X1 FILLER_129_659 ();
 FILLCELL_X1 FILLER_129_680 ();
 FILLCELL_X4 FILLER_129_697 ();
 FILLCELL_X2 FILLER_129_701 ();
 FILLCELL_X1 FILLER_129_703 ();
 FILLCELL_X2 FILLER_129_717 ();
 FILLCELL_X2 FILLER_129_737 ();
 FILLCELL_X1 FILLER_129_739 ();
 FILLCELL_X2 FILLER_129_755 ();
 FILLCELL_X4 FILLER_129_761 ();
 FILLCELL_X4 FILLER_129_768 ();
 FILLCELL_X2 FILLER_129_772 ();
 FILLCELL_X4 FILLER_129_798 ();
 FILLCELL_X2 FILLER_129_819 ();
 FILLCELL_X1 FILLER_129_821 ();
 FILLCELL_X8 FILLER_129_847 ();
 FILLCELL_X2 FILLER_129_855 ();
 FILLCELL_X4 FILLER_129_892 ();
 FILLCELL_X1 FILLER_129_901 ();
 FILLCELL_X4 FILLER_129_905 ();
 FILLCELL_X2 FILLER_129_909 ();
 FILLCELL_X2 FILLER_129_916 ();
 FILLCELL_X4 FILLER_129_932 ();
 FILLCELL_X2 FILLER_129_936 ();
 FILLCELL_X1 FILLER_129_938 ();
 FILLCELL_X8 FILLER_129_949 ();
 FILLCELL_X2 FILLER_129_957 ();
 FILLCELL_X8 FILLER_129_966 ();
 FILLCELL_X4 FILLER_129_974 ();
 FILLCELL_X4 FILLER_129_987 ();
 FILLCELL_X8 FILLER_129_996 ();
 FILLCELL_X8 FILLER_129_1008 ();
 FILLCELL_X2 FILLER_129_1016 ();
 FILLCELL_X1 FILLER_129_1022 ();
 FILLCELL_X4 FILLER_129_1040 ();
 FILLCELL_X2 FILLER_129_1044 ();
 FILLCELL_X1 FILLER_129_1046 ();
 FILLCELL_X1 FILLER_129_1060 ();
 FILLCELL_X16 FILLER_129_1078 ();
 FILLCELL_X8 FILLER_129_1094 ();
 FILLCELL_X4 FILLER_129_1102 ();
 FILLCELL_X1 FILLER_129_1106 ();
 FILLCELL_X16 FILLER_129_1139 ();
 FILLCELL_X2 FILLER_129_1155 ();
 FILLCELL_X1 FILLER_129_1157 ();
 FILLCELL_X4 FILLER_129_1173 ();
 FILLCELL_X2 FILLER_129_1177 ();
 FILLCELL_X1 FILLER_129_1179 ();
 FILLCELL_X8 FILLER_129_1187 ();
 FILLCELL_X2 FILLER_129_1195 ();
 FILLCELL_X32 FILLER_129_1211 ();
 FILLCELL_X16 FILLER_129_1243 ();
 FILLCELL_X1 FILLER_129_1259 ();
 FILLCELL_X4 FILLER_130_1 ();
 FILLCELL_X2 FILLER_130_5 ();
 FILLCELL_X1 FILLER_130_7 ();
 FILLCELL_X8 FILLER_130_49 ();
 FILLCELL_X1 FILLER_130_57 ();
 FILLCELL_X8 FILLER_130_105 ();
 FILLCELL_X1 FILLER_130_113 ();
 FILLCELL_X4 FILLER_130_121 ();
 FILLCELL_X2 FILLER_130_152 ();
 FILLCELL_X8 FILLER_130_163 ();
 FILLCELL_X2 FILLER_130_171 ();
 FILLCELL_X1 FILLER_130_173 ();
 FILLCELL_X1 FILLER_130_191 ();
 FILLCELL_X4 FILLER_130_244 ();
 FILLCELL_X2 FILLER_130_248 ();
 FILLCELL_X2 FILLER_130_277 ();
 FILLCELL_X1 FILLER_130_279 ();
 FILLCELL_X2 FILLER_130_300 ();
 FILLCELL_X8 FILLER_130_312 ();
 FILLCELL_X2 FILLER_130_327 ();
 FILLCELL_X1 FILLER_130_329 ();
 FILLCELL_X8 FILLER_130_350 ();
 FILLCELL_X4 FILLER_130_358 ();
 FILLCELL_X2 FILLER_130_362 ();
 FILLCELL_X4 FILLER_130_374 ();
 FILLCELL_X2 FILLER_130_378 ();
 FILLCELL_X1 FILLER_130_380 ();
 FILLCELL_X1 FILLER_130_417 ();
 FILLCELL_X4 FILLER_130_445 ();
 FILLCELL_X1 FILLER_130_449 ();
 FILLCELL_X8 FILLER_130_457 ();
 FILLCELL_X2 FILLER_130_465 ();
 FILLCELL_X16 FILLER_130_471 ();
 FILLCELL_X8 FILLER_130_487 ();
 FILLCELL_X2 FILLER_130_495 ();
 FILLCELL_X2 FILLER_130_517 ();
 FILLCELL_X8 FILLER_130_533 ();
 FILLCELL_X2 FILLER_130_541 ();
 FILLCELL_X4 FILLER_130_561 ();
 FILLCELL_X2 FILLER_130_568 ();
 FILLCELL_X1 FILLER_130_570 ();
 FILLCELL_X8 FILLER_130_578 ();
 FILLCELL_X4 FILLER_130_586 ();
 FILLCELL_X2 FILLER_130_594 ();
 FILLCELL_X1 FILLER_130_596 ();
 FILLCELL_X4 FILLER_130_600 ();
 FILLCELL_X2 FILLER_130_632 ();
 FILLCELL_X1 FILLER_130_634 ();
 FILLCELL_X2 FILLER_130_642 ();
 FILLCELL_X8 FILLER_130_664 ();
 FILLCELL_X4 FILLER_130_684 ();
 FILLCELL_X4 FILLER_130_699 ();
 FILLCELL_X2 FILLER_130_703 ();
 FILLCELL_X16 FILLER_130_712 ();
 FILLCELL_X4 FILLER_130_761 ();
 FILLCELL_X1 FILLER_130_765 ();
 FILLCELL_X4 FILLER_130_793 ();
 FILLCELL_X1 FILLER_130_797 ();
 FILLCELL_X4 FILLER_130_805 ();
 FILLCELL_X1 FILLER_130_809 ();
 FILLCELL_X4 FILLER_130_838 ();
 FILLCELL_X2 FILLER_130_842 ();
 FILLCELL_X1 FILLER_130_844 ();
 FILLCELL_X2 FILLER_130_853 ();
 FILLCELL_X1 FILLER_130_863 ();
 FILLCELL_X4 FILLER_130_879 ();
 FILLCELL_X1 FILLER_130_890 ();
 FILLCELL_X2 FILLER_130_933 ();
 FILLCELL_X1 FILLER_130_935 ();
 FILLCELL_X8 FILLER_130_970 ();
 FILLCELL_X4 FILLER_130_978 ();
 FILLCELL_X2 FILLER_130_982 ();
 FILLCELL_X1 FILLER_130_984 ();
 FILLCELL_X4 FILLER_130_993 ();
 FILLCELL_X2 FILLER_130_1010 ();
 FILLCELL_X4 FILLER_130_1021 ();
 FILLCELL_X2 FILLER_130_1025 ();
 FILLCELL_X16 FILLER_130_1043 ();
 FILLCELL_X2 FILLER_130_1059 ();
 FILLCELL_X2 FILLER_130_1078 ();
 FILLCELL_X16 FILLER_130_1089 ();
 FILLCELL_X2 FILLER_130_1105 ();
 FILLCELL_X16 FILLER_130_1112 ();
 FILLCELL_X1 FILLER_130_1128 ();
 FILLCELL_X1 FILLER_130_1183 ();
 FILLCELL_X32 FILLER_130_1211 ();
 FILLCELL_X16 FILLER_130_1243 ();
 FILLCELL_X1 FILLER_130_1259 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X2 FILLER_131_33 ();
 FILLCELL_X1 FILLER_131_35 ();
 FILLCELL_X16 FILLER_131_43 ();
 FILLCELL_X8 FILLER_131_59 ();
 FILLCELL_X2 FILLER_131_67 ();
 FILLCELL_X16 FILLER_131_96 ();
 FILLCELL_X2 FILLER_131_112 ();
 FILLCELL_X1 FILLER_131_114 ();
 FILLCELL_X1 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_137 ();
 FILLCELL_X4 FILLER_131_169 ();
 FILLCELL_X2 FILLER_131_173 ();
 FILLCELL_X1 FILLER_131_175 ();
 FILLCELL_X4 FILLER_131_191 ();
 FILLCELL_X2 FILLER_131_195 ();
 FILLCELL_X4 FILLER_131_204 ();
 FILLCELL_X2 FILLER_131_208 ();
 FILLCELL_X1 FILLER_131_210 ();
 FILLCELL_X1 FILLER_131_223 ();
 FILLCELL_X2 FILLER_131_231 ();
 FILLCELL_X16 FILLER_131_240 ();
 FILLCELL_X4 FILLER_131_256 ();
 FILLCELL_X2 FILLER_131_260 ();
 FILLCELL_X2 FILLER_131_286 ();
 FILLCELL_X1 FILLER_131_291 ();
 FILLCELL_X1 FILLER_131_312 ();
 FILLCELL_X1 FILLER_131_336 ();
 FILLCELL_X8 FILLER_131_344 ();
 FILLCELL_X4 FILLER_131_352 ();
 FILLCELL_X2 FILLER_131_356 ();
 FILLCELL_X4 FILLER_131_376 ();
 FILLCELL_X2 FILLER_131_380 ();
 FILLCELL_X2 FILLER_131_386 ();
 FILLCELL_X2 FILLER_131_392 ();
 FILLCELL_X2 FILLER_131_397 ();
 FILLCELL_X1 FILLER_131_402 ();
 FILLCELL_X1 FILLER_131_407 ();
 FILLCELL_X2 FILLER_131_411 ();
 FILLCELL_X4 FILLER_131_436 ();
 FILLCELL_X1 FILLER_131_440 ();
 FILLCELL_X4 FILLER_131_448 ();
 FILLCELL_X1 FILLER_131_452 ();
 FILLCELL_X1 FILLER_131_473 ();
 FILLCELL_X2 FILLER_131_497 ();
 FILLCELL_X2 FILLER_131_506 ();
 FILLCELL_X2 FILLER_131_616 ();
 FILLCELL_X1 FILLER_131_618 ();
 FILLCELL_X2 FILLER_131_656 ();
 FILLCELL_X1 FILLER_131_658 ();
 FILLCELL_X4 FILLER_131_662 ();
 FILLCELL_X8 FILLER_131_693 ();
 FILLCELL_X2 FILLER_131_701 ();
 FILLCELL_X16 FILLER_131_730 ();
 FILLCELL_X8 FILLER_131_746 ();
 FILLCELL_X1 FILLER_131_754 ();
 FILLCELL_X2 FILLER_131_779 ();
 FILLCELL_X1 FILLER_131_781 ();
 FILLCELL_X16 FILLER_131_785 ();
 FILLCELL_X8 FILLER_131_801 ();
 FILLCELL_X2 FILLER_131_809 ();
 FILLCELL_X1 FILLER_131_811 ();
 FILLCELL_X2 FILLER_131_819 ();
 FILLCELL_X1 FILLER_131_821 ();
 FILLCELL_X2 FILLER_131_825 ();
 FILLCELL_X1 FILLER_131_827 ();
 FILLCELL_X4 FILLER_131_840 ();
 FILLCELL_X1 FILLER_131_844 ();
 FILLCELL_X4 FILLER_131_850 ();
 FILLCELL_X1 FILLER_131_854 ();
 FILLCELL_X1 FILLER_131_865 ();
 FILLCELL_X2 FILLER_131_873 ();
 FILLCELL_X2 FILLER_131_884 ();
 FILLCELL_X2 FILLER_131_893 ();
 FILLCELL_X16 FILLER_131_902 ();
 FILLCELL_X2 FILLER_131_918 ();
 FILLCELL_X1 FILLER_131_920 ();
 FILLCELL_X2 FILLER_131_927 ();
 FILLCELL_X2 FILLER_131_956 ();
 FILLCELL_X1 FILLER_131_958 ();
 FILLCELL_X1 FILLER_131_983 ();
 FILLCELL_X1 FILLER_131_994 ();
 FILLCELL_X1 FILLER_131_1000 ();
 FILLCELL_X4 FILLER_131_1008 ();
 FILLCELL_X2 FILLER_131_1012 ();
 FILLCELL_X1 FILLER_131_1026 ();
 FILLCELL_X1 FILLER_131_1031 ();
 FILLCELL_X4 FILLER_131_1039 ();
 FILLCELL_X1 FILLER_131_1043 ();
 FILLCELL_X1 FILLER_131_1066 ();
 FILLCELL_X2 FILLER_131_1072 ();
 FILLCELL_X1 FILLER_131_1074 ();
 FILLCELL_X2 FILLER_131_1084 ();
 FILLCELL_X2 FILLER_131_1108 ();
 FILLCELL_X8 FILLER_131_1114 ();
 FILLCELL_X4 FILLER_131_1122 ();
 FILLCELL_X1 FILLER_131_1126 ();
 FILLCELL_X32 FILLER_131_1146 ();
 FILLCELL_X32 FILLER_131_1178 ();
 FILLCELL_X32 FILLER_131_1210 ();
 FILLCELL_X16 FILLER_131_1242 ();
 FILLCELL_X2 FILLER_131_1258 ();
 FILLCELL_X16 FILLER_132_1 ();
 FILLCELL_X4 FILLER_132_44 ();
 FILLCELL_X2 FILLER_132_48 ();
 FILLCELL_X8 FILLER_132_57 ();
 FILLCELL_X1 FILLER_132_65 ();
 FILLCELL_X2 FILLER_132_113 ();
 FILLCELL_X2 FILLER_132_132 ();
 FILLCELL_X2 FILLER_132_138 ();
 FILLCELL_X1 FILLER_132_140 ();
 FILLCELL_X2 FILLER_132_148 ();
 FILLCELL_X1 FILLER_132_150 ();
 FILLCELL_X8 FILLER_132_160 ();
 FILLCELL_X4 FILLER_132_168 ();
 FILLCELL_X2 FILLER_132_172 ();
 FILLCELL_X2 FILLER_132_223 ();
 FILLCELL_X2 FILLER_132_245 ();
 FILLCELL_X1 FILLER_132_247 ();
 FILLCELL_X1 FILLER_132_268 ();
 FILLCELL_X2 FILLER_132_276 ();
 FILLCELL_X1 FILLER_132_278 ();
 FILLCELL_X1 FILLER_132_282 ();
 FILLCELL_X2 FILLER_132_291 ();
 FILLCELL_X8 FILLER_132_302 ();
 FILLCELL_X2 FILLER_132_310 ();
 FILLCELL_X1 FILLER_132_312 ();
 FILLCELL_X1 FILLER_132_327 ();
 FILLCELL_X2 FILLER_132_335 ();
 FILLCELL_X1 FILLER_132_337 ();
 FILLCELL_X2 FILLER_132_370 ();
 FILLCELL_X2 FILLER_132_376 ();
 FILLCELL_X1 FILLER_132_378 ();
 FILLCELL_X1 FILLER_132_390 ();
 FILLCELL_X2 FILLER_132_401 ();
 FILLCELL_X1 FILLER_132_425 ();
 FILLCELL_X4 FILLER_132_429 ();
 FILLCELL_X16 FILLER_132_436 ();
 FILLCELL_X1 FILLER_132_452 ();
 FILLCELL_X8 FILLER_132_456 ();
 FILLCELL_X2 FILLER_132_464 ();
 FILLCELL_X4 FILLER_132_473 ();
 FILLCELL_X2 FILLER_132_477 ();
 FILLCELL_X2 FILLER_132_496 ();
 FILLCELL_X8 FILLER_132_521 ();
 FILLCELL_X2 FILLER_132_536 ();
 FILLCELL_X1 FILLER_132_538 ();
 FILLCELL_X2 FILLER_132_553 ();
 FILLCELL_X1 FILLER_132_555 ();
 FILLCELL_X1 FILLER_132_560 ();
 FILLCELL_X16 FILLER_132_564 ();
 FILLCELL_X4 FILLER_132_580 ();
 FILLCELL_X2 FILLER_132_584 ();
 FILLCELL_X1 FILLER_132_586 ();
 FILLCELL_X4 FILLER_132_600 ();
 FILLCELL_X1 FILLER_132_604 ();
 FILLCELL_X2 FILLER_132_619 ();
 FILLCELL_X1 FILLER_132_621 ();
 FILLCELL_X4 FILLER_132_626 ();
 FILLCELL_X1 FILLER_132_630 ();
 FILLCELL_X1 FILLER_132_662 ();
 FILLCELL_X8 FILLER_132_667 ();
 FILLCELL_X1 FILLER_132_675 ();
 FILLCELL_X2 FILLER_132_730 ();
 FILLCELL_X1 FILLER_132_739 ();
 FILLCELL_X8 FILLER_132_743 ();
 FILLCELL_X2 FILLER_132_751 ();
 FILLCELL_X1 FILLER_132_753 ();
 FILLCELL_X4 FILLER_132_770 ();
 FILLCELL_X2 FILLER_132_774 ();
 FILLCELL_X1 FILLER_132_804 ();
 FILLCELL_X16 FILLER_132_822 ();
 FILLCELL_X8 FILLER_132_838 ();
 FILLCELL_X2 FILLER_132_846 ();
 FILLCELL_X1 FILLER_132_848 ();
 FILLCELL_X1 FILLER_132_889 ();
 FILLCELL_X1 FILLER_132_897 ();
 FILLCELL_X4 FILLER_132_942 ();
 FILLCELL_X1 FILLER_132_966 ();
 FILLCELL_X4 FILLER_132_974 ();
 FILLCELL_X2 FILLER_132_978 ();
 FILLCELL_X1 FILLER_132_980 ();
 FILLCELL_X2 FILLER_132_989 ();
 FILLCELL_X1 FILLER_132_991 ();
 FILLCELL_X4 FILLER_132_1038 ();
 FILLCELL_X2 FILLER_132_1042 ();
 FILLCELL_X4 FILLER_132_1054 ();
 FILLCELL_X2 FILLER_132_1058 ();
 FILLCELL_X1 FILLER_132_1060 ();
 FILLCELL_X1 FILLER_132_1071 ();
 FILLCELL_X8 FILLER_132_1076 ();
 FILLCELL_X4 FILLER_132_1084 ();
 FILLCELL_X4 FILLER_132_1095 ();
 FILLCELL_X1 FILLER_132_1099 ();
 FILLCELL_X1 FILLER_132_1102 ();
 FILLCELL_X4 FILLER_132_1113 ();
 FILLCELL_X2 FILLER_132_1117 ();
 FILLCELL_X1 FILLER_132_1119 ();
 FILLCELL_X4 FILLER_132_1136 ();
 FILLCELL_X2 FILLER_132_1140 ();
 FILLCELL_X1 FILLER_132_1142 ();
 FILLCELL_X32 FILLER_132_1164 ();
 FILLCELL_X32 FILLER_132_1196 ();
 FILLCELL_X32 FILLER_132_1228 ();
 FILLCELL_X4 FILLER_133_28 ();
 FILLCELL_X1 FILLER_133_32 ();
 FILLCELL_X1 FILLER_133_47 ();
 FILLCELL_X4 FILLER_133_89 ();
 FILLCELL_X1 FILLER_133_93 ();
 FILLCELL_X2 FILLER_133_127 ();
 FILLCELL_X1 FILLER_133_173 ();
 FILLCELL_X2 FILLER_133_195 ();
 FILLCELL_X1 FILLER_133_204 ();
 FILLCELL_X2 FILLER_133_225 ();
 FILLCELL_X4 FILLER_133_244 ();
 FILLCELL_X1 FILLER_133_248 ();
 FILLCELL_X1 FILLER_133_256 ();
 FILLCELL_X2 FILLER_133_264 ();
 FILLCELL_X1 FILLER_133_297 ();
 FILLCELL_X1 FILLER_133_302 ();
 FILLCELL_X1 FILLER_133_326 ();
 FILLCELL_X4 FILLER_133_337 ();
 FILLCELL_X2 FILLER_133_341 ();
 FILLCELL_X1 FILLER_133_343 ();
 FILLCELL_X2 FILLER_133_347 ();
 FILLCELL_X4 FILLER_133_353 ();
 FILLCELL_X2 FILLER_133_357 ();
 FILLCELL_X2 FILLER_133_370 ();
 FILLCELL_X1 FILLER_133_372 ();
 FILLCELL_X4 FILLER_133_384 ();
 FILLCELL_X2 FILLER_133_388 ();
 FILLCELL_X1 FILLER_133_390 ();
 FILLCELL_X4 FILLER_133_413 ();
 FILLCELL_X8 FILLER_133_436 ();
 FILLCELL_X1 FILLER_133_444 ();
 FILLCELL_X4 FILLER_133_517 ();
 FILLCELL_X1 FILLER_133_521 ();
 FILLCELL_X2 FILLER_133_542 ();
 FILLCELL_X1 FILLER_133_544 ();
 FILLCELL_X1 FILLER_133_572 ();
 FILLCELL_X16 FILLER_133_607 ();
 FILLCELL_X4 FILLER_133_623 ();
 FILLCELL_X1 FILLER_133_627 ();
 FILLCELL_X8 FILLER_133_642 ();
 FILLCELL_X2 FILLER_133_650 ();
 FILLCELL_X16 FILLER_133_659 ();
 FILLCELL_X8 FILLER_133_675 ();
 FILLCELL_X4 FILLER_133_683 ();
 FILLCELL_X1 FILLER_133_687 ();
 FILLCELL_X8 FILLER_133_691 ();
 FILLCELL_X4 FILLER_133_699 ();
 FILLCELL_X1 FILLER_133_730 ();
 FILLCELL_X1 FILLER_133_751 ();
 FILLCELL_X2 FILLER_133_759 ();
 FILLCELL_X2 FILLER_133_807 ();
 FILLCELL_X1 FILLER_133_809 ();
 FILLCELL_X4 FILLER_133_817 ();
 FILLCELL_X1 FILLER_133_821 ();
 FILLCELL_X1 FILLER_133_836 ();
 FILLCELL_X4 FILLER_133_853 ();
 FILLCELL_X2 FILLER_133_857 ();
 FILLCELL_X1 FILLER_133_859 ();
 FILLCELL_X8 FILLER_133_867 ();
 FILLCELL_X4 FILLER_133_875 ();
 FILLCELL_X2 FILLER_133_879 ();
 FILLCELL_X8 FILLER_133_896 ();
 FILLCELL_X4 FILLER_133_915 ();
 FILLCELL_X1 FILLER_133_919 ();
 FILLCELL_X1 FILLER_133_932 ();
 FILLCELL_X16 FILLER_133_940 ();
 FILLCELL_X1 FILLER_133_960 ();
 FILLCELL_X8 FILLER_133_968 ();
 FILLCELL_X2 FILLER_133_976 ();
 FILLCELL_X1 FILLER_133_978 ();
 FILLCELL_X2 FILLER_133_983 ();
 FILLCELL_X4 FILLER_133_989 ();
 FILLCELL_X2 FILLER_133_993 ();
 FILLCELL_X8 FILLER_133_1000 ();
 FILLCELL_X1 FILLER_133_1023 ();
 FILLCELL_X4 FILLER_133_1041 ();
 FILLCELL_X2 FILLER_133_1055 ();
 FILLCELL_X1 FILLER_133_1057 ();
 FILLCELL_X2 FILLER_133_1078 ();
 FILLCELL_X1 FILLER_133_1080 ();
 FILLCELL_X4 FILLER_133_1103 ();
 FILLCELL_X1 FILLER_133_1107 ();
 FILLCELL_X8 FILLER_133_1128 ();
 FILLCELL_X4 FILLER_133_1136 ();
 FILLCELL_X1 FILLER_133_1152 ();
 FILLCELL_X32 FILLER_133_1171 ();
 FILLCELL_X16 FILLER_133_1203 ();
 FILLCELL_X8 FILLER_133_1219 ();
 FILLCELL_X4 FILLER_133_1227 ();
 FILLCELL_X1 FILLER_133_1231 ();
 FILLCELL_X16 FILLER_133_1235 ();
 FILLCELL_X8 FILLER_133_1251 ();
 FILLCELL_X1 FILLER_133_1259 ();
 FILLCELL_X2 FILLER_134_1 ();
 FILLCELL_X2 FILLER_134_23 ();
 FILLCELL_X1 FILLER_134_25 ();
 FILLCELL_X1 FILLER_134_33 ();
 FILLCELL_X16 FILLER_134_41 ();
 FILLCELL_X4 FILLER_134_57 ();
 FILLCELL_X2 FILLER_134_61 ();
 FILLCELL_X1 FILLER_134_63 ();
 FILLCELL_X1 FILLER_134_125 ();
 FILLCELL_X1 FILLER_134_133 ();
 FILLCELL_X16 FILLER_134_145 ();
 FILLCELL_X8 FILLER_134_161 ();
 FILLCELL_X8 FILLER_134_176 ();
 FILLCELL_X16 FILLER_134_188 ();
 FILLCELL_X8 FILLER_134_204 ();
 FILLCELL_X4 FILLER_134_212 ();
 FILLCELL_X2 FILLER_134_216 ();
 FILLCELL_X4 FILLER_134_225 ();
 FILLCELL_X2 FILLER_134_243 ();
 FILLCELL_X4 FILLER_134_265 ();
 FILLCELL_X8 FILLER_134_300 ();
 FILLCELL_X8 FILLER_134_311 ();
 FILLCELL_X2 FILLER_134_319 ();
 FILLCELL_X2 FILLER_134_325 ();
 FILLCELL_X8 FILLER_134_330 ();
 FILLCELL_X2 FILLER_134_338 ();
 FILLCELL_X1 FILLER_134_340 ();
 FILLCELL_X4 FILLER_134_345 ();
 FILLCELL_X2 FILLER_134_349 ();
 FILLCELL_X1 FILLER_134_351 ();
 FILLCELL_X1 FILLER_134_356 ();
 FILLCELL_X8 FILLER_134_360 ();
 FILLCELL_X2 FILLER_134_368 ();
 FILLCELL_X8 FILLER_134_391 ();
 FILLCELL_X4 FILLER_134_399 ();
 FILLCELL_X2 FILLER_134_403 ();
 FILLCELL_X2 FILLER_134_407 ();
 FILLCELL_X1 FILLER_134_420 ();
 FILLCELL_X1 FILLER_134_424 ();
 FILLCELL_X8 FILLER_134_450 ();
 FILLCELL_X4 FILLER_134_458 ();
 FILLCELL_X2 FILLER_134_462 ();
 FILLCELL_X4 FILLER_134_467 ();
 FILLCELL_X2 FILLER_134_471 ();
 FILLCELL_X1 FILLER_134_473 ();
 FILLCELL_X4 FILLER_134_506 ();
 FILLCELL_X1 FILLER_134_510 ();
 FILLCELL_X8 FILLER_134_516 ();
 FILLCELL_X2 FILLER_134_524 ();
 FILLCELL_X1 FILLER_134_526 ();
 FILLCELL_X1 FILLER_134_535 ();
 FILLCELL_X4 FILLER_134_539 ();
 FILLCELL_X2 FILLER_134_543 ();
 FILLCELL_X8 FILLER_134_548 ();
 FILLCELL_X4 FILLER_134_556 ();
 FILLCELL_X2 FILLER_134_560 ();
 FILLCELL_X1 FILLER_134_562 ();
 FILLCELL_X4 FILLER_134_591 ();
 FILLCELL_X1 FILLER_134_595 ();
 FILLCELL_X4 FILLER_134_610 ();
 FILLCELL_X2 FILLER_134_614 ();
 FILLCELL_X1 FILLER_134_616 ();
 FILLCELL_X4 FILLER_134_624 ();
 FILLCELL_X2 FILLER_134_628 ();
 FILLCELL_X1 FILLER_134_630 ();
 FILLCELL_X4 FILLER_134_632 ();
 FILLCELL_X2 FILLER_134_636 ();
 FILLCELL_X1 FILLER_134_638 ();
 FILLCELL_X1 FILLER_134_659 ();
 FILLCELL_X8 FILLER_134_667 ();
 FILLCELL_X4 FILLER_134_675 ();
 FILLCELL_X32 FILLER_134_693 ();
 FILLCELL_X2 FILLER_134_725 ();
 FILLCELL_X8 FILLER_134_761 ();
 FILLCELL_X4 FILLER_134_769 ();
 FILLCELL_X8 FILLER_134_780 ();
 FILLCELL_X2 FILLER_134_795 ();
 FILLCELL_X2 FILLER_134_818 ();
 FILLCELL_X4 FILLER_134_830 ();
 FILLCELL_X2 FILLER_134_844 ();
 FILLCELL_X2 FILLER_134_852 ();
 FILLCELL_X1 FILLER_134_858 ();
 FILLCELL_X8 FILLER_134_869 ();
 FILLCELL_X4 FILLER_134_877 ();
 FILLCELL_X1 FILLER_134_881 ();
 FILLCELL_X4 FILLER_134_887 ();
 FILLCELL_X4 FILLER_134_895 ();
 FILLCELL_X2 FILLER_134_899 ();
 FILLCELL_X4 FILLER_134_904 ();
 FILLCELL_X4 FILLER_134_917 ();
 FILLCELL_X1 FILLER_134_928 ();
 FILLCELL_X1 FILLER_134_938 ();
 FILLCELL_X1 FILLER_134_946 ();
 FILLCELL_X4 FILLER_134_950 ();
 FILLCELL_X2 FILLER_134_954 ();
 FILLCELL_X1 FILLER_134_956 ();
 FILLCELL_X8 FILLER_134_970 ();
 FILLCELL_X8 FILLER_134_982 ();
 FILLCELL_X4 FILLER_134_990 ();
 FILLCELL_X1 FILLER_134_994 ();
 FILLCELL_X16 FILLER_134_997 ();
 FILLCELL_X2 FILLER_134_1013 ();
 FILLCELL_X4 FILLER_134_1019 ();
 FILLCELL_X2 FILLER_134_1023 ();
 FILLCELL_X1 FILLER_134_1071 ();
 FILLCELL_X1 FILLER_134_1094 ();
 FILLCELL_X1 FILLER_134_1097 ();
 FILLCELL_X4 FILLER_134_1112 ();
 FILLCELL_X1 FILLER_134_1116 ();
 FILLCELL_X8 FILLER_134_1129 ();
 FILLCELL_X1 FILLER_134_1137 ();
 FILLCELL_X4 FILLER_134_1140 ();
 FILLCELL_X2 FILLER_134_1144 ();
 FILLCELL_X8 FILLER_134_1148 ();
 FILLCELL_X2 FILLER_134_1156 ();
 FILLCELL_X2 FILLER_134_1161 ();
 FILLCELL_X1 FILLER_134_1163 ();
 FILLCELL_X32 FILLER_134_1181 ();
 FILLCELL_X32 FILLER_134_1213 ();
 FILLCELL_X8 FILLER_134_1245 ();
 FILLCELL_X4 FILLER_134_1253 ();
 FILLCELL_X2 FILLER_134_1257 ();
 FILLCELL_X1 FILLER_134_1259 ();
 FILLCELL_X4 FILLER_135_1 ();
 FILLCELL_X2 FILLER_135_5 ();
 FILLCELL_X2 FILLER_135_41 ();
 FILLCELL_X16 FILLER_135_50 ();
 FILLCELL_X8 FILLER_135_66 ();
 FILLCELL_X8 FILLER_135_79 ();
 FILLCELL_X2 FILLER_135_87 ();
 FILLCELL_X1 FILLER_135_103 ();
 FILLCELL_X1 FILLER_135_148 ();
 FILLCELL_X2 FILLER_135_183 ();
 FILLCELL_X16 FILLER_135_251 ();
 FILLCELL_X1 FILLER_135_267 ();
 FILLCELL_X4 FILLER_135_275 ();
 FILLCELL_X2 FILLER_135_279 ();
 FILLCELL_X8 FILLER_135_295 ();
 FILLCELL_X1 FILLER_135_303 ();
 FILLCELL_X1 FILLER_135_308 ();
 FILLCELL_X2 FILLER_135_329 ();
 FILLCELL_X1 FILLER_135_338 ();
 FILLCELL_X4 FILLER_135_369 ();
 FILLCELL_X2 FILLER_135_373 ();
 FILLCELL_X1 FILLER_135_378 ();
 FILLCELL_X4 FILLER_135_425 ();
 FILLCELL_X2 FILLER_135_429 ();
 FILLCELL_X1 FILLER_135_433 ();
 FILLCELL_X2 FILLER_135_440 ();
 FILLCELL_X1 FILLER_135_442 ();
 FILLCELL_X2 FILLER_135_450 ();
 FILLCELL_X4 FILLER_135_473 ();
 FILLCELL_X2 FILLER_135_477 ();
 FILLCELL_X2 FILLER_135_500 ();
 FILLCELL_X8 FILLER_135_507 ();
 FILLCELL_X1 FILLER_135_515 ();
 FILLCELL_X2 FILLER_135_584 ();
 FILLCELL_X2 FILLER_135_621 ();
 FILLCELL_X16 FILLER_135_630 ();
 FILLCELL_X2 FILLER_135_646 ();
 FILLCELL_X1 FILLER_135_648 ();
 FILLCELL_X4 FILLER_135_672 ();
 FILLCELL_X1 FILLER_135_676 ();
 FILLCELL_X8 FILLER_135_684 ();
 FILLCELL_X4 FILLER_135_692 ();
 FILLCELL_X1 FILLER_135_696 ();
 FILLCELL_X2 FILLER_135_701 ();
 FILLCELL_X16 FILLER_135_706 ();
 FILLCELL_X1 FILLER_135_753 ();
 FILLCELL_X1 FILLER_135_757 ();
 FILLCELL_X8 FILLER_135_793 ();
 FILLCELL_X4 FILLER_135_801 ();
 FILLCELL_X1 FILLER_135_805 ();
 FILLCELL_X2 FILLER_135_820 ();
 FILLCELL_X8 FILLER_135_836 ();
 FILLCELL_X4 FILLER_135_844 ();
 FILLCELL_X8 FILLER_135_866 ();
 FILLCELL_X4 FILLER_135_924 ();
 FILLCELL_X2 FILLER_135_933 ();
 FILLCELL_X2 FILLER_135_942 ();
 FILLCELL_X1 FILLER_135_944 ();
 FILLCELL_X1 FILLER_135_954 ();
 FILLCELL_X2 FILLER_135_959 ();
 FILLCELL_X1 FILLER_135_970 ();
 FILLCELL_X1 FILLER_135_985 ();
 FILLCELL_X2 FILLER_135_993 ();
 FILLCELL_X1 FILLER_135_995 ();
 FILLCELL_X4 FILLER_135_1006 ();
 FILLCELL_X2 FILLER_135_1010 ();
 FILLCELL_X16 FILLER_135_1022 ();
 FILLCELL_X8 FILLER_135_1038 ();
 FILLCELL_X4 FILLER_135_1046 ();
 FILLCELL_X2 FILLER_135_1050 ();
 FILLCELL_X8 FILLER_135_1066 ();
 FILLCELL_X8 FILLER_135_1084 ();
 FILLCELL_X4 FILLER_135_1092 ();
 FILLCELL_X2 FILLER_135_1096 ();
 FILLCELL_X2 FILLER_135_1130 ();
 FILLCELL_X1 FILLER_135_1132 ();
 FILLCELL_X2 FILLER_135_1149 ();
 FILLCELL_X2 FILLER_135_1153 ();
 FILLCELL_X1 FILLER_135_1176 ();
 FILLCELL_X32 FILLER_135_1193 ();
 FILLCELL_X32 FILLER_135_1225 ();
 FILLCELL_X2 FILLER_135_1257 ();
 FILLCELL_X1 FILLER_135_1259 ();
 FILLCELL_X8 FILLER_136_1 ();
 FILLCELL_X2 FILLER_136_9 ();
 FILLCELL_X4 FILLER_136_19 ();
 FILLCELL_X2 FILLER_136_23 ();
 FILLCELL_X1 FILLER_136_25 ();
 FILLCELL_X1 FILLER_136_47 ();
 FILLCELL_X4 FILLER_136_55 ();
 FILLCELL_X2 FILLER_136_59 ();
 FILLCELL_X1 FILLER_136_61 ();
 FILLCELL_X2 FILLER_136_123 ();
 FILLCELL_X4 FILLER_136_158 ();
 FILLCELL_X2 FILLER_136_162 ();
 FILLCELL_X2 FILLER_136_171 ();
 FILLCELL_X1 FILLER_136_173 ();
 FILLCELL_X8 FILLER_136_184 ();
 FILLCELL_X4 FILLER_136_192 ();
 FILLCELL_X1 FILLER_136_196 ();
 FILLCELL_X8 FILLER_136_217 ();
 FILLCELL_X1 FILLER_136_225 ();
 FILLCELL_X4 FILLER_136_233 ();
 FILLCELL_X2 FILLER_136_237 ();
 FILLCELL_X1 FILLER_136_239 ();
 FILLCELL_X1 FILLER_136_267 ();
 FILLCELL_X1 FILLER_136_275 ();
 FILLCELL_X1 FILLER_136_318 ();
 FILLCELL_X1 FILLER_136_322 ();
 FILLCELL_X1 FILLER_136_327 ();
 FILLCELL_X2 FILLER_136_338 ();
 FILLCELL_X8 FILLER_136_343 ();
 FILLCELL_X4 FILLER_136_351 ();
 FILLCELL_X1 FILLER_136_355 ();
 FILLCELL_X2 FILLER_136_370 ();
 FILLCELL_X1 FILLER_136_372 ();
 FILLCELL_X2 FILLER_136_376 ();
 FILLCELL_X1 FILLER_136_378 ();
 FILLCELL_X2 FILLER_136_386 ();
 FILLCELL_X2 FILLER_136_397 ();
 FILLCELL_X4 FILLER_136_403 ();
 FILLCELL_X4 FILLER_136_410 ();
 FILLCELL_X1 FILLER_136_414 ();
 FILLCELL_X2 FILLER_136_455 ();
 FILLCELL_X1 FILLER_136_457 ();
 FILLCELL_X4 FILLER_136_461 ();
 FILLCELL_X1 FILLER_136_465 ();
 FILLCELL_X4 FILLER_136_480 ();
 FILLCELL_X1 FILLER_136_484 ();
 FILLCELL_X8 FILLER_136_495 ();
 FILLCELL_X2 FILLER_136_503 ();
 FILLCELL_X2 FILLER_136_535 ();
 FILLCELL_X1 FILLER_136_537 ();
 FILLCELL_X8 FILLER_136_558 ();
 FILLCELL_X2 FILLER_136_566 ();
 FILLCELL_X16 FILLER_136_598 ();
 FILLCELL_X1 FILLER_136_614 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X1 FILLER_136_632 ();
 FILLCELL_X1 FILLER_136_636 ();
 FILLCELL_X8 FILLER_136_644 ();
 FILLCELL_X1 FILLER_136_652 ();
 FILLCELL_X1 FILLER_136_658 ();
 FILLCELL_X2 FILLER_136_691 ();
 FILLCELL_X4 FILLER_136_722 ();
 FILLCELL_X8 FILLER_136_733 ();
 FILLCELL_X4 FILLER_136_741 ();
 FILLCELL_X2 FILLER_136_745 ();
 FILLCELL_X8 FILLER_136_750 ();
 FILLCELL_X2 FILLER_136_758 ();
 FILLCELL_X2 FILLER_136_784 ();
 FILLCELL_X1 FILLER_136_786 ();
 FILLCELL_X2 FILLER_136_804 ();
 FILLCELL_X4 FILLER_136_816 ();
 FILLCELL_X1 FILLER_136_820 ();
 FILLCELL_X1 FILLER_136_837 ();
 FILLCELL_X2 FILLER_136_848 ();
 FILLCELL_X1 FILLER_136_850 ();
 FILLCELL_X2 FILLER_136_882 ();
 FILLCELL_X4 FILLER_136_916 ();
 FILLCELL_X2 FILLER_136_929 ();
 FILLCELL_X1 FILLER_136_931 ();
 FILLCELL_X8 FILLER_136_949 ();
 FILLCELL_X2 FILLER_136_970 ();
 FILLCELL_X1 FILLER_136_972 ();
 FILLCELL_X4 FILLER_136_978 ();
 FILLCELL_X1 FILLER_136_982 ();
 FILLCELL_X1 FILLER_136_999 ();
 FILLCELL_X2 FILLER_136_1007 ();
 FILLCELL_X1 FILLER_136_1009 ();
 FILLCELL_X4 FILLER_136_1013 ();
 FILLCELL_X1 FILLER_136_1017 ();
 FILLCELL_X2 FILLER_136_1038 ();
 FILLCELL_X1 FILLER_136_1040 ();
 FILLCELL_X2 FILLER_136_1051 ();
 FILLCELL_X4 FILLER_136_1055 ();
 FILLCELL_X1 FILLER_136_1059 ();
 FILLCELL_X8 FILLER_136_1076 ();
 FILLCELL_X1 FILLER_136_1084 ();
 FILLCELL_X2 FILLER_136_1103 ();
 FILLCELL_X1 FILLER_136_1105 ();
 FILLCELL_X2 FILLER_136_1108 ();
 FILLCELL_X2 FILLER_136_1120 ();
 FILLCELL_X1 FILLER_136_1122 ();
 FILLCELL_X2 FILLER_136_1125 ();
 FILLCELL_X4 FILLER_136_1131 ();
 FILLCELL_X2 FILLER_136_1135 ();
 FILLCELL_X1 FILLER_136_1147 ();
 FILLCELL_X1 FILLER_136_1164 ();
 FILLCELL_X32 FILLER_136_1192 ();
 FILLCELL_X32 FILLER_136_1224 ();
 FILLCELL_X4 FILLER_136_1256 ();
 FILLCELL_X8 FILLER_137_1 ();
 FILLCELL_X2 FILLER_137_9 ();
 FILLCELL_X1 FILLER_137_11 ();
 FILLCELL_X4 FILLER_137_32 ();
 FILLCELL_X1 FILLER_137_36 ();
 FILLCELL_X2 FILLER_137_44 ();
 FILLCELL_X16 FILLER_137_53 ();
 FILLCELL_X8 FILLER_137_69 ();
 FILLCELL_X1 FILLER_137_77 ();
 FILLCELL_X1 FILLER_137_126 ();
 FILLCELL_X1 FILLER_137_134 ();
 FILLCELL_X4 FILLER_137_176 ();
 FILLCELL_X1 FILLER_137_180 ();
 FILLCELL_X1 FILLER_137_195 ();
 FILLCELL_X1 FILLER_137_200 ();
 FILLCELL_X1 FILLER_137_205 ();
 FILLCELL_X8 FILLER_137_220 ();
 FILLCELL_X1 FILLER_137_228 ();
 FILLCELL_X8 FILLER_137_236 ();
 FILLCELL_X1 FILLER_137_244 ();
 FILLCELL_X4 FILLER_137_252 ();
 FILLCELL_X1 FILLER_137_263 ();
 FILLCELL_X2 FILLER_137_271 ();
 FILLCELL_X1 FILLER_137_280 ();
 FILLCELL_X2 FILLER_137_284 ();
 FILLCELL_X2 FILLER_137_289 ();
 FILLCELL_X8 FILLER_137_296 ();
 FILLCELL_X2 FILLER_137_304 ();
 FILLCELL_X1 FILLER_137_306 ();
 FILLCELL_X4 FILLER_137_314 ();
 FILLCELL_X1 FILLER_137_331 ();
 FILLCELL_X2 FILLER_137_371 ();
 FILLCELL_X1 FILLER_137_373 ();
 FILLCELL_X2 FILLER_137_388 ();
 FILLCELL_X2 FILLER_137_412 ();
 FILLCELL_X16 FILLER_137_445 ();
 FILLCELL_X2 FILLER_137_461 ();
 FILLCELL_X1 FILLER_137_463 ();
 FILLCELL_X8 FILLER_137_481 ();
 FILLCELL_X2 FILLER_137_489 ();
 FILLCELL_X1 FILLER_137_491 ();
 FILLCELL_X8 FILLER_137_503 ();
 FILLCELL_X4 FILLER_137_511 ();
 FILLCELL_X1 FILLER_137_522 ();
 FILLCELL_X1 FILLER_137_530 ();
 FILLCELL_X2 FILLER_137_535 ();
 FILLCELL_X1 FILLER_137_537 ();
 FILLCELL_X2 FILLER_137_558 ();
 FILLCELL_X2 FILLER_137_567 ();
 FILLCELL_X1 FILLER_137_587 ();
 FILLCELL_X2 FILLER_137_602 ();
 FILLCELL_X2 FILLER_137_611 ();
 FILLCELL_X4 FILLER_137_626 ();
 FILLCELL_X1 FILLER_137_630 ();
 FILLCELL_X4 FILLER_137_702 ();
 FILLCELL_X2 FILLER_137_706 ();
 FILLCELL_X2 FILLER_137_717 ();
 FILLCELL_X2 FILLER_137_750 ();
 FILLCELL_X1 FILLER_137_762 ();
 FILLCELL_X1 FILLER_137_777 ();
 FILLCELL_X2 FILLER_137_799 ();
 FILLCELL_X1 FILLER_137_801 ();
 FILLCELL_X2 FILLER_137_809 ();
 FILLCELL_X1 FILLER_137_811 ();
 FILLCELL_X8 FILLER_137_835 ();
 FILLCELL_X4 FILLER_137_843 ();
 FILLCELL_X2 FILLER_137_847 ();
 FILLCELL_X1 FILLER_137_849 ();
 FILLCELL_X2 FILLER_137_854 ();
 FILLCELL_X2 FILLER_137_873 ();
 FILLCELL_X2 FILLER_137_888 ();
 FILLCELL_X1 FILLER_137_890 ();
 FILLCELL_X4 FILLER_137_923 ();
 FILLCELL_X4 FILLER_137_934 ();
 FILLCELL_X1 FILLER_137_942 ();
 FILLCELL_X2 FILLER_137_947 ();
 FILLCELL_X1 FILLER_137_949 ();
 FILLCELL_X2 FILLER_137_954 ();
 FILLCELL_X2 FILLER_137_975 ();
 FILLCELL_X2 FILLER_137_989 ();
 FILLCELL_X8 FILLER_137_996 ();
 FILLCELL_X1 FILLER_137_1004 ();
 FILLCELL_X2 FILLER_137_1021 ();
 FILLCELL_X1 FILLER_137_1025 ();
 FILLCELL_X1 FILLER_137_1029 ();
 FILLCELL_X1 FILLER_137_1033 ();
 FILLCELL_X1 FILLER_137_1037 ();
 FILLCELL_X1 FILLER_137_1054 ();
 FILLCELL_X1 FILLER_137_1094 ();
 FILLCELL_X1 FILLER_137_1098 ();
 FILLCELL_X1 FILLER_137_1109 ();
 FILLCELL_X2 FILLER_137_1112 ();
 FILLCELL_X4 FILLER_137_1142 ();
 FILLCELL_X16 FILLER_137_1148 ();
 FILLCELL_X4 FILLER_137_1164 ();
 FILLCELL_X2 FILLER_137_1168 ();
 FILLCELL_X1 FILLER_137_1187 ();
 FILLCELL_X32 FILLER_137_1191 ();
 FILLCELL_X32 FILLER_137_1223 ();
 FILLCELL_X4 FILLER_137_1255 ();
 FILLCELL_X1 FILLER_137_1259 ();
 FILLCELL_X16 FILLER_138_49 ();
 FILLCELL_X1 FILLER_138_65 ();
 FILLCELL_X16 FILLER_138_93 ();
 FILLCELL_X2 FILLER_138_109 ();
 FILLCELL_X8 FILLER_138_120 ();
 FILLCELL_X1 FILLER_138_128 ();
 FILLCELL_X8 FILLER_138_139 ();
 FILLCELL_X2 FILLER_138_154 ();
 FILLCELL_X1 FILLER_138_156 ();
 FILLCELL_X2 FILLER_138_182 ();
 FILLCELL_X1 FILLER_138_184 ();
 FILLCELL_X8 FILLER_138_198 ();
 FILLCELL_X2 FILLER_138_206 ();
 FILLCELL_X4 FILLER_138_221 ();
 FILLCELL_X2 FILLER_138_225 ();
 FILLCELL_X2 FILLER_138_234 ();
 FILLCELL_X1 FILLER_138_236 ();
 FILLCELL_X8 FILLER_138_284 ();
 FILLCELL_X4 FILLER_138_292 ();
 FILLCELL_X2 FILLER_138_371 ();
 FILLCELL_X1 FILLER_138_373 ();
 FILLCELL_X2 FILLER_138_402 ();
 FILLCELL_X1 FILLER_138_404 ();
 FILLCELL_X2 FILLER_138_412 ();
 FILLCELL_X1 FILLER_138_414 ();
 FILLCELL_X2 FILLER_138_418 ();
 FILLCELL_X1 FILLER_138_420 ();
 FILLCELL_X4 FILLER_138_435 ();
 FILLCELL_X2 FILLER_138_439 ();
 FILLCELL_X1 FILLER_138_441 ();
 FILLCELL_X16 FILLER_138_456 ();
 FILLCELL_X2 FILLER_138_472 ();
 FILLCELL_X1 FILLER_138_474 ();
 FILLCELL_X2 FILLER_138_482 ();
 FILLCELL_X1 FILLER_138_484 ();
 FILLCELL_X2 FILLER_138_505 ();
 FILLCELL_X2 FILLER_138_514 ();
 FILLCELL_X1 FILLER_138_516 ();
 FILLCELL_X1 FILLER_138_524 ();
 FILLCELL_X2 FILLER_138_532 ();
 FILLCELL_X2 FILLER_138_615 ();
 FILLCELL_X1 FILLER_138_617 ();
 FILLCELL_X1 FILLER_138_632 ();
 FILLCELL_X2 FILLER_138_646 ();
 FILLCELL_X2 FILLER_138_655 ();
 FILLCELL_X2 FILLER_138_664 ();
 FILLCELL_X2 FILLER_138_670 ();
 FILLCELL_X16 FILLER_138_675 ();
 FILLCELL_X1 FILLER_138_691 ();
 FILLCELL_X16 FILLER_138_699 ();
 FILLCELL_X8 FILLER_138_715 ();
 FILLCELL_X4 FILLER_138_733 ();
 FILLCELL_X2 FILLER_138_737 ();
 FILLCELL_X4 FILLER_138_749 ();
 FILLCELL_X1 FILLER_138_787 ();
 FILLCELL_X4 FILLER_138_802 ();
 FILLCELL_X1 FILLER_138_825 ();
 FILLCELL_X1 FILLER_138_838 ();
 FILLCELL_X4 FILLER_138_849 ();
 FILLCELL_X2 FILLER_138_853 ();
 FILLCELL_X1 FILLER_138_855 ();
 FILLCELL_X4 FILLER_138_870 ();
 FILLCELL_X2 FILLER_138_874 ();
 FILLCELL_X1 FILLER_138_876 ();
 FILLCELL_X1 FILLER_138_889 ();
 FILLCELL_X2 FILLER_138_931 ();
 FILLCELL_X1 FILLER_138_949 ();
 FILLCELL_X2 FILLER_138_963 ();
 FILLCELL_X1 FILLER_138_965 ();
 FILLCELL_X2 FILLER_138_979 ();
 FILLCELL_X1 FILLER_138_981 ();
 FILLCELL_X4 FILLER_138_1001 ();
 FILLCELL_X1 FILLER_138_1005 ();
 FILLCELL_X2 FILLER_138_1017 ();
 FILLCELL_X4 FILLER_138_1038 ();
 FILLCELL_X2 FILLER_138_1042 ();
 FILLCELL_X1 FILLER_138_1050 ();
 FILLCELL_X2 FILLER_138_1061 ();
 FILLCELL_X4 FILLER_138_1066 ();
 FILLCELL_X2 FILLER_138_1070 ();
 FILLCELL_X8 FILLER_138_1107 ();
 FILLCELL_X4 FILLER_138_1117 ();
 FILLCELL_X2 FILLER_138_1121 ();
 FILLCELL_X1 FILLER_138_1123 ();
 FILLCELL_X2 FILLER_138_1134 ();
 FILLCELL_X1 FILLER_138_1136 ();
 FILLCELL_X1 FILLER_138_1141 ();
 FILLCELL_X8 FILLER_138_1144 ();
 FILLCELL_X4 FILLER_138_1152 ();
 FILLCELL_X32 FILLER_138_1182 ();
 FILLCELL_X32 FILLER_138_1214 ();
 FILLCELL_X8 FILLER_138_1246 ();
 FILLCELL_X4 FILLER_138_1254 ();
 FILLCELL_X2 FILLER_138_1258 ();
 FILLCELL_X16 FILLER_139_1 ();
 FILLCELL_X2 FILLER_139_44 ();
 FILLCELL_X1 FILLER_139_46 ();
 FILLCELL_X1 FILLER_139_74 ();
 FILLCELL_X4 FILLER_139_82 ();
 FILLCELL_X2 FILLER_139_86 ();
 FILLCELL_X1 FILLER_139_88 ();
 FILLCELL_X4 FILLER_139_117 ();
 FILLCELL_X2 FILLER_139_121 ();
 FILLCELL_X1 FILLER_139_123 ();
 FILLCELL_X4 FILLER_139_131 ();
 FILLCELL_X2 FILLER_139_135 ();
 FILLCELL_X16 FILLER_139_144 ();
 FILLCELL_X4 FILLER_139_160 ();
 FILLCELL_X16 FILLER_139_171 ();
 FILLCELL_X4 FILLER_139_187 ();
 FILLCELL_X2 FILLER_139_211 ();
 FILLCELL_X1 FILLER_139_213 ();
 FILLCELL_X4 FILLER_139_221 ();
 FILLCELL_X4 FILLER_139_239 ();
 FILLCELL_X1 FILLER_139_243 ();
 FILLCELL_X4 FILLER_139_251 ();
 FILLCELL_X2 FILLER_139_255 ();
 FILLCELL_X2 FILLER_139_264 ();
 FILLCELL_X1 FILLER_139_266 ();
 FILLCELL_X8 FILLER_139_274 ();
 FILLCELL_X4 FILLER_139_282 ();
 FILLCELL_X2 FILLER_139_286 ();
 FILLCELL_X1 FILLER_139_288 ();
 FILLCELL_X1 FILLER_139_316 ();
 FILLCELL_X4 FILLER_139_320 ();
 FILLCELL_X2 FILLER_139_328 ();
 FILLCELL_X8 FILLER_139_334 ();
 FILLCELL_X2 FILLER_139_342 ();
 FILLCELL_X1 FILLER_139_344 ();
 FILLCELL_X1 FILLER_139_352 ();
 FILLCELL_X1 FILLER_139_356 ();
 FILLCELL_X2 FILLER_139_368 ();
 FILLCELL_X8 FILLER_139_373 ();
 FILLCELL_X1 FILLER_139_385 ();
 FILLCELL_X4 FILLER_139_406 ();
 FILLCELL_X2 FILLER_139_410 ();
 FILLCELL_X1 FILLER_139_412 ();
 FILLCELL_X1 FILLER_139_426 ();
 FILLCELL_X2 FILLER_139_435 ();
 FILLCELL_X1 FILLER_139_437 ();
 FILLCELL_X2 FILLER_139_459 ();
 FILLCELL_X4 FILLER_139_495 ();
 FILLCELL_X1 FILLER_139_499 ();
 FILLCELL_X2 FILLER_139_503 ();
 FILLCELL_X2 FILLER_139_525 ();
 FILLCELL_X2 FILLER_139_534 ();
 FILLCELL_X1 FILLER_139_536 ();
 FILLCELL_X1 FILLER_139_544 ();
 FILLCELL_X4 FILLER_139_557 ();
 FILLCELL_X2 FILLER_139_561 ();
 FILLCELL_X1 FILLER_139_563 ();
 FILLCELL_X2 FILLER_139_604 ();
 FILLCELL_X16 FILLER_139_633 ();
 FILLCELL_X2 FILLER_139_649 ();
 FILLCELL_X2 FILLER_139_678 ();
 FILLCELL_X8 FILLER_139_700 ();
 FILLCELL_X4 FILLER_139_708 ();
 FILLCELL_X1 FILLER_139_712 ();
 FILLCELL_X1 FILLER_139_755 ();
 FILLCELL_X1 FILLER_139_770 ();
 FILLCELL_X8 FILLER_139_791 ();
 FILLCELL_X4 FILLER_139_799 ();
 FILLCELL_X2 FILLER_139_803 ();
 FILLCELL_X1 FILLER_139_823 ();
 FILLCELL_X1 FILLER_139_826 ();
 FILLCELL_X1 FILLER_139_843 ();
 FILLCELL_X1 FILLER_139_866 ();
 FILLCELL_X4 FILLER_139_869 ();
 FILLCELL_X1 FILLER_139_913 ();
 FILLCELL_X2 FILLER_139_918 ();
 FILLCELL_X1 FILLER_139_920 ();
 FILLCELL_X1 FILLER_139_930 ();
 FILLCELL_X2 FILLER_139_940 ();
 FILLCELL_X1 FILLER_139_949 ();
 FILLCELL_X4 FILLER_139_968 ();
 FILLCELL_X2 FILLER_139_972 ();
 FILLCELL_X8 FILLER_139_980 ();
 FILLCELL_X2 FILLER_139_988 ();
 FILLCELL_X1 FILLER_139_990 ();
 FILLCELL_X2 FILLER_139_1000 ();
 FILLCELL_X1 FILLER_139_1002 ();
 FILLCELL_X16 FILLER_139_1008 ();
 FILLCELL_X1 FILLER_139_1043 ();
 FILLCELL_X4 FILLER_139_1091 ();
 FILLCELL_X8 FILLER_139_1099 ();
 FILLCELL_X1 FILLER_139_1107 ();
 FILLCELL_X4 FILLER_139_1111 ();
 FILLCELL_X4 FILLER_139_1125 ();
 FILLCELL_X2 FILLER_139_1129 ();
 FILLCELL_X1 FILLER_139_1131 ();
 FILLCELL_X8 FILLER_139_1162 ();
 FILLCELL_X1 FILLER_139_1170 ();
 FILLCELL_X32 FILLER_139_1178 ();
 FILLCELL_X32 FILLER_139_1210 ();
 FILLCELL_X16 FILLER_139_1242 ();
 FILLCELL_X2 FILLER_139_1258 ();
 FILLCELL_X16 FILLER_140_1 ();
 FILLCELL_X2 FILLER_140_44 ();
 FILLCELL_X1 FILLER_140_46 ();
 FILLCELL_X1 FILLER_140_67 ();
 FILLCELL_X4 FILLER_140_115 ();
 FILLCELL_X4 FILLER_140_126 ();
 FILLCELL_X1 FILLER_140_160 ();
 FILLCELL_X4 FILLER_140_188 ();
 FILLCELL_X2 FILLER_140_192 ();
 FILLCELL_X1 FILLER_140_194 ();
 FILLCELL_X4 FILLER_140_202 ();
 FILLCELL_X2 FILLER_140_206 ();
 FILLCELL_X1 FILLER_140_208 ();
 FILLCELL_X1 FILLER_140_236 ();
 FILLCELL_X8 FILLER_140_257 ();
 FILLCELL_X2 FILLER_140_265 ();
 FILLCELL_X1 FILLER_140_267 ();
 FILLCELL_X2 FILLER_140_275 ();
 FILLCELL_X1 FILLER_140_280 ();
 FILLCELL_X1 FILLER_140_288 ();
 FILLCELL_X2 FILLER_140_310 ();
 FILLCELL_X1 FILLER_140_312 ();
 FILLCELL_X4 FILLER_140_317 ();
 FILLCELL_X1 FILLER_140_354 ();
 FILLCELL_X2 FILLER_140_358 ();
 FILLCELL_X1 FILLER_140_367 ();
 FILLCELL_X2 FILLER_140_375 ();
 FILLCELL_X1 FILLER_140_397 ();
 FILLCELL_X1 FILLER_140_412 ();
 FILLCELL_X2 FILLER_140_436 ();
 FILLCELL_X1 FILLER_140_438 ();
 FILLCELL_X4 FILLER_140_457 ();
 FILLCELL_X1 FILLER_140_464 ();
 FILLCELL_X4 FILLER_140_468 ();
 FILLCELL_X4 FILLER_140_479 ();
 FILLCELL_X1 FILLER_140_497 ();
 FILLCELL_X2 FILLER_140_505 ();
 FILLCELL_X1 FILLER_140_514 ();
 FILLCELL_X8 FILLER_140_522 ();
 FILLCELL_X1 FILLER_140_544 ();
 FILLCELL_X8 FILLER_140_555 ();
 FILLCELL_X2 FILLER_140_563 ();
 FILLCELL_X2 FILLER_140_614 ();
 FILLCELL_X1 FILLER_140_616 ();
 FILLCELL_X4 FILLER_140_639 ();
 FILLCELL_X4 FILLER_140_671 ();
 FILLCELL_X2 FILLER_140_675 ();
 FILLCELL_X4 FILLER_140_684 ();
 FILLCELL_X2 FILLER_140_688 ();
 FILLCELL_X1 FILLER_140_690 ();
 FILLCELL_X8 FILLER_140_705 ();
 FILLCELL_X2 FILLER_140_713 ();
 FILLCELL_X1 FILLER_140_715 ();
 FILLCELL_X2 FILLER_140_726 ();
 FILLCELL_X1 FILLER_140_728 ();
 FILLCELL_X8 FILLER_140_732 ();
 FILLCELL_X2 FILLER_140_747 ();
 FILLCELL_X2 FILLER_140_752 ();
 FILLCELL_X1 FILLER_140_754 ();
 FILLCELL_X4 FILLER_140_769 ();
 FILLCELL_X2 FILLER_140_773 ();
 FILLCELL_X1 FILLER_140_775 ();
 FILLCELL_X4 FILLER_140_783 ();
 FILLCELL_X2 FILLER_140_787 ();
 FILLCELL_X1 FILLER_140_789 ();
 FILLCELL_X8 FILLER_140_797 ();
 FILLCELL_X1 FILLER_140_805 ();
 FILLCELL_X8 FILLER_140_808 ();
 FILLCELL_X4 FILLER_140_816 ();
 FILLCELL_X8 FILLER_140_854 ();
 FILLCELL_X1 FILLER_140_862 ();
 FILLCELL_X1 FILLER_140_881 ();
 FILLCELL_X1 FILLER_140_886 ();
 FILLCELL_X8 FILLER_140_906 ();
 FILLCELL_X4 FILLER_140_914 ();
 FILLCELL_X4 FILLER_140_920 ();
 FILLCELL_X2 FILLER_140_924 ();
 FILLCELL_X2 FILLER_140_946 ();
 FILLCELL_X1 FILLER_140_950 ();
 FILLCELL_X2 FILLER_140_966 ();
 FILLCELL_X2 FILLER_140_985 ();
 FILLCELL_X2 FILLER_140_993 ();
 FILLCELL_X1 FILLER_140_995 ();
 FILLCELL_X2 FILLER_140_1000 ();
 FILLCELL_X8 FILLER_140_1005 ();
 FILLCELL_X2 FILLER_140_1013 ();
 FILLCELL_X1 FILLER_140_1015 ();
 FILLCELL_X4 FILLER_140_1024 ();
 FILLCELL_X1 FILLER_140_1028 ();
 FILLCELL_X1 FILLER_140_1032 ();
 FILLCELL_X1 FILLER_140_1035 ();
 FILLCELL_X1 FILLER_140_1039 ();
 FILLCELL_X1 FILLER_140_1056 ();
 FILLCELL_X1 FILLER_140_1060 ();
 FILLCELL_X4 FILLER_140_1066 ();
 FILLCELL_X2 FILLER_140_1070 ();
 FILLCELL_X8 FILLER_140_1093 ();
 FILLCELL_X2 FILLER_140_1101 ();
 FILLCELL_X1 FILLER_140_1103 ();
 FILLCELL_X1 FILLER_140_1114 ();
 FILLCELL_X2 FILLER_140_1125 ();
 FILLCELL_X4 FILLER_140_1129 ();
 FILLCELL_X2 FILLER_140_1133 ();
 FILLCELL_X1 FILLER_140_1135 ();
 FILLCELL_X1 FILLER_140_1146 ();
 FILLCELL_X1 FILLER_140_1149 ();
 FILLCELL_X32 FILLER_140_1176 ();
 FILLCELL_X32 FILLER_140_1208 ();
 FILLCELL_X16 FILLER_140_1240 ();
 FILLCELL_X4 FILLER_140_1256 ();
 FILLCELL_X8 FILLER_141_35 ();
 FILLCELL_X2 FILLER_141_43 ();
 FILLCELL_X2 FILLER_141_72 ();
 FILLCELL_X1 FILLER_141_74 ();
 FILLCELL_X8 FILLER_141_80 ();
 FILLCELL_X2 FILLER_141_88 ();
 FILLCELL_X1 FILLER_141_90 ();
 FILLCELL_X4 FILLER_141_98 ();
 FILLCELL_X1 FILLER_141_102 ();
 FILLCELL_X8 FILLER_141_117 ();
 FILLCELL_X4 FILLER_141_125 ();
 FILLCELL_X16 FILLER_141_136 ();
 FILLCELL_X2 FILLER_141_152 ();
 FILLCELL_X2 FILLER_141_161 ();
 FILLCELL_X4 FILLER_141_177 ();
 FILLCELL_X2 FILLER_141_181 ();
 FILLCELL_X1 FILLER_141_183 ();
 FILLCELL_X4 FILLER_141_191 ();
 FILLCELL_X2 FILLER_141_195 ();
 FILLCELL_X8 FILLER_141_231 ();
 FILLCELL_X4 FILLER_141_239 ();
 FILLCELL_X2 FILLER_141_243 ();
 FILLCELL_X8 FILLER_141_286 ();
 FILLCELL_X1 FILLER_141_294 ();
 FILLCELL_X8 FILLER_141_328 ();
 FILLCELL_X2 FILLER_141_336 ();
 FILLCELL_X8 FILLER_141_341 ();
 FILLCELL_X1 FILLER_141_349 ();
 FILLCELL_X1 FILLER_141_357 ();
 FILLCELL_X2 FILLER_141_362 ();
 FILLCELL_X2 FILLER_141_367 ();
 FILLCELL_X1 FILLER_141_369 ();
 FILLCELL_X8 FILLER_141_377 ();
 FILLCELL_X1 FILLER_141_385 ();
 FILLCELL_X1 FILLER_141_457 ();
 FILLCELL_X1 FILLER_141_465 ();
 FILLCELL_X2 FILLER_141_493 ();
 FILLCELL_X1 FILLER_141_495 ();
 FILLCELL_X4 FILLER_141_503 ();
 FILLCELL_X2 FILLER_141_507 ();
 FILLCELL_X8 FILLER_141_513 ();
 FILLCELL_X2 FILLER_141_521 ();
 FILLCELL_X2 FILLER_141_533 ();
 FILLCELL_X2 FILLER_141_555 ();
 FILLCELL_X1 FILLER_141_557 ();
 FILLCELL_X2 FILLER_141_608 ();
 FILLCELL_X2 FILLER_141_617 ();
 FILLCELL_X2 FILLER_141_654 ();
 FILLCELL_X1 FILLER_141_663 ();
 FILLCELL_X16 FILLER_141_713 ();
 FILLCELL_X32 FILLER_141_736 ();
 FILLCELL_X4 FILLER_141_768 ();
 FILLCELL_X1 FILLER_141_788 ();
 FILLCELL_X4 FILLER_141_807 ();
 FILLCELL_X1 FILLER_141_811 ();
 FILLCELL_X4 FILLER_141_814 ();
 FILLCELL_X2 FILLER_141_818 ();
 FILLCELL_X1 FILLER_141_820 ();
 FILLCELL_X8 FILLER_141_823 ();
 FILLCELL_X8 FILLER_141_845 ();
 FILLCELL_X1 FILLER_141_853 ();
 FILLCELL_X8 FILLER_141_868 ();
 FILLCELL_X4 FILLER_141_876 ();
 FILLCELL_X8 FILLER_141_892 ();
 FILLCELL_X1 FILLER_141_914 ();
 FILLCELL_X4 FILLER_141_931 ();
 FILLCELL_X1 FILLER_141_951 ();
 FILLCELL_X1 FILLER_141_956 ();
 FILLCELL_X1 FILLER_141_977 ();
 FILLCELL_X2 FILLER_141_996 ();
 FILLCELL_X1 FILLER_141_998 ();
 FILLCELL_X8 FILLER_141_1009 ();
 FILLCELL_X4 FILLER_141_1017 ();
 FILLCELL_X2 FILLER_141_1021 ();
 FILLCELL_X1 FILLER_141_1023 ();
 FILLCELL_X2 FILLER_141_1049 ();
 FILLCELL_X2 FILLER_141_1067 ();
 FILLCELL_X8 FILLER_141_1088 ();
 FILLCELL_X2 FILLER_141_1096 ();
 FILLCELL_X2 FILLER_141_1142 ();
 FILLCELL_X1 FILLER_141_1144 ();
 FILLCELL_X2 FILLER_141_1161 ();
 FILLCELL_X1 FILLER_141_1163 ();
 FILLCELL_X32 FILLER_141_1182 ();
 FILLCELL_X32 FILLER_141_1214 ();
 FILLCELL_X8 FILLER_141_1246 ();
 FILLCELL_X4 FILLER_141_1254 ();
 FILLCELL_X2 FILLER_141_1258 ();
 FILLCELL_X16 FILLER_142_1 ();
 FILLCELL_X1 FILLER_142_17 ();
 FILLCELL_X2 FILLER_142_38 ();
 FILLCELL_X4 FILLER_142_47 ();
 FILLCELL_X2 FILLER_142_58 ();
 FILLCELL_X1 FILLER_142_60 ();
 FILLCELL_X16 FILLER_142_101 ();
 FILLCELL_X4 FILLER_142_117 ();
 FILLCELL_X2 FILLER_142_121 ();
 FILLCELL_X1 FILLER_142_123 ();
 FILLCELL_X2 FILLER_142_131 ();
 FILLCELL_X2 FILLER_142_160 ();
 FILLCELL_X1 FILLER_142_162 ();
 FILLCELL_X4 FILLER_142_183 ();
 FILLCELL_X1 FILLER_142_187 ();
 FILLCELL_X1 FILLER_142_216 ();
 FILLCELL_X8 FILLER_142_238 ();
 FILLCELL_X2 FILLER_142_246 ();
 FILLCELL_X1 FILLER_142_255 ();
 FILLCELL_X4 FILLER_142_263 ();
 FILLCELL_X2 FILLER_142_267 ();
 FILLCELL_X1 FILLER_142_269 ();
 FILLCELL_X2 FILLER_142_277 ();
 FILLCELL_X4 FILLER_142_286 ();
 FILLCELL_X2 FILLER_142_308 ();
 FILLCELL_X1 FILLER_142_310 ();
 FILLCELL_X2 FILLER_142_325 ();
 FILLCELL_X1 FILLER_142_327 ();
 FILLCELL_X2 FILLER_142_332 ();
 FILLCELL_X1 FILLER_142_334 ();
 FILLCELL_X2 FILLER_142_389 ();
 FILLCELL_X1 FILLER_142_391 ();
 FILLCELL_X2 FILLER_142_399 ();
 FILLCELL_X1 FILLER_142_401 ();
 FILLCELL_X16 FILLER_142_434 ();
 FILLCELL_X4 FILLER_142_450 ();
 FILLCELL_X1 FILLER_142_454 ();
 FILLCELL_X1 FILLER_142_460 ();
 FILLCELL_X8 FILLER_142_468 ();
 FILLCELL_X4 FILLER_142_476 ();
 FILLCELL_X2 FILLER_142_480 ();
 FILLCELL_X4 FILLER_142_502 ();
 FILLCELL_X1 FILLER_142_506 ();
 FILLCELL_X4 FILLER_142_527 ();
 FILLCELL_X2 FILLER_142_531 ();
 FILLCELL_X1 FILLER_142_533 ();
 FILLCELL_X2 FILLER_142_541 ();
 FILLCELL_X2 FILLER_142_547 ();
 FILLCELL_X8 FILLER_142_552 ();
 FILLCELL_X8 FILLER_142_564 ();
 FILLCELL_X2 FILLER_142_572 ();
 FILLCELL_X1 FILLER_142_585 ();
 FILLCELL_X2 FILLER_142_610 ();
 FILLCELL_X1 FILLER_142_612 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X4 FILLER_142_652 ();
 FILLCELL_X2 FILLER_142_656 ();
 FILLCELL_X1 FILLER_142_658 ();
 FILLCELL_X8 FILLER_142_682 ();
 FILLCELL_X1 FILLER_142_690 ();
 FILLCELL_X32 FILLER_142_711 ();
 FILLCELL_X32 FILLER_142_743 ();
 FILLCELL_X8 FILLER_142_775 ();
 FILLCELL_X2 FILLER_142_783 ();
 FILLCELL_X1 FILLER_142_787 ();
 FILLCELL_X4 FILLER_142_790 ();
 FILLCELL_X2 FILLER_142_794 ();
 FILLCELL_X1 FILLER_142_796 ();
 FILLCELL_X8 FILLER_142_823 ();
 FILLCELL_X1 FILLER_142_831 ();
 FILLCELL_X4 FILLER_142_850 ();
 FILLCELL_X4 FILLER_142_872 ();
 FILLCELL_X2 FILLER_142_876 ();
 FILLCELL_X8 FILLER_142_896 ();
 FILLCELL_X2 FILLER_142_904 ();
 FILLCELL_X16 FILLER_142_910 ();
 FILLCELL_X4 FILLER_142_926 ();
 FILLCELL_X1 FILLER_142_930 ();
 FILLCELL_X2 FILLER_142_933 ();
 FILLCELL_X8 FILLER_142_937 ();
 FILLCELL_X4 FILLER_142_945 ();
 FILLCELL_X2 FILLER_142_959 ();
 FILLCELL_X1 FILLER_142_961 ();
 FILLCELL_X4 FILLER_142_1008 ();
 FILLCELL_X2 FILLER_142_1012 ();
 FILLCELL_X1 FILLER_142_1014 ();
 FILLCELL_X2 FILLER_142_1049 ();
 FILLCELL_X1 FILLER_142_1051 ();
 FILLCELL_X2 FILLER_142_1055 ();
 FILLCELL_X1 FILLER_142_1057 ();
 FILLCELL_X8 FILLER_142_1063 ();
 FILLCELL_X4 FILLER_142_1071 ();
 FILLCELL_X1 FILLER_142_1075 ();
 FILLCELL_X8 FILLER_142_1092 ();
 FILLCELL_X4 FILLER_142_1100 ();
 FILLCELL_X2 FILLER_142_1104 ();
 FILLCELL_X4 FILLER_142_1108 ();
 FILLCELL_X1 FILLER_142_1112 ();
 FILLCELL_X1 FILLER_142_1123 ();
 FILLCELL_X4 FILLER_142_1146 ();
 FILLCELL_X1 FILLER_142_1150 ();
 FILLCELL_X8 FILLER_142_1161 ();
 FILLCELL_X2 FILLER_142_1169 ();
 FILLCELL_X2 FILLER_142_1183 ();
 FILLCELL_X1 FILLER_142_1185 ();
 FILLCELL_X32 FILLER_142_1189 ();
 FILLCELL_X32 FILLER_142_1221 ();
 FILLCELL_X4 FILLER_142_1253 ();
 FILLCELL_X2 FILLER_142_1257 ();
 FILLCELL_X1 FILLER_142_1259 ();
 FILLCELL_X16 FILLER_143_1 ();
 FILLCELL_X2 FILLER_143_17 ();
 FILLCELL_X1 FILLER_143_19 ();
 FILLCELL_X8 FILLER_143_54 ();
 FILLCELL_X8 FILLER_143_69 ();
 FILLCELL_X2 FILLER_143_77 ();
 FILLCELL_X4 FILLER_143_86 ();
 FILLCELL_X1 FILLER_143_90 ();
 FILLCELL_X1 FILLER_143_111 ();
 FILLCELL_X2 FILLER_143_119 ();
 FILLCELL_X4 FILLER_143_128 ();
 FILLCELL_X2 FILLER_143_132 ();
 FILLCELL_X1 FILLER_143_134 ();
 FILLCELL_X8 FILLER_143_142 ();
 FILLCELL_X2 FILLER_143_150 ();
 FILLCELL_X4 FILLER_143_171 ();
 FILLCELL_X2 FILLER_143_175 ();
 FILLCELL_X16 FILLER_143_220 ();
 FILLCELL_X2 FILLER_143_236 ();
 FILLCELL_X4 FILLER_143_245 ();
 FILLCELL_X2 FILLER_143_249 ();
 FILLCELL_X8 FILLER_143_286 ();
 FILLCELL_X1 FILLER_143_294 ();
 FILLCELL_X4 FILLER_143_352 ();
 FILLCELL_X1 FILLER_143_356 ();
 FILLCELL_X4 FILLER_143_371 ();
 FILLCELL_X1 FILLER_143_375 ();
 FILLCELL_X2 FILLER_143_380 ();
 FILLCELL_X1 FILLER_143_382 ();
 FILLCELL_X4 FILLER_143_407 ();
 FILLCELL_X2 FILLER_143_411 ();
 FILLCELL_X1 FILLER_143_413 ();
 FILLCELL_X2 FILLER_143_421 ();
 FILLCELL_X1 FILLER_143_423 ();
 FILLCELL_X2 FILLER_143_445 ();
 FILLCELL_X1 FILLER_143_450 ();
 FILLCELL_X8 FILLER_143_461 ();
 FILLCELL_X4 FILLER_143_469 ();
 FILLCELL_X1 FILLER_143_473 ();
 FILLCELL_X4 FILLER_143_479 ();
 FILLCELL_X2 FILLER_143_483 ();
 FILLCELL_X4 FILLER_143_499 ();
 FILLCELL_X1 FILLER_143_518 ();
 FILLCELL_X2 FILLER_143_533 ();
 FILLCELL_X4 FILLER_143_555 ();
 FILLCELL_X2 FILLER_143_572 ();
 FILLCELL_X4 FILLER_143_594 ();
 FILLCELL_X1 FILLER_143_605 ();
 FILLCELL_X8 FILLER_143_613 ();
 FILLCELL_X4 FILLER_143_621 ();
 FILLCELL_X1 FILLER_143_632 ();
 FILLCELL_X8 FILLER_143_637 ();
 FILLCELL_X1 FILLER_143_645 ();
 FILLCELL_X8 FILLER_143_656 ();
 FILLCELL_X32 FILLER_143_685 ();
 FILLCELL_X32 FILLER_143_717 ();
 FILLCELL_X16 FILLER_143_749 ();
 FILLCELL_X8 FILLER_143_765 ();
 FILLCELL_X2 FILLER_143_773 ();
 FILLCELL_X1 FILLER_143_775 ();
 FILLCELL_X1 FILLER_143_794 ();
 FILLCELL_X2 FILLER_143_797 ();
 FILLCELL_X1 FILLER_143_799 ();
 FILLCELL_X8 FILLER_143_802 ();
 FILLCELL_X2 FILLER_143_810 ();
 FILLCELL_X1 FILLER_143_812 ();
 FILLCELL_X1 FILLER_143_849 ();
 FILLCELL_X2 FILLER_143_852 ();
 FILLCELL_X1 FILLER_143_870 ();
 FILLCELL_X1 FILLER_143_875 ();
 FILLCELL_X8 FILLER_143_892 ();
 FILLCELL_X2 FILLER_143_930 ();
 FILLCELL_X1 FILLER_143_932 ();
 FILLCELL_X2 FILLER_143_965 ();
 FILLCELL_X1 FILLER_143_967 ();
 FILLCELL_X16 FILLER_143_1000 ();
 FILLCELL_X1 FILLER_143_1016 ();
 FILLCELL_X2 FILLER_143_1026 ();
 FILLCELL_X1 FILLER_143_1028 ();
 FILLCELL_X1 FILLER_143_1038 ();
 FILLCELL_X4 FILLER_143_1046 ();
 FILLCELL_X1 FILLER_143_1050 ();
 FILLCELL_X4 FILLER_143_1088 ();
 FILLCELL_X1 FILLER_143_1092 ();
 FILLCELL_X1 FILLER_143_1096 ();
 FILLCELL_X4 FILLER_143_1131 ();
 FILLCELL_X4 FILLER_143_1137 ();
 FILLCELL_X2 FILLER_143_1141 ();
 FILLCELL_X4 FILLER_143_1147 ();
 FILLCELL_X2 FILLER_143_1169 ();
 FILLCELL_X1 FILLER_143_1171 ();
 FILLCELL_X32 FILLER_143_1186 ();
 FILLCELL_X32 FILLER_143_1218 ();
 FILLCELL_X8 FILLER_143_1250 ();
 FILLCELL_X2 FILLER_143_1258 ();
 FILLCELL_X16 FILLER_144_1 ();
 FILLCELL_X4 FILLER_144_17 ();
 FILLCELL_X1 FILLER_144_33 ();
 FILLCELL_X4 FILLER_144_62 ();
 FILLCELL_X2 FILLER_144_66 ();
 FILLCELL_X1 FILLER_144_68 ();
 FILLCELL_X4 FILLER_144_76 ();
 FILLCELL_X2 FILLER_144_80 ();
 FILLCELL_X2 FILLER_144_109 ();
 FILLCELL_X1 FILLER_144_111 ();
 FILLCELL_X2 FILLER_144_126 ();
 FILLCELL_X4 FILLER_144_151 ();
 FILLCELL_X1 FILLER_144_155 ();
 FILLCELL_X8 FILLER_144_163 ();
 FILLCELL_X4 FILLER_144_171 ();
 FILLCELL_X2 FILLER_144_202 ();
 FILLCELL_X4 FILLER_144_232 ();
 FILLCELL_X2 FILLER_144_236 ();
 FILLCELL_X1 FILLER_144_238 ();
 FILLCELL_X4 FILLER_144_252 ();
 FILLCELL_X1 FILLER_144_256 ();
 FILLCELL_X32 FILLER_144_284 ();
 FILLCELL_X2 FILLER_144_316 ();
 FILLCELL_X16 FILLER_144_328 ();
 FILLCELL_X4 FILLER_144_344 ();
 FILLCELL_X1 FILLER_144_348 ();
 FILLCELL_X4 FILLER_144_362 ();
 FILLCELL_X4 FILLER_144_369 ();
 FILLCELL_X2 FILLER_144_373 ();
 FILLCELL_X1 FILLER_144_375 ();
 FILLCELL_X4 FILLER_144_399 ();
 FILLCELL_X2 FILLER_144_403 ();
 FILLCELL_X1 FILLER_144_405 ();
 FILLCELL_X8 FILLER_144_413 ();
 FILLCELL_X1 FILLER_144_421 ();
 FILLCELL_X2 FILLER_144_426 ();
 FILLCELL_X1 FILLER_144_501 ();
 FILLCELL_X8 FILLER_144_516 ();
 FILLCELL_X4 FILLER_144_524 ();
 FILLCELL_X1 FILLER_144_528 ();
 FILLCELL_X2 FILLER_144_562 ();
 FILLCELL_X1 FILLER_144_564 ();
 FILLCELL_X4 FILLER_144_573 ();
 FILLCELL_X2 FILLER_144_577 ();
 FILLCELL_X4 FILLER_144_606 ();
 FILLCELL_X1 FILLER_144_610 ();
 FILLCELL_X4 FILLER_144_632 ();
 FILLCELL_X1 FILLER_144_636 ();
 FILLCELL_X4 FILLER_144_657 ();
 FILLCELL_X1 FILLER_144_668 ();
 FILLCELL_X1 FILLER_144_683 ();
 FILLCELL_X32 FILLER_144_704 ();
 FILLCELL_X16 FILLER_144_736 ();
 FILLCELL_X8 FILLER_144_752 ();
 FILLCELL_X4 FILLER_144_760 ();
 FILLCELL_X1 FILLER_144_764 ();
 FILLCELL_X1 FILLER_144_793 ();
 FILLCELL_X2 FILLER_144_804 ();
 FILLCELL_X2 FILLER_144_827 ();
 FILLCELL_X1 FILLER_144_829 ();
 FILLCELL_X4 FILLER_144_832 ();
 FILLCELL_X4 FILLER_144_838 ();
 FILLCELL_X2 FILLER_144_842 ();
 FILLCELL_X4 FILLER_144_860 ();
 FILLCELL_X8 FILLER_144_882 ();
 FILLCELL_X2 FILLER_144_890 ();
 FILLCELL_X2 FILLER_144_910 ();
 FILLCELL_X1 FILLER_144_912 ();
 FILLCELL_X2 FILLER_144_931 ();
 FILLCELL_X4 FILLER_144_935 ();
 FILLCELL_X4 FILLER_144_941 ();
 FILLCELL_X1 FILLER_144_945 ();
 FILLCELL_X2 FILLER_144_948 ();
 FILLCELL_X16 FILLER_144_952 ();
 FILLCELL_X1 FILLER_144_984 ();
 FILLCELL_X16 FILLER_144_992 ();
 FILLCELL_X2 FILLER_144_1027 ();
 FILLCELL_X8 FILLER_144_1038 ();
 FILLCELL_X2 FILLER_144_1052 ();
 FILLCELL_X8 FILLER_144_1060 ();
 FILLCELL_X4 FILLER_144_1068 ();
 FILLCELL_X8 FILLER_144_1081 ();
 FILLCELL_X4 FILLER_144_1089 ();
 FILLCELL_X1 FILLER_144_1093 ();
 FILLCELL_X4 FILLER_144_1110 ();
 FILLCELL_X2 FILLER_144_1114 ();
 FILLCELL_X4 FILLER_144_1118 ();
 FILLCELL_X4 FILLER_144_1152 ();
 FILLCELL_X2 FILLER_144_1156 ();
 FILLCELL_X8 FILLER_144_1160 ();
 FILLCELL_X1 FILLER_144_1168 ();
 FILLCELL_X32 FILLER_144_1188 ();
 FILLCELL_X32 FILLER_144_1220 ();
 FILLCELL_X8 FILLER_144_1252 ();
 FILLCELL_X16 FILLER_145_1 ();
 FILLCELL_X2 FILLER_145_17 ();
 FILLCELL_X8 FILLER_145_39 ();
 FILLCELL_X4 FILLER_145_54 ();
 FILLCELL_X2 FILLER_145_58 ();
 FILLCELL_X1 FILLER_145_60 ();
 FILLCELL_X4 FILLER_145_81 ();
 FILLCELL_X1 FILLER_145_85 ();
 FILLCELL_X4 FILLER_145_93 ();
 FILLCELL_X1 FILLER_145_97 ();
 FILLCELL_X2 FILLER_145_152 ();
 FILLCELL_X1 FILLER_145_154 ();
 FILLCELL_X4 FILLER_145_162 ();
 FILLCELL_X2 FILLER_145_166 ();
 FILLCELL_X32 FILLER_145_175 ();
 FILLCELL_X2 FILLER_145_207 ();
 FILLCELL_X1 FILLER_145_209 ();
 FILLCELL_X16 FILLER_145_217 ();
 FILLCELL_X8 FILLER_145_243 ();
 FILLCELL_X4 FILLER_145_251 ();
 FILLCELL_X1 FILLER_145_255 ();
 FILLCELL_X1 FILLER_145_263 ();
 FILLCELL_X2 FILLER_145_268 ();
 FILLCELL_X8 FILLER_145_297 ();
 FILLCELL_X4 FILLER_145_305 ();
 FILLCELL_X2 FILLER_145_309 ();
 FILLCELL_X1 FILLER_145_331 ();
 FILLCELL_X2 FILLER_145_341 ();
 FILLCELL_X1 FILLER_145_346 ();
 FILLCELL_X1 FILLER_145_355 ();
 FILLCELL_X8 FILLER_145_360 ();
 FILLCELL_X2 FILLER_145_368 ();
 FILLCELL_X1 FILLER_145_370 ();
 FILLCELL_X1 FILLER_145_380 ();
 FILLCELL_X16 FILLER_145_384 ();
 FILLCELL_X2 FILLER_145_414 ();
 FILLCELL_X2 FILLER_145_436 ();
 FILLCELL_X2 FILLER_145_454 ();
 FILLCELL_X4 FILLER_145_482 ();
 FILLCELL_X1 FILLER_145_490 ();
 FILLCELL_X8 FILLER_145_498 ();
 FILLCELL_X2 FILLER_145_506 ();
 FILLCELL_X1 FILLER_145_535 ();
 FILLCELL_X2 FILLER_145_540 ();
 FILLCELL_X2 FILLER_145_558 ();
 FILLCELL_X1 FILLER_145_560 ();
 FILLCELL_X4 FILLER_145_568 ();
 FILLCELL_X1 FILLER_145_572 ();
 FILLCELL_X1 FILLER_145_579 ();
 FILLCELL_X2 FILLER_145_592 ();
 FILLCELL_X1 FILLER_145_594 ();
 FILLCELL_X1 FILLER_145_616 ();
 FILLCELL_X8 FILLER_145_624 ();
 FILLCELL_X4 FILLER_145_632 ();
 FILLCELL_X2 FILLER_145_636 ();
 FILLCELL_X4 FILLER_145_645 ();
 FILLCELL_X1 FILLER_145_653 ();
 FILLCELL_X4 FILLER_145_664 ();
 FILLCELL_X2 FILLER_145_668 ();
 FILLCELL_X1 FILLER_145_670 ();
 FILLCELL_X4 FILLER_145_678 ();
 FILLCELL_X2 FILLER_145_682 ();
 FILLCELL_X1 FILLER_145_684 ();
 FILLCELL_X2 FILLER_145_689 ();
 FILLCELL_X1 FILLER_145_691 ();
 FILLCELL_X32 FILLER_145_695 ();
 FILLCELL_X32 FILLER_145_727 ();
 FILLCELL_X4 FILLER_145_759 ();
 FILLCELL_X2 FILLER_145_763 ();
 FILLCELL_X1 FILLER_145_765 ();
 FILLCELL_X1 FILLER_145_788 ();
 FILLCELL_X1 FILLER_145_791 ();
 FILLCELL_X1 FILLER_145_824 ();
 FILLCELL_X16 FILLER_145_841 ();
 FILLCELL_X4 FILLER_145_857 ();
 FILLCELL_X2 FILLER_145_861 ();
 FILLCELL_X1 FILLER_145_863 ();
 FILLCELL_X16 FILLER_145_866 ();
 FILLCELL_X1 FILLER_145_882 ();
 FILLCELL_X8 FILLER_145_917 ();
 FILLCELL_X2 FILLER_145_925 ();
 FILLCELL_X1 FILLER_145_927 ();
 FILLCELL_X2 FILLER_145_930 ();
 FILLCELL_X4 FILLER_145_962 ();
 FILLCELL_X1 FILLER_145_966 ();
 FILLCELL_X8 FILLER_145_969 ();
 FILLCELL_X4 FILLER_145_977 ();
 FILLCELL_X4 FILLER_145_983 ();
 FILLCELL_X1 FILLER_145_1025 ();
 FILLCELL_X2 FILLER_145_1042 ();
 FILLCELL_X1 FILLER_145_1044 ();
 FILLCELL_X1 FILLER_145_1122 ();
 FILLCELL_X16 FILLER_145_1133 ();
 FILLCELL_X2 FILLER_145_1149 ();
 FILLCELL_X1 FILLER_145_1151 ();
 FILLCELL_X1 FILLER_145_1183 ();
 FILLCELL_X32 FILLER_145_1195 ();
 FILLCELL_X32 FILLER_145_1227 ();
 FILLCELL_X1 FILLER_145_1259 ();
 FILLCELL_X16 FILLER_146_1 ();
 FILLCELL_X1 FILLER_146_17 ();
 FILLCELL_X2 FILLER_146_25 ();
 FILLCELL_X1 FILLER_146_27 ();
 FILLCELL_X2 FILLER_146_35 ();
 FILLCELL_X1 FILLER_146_37 ();
 FILLCELL_X8 FILLER_146_52 ();
 FILLCELL_X1 FILLER_146_60 ();
 FILLCELL_X8 FILLER_146_88 ();
 FILLCELL_X4 FILLER_146_96 ();
 FILLCELL_X2 FILLER_146_100 ();
 FILLCELL_X1 FILLER_146_102 ();
 FILLCELL_X1 FILLER_146_110 ();
 FILLCELL_X4 FILLER_146_118 ();
 FILLCELL_X2 FILLER_146_122 ();
 FILLCELL_X8 FILLER_146_138 ();
 FILLCELL_X1 FILLER_146_146 ();
 FILLCELL_X1 FILLER_146_167 ();
 FILLCELL_X2 FILLER_146_195 ();
 FILLCELL_X1 FILLER_146_197 ();
 FILLCELL_X8 FILLER_146_218 ();
 FILLCELL_X2 FILLER_146_226 ();
 FILLCELL_X1 FILLER_146_228 ();
 FILLCELL_X2 FILLER_146_270 ();
 FILLCELL_X4 FILLER_146_279 ();
 FILLCELL_X8 FILLER_146_287 ();
 FILLCELL_X2 FILLER_146_295 ();
 FILLCELL_X1 FILLER_146_297 ();
 FILLCELL_X1 FILLER_146_318 ();
 FILLCELL_X1 FILLER_146_348 ();
 FILLCELL_X2 FILLER_146_372 ();
 FILLCELL_X1 FILLER_146_374 ();
 FILLCELL_X2 FILLER_146_400 ();
 FILLCELL_X1 FILLER_146_409 ();
 FILLCELL_X8 FILLER_146_520 ();
 FILLCELL_X4 FILLER_146_528 ();
 FILLCELL_X2 FILLER_146_532 ();
 FILLCELL_X1 FILLER_146_534 ();
 FILLCELL_X1 FILLER_146_539 ();
 FILLCELL_X16 FILLER_146_543 ();
 FILLCELL_X8 FILLER_146_559 ();
 FILLCELL_X2 FILLER_146_567 ();
 FILLCELL_X1 FILLER_146_569 ();
 FILLCELL_X4 FILLER_146_610 ();
 FILLCELL_X2 FILLER_146_632 ();
 FILLCELL_X1 FILLER_146_634 ();
 FILLCELL_X1 FILLER_146_655 ();
 FILLCELL_X8 FILLER_146_670 ();
 FILLCELL_X32 FILLER_146_702 ();
 FILLCELL_X16 FILLER_146_734 ();
 FILLCELL_X8 FILLER_146_750 ();
 FILLCELL_X4 FILLER_146_758 ();
 FILLCELL_X1 FILLER_146_762 ();
 FILLCELL_X2 FILLER_146_781 ();
 FILLCELL_X16 FILLER_146_785 ();
 FILLCELL_X4 FILLER_146_801 ();
 FILLCELL_X2 FILLER_146_805 ();
 FILLCELL_X16 FILLER_146_825 ();
 FILLCELL_X4 FILLER_146_841 ();
 FILLCELL_X2 FILLER_146_895 ();
 FILLCELL_X2 FILLER_146_899 ();
 FILLCELL_X1 FILLER_146_901 ();
 FILLCELL_X1 FILLER_146_918 ();
 FILLCELL_X4 FILLER_146_951 ();
 FILLCELL_X1 FILLER_146_955 ();
 FILLCELL_X2 FILLER_146_974 ();
 FILLCELL_X1 FILLER_146_976 ();
 FILLCELL_X4 FILLER_146_997 ();
 FILLCELL_X8 FILLER_146_1003 ();
 FILLCELL_X1 FILLER_146_1013 ();
 FILLCELL_X1 FILLER_146_1017 ();
 FILLCELL_X4 FILLER_146_1020 ();
 FILLCELL_X4 FILLER_146_1026 ();
 FILLCELL_X2 FILLER_146_1030 ();
 FILLCELL_X1 FILLER_146_1034 ();
 FILLCELL_X2 FILLER_146_1038 ();
 FILLCELL_X1 FILLER_146_1053 ();
 FILLCELL_X4 FILLER_146_1070 ();
 FILLCELL_X2 FILLER_146_1090 ();
 FILLCELL_X8 FILLER_146_1094 ();
 FILLCELL_X2 FILLER_146_1102 ();
 FILLCELL_X1 FILLER_146_1104 ();
 FILLCELL_X1 FILLER_146_1109 ();
 FILLCELL_X8 FILLER_146_1112 ();
 FILLCELL_X2 FILLER_146_1120 ();
 FILLCELL_X4 FILLER_146_1140 ();
 FILLCELL_X2 FILLER_146_1144 ();
 FILLCELL_X4 FILLER_146_1148 ();
 FILLCELL_X1 FILLER_146_1152 ();
 FILLCELL_X4 FILLER_146_1155 ();
 FILLCELL_X2 FILLER_146_1159 ();
 FILLCELL_X4 FILLER_146_1163 ();
 FILLCELL_X2 FILLER_146_1167 ();
 FILLCELL_X32 FILLER_146_1202 ();
 FILLCELL_X16 FILLER_146_1234 ();
 FILLCELL_X8 FILLER_146_1250 ();
 FILLCELL_X2 FILLER_146_1258 ();
 FILLCELL_X4 FILLER_147_1 ();
 FILLCELL_X1 FILLER_147_45 ();
 FILLCELL_X8 FILLER_147_53 ();
 FILLCELL_X1 FILLER_147_61 ();
 FILLCELL_X2 FILLER_147_97 ();
 FILLCELL_X4 FILLER_147_113 ();
 FILLCELL_X4 FILLER_147_121 ();
 FILLCELL_X1 FILLER_147_125 ();
 FILLCELL_X1 FILLER_147_153 ();
 FILLCELL_X2 FILLER_147_168 ();
 FILLCELL_X1 FILLER_147_170 ();
 FILLCELL_X1 FILLER_147_211 ();
 FILLCELL_X4 FILLER_147_232 ();
 FILLCELL_X1 FILLER_147_236 ();
 FILLCELL_X2 FILLER_147_268 ();
 FILLCELL_X16 FILLER_147_297 ();
 FILLCELL_X2 FILLER_147_320 ();
 FILLCELL_X1 FILLER_147_326 ();
 FILLCELL_X32 FILLER_147_335 ();
 FILLCELL_X1 FILLER_147_367 ();
 FILLCELL_X1 FILLER_147_380 ();
 FILLCELL_X1 FILLER_147_401 ();
 FILLCELL_X4 FILLER_147_405 ();
 FILLCELL_X2 FILLER_147_409 ();
 FILLCELL_X1 FILLER_147_411 ();
 FILLCELL_X2 FILLER_147_416 ();
 FILLCELL_X1 FILLER_147_434 ();
 FILLCELL_X1 FILLER_147_449 ();
 FILLCELL_X8 FILLER_147_464 ();
 FILLCELL_X4 FILLER_147_472 ();
 FILLCELL_X4 FILLER_147_481 ();
 FILLCELL_X1 FILLER_147_485 ();
 FILLCELL_X4 FILLER_147_490 ();
 FILLCELL_X2 FILLER_147_501 ();
 FILLCELL_X1 FILLER_147_506 ();
 FILLCELL_X1 FILLER_147_532 ();
 FILLCELL_X2 FILLER_147_560 ();
 FILLCELL_X2 FILLER_147_582 ();
 FILLCELL_X8 FILLER_147_601 ();
 FILLCELL_X4 FILLER_147_609 ();
 FILLCELL_X8 FILLER_147_617 ();
 FILLCELL_X4 FILLER_147_631 ();
 FILLCELL_X1 FILLER_147_635 ();
 FILLCELL_X2 FILLER_147_640 ();
 FILLCELL_X1 FILLER_147_642 ();
 FILLCELL_X16 FILLER_147_646 ();
 FILLCELL_X8 FILLER_147_662 ();
 FILLCELL_X1 FILLER_147_670 ();
 FILLCELL_X8 FILLER_147_685 ();
 FILLCELL_X32 FILLER_147_696 ();
 FILLCELL_X32 FILLER_147_728 ();
 FILLCELL_X4 FILLER_147_760 ();
 FILLCELL_X1 FILLER_147_764 ();
 FILLCELL_X4 FILLER_147_783 ();
 FILLCELL_X1 FILLER_147_805 ();
 FILLCELL_X1 FILLER_147_826 ();
 FILLCELL_X8 FILLER_147_843 ();
 FILLCELL_X2 FILLER_147_851 ();
 FILLCELL_X16 FILLER_147_885 ();
 FILLCELL_X4 FILLER_147_901 ();
 FILLCELL_X2 FILLER_147_905 ();
 FILLCELL_X1 FILLER_147_907 ();
 FILLCELL_X4 FILLER_147_911 ();
 FILLCELL_X2 FILLER_147_915 ();
 FILLCELL_X8 FILLER_147_920 ();
 FILLCELL_X4 FILLER_147_928 ();
 FILLCELL_X2 FILLER_147_932 ();
 FILLCELL_X1 FILLER_147_934 ();
 FILLCELL_X4 FILLER_147_937 ();
 FILLCELL_X2 FILLER_147_941 ();
 FILLCELL_X1 FILLER_147_943 ();
 FILLCELL_X1 FILLER_147_946 ();
 FILLCELL_X4 FILLER_147_963 ();
 FILLCELL_X2 FILLER_147_967 ();
 FILLCELL_X1 FILLER_147_969 ();
 FILLCELL_X1 FILLER_147_1023 ();
 FILLCELL_X4 FILLER_147_1043 ();
 FILLCELL_X8 FILLER_147_1063 ();
 FILLCELL_X4 FILLER_147_1071 ();
 FILLCELL_X8 FILLER_147_1077 ();
 FILLCELL_X4 FILLER_147_1085 ();
 FILLCELL_X1 FILLER_147_1091 ();
 FILLCELL_X4 FILLER_147_1105 ();
 FILLCELL_X2 FILLER_147_1109 ();
 FILLCELL_X4 FILLER_147_1121 ();
 FILLCELL_X1 FILLER_147_1125 ();
 FILLCELL_X4 FILLER_147_1166 ();
 FILLCELL_X1 FILLER_147_1170 ();
 FILLCELL_X4 FILLER_147_1174 ();
 FILLCELL_X1 FILLER_147_1178 ();
 FILLCELL_X32 FILLER_147_1197 ();
 FILLCELL_X16 FILLER_147_1229 ();
 FILLCELL_X8 FILLER_147_1245 ();
 FILLCELL_X4 FILLER_147_1253 ();
 FILLCELL_X2 FILLER_147_1257 ();
 FILLCELL_X1 FILLER_147_1259 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X4 FILLER_148_40 ();
 FILLCELL_X2 FILLER_148_44 ();
 FILLCELL_X1 FILLER_148_46 ();
 FILLCELL_X4 FILLER_148_61 ();
 FILLCELL_X8 FILLER_148_72 ();
 FILLCELL_X4 FILLER_148_80 ();
 FILLCELL_X1 FILLER_148_84 ();
 FILLCELL_X4 FILLER_148_123 ();
 FILLCELL_X1 FILLER_148_127 ();
 FILLCELL_X4 FILLER_148_154 ();
 FILLCELL_X2 FILLER_148_158 ();
 FILLCELL_X4 FILLER_148_167 ();
 FILLCELL_X1 FILLER_148_171 ();
 FILLCELL_X4 FILLER_148_179 ();
 FILLCELL_X1 FILLER_148_201 ();
 FILLCELL_X8 FILLER_148_209 ();
 FILLCELL_X1 FILLER_148_217 ();
 FILLCELL_X4 FILLER_148_222 ();
 FILLCELL_X2 FILLER_148_226 ();
 FILLCELL_X1 FILLER_148_228 ();
 FILLCELL_X4 FILLER_148_236 ();
 FILLCELL_X2 FILLER_148_240 ();
 FILLCELL_X4 FILLER_148_249 ();
 FILLCELL_X2 FILLER_148_253 ();
 FILLCELL_X1 FILLER_148_269 ();
 FILLCELL_X1 FILLER_148_298 ();
 FILLCELL_X4 FILLER_148_360 ();
 FILLCELL_X4 FILLER_148_404 ();
 FILLCELL_X2 FILLER_148_408 ();
 FILLCELL_X1 FILLER_148_410 ();
 FILLCELL_X4 FILLER_148_418 ();
 FILLCELL_X2 FILLER_148_445 ();
 FILLCELL_X1 FILLER_148_447 ();
 FILLCELL_X8 FILLER_148_455 ();
 FILLCELL_X8 FILLER_148_474 ();
 FILLCELL_X4 FILLER_148_482 ();
 FILLCELL_X4 FILLER_148_513 ();
 FILLCELL_X1 FILLER_148_517 ();
 FILLCELL_X8 FILLER_148_525 ();
 FILLCELL_X1 FILLER_148_537 ();
 FILLCELL_X2 FILLER_148_541 ();
 FILLCELL_X2 FILLER_148_550 ();
 FILLCELL_X4 FILLER_148_559 ();
 FILLCELL_X2 FILLER_148_563 ();
 FILLCELL_X2 FILLER_148_572 ();
 FILLCELL_X1 FILLER_148_574 ();
 FILLCELL_X4 FILLER_148_578 ();
 FILLCELL_X2 FILLER_148_582 ();
 FILLCELL_X1 FILLER_148_588 ();
 FILLCELL_X4 FILLER_148_603 ();
 FILLCELL_X2 FILLER_148_607 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X4 FILLER_148_632 ();
 FILLCELL_X2 FILLER_148_636 ();
 FILLCELL_X1 FILLER_148_638 ();
 FILLCELL_X1 FILLER_148_659 ();
 FILLCELL_X2 FILLER_148_681 ();
 FILLCELL_X1 FILLER_148_683 ();
 FILLCELL_X32 FILLER_148_691 ();
 FILLCELL_X32 FILLER_148_723 ();
 FILLCELL_X8 FILLER_148_755 ();
 FILLCELL_X8 FILLER_148_765 ();
 FILLCELL_X4 FILLER_148_773 ();
 FILLCELL_X1 FILLER_148_777 ();
 FILLCELL_X4 FILLER_148_788 ();
 FILLCELL_X2 FILLER_148_792 ();
 FILLCELL_X2 FILLER_148_796 ();
 FILLCELL_X4 FILLER_148_814 ();
 FILLCELL_X8 FILLER_148_882 ();
 FILLCELL_X2 FILLER_148_890 ();
 FILLCELL_X1 FILLER_148_892 ();
 FILLCELL_X2 FILLER_148_928 ();
 FILLCELL_X4 FILLER_148_954 ();
 FILLCELL_X1 FILLER_148_967 ();
 FILLCELL_X1 FILLER_148_980 ();
 FILLCELL_X4 FILLER_148_983 ();
 FILLCELL_X4 FILLER_148_989 ();
 FILLCELL_X2 FILLER_148_993 ();
 FILLCELL_X1 FILLER_148_995 ();
 FILLCELL_X4 FILLER_148_1014 ();
 FILLCELL_X2 FILLER_148_1018 ();
 FILLCELL_X4 FILLER_148_1036 ();
 FILLCELL_X2 FILLER_148_1040 ();
 FILLCELL_X2 FILLER_148_1074 ();
 FILLCELL_X4 FILLER_148_1078 ();
 FILLCELL_X1 FILLER_148_1082 ();
 FILLCELL_X4 FILLER_148_1085 ();
 FILLCELL_X1 FILLER_148_1089 ();
 FILLCELL_X1 FILLER_148_1095 ();
 FILLCELL_X8 FILLER_148_1114 ();
 FILLCELL_X2 FILLER_148_1122 ();
 FILLCELL_X1 FILLER_148_1124 ();
 FILLCELL_X8 FILLER_148_1127 ();
 FILLCELL_X4 FILLER_148_1135 ();
 FILLCELL_X1 FILLER_148_1141 ();
 FILLCELL_X1 FILLER_148_1144 ();
 FILLCELL_X1 FILLER_148_1155 ();
 FILLCELL_X8 FILLER_148_1174 ();
 FILLCELL_X4 FILLER_148_1182 ();
 FILLCELL_X32 FILLER_148_1189 ();
 FILLCELL_X32 FILLER_148_1221 ();
 FILLCELL_X4 FILLER_148_1253 ();
 FILLCELL_X2 FILLER_148_1257 ();
 FILLCELL_X1 FILLER_148_1259 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X2 FILLER_149_33 ();
 FILLCELL_X1 FILLER_149_62 ();
 FILLCELL_X8 FILLER_149_83 ();
 FILLCELL_X4 FILLER_149_112 ();
 FILLCELL_X1 FILLER_149_116 ();
 FILLCELL_X4 FILLER_149_131 ();
 FILLCELL_X8 FILLER_149_142 ();
 FILLCELL_X4 FILLER_149_150 ();
 FILLCELL_X2 FILLER_149_154 ();
 FILLCELL_X2 FILLER_149_183 ();
 FILLCELL_X1 FILLER_149_185 ();
 FILLCELL_X16 FILLER_149_200 ();
 FILLCELL_X16 FILLER_149_223 ();
 FILLCELL_X4 FILLER_149_239 ();
 FILLCELL_X2 FILLER_149_243 ();
 FILLCELL_X2 FILLER_149_252 ();
 FILLCELL_X4 FILLER_149_280 ();
 FILLCELL_X2 FILLER_149_284 ();
 FILLCELL_X2 FILLER_149_293 ();
 FILLCELL_X1 FILLER_149_295 ();
 FILLCELL_X8 FILLER_149_310 ();
 FILLCELL_X4 FILLER_149_318 ();
 FILLCELL_X1 FILLER_149_322 ();
 FILLCELL_X1 FILLER_149_354 ();
 FILLCELL_X2 FILLER_149_362 ();
 FILLCELL_X1 FILLER_149_364 ();
 FILLCELL_X4 FILLER_149_381 ();
 FILLCELL_X2 FILLER_149_385 ();
 FILLCELL_X2 FILLER_149_397 ();
 FILLCELL_X2 FILLER_149_410 ();
 FILLCELL_X1 FILLER_149_412 ();
 FILLCELL_X4 FILLER_149_482 ();
 FILLCELL_X2 FILLER_149_486 ();
 FILLCELL_X8 FILLER_149_492 ();
 FILLCELL_X2 FILLER_149_503 ();
 FILLCELL_X1 FILLER_149_505 ();
 FILLCELL_X4 FILLER_149_513 ();
 FILLCELL_X2 FILLER_149_517 ();
 FILLCELL_X1 FILLER_149_519 ();
 FILLCELL_X4 FILLER_149_527 ();
 FILLCELL_X1 FILLER_149_558 ();
 FILLCELL_X2 FILLER_149_602 ();
 FILLCELL_X4 FILLER_149_608 ();
 FILLCELL_X2 FILLER_149_612 ();
 FILLCELL_X1 FILLER_149_614 ();
 FILLCELL_X2 FILLER_149_618 ();
 FILLCELL_X1 FILLER_149_620 ();
 FILLCELL_X4 FILLER_149_635 ();
 FILLCELL_X1 FILLER_149_639 ();
 FILLCELL_X8 FILLER_149_647 ();
 FILLCELL_X4 FILLER_149_655 ();
 FILLCELL_X2 FILLER_149_659 ();
 FILLCELL_X1 FILLER_149_661 ();
 FILLCELL_X1 FILLER_149_669 ();
 FILLCELL_X2 FILLER_149_677 ();
 FILLCELL_X1 FILLER_149_679 ();
 FILLCELL_X32 FILLER_149_700 ();
 FILLCELL_X32 FILLER_149_732 ();
 FILLCELL_X4 FILLER_149_764 ();
 FILLCELL_X2 FILLER_149_768 ();
 FILLCELL_X16 FILLER_149_780 ();
 FILLCELL_X2 FILLER_149_796 ();
 FILLCELL_X8 FILLER_149_814 ();
 FILLCELL_X4 FILLER_149_822 ();
 FILLCELL_X2 FILLER_149_826 ();
 FILLCELL_X16 FILLER_149_860 ();
 FILLCELL_X4 FILLER_149_876 ();
 FILLCELL_X16 FILLER_149_896 ();
 FILLCELL_X4 FILLER_149_912 ();
 FILLCELL_X2 FILLER_149_916 ();
 FILLCELL_X8 FILLER_149_937 ();
 FILLCELL_X2 FILLER_149_945 ();
 FILLCELL_X16 FILLER_149_963 ();
 FILLCELL_X2 FILLER_149_979 ();
 FILLCELL_X2 FILLER_149_997 ();
 FILLCELL_X4 FILLER_149_1001 ();
 FILLCELL_X2 FILLER_149_1005 ();
 FILLCELL_X4 FILLER_149_1009 ();
 FILLCELL_X16 FILLER_149_1015 ();
 FILLCELL_X1 FILLER_149_1031 ();
 FILLCELL_X4 FILLER_149_1067 ();
 FILLCELL_X8 FILLER_149_1073 ();
 FILLCELL_X2 FILLER_149_1110 ();
 FILLCELL_X2 FILLER_149_1144 ();
 FILLCELL_X1 FILLER_149_1148 ();
 FILLCELL_X4 FILLER_149_1168 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X2 FILLER_149_1257 ();
 FILLCELL_X1 FILLER_149_1259 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X1 FILLER_150_33 ();
 FILLCELL_X8 FILLER_150_61 ();
 FILLCELL_X4 FILLER_150_69 ();
 FILLCELL_X1 FILLER_150_73 ();
 FILLCELL_X2 FILLER_150_115 ();
 FILLCELL_X4 FILLER_150_138 ();
 FILLCELL_X2 FILLER_150_142 ();
 FILLCELL_X1 FILLER_150_144 ();
 FILLCELL_X1 FILLER_150_185 ();
 FILLCELL_X4 FILLER_150_200 ();
 FILLCELL_X2 FILLER_150_204 ();
 FILLCELL_X2 FILLER_150_226 ();
 FILLCELL_X1 FILLER_150_228 ();
 FILLCELL_X1 FILLER_150_234 ();
 FILLCELL_X4 FILLER_150_262 ();
 FILLCELL_X1 FILLER_150_266 ();
 FILLCELL_X1 FILLER_150_270 ();
 FILLCELL_X4 FILLER_150_278 ();
 FILLCELL_X8 FILLER_150_302 ();
 FILLCELL_X4 FILLER_150_310 ();
 FILLCELL_X2 FILLER_150_314 ();
 FILLCELL_X2 FILLER_150_323 ();
 FILLCELL_X1 FILLER_150_325 ();
 FILLCELL_X1 FILLER_150_330 ();
 FILLCELL_X4 FILLER_150_334 ();
 FILLCELL_X2 FILLER_150_338 ();
 FILLCELL_X2 FILLER_150_344 ();
 FILLCELL_X1 FILLER_150_349 ();
 FILLCELL_X2 FILLER_150_357 ();
 FILLCELL_X1 FILLER_150_359 ();
 FILLCELL_X4 FILLER_150_380 ();
 FILLCELL_X2 FILLER_150_397 ();
 FILLCELL_X4 FILLER_150_420 ();
 FILLCELL_X8 FILLER_150_431 ();
 FILLCELL_X2 FILLER_150_439 ();
 FILLCELL_X1 FILLER_150_455 ();
 FILLCELL_X16 FILLER_150_470 ();
 FILLCELL_X4 FILLER_150_506 ();
 FILLCELL_X2 FILLER_150_510 ();
 FILLCELL_X1 FILLER_150_526 ();
 FILLCELL_X4 FILLER_150_534 ();
 FILLCELL_X1 FILLER_150_538 ();
 FILLCELL_X1 FILLER_150_546 ();
 FILLCELL_X16 FILLER_150_561 ();
 FILLCELL_X1 FILLER_150_577 ();
 FILLCELL_X4 FILLER_150_583 ();
 FILLCELL_X4 FILLER_150_591 ();
 FILLCELL_X2 FILLER_150_595 ();
 FILLCELL_X2 FILLER_150_620 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X1 FILLER_150_639 ();
 FILLCELL_X4 FILLER_150_647 ();
 FILLCELL_X1 FILLER_150_651 ();
 FILLCELL_X4 FILLER_150_659 ();
 FILLCELL_X32 FILLER_150_683 ();
 FILLCELL_X32 FILLER_150_715 ();
 FILLCELL_X16 FILLER_150_747 ();
 FILLCELL_X8 FILLER_150_763 ();
 FILLCELL_X2 FILLER_150_803 ();
 FILLCELL_X1 FILLER_150_805 ();
 FILLCELL_X16 FILLER_150_827 ();
 FILLCELL_X4 FILLER_150_843 ();
 FILLCELL_X16 FILLER_150_853 ();
 FILLCELL_X2 FILLER_150_869 ();
 FILLCELL_X2 FILLER_150_873 ();
 FILLCELL_X2 FILLER_150_883 ();
 FILLCELL_X2 FILLER_150_904 ();
 FILLCELL_X1 FILLER_150_906 ();
 FILLCELL_X1 FILLER_150_926 ();
 FILLCELL_X1 FILLER_150_946 ();
 FILLCELL_X4 FILLER_150_960 ();
 FILLCELL_X1 FILLER_150_966 ();
 FILLCELL_X4 FILLER_150_978 ();
 FILLCELL_X4 FILLER_150_984 ();
 FILLCELL_X2 FILLER_150_988 ();
 FILLCELL_X1 FILLER_150_993 ();
 FILLCELL_X4 FILLER_150_996 ();
 FILLCELL_X2 FILLER_150_1008 ();
 FILLCELL_X4 FILLER_150_1035 ();
 FILLCELL_X1 FILLER_150_1039 ();
 FILLCELL_X4 FILLER_150_1045 ();
 FILLCELL_X8 FILLER_150_1068 ();
 FILLCELL_X2 FILLER_150_1105 ();
 FILLCELL_X2 FILLER_150_1112 ();
 FILLCELL_X8 FILLER_150_1148 ();
 FILLCELL_X1 FILLER_150_1187 ();
 FILLCELL_X32 FILLER_150_1191 ();
 FILLCELL_X32 FILLER_150_1223 ();
 FILLCELL_X4 FILLER_150_1255 ();
 FILLCELL_X1 FILLER_150_1259 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X8 FILLER_151_65 ();
 FILLCELL_X2 FILLER_151_73 ();
 FILLCELL_X1 FILLER_151_82 ();
 FILLCELL_X32 FILLER_151_110 ();
 FILLCELL_X16 FILLER_151_142 ();
 FILLCELL_X2 FILLER_151_158 ();
 FILLCELL_X1 FILLER_151_160 ();
 FILLCELL_X8 FILLER_151_175 ();
 FILLCELL_X4 FILLER_151_183 ();
 FILLCELL_X4 FILLER_151_208 ();
 FILLCELL_X4 FILLER_151_233 ();
 FILLCELL_X2 FILLER_151_237 ();
 FILLCELL_X4 FILLER_151_259 ();
 FILLCELL_X8 FILLER_151_303 ();
 FILLCELL_X2 FILLER_151_311 ();
 FILLCELL_X1 FILLER_151_313 ();
 FILLCELL_X8 FILLER_151_354 ();
 FILLCELL_X4 FILLER_151_362 ();
 FILLCELL_X2 FILLER_151_366 ();
 FILLCELL_X4 FILLER_151_404 ();
 FILLCELL_X8 FILLER_151_415 ();
 FILLCELL_X1 FILLER_151_423 ();
 FILLCELL_X1 FILLER_151_448 ();
 FILLCELL_X1 FILLER_151_452 ();
 FILLCELL_X2 FILLER_151_460 ();
 FILLCELL_X1 FILLER_151_462 ();
 FILLCELL_X8 FILLER_151_475 ();
 FILLCELL_X2 FILLER_151_483 ();
 FILLCELL_X2 FILLER_151_489 ();
 FILLCELL_X4 FILLER_151_521 ();
 FILLCELL_X8 FILLER_151_532 ();
 FILLCELL_X2 FILLER_151_540 ();
 FILLCELL_X1 FILLER_151_542 ();
 FILLCELL_X1 FILLER_151_547 ();
 FILLCELL_X2 FILLER_151_551 ();
 FILLCELL_X1 FILLER_151_553 ();
 FILLCELL_X2 FILLER_151_558 ();
 FILLCELL_X8 FILLER_151_563 ();
 FILLCELL_X8 FILLER_151_603 ();
 FILLCELL_X4 FILLER_151_611 ();
 FILLCELL_X1 FILLER_151_615 ();
 FILLCELL_X1 FILLER_151_675 ();
 FILLCELL_X32 FILLER_151_682 ();
 FILLCELL_X32 FILLER_151_714 ();
 FILLCELL_X8 FILLER_151_746 ();
 FILLCELL_X4 FILLER_151_754 ();
 FILLCELL_X1 FILLER_151_758 ();
 FILLCELL_X1 FILLER_151_775 ();
 FILLCELL_X2 FILLER_151_792 ();
 FILLCELL_X1 FILLER_151_794 ();
 FILLCELL_X2 FILLER_151_799 ();
 FILLCELL_X2 FILLER_151_817 ();
 FILLCELL_X1 FILLER_151_819 ();
 FILLCELL_X2 FILLER_151_868 ();
 FILLCELL_X8 FILLER_151_886 ();
 FILLCELL_X4 FILLER_151_918 ();
 FILLCELL_X2 FILLER_151_922 ();
 FILLCELL_X1 FILLER_151_924 ();
 FILLCELL_X1 FILLER_151_928 ();
 FILLCELL_X1 FILLER_151_932 ();
 FILLCELL_X1 FILLER_151_936 ();
 FILLCELL_X2 FILLER_151_940 ();
 FILLCELL_X2 FILLER_151_947 ();
 FILLCELL_X1 FILLER_151_949 ();
 FILLCELL_X2 FILLER_151_1041 ();
 FILLCELL_X8 FILLER_151_1049 ();
 FILLCELL_X1 FILLER_151_1057 ();
 FILLCELL_X4 FILLER_151_1061 ();
 FILLCELL_X8 FILLER_151_1083 ();
 FILLCELL_X2 FILLER_151_1091 ();
 FILLCELL_X2 FILLER_151_1096 ();
 FILLCELL_X1 FILLER_151_1098 ();
 FILLCELL_X4 FILLER_151_1118 ();
 FILLCELL_X2 FILLER_151_1122 ();
 FILLCELL_X1 FILLER_151_1124 ();
 FILLCELL_X4 FILLER_151_1127 ();
 FILLCELL_X1 FILLER_151_1131 ();
 FILLCELL_X8 FILLER_151_1168 ();
 FILLCELL_X2 FILLER_151_1176 ();
 FILLCELL_X1 FILLER_151_1178 ();
 FILLCELL_X32 FILLER_151_1196 ();
 FILLCELL_X32 FILLER_151_1228 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X4 FILLER_152_65 ();
 FILLCELL_X2 FILLER_152_69 ();
 FILLCELL_X1 FILLER_152_71 ();
 FILLCELL_X16 FILLER_152_80 ();
 FILLCELL_X2 FILLER_152_96 ();
 FILLCELL_X1 FILLER_152_132 ();
 FILLCELL_X4 FILLER_152_140 ();
 FILLCELL_X1 FILLER_152_235 ();
 FILLCELL_X4 FILLER_152_243 ();
 FILLCELL_X1 FILLER_152_247 ();
 FILLCELL_X8 FILLER_152_255 ();
 FILLCELL_X8 FILLER_152_270 ();
 FILLCELL_X1 FILLER_152_278 ();
 FILLCELL_X1 FILLER_152_286 ();
 FILLCELL_X2 FILLER_152_294 ();
 FILLCELL_X1 FILLER_152_303 ();
 FILLCELL_X1 FILLER_152_324 ();
 FILLCELL_X8 FILLER_152_332 ();
 FILLCELL_X2 FILLER_152_340 ();
 FILLCELL_X4 FILLER_152_349 ();
 FILLCELL_X2 FILLER_152_360 ();
 FILLCELL_X2 FILLER_152_389 ();
 FILLCELL_X1 FILLER_152_391 ();
 FILLCELL_X2 FILLER_152_412 ();
 FILLCELL_X1 FILLER_152_414 ();
 FILLCELL_X8 FILLER_152_427 ();
 FILLCELL_X1 FILLER_152_435 ();
 FILLCELL_X8 FILLER_152_443 ();
 FILLCELL_X2 FILLER_152_451 ();
 FILLCELL_X4 FILLER_152_473 ();
 FILLCELL_X8 FILLER_152_497 ();
 FILLCELL_X4 FILLER_152_505 ();
 FILLCELL_X1 FILLER_152_509 ();
 FILLCELL_X4 FILLER_152_590 ();
 FILLCELL_X1 FILLER_152_594 ();
 FILLCELL_X4 FILLER_152_602 ();
 FILLCELL_X2 FILLER_152_606 ();
 FILLCELL_X1 FILLER_152_608 ();
 FILLCELL_X2 FILLER_152_622 ();
 FILLCELL_X4 FILLER_152_635 ();
 FILLCELL_X1 FILLER_152_639 ();
 FILLCELL_X4 FILLER_152_647 ();
 FILLCELL_X2 FILLER_152_651 ();
 FILLCELL_X1 FILLER_152_672 ();
 FILLCELL_X32 FILLER_152_697 ();
 FILLCELL_X32 FILLER_152_729 ();
 FILLCELL_X4 FILLER_152_761 ();
 FILLCELL_X1 FILLER_152_771 ();
 FILLCELL_X32 FILLER_152_778 ();
 FILLCELL_X4 FILLER_152_813 ();
 FILLCELL_X2 FILLER_152_833 ();
 FILLCELL_X8 FILLER_152_854 ();
 FILLCELL_X4 FILLER_152_862 ();
 FILLCELL_X1 FILLER_152_866 ();
 FILLCELL_X1 FILLER_152_879 ();
 FILLCELL_X2 FILLER_152_898 ();
 FILLCELL_X1 FILLER_152_900 ();
 FILLCELL_X1 FILLER_152_904 ();
 FILLCELL_X1 FILLER_152_937 ();
 FILLCELL_X2 FILLER_152_940 ();
 FILLCELL_X1 FILLER_152_942 ();
 FILLCELL_X1 FILLER_152_950 ();
 FILLCELL_X8 FILLER_152_957 ();
 FILLCELL_X4 FILLER_152_965 ();
 FILLCELL_X1 FILLER_152_969 ();
 FILLCELL_X2 FILLER_152_976 ();
 FILLCELL_X1 FILLER_152_978 ();
 FILLCELL_X8 FILLER_152_981 ();
 FILLCELL_X1 FILLER_152_989 ();
 FILLCELL_X2 FILLER_152_993 ();
 FILLCELL_X1 FILLER_152_995 ();
 FILLCELL_X4 FILLER_152_998 ();
 FILLCELL_X1 FILLER_152_1002 ();
 FILLCELL_X4 FILLER_152_1009 ();
 FILLCELL_X4 FILLER_152_1030 ();
 FILLCELL_X1 FILLER_152_1034 ();
 FILLCELL_X2 FILLER_152_1054 ();
 FILLCELL_X1 FILLER_152_1056 ();
 FILLCELL_X8 FILLER_152_1060 ();
 FILLCELL_X2 FILLER_152_1068 ();
 FILLCELL_X2 FILLER_152_1072 ();
 FILLCELL_X1 FILLER_152_1074 ();
 FILLCELL_X1 FILLER_152_1077 ();
 FILLCELL_X8 FILLER_152_1112 ();
 FILLCELL_X1 FILLER_152_1120 ();
 FILLCELL_X8 FILLER_152_1123 ();
 FILLCELL_X4 FILLER_152_1131 ();
 FILLCELL_X2 FILLER_152_1135 ();
 FILLCELL_X1 FILLER_152_1137 ();
 FILLCELL_X1 FILLER_152_1158 ();
 FILLCELL_X4 FILLER_152_1164 ();
 FILLCELL_X2 FILLER_152_1181 ();
 FILLCELL_X1 FILLER_152_1183 ();
 FILLCELL_X32 FILLER_152_1191 ();
 FILLCELL_X32 FILLER_152_1223 ();
 FILLCELL_X4 FILLER_152_1255 ();
 FILLCELL_X1 FILLER_152_1259 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X16 FILLER_153_65 ();
 FILLCELL_X8 FILLER_153_81 ();
 FILLCELL_X4 FILLER_153_89 ();
 FILLCELL_X2 FILLER_153_93 ();
 FILLCELL_X1 FILLER_153_95 ();
 FILLCELL_X4 FILLER_153_116 ();
 FILLCELL_X2 FILLER_153_120 ();
 FILLCELL_X8 FILLER_153_142 ();
 FILLCELL_X4 FILLER_153_150 ();
 FILLCELL_X4 FILLER_153_166 ();
 FILLCELL_X1 FILLER_153_170 ();
 FILLCELL_X4 FILLER_153_178 ();
 FILLCELL_X2 FILLER_153_182 ();
 FILLCELL_X1 FILLER_153_184 ();
 FILLCELL_X2 FILLER_153_192 ();
 FILLCELL_X1 FILLER_153_194 ();
 FILLCELL_X8 FILLER_153_215 ();
 FILLCELL_X2 FILLER_153_223 ();
 FILLCELL_X1 FILLER_153_225 ();
 FILLCELL_X4 FILLER_153_240 ();
 FILLCELL_X2 FILLER_153_244 ();
 FILLCELL_X1 FILLER_153_246 ();
 FILLCELL_X8 FILLER_153_254 ();
 FILLCELL_X2 FILLER_153_296 ();
 FILLCELL_X2 FILLER_153_305 ();
 FILLCELL_X1 FILLER_153_310 ();
 FILLCELL_X2 FILLER_153_316 ();
 FILLCELL_X1 FILLER_153_318 ();
 FILLCELL_X1 FILLER_153_326 ();
 FILLCELL_X8 FILLER_153_334 ();
 FILLCELL_X4 FILLER_153_342 ();
 FILLCELL_X2 FILLER_153_346 ();
 FILLCELL_X1 FILLER_153_348 ();
 FILLCELL_X2 FILLER_153_372 ();
 FILLCELL_X2 FILLER_153_384 ();
 FILLCELL_X1 FILLER_153_386 ();
 FILLCELL_X1 FILLER_153_391 ();
 FILLCELL_X1 FILLER_153_408 ();
 FILLCELL_X16 FILLER_153_423 ();
 FILLCELL_X4 FILLER_153_439 ();
 FILLCELL_X8 FILLER_153_457 ();
 FILLCELL_X4 FILLER_153_465 ();
 FILLCELL_X1 FILLER_153_469 ();
 FILLCELL_X4 FILLER_153_477 ();
 FILLCELL_X2 FILLER_153_481 ();
 FILLCELL_X1 FILLER_153_483 ();
 FILLCELL_X16 FILLER_153_502 ();
 FILLCELL_X2 FILLER_153_518 ();
 FILLCELL_X1 FILLER_153_529 ();
 FILLCELL_X4 FILLER_153_533 ();
 FILLCELL_X2 FILLER_153_537 ();
 FILLCELL_X2 FILLER_153_543 ();
 FILLCELL_X1 FILLER_153_545 ();
 FILLCELL_X8 FILLER_153_549 ();
 FILLCELL_X2 FILLER_153_557 ();
 FILLCELL_X4 FILLER_153_563 ();
 FILLCELL_X1 FILLER_153_567 ();
 FILLCELL_X4 FILLER_153_571 ();
 FILLCELL_X4 FILLER_153_578 ();
 FILLCELL_X4 FILLER_153_586 ();
 FILLCELL_X2 FILLER_153_590 ();
 FILLCELL_X1 FILLER_153_592 ();
 FILLCELL_X2 FILLER_153_603 ();
 FILLCELL_X2 FILLER_153_612 ();
 FILLCELL_X1 FILLER_153_614 ();
 FILLCELL_X2 FILLER_153_635 ();
 FILLCELL_X1 FILLER_153_637 ();
 FILLCELL_X2 FILLER_153_645 ();
 FILLCELL_X1 FILLER_153_654 ();
 FILLCELL_X2 FILLER_153_662 ();
 FILLCELL_X1 FILLER_153_664 ();
 FILLCELL_X32 FILLER_153_687 ();
 FILLCELL_X32 FILLER_153_719 ();
 FILLCELL_X8 FILLER_153_751 ();
 FILLCELL_X4 FILLER_153_759 ();
 FILLCELL_X2 FILLER_153_763 ();
 FILLCELL_X4 FILLER_153_767 ();
 FILLCELL_X2 FILLER_153_771 ();
 FILLCELL_X8 FILLER_153_785 ();
 FILLCELL_X2 FILLER_153_793 ();
 FILLCELL_X1 FILLER_153_811 ();
 FILLCELL_X8 FILLER_153_875 ();
 FILLCELL_X4 FILLER_153_883 ();
 FILLCELL_X2 FILLER_153_966 ();
 FILLCELL_X4 FILLER_153_979 ();
 FILLCELL_X2 FILLER_153_983 ();
 FILLCELL_X1 FILLER_153_985 ();
 FILLCELL_X2 FILLER_153_989 ();
 FILLCELL_X1 FILLER_153_991 ();
 FILLCELL_X2 FILLER_153_1014 ();
 FILLCELL_X1 FILLER_153_1018 ();
 FILLCELL_X2 FILLER_153_1022 ();
 FILLCELL_X1 FILLER_153_1056 ();
 FILLCELL_X1 FILLER_153_1073 ();
 FILLCELL_X2 FILLER_153_1092 ();
 FILLCELL_X1 FILLER_153_1094 ();
 FILLCELL_X2 FILLER_153_1098 ();
 FILLCELL_X1 FILLER_153_1126 ();
 FILLCELL_X1 FILLER_153_1137 ();
 FILLCELL_X1 FILLER_153_1148 ();
 FILLCELL_X2 FILLER_153_1152 ();
 FILLCELL_X1 FILLER_153_1154 ();
 FILLCELL_X32 FILLER_153_1199 ();
 FILLCELL_X16 FILLER_153_1231 ();
 FILLCELL_X8 FILLER_153_1247 ();
 FILLCELL_X4 FILLER_153_1255 ();
 FILLCELL_X1 FILLER_153_1259 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X4 FILLER_154_97 ();
 FILLCELL_X2 FILLER_154_101 ();
 FILLCELL_X1 FILLER_154_103 ();
 FILLCELL_X32 FILLER_154_131 ();
 FILLCELL_X4 FILLER_154_203 ();
 FILLCELL_X2 FILLER_154_207 ();
 FILLCELL_X4 FILLER_154_237 ();
 FILLCELL_X1 FILLER_154_241 ();
 FILLCELL_X1 FILLER_154_269 ();
 FILLCELL_X4 FILLER_154_277 ();
 FILLCELL_X1 FILLER_154_281 ();
 FILLCELL_X16 FILLER_154_289 ();
 FILLCELL_X4 FILLER_154_309 ();
 FILLCELL_X2 FILLER_154_313 ();
 FILLCELL_X1 FILLER_154_315 ();
 FILLCELL_X1 FILLER_154_343 ();
 FILLCELL_X2 FILLER_154_351 ();
 FILLCELL_X1 FILLER_154_353 ();
 FILLCELL_X4 FILLER_154_358 ();
 FILLCELL_X2 FILLER_154_362 ();
 FILLCELL_X1 FILLER_154_364 ();
 FILLCELL_X4 FILLER_154_405 ();
 FILLCELL_X8 FILLER_154_416 ();
 FILLCELL_X8 FILLER_154_431 ();
 FILLCELL_X4 FILLER_154_439 ();
 FILLCELL_X4 FILLER_154_450 ();
 FILLCELL_X2 FILLER_154_454 ();
 FILLCELL_X1 FILLER_154_456 ();
 FILLCELL_X2 FILLER_154_532 ();
 FILLCELL_X2 FILLER_154_574 ();
 FILLCELL_X1 FILLER_154_576 ();
 FILLCELL_X2 FILLER_154_597 ();
 FILLCELL_X1 FILLER_154_599 ();
 FILLCELL_X4 FILLER_154_607 ();
 FILLCELL_X2 FILLER_154_611 ();
 FILLCELL_X8 FILLER_154_620 ();
 FILLCELL_X2 FILLER_154_628 ();
 FILLCELL_X1 FILLER_154_630 ();
 FILLCELL_X16 FILLER_154_632 ();
 FILLCELL_X4 FILLER_154_648 ();
 FILLCELL_X4 FILLER_154_666 ();
 FILLCELL_X2 FILLER_154_670 ();
 FILLCELL_X1 FILLER_154_672 ();
 FILLCELL_X8 FILLER_154_677 ();
 FILLCELL_X1 FILLER_154_685 ();
 FILLCELL_X32 FILLER_154_689 ();
 FILLCELL_X32 FILLER_154_721 ();
 FILLCELL_X8 FILLER_154_753 ();
 FILLCELL_X2 FILLER_154_761 ();
 FILLCELL_X2 FILLER_154_765 ();
 FILLCELL_X4 FILLER_154_777 ();
 FILLCELL_X2 FILLER_154_799 ();
 FILLCELL_X1 FILLER_154_801 ();
 FILLCELL_X4 FILLER_154_804 ();
 FILLCELL_X2 FILLER_154_808 ();
 FILLCELL_X4 FILLER_154_812 ();
 FILLCELL_X2 FILLER_154_816 ();
 FILLCELL_X4 FILLER_154_834 ();
 FILLCELL_X1 FILLER_154_838 ();
 FILLCELL_X1 FILLER_154_877 ();
 FILLCELL_X8 FILLER_154_884 ();
 FILLCELL_X4 FILLER_154_892 ();
 FILLCELL_X2 FILLER_154_896 ();
 FILLCELL_X2 FILLER_154_904 ();
 FILLCELL_X8 FILLER_154_909 ();
 FILLCELL_X2 FILLER_154_917 ();
 FILLCELL_X1 FILLER_154_919 ();
 FILLCELL_X1 FILLER_154_923 ();
 FILLCELL_X1 FILLER_154_929 ();
 FILLCELL_X1 FILLER_154_933 ();
 FILLCELL_X16 FILLER_154_937 ();
 FILLCELL_X1 FILLER_154_978 ();
 FILLCELL_X4 FILLER_154_995 ();
 FILLCELL_X2 FILLER_154_999 ();
 FILLCELL_X1 FILLER_154_1001 ();
 FILLCELL_X4 FILLER_154_1008 ();
 FILLCELL_X1 FILLER_154_1015 ();
 FILLCELL_X4 FILLER_154_1032 ();
 FILLCELL_X1 FILLER_154_1036 ();
 FILLCELL_X1 FILLER_154_1039 ();
 FILLCELL_X8 FILLER_154_1055 ();
 FILLCELL_X2 FILLER_154_1063 ();
 FILLCELL_X1 FILLER_154_1065 ();
 FILLCELL_X2 FILLER_154_1083 ();
 FILLCELL_X2 FILLER_154_1095 ();
 FILLCELL_X1 FILLER_154_1097 ();
 FILLCELL_X2 FILLER_154_1100 ();
 FILLCELL_X1 FILLER_154_1102 ();
 FILLCELL_X2 FILLER_154_1108 ();
 FILLCELL_X1 FILLER_154_1110 ();
 FILLCELL_X4 FILLER_154_1114 ();
 FILLCELL_X1 FILLER_154_1118 ();
 FILLCELL_X1 FILLER_154_1121 ();
 FILLCELL_X4 FILLER_154_1134 ();
 FILLCELL_X2 FILLER_154_1138 ();
 FILLCELL_X1 FILLER_154_1140 ();
 FILLCELL_X8 FILLER_154_1151 ();
 FILLCELL_X1 FILLER_154_1159 ();
 FILLCELL_X2 FILLER_154_1162 ();
 FILLCELL_X1 FILLER_154_1164 ();
 FILLCELL_X1 FILLER_154_1175 ();
 FILLCELL_X32 FILLER_154_1189 ();
 FILLCELL_X32 FILLER_154_1221 ();
 FILLCELL_X4 FILLER_154_1253 ();
 FILLCELL_X2 FILLER_154_1257 ();
 FILLCELL_X1 FILLER_154_1259 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X4 FILLER_155_161 ();
 FILLCELL_X1 FILLER_155_165 ();
 FILLCELL_X8 FILLER_155_173 ();
 FILLCELL_X4 FILLER_155_181 ();
 FILLCELL_X4 FILLER_155_212 ();
 FILLCELL_X2 FILLER_155_216 ();
 FILLCELL_X1 FILLER_155_218 ();
 FILLCELL_X8 FILLER_155_226 ();
 FILLCELL_X4 FILLER_155_234 ();
 FILLCELL_X2 FILLER_155_238 ();
 FILLCELL_X4 FILLER_155_247 ();
 FILLCELL_X1 FILLER_155_251 ();
 FILLCELL_X2 FILLER_155_271 ();
 FILLCELL_X8 FILLER_155_293 ();
 FILLCELL_X4 FILLER_155_301 ();
 FILLCELL_X8 FILLER_155_312 ();
 FILLCELL_X4 FILLER_155_320 ();
 FILLCELL_X1 FILLER_155_324 ();
 FILLCELL_X4 FILLER_155_343 ();
 FILLCELL_X2 FILLER_155_347 ();
 FILLCELL_X2 FILLER_155_353 ();
 FILLCELL_X4 FILLER_155_362 ();
 FILLCELL_X4 FILLER_155_373 ();
 FILLCELL_X2 FILLER_155_397 ();
 FILLCELL_X1 FILLER_155_399 ();
 FILLCELL_X2 FILLER_155_404 ();
 FILLCELL_X4 FILLER_155_420 ();
 FILLCELL_X4 FILLER_155_458 ();
 FILLCELL_X1 FILLER_155_462 ();
 FILLCELL_X16 FILLER_155_470 ();
 FILLCELL_X2 FILLER_155_489 ();
 FILLCELL_X2 FILLER_155_498 ();
 FILLCELL_X1 FILLER_155_507 ();
 FILLCELL_X4 FILLER_155_535 ();
 FILLCELL_X2 FILLER_155_539 ();
 FILLCELL_X1 FILLER_155_541 ();
 FILLCELL_X2 FILLER_155_546 ();
 FILLCELL_X2 FILLER_155_572 ();
 FILLCELL_X1 FILLER_155_579 ();
 FILLCELL_X2 FILLER_155_587 ();
 FILLCELL_X1 FILLER_155_589 ();
 FILLCELL_X4 FILLER_155_611 ();
 FILLCELL_X2 FILLER_155_615 ();
 FILLCELL_X2 FILLER_155_644 ();
 FILLCELL_X1 FILLER_155_646 ();
 FILLCELL_X2 FILLER_155_661 ();
 FILLCELL_X4 FILLER_155_667 ();
 FILLCELL_X2 FILLER_155_671 ();
 FILLCELL_X1 FILLER_155_680 ();
 FILLCELL_X32 FILLER_155_684 ();
 FILLCELL_X32 FILLER_155_716 ();
 FILLCELL_X16 FILLER_155_748 ();
 FILLCELL_X1 FILLER_155_764 ();
 FILLCELL_X8 FILLER_155_783 ();
 FILLCELL_X1 FILLER_155_858 ();
 FILLCELL_X1 FILLER_155_862 ();
 FILLCELL_X2 FILLER_155_870 ();
 FILLCELL_X1 FILLER_155_872 ();
 FILLCELL_X1 FILLER_155_892 ();
 FILLCELL_X1 FILLER_155_912 ();
 FILLCELL_X2 FILLER_155_916 ();
 FILLCELL_X1 FILLER_155_918 ();
 FILLCELL_X2 FILLER_155_922 ();
 FILLCELL_X1 FILLER_155_924 ();
 FILLCELL_X4 FILLER_155_964 ();
 FILLCELL_X2 FILLER_155_968 ();
 FILLCELL_X2 FILLER_155_973 ();
 FILLCELL_X1 FILLER_155_975 ();
 FILLCELL_X1 FILLER_155_979 ();
 FILLCELL_X1 FILLER_155_983 ();
 FILLCELL_X1 FILLER_155_990 ();
 FILLCELL_X1 FILLER_155_994 ();
 FILLCELL_X2 FILLER_155_1011 ();
 FILLCELL_X4 FILLER_155_1016 ();
 FILLCELL_X2 FILLER_155_1023 ();
 FILLCELL_X1 FILLER_155_1025 ();
 FILLCELL_X4 FILLER_155_1028 ();
 FILLCELL_X1 FILLER_155_1032 ();
 FILLCELL_X2 FILLER_155_1061 ();
 FILLCELL_X1 FILLER_155_1063 ();
 FILLCELL_X4 FILLER_155_1086 ();
 FILLCELL_X2 FILLER_155_1090 ();
 FILLCELL_X1 FILLER_155_1124 ();
 FILLCELL_X2 FILLER_155_1141 ();
 FILLCELL_X16 FILLER_155_1159 ();
 FILLCELL_X2 FILLER_155_1175 ();
 FILLCELL_X32 FILLER_155_1190 ();
 FILLCELL_X32 FILLER_155_1222 ();
 FILLCELL_X4 FILLER_155_1254 ();
 FILLCELL_X2 FILLER_155_1258 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X4 FILLER_156_161 ();
 FILLCELL_X2 FILLER_156_165 ();
 FILLCELL_X16 FILLER_156_187 ();
 FILLCELL_X4 FILLER_156_230 ();
 FILLCELL_X2 FILLER_156_234 ();
 FILLCELL_X4 FILLER_156_256 ();
 FILLCELL_X2 FILLER_156_267 ();
 FILLCELL_X4 FILLER_156_289 ();
 FILLCELL_X1 FILLER_156_336 ();
 FILLCELL_X8 FILLER_156_379 ();
 FILLCELL_X1 FILLER_156_434 ();
 FILLCELL_X2 FILLER_156_455 ();
 FILLCELL_X4 FILLER_156_477 ();
 FILLCELL_X2 FILLER_156_481 ();
 FILLCELL_X1 FILLER_156_483 ();
 FILLCELL_X2 FILLER_156_512 ();
 FILLCELL_X1 FILLER_156_514 ();
 FILLCELL_X16 FILLER_156_522 ();
 FILLCELL_X1 FILLER_156_558 ();
 FILLCELL_X1 FILLER_156_566 ();
 FILLCELL_X1 FILLER_156_574 ();
 FILLCELL_X2 FILLER_156_595 ();
 FILLCELL_X2 FILLER_156_604 ();
 FILLCELL_X2 FILLER_156_613 ();
 FILLCELL_X1 FILLER_156_615 ();
 FILLCELL_X2 FILLER_156_620 ();
 FILLCELL_X1 FILLER_156_622 ();
 FILLCELL_X4 FILLER_156_626 ();
 FILLCELL_X1 FILLER_156_630 ();
 FILLCELL_X4 FILLER_156_632 ();
 FILLCELL_X2 FILLER_156_636 ();
 FILLCELL_X1 FILLER_156_638 ();
 FILLCELL_X2 FILLER_156_657 ();
 FILLCELL_X1 FILLER_156_659 ();
 FILLCELL_X32 FILLER_156_700 ();
 FILLCELL_X32 FILLER_156_732 ();
 FILLCELL_X4 FILLER_156_764 ();
 FILLCELL_X2 FILLER_156_778 ();
 FILLCELL_X2 FILLER_156_782 ();
 FILLCELL_X32 FILLER_156_800 ();
 FILLCELL_X4 FILLER_156_832 ();
 FILLCELL_X4 FILLER_156_838 ();
 FILLCELL_X2 FILLER_156_842 ();
 FILLCELL_X8 FILLER_156_846 ();
 FILLCELL_X4 FILLER_156_854 ();
 FILLCELL_X2 FILLER_156_858 ();
 FILLCELL_X2 FILLER_156_871 ();
 FILLCELL_X8 FILLER_156_901 ();
 FILLCELL_X2 FILLER_156_909 ();
 FILLCELL_X4 FILLER_156_929 ();
 FILLCELL_X2 FILLER_156_933 ();
 FILLCELL_X1 FILLER_156_935 ();
 FILLCELL_X8 FILLER_156_939 ();
 FILLCELL_X2 FILLER_156_947 ();
 FILLCELL_X1 FILLER_156_949 ();
 FILLCELL_X2 FILLER_156_966 ();
 FILLCELL_X1 FILLER_156_1005 ();
 FILLCELL_X1 FILLER_156_1043 ();
 FILLCELL_X4 FILLER_156_1046 ();
 FILLCELL_X1 FILLER_156_1050 ();
 FILLCELL_X8 FILLER_156_1061 ();
 FILLCELL_X2 FILLER_156_1069 ();
 FILLCELL_X8 FILLER_156_1082 ();
 FILLCELL_X4 FILLER_156_1090 ();
 FILLCELL_X1 FILLER_156_1097 ();
 FILLCELL_X1 FILLER_156_1101 ();
 FILLCELL_X32 FILLER_156_1155 ();
 FILLCELL_X32 FILLER_156_1187 ();
 FILLCELL_X32 FILLER_156_1219 ();
 FILLCELL_X8 FILLER_156_1251 ();
 FILLCELL_X1 FILLER_156_1259 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X4 FILLER_157_161 ();
 FILLCELL_X2 FILLER_157_165 ();
 FILLCELL_X8 FILLER_157_209 ();
 FILLCELL_X4 FILLER_157_238 ();
 FILLCELL_X1 FILLER_157_242 ();
 FILLCELL_X2 FILLER_157_250 ();
 FILLCELL_X1 FILLER_157_252 ();
 FILLCELL_X16 FILLER_157_274 ();
 FILLCELL_X8 FILLER_157_290 ();
 FILLCELL_X4 FILLER_157_298 ();
 FILLCELL_X2 FILLER_157_302 ();
 FILLCELL_X4 FILLER_157_314 ();
 FILLCELL_X2 FILLER_157_318 ();
 FILLCELL_X1 FILLER_157_327 ();
 FILLCELL_X1 FILLER_157_345 ();
 FILLCELL_X2 FILLER_157_353 ();
 FILLCELL_X1 FILLER_157_385 ();
 FILLCELL_X2 FILLER_157_390 ();
 FILLCELL_X1 FILLER_157_392 ();
 FILLCELL_X4 FILLER_157_396 ();
 FILLCELL_X2 FILLER_157_400 ();
 FILLCELL_X8 FILLER_157_405 ();
 FILLCELL_X4 FILLER_157_413 ();
 FILLCELL_X8 FILLER_157_431 ();
 FILLCELL_X4 FILLER_157_439 ();
 FILLCELL_X1 FILLER_157_443 ();
 FILLCELL_X4 FILLER_157_455 ();
 FILLCELL_X1 FILLER_157_459 ();
 FILLCELL_X4 FILLER_157_463 ();
 FILLCELL_X1 FILLER_157_467 ();
 FILLCELL_X2 FILLER_157_475 ();
 FILLCELL_X1 FILLER_157_477 ();
 FILLCELL_X1 FILLER_157_485 ();
 FILLCELL_X8 FILLER_157_500 ();
 FILLCELL_X4 FILLER_157_508 ();
 FILLCELL_X2 FILLER_157_519 ();
 FILLCELL_X1 FILLER_157_521 ();
 FILLCELL_X8 FILLER_157_549 ();
 FILLCELL_X2 FILLER_157_557 ();
 FILLCELL_X2 FILLER_157_573 ();
 FILLCELL_X1 FILLER_157_575 ();
 FILLCELL_X8 FILLER_157_583 ();
 FILLCELL_X2 FILLER_157_591 ();
 FILLCELL_X1 FILLER_157_593 ();
 FILLCELL_X2 FILLER_157_608 ();
 FILLCELL_X1 FILLER_157_610 ();
 FILLCELL_X4 FILLER_157_631 ();
 FILLCELL_X1 FILLER_157_635 ();
 FILLCELL_X32 FILLER_157_663 ();
 FILLCELL_X32 FILLER_157_695 ();
 FILLCELL_X32 FILLER_157_727 ();
 FILLCELL_X8 FILLER_157_759 ();
 FILLCELL_X4 FILLER_157_767 ();
 FILLCELL_X1 FILLER_157_771 ();
 FILLCELL_X16 FILLER_157_794 ();
 FILLCELL_X4 FILLER_157_810 ();
 FILLCELL_X4 FILLER_157_878 ();
 FILLCELL_X2 FILLER_157_882 ();
 FILLCELL_X8 FILLER_157_900 ();
 FILLCELL_X2 FILLER_157_908 ();
 FILLCELL_X1 FILLER_157_910 ();
 FILLCELL_X8 FILLER_157_913 ();
 FILLCELL_X4 FILLER_157_921 ();
 FILLCELL_X2 FILLER_157_925 ();
 FILLCELL_X1 FILLER_157_927 ();
 FILLCELL_X16 FILLER_157_944 ();
 FILLCELL_X2 FILLER_157_960 ();
 FILLCELL_X1 FILLER_157_964 ();
 FILLCELL_X1 FILLER_157_981 ();
 FILLCELL_X2 FILLER_157_998 ();
 FILLCELL_X2 FILLER_157_1003 ();
 FILLCELL_X2 FILLER_157_1021 ();
 FILLCELL_X4 FILLER_157_1026 ();
 FILLCELL_X2 FILLER_157_1030 ();
 FILLCELL_X1 FILLER_157_1032 ();
 FILLCELL_X2 FILLER_157_1038 ();
 FILLCELL_X1 FILLER_157_1040 ();
 FILLCELL_X2 FILLER_157_1051 ();
 FILLCELL_X1 FILLER_157_1053 ();
 FILLCELL_X4 FILLER_157_1064 ();
 FILLCELL_X8 FILLER_157_1103 ();
 FILLCELL_X1 FILLER_157_1111 ();
 FILLCELL_X4 FILLER_157_1118 ();
 FILLCELL_X2 FILLER_157_1122 ();
 FILLCELL_X1 FILLER_157_1142 ();
 FILLCELL_X16 FILLER_157_1147 ();
 FILLCELL_X2 FILLER_157_1163 ();
 FILLCELL_X1 FILLER_157_1165 ();
 FILLCELL_X32 FILLER_157_1168 ();
 FILLCELL_X32 FILLER_157_1200 ();
 FILLCELL_X16 FILLER_157_1232 ();
 FILLCELL_X8 FILLER_157_1248 ();
 FILLCELL_X4 FILLER_157_1256 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X8 FILLER_158_193 ();
 FILLCELL_X1 FILLER_158_201 ();
 FILLCELL_X4 FILLER_158_209 ();
 FILLCELL_X1 FILLER_158_213 ();
 FILLCELL_X1 FILLER_158_268 ();
 FILLCELL_X2 FILLER_158_289 ();
 FILLCELL_X1 FILLER_158_291 ();
 FILLCELL_X1 FILLER_158_312 ();
 FILLCELL_X16 FILLER_158_340 ();
 FILLCELL_X8 FILLER_158_356 ();
 FILLCELL_X2 FILLER_158_364 ();
 FILLCELL_X8 FILLER_158_373 ();
 FILLCELL_X2 FILLER_158_381 ();
 FILLCELL_X1 FILLER_158_383 ();
 FILLCELL_X1 FILLER_158_388 ();
 FILLCELL_X8 FILLER_158_392 ();
 FILLCELL_X2 FILLER_158_400 ();
 FILLCELL_X4 FILLER_158_443 ();
 FILLCELL_X1 FILLER_158_447 ();
 FILLCELL_X16 FILLER_158_468 ();
 FILLCELL_X4 FILLER_158_484 ();
 FILLCELL_X4 FILLER_158_491 ();
 FILLCELL_X1 FILLER_158_495 ();
 FILLCELL_X8 FILLER_158_503 ();
 FILLCELL_X1 FILLER_158_511 ();
 FILLCELL_X2 FILLER_158_519 ();
 FILLCELL_X1 FILLER_158_521 ();
 FILLCELL_X4 FILLER_158_529 ();
 FILLCELL_X2 FILLER_158_533 ();
 FILLCELL_X2 FILLER_158_542 ();
 FILLCELL_X1 FILLER_158_544 ();
 FILLCELL_X2 FILLER_158_552 ();
 FILLCELL_X1 FILLER_158_554 ();
 FILLCELL_X1 FILLER_158_565 ();
 FILLCELL_X4 FILLER_158_573 ();
 FILLCELL_X1 FILLER_158_577 ();
 FILLCELL_X1 FILLER_158_585 ();
 FILLCELL_X2 FILLER_158_599 ();
 FILLCELL_X8 FILLER_158_608 ();
 FILLCELL_X1 FILLER_158_616 ();
 FILLCELL_X32 FILLER_158_657 ();
 FILLCELL_X32 FILLER_158_689 ();
 FILLCELL_X32 FILLER_158_721 ();
 FILLCELL_X16 FILLER_158_753 ();
 FILLCELL_X2 FILLER_158_769 ();
 FILLCELL_X2 FILLER_158_781 ();
 FILLCELL_X1 FILLER_158_783 ();
 FILLCELL_X16 FILLER_158_828 ();
 FILLCELL_X8 FILLER_158_844 ();
 FILLCELL_X4 FILLER_158_860 ();
 FILLCELL_X4 FILLER_158_885 ();
 FILLCELL_X4 FILLER_158_892 ();
 FILLCELL_X1 FILLER_158_896 ();
 FILLCELL_X8 FILLER_158_900 ();
 FILLCELL_X4 FILLER_158_908 ();
 FILLCELL_X2 FILLER_158_912 ();
 FILLCELL_X1 FILLER_158_914 ();
 FILLCELL_X4 FILLER_158_979 ();
 FILLCELL_X2 FILLER_158_983 ();
 FILLCELL_X1 FILLER_158_985 ();
 FILLCELL_X2 FILLER_158_988 ();
 FILLCELL_X1 FILLER_158_990 ();
 FILLCELL_X8 FILLER_158_1009 ();
 FILLCELL_X4 FILLER_158_1017 ();
 FILLCELL_X2 FILLER_158_1021 ();
 FILLCELL_X1 FILLER_158_1023 ();
 FILLCELL_X4 FILLER_158_1026 ();
 FILLCELL_X2 FILLER_158_1030 ();
 FILLCELL_X1 FILLER_158_1032 ();
 FILLCELL_X2 FILLER_158_1051 ();
 FILLCELL_X8 FILLER_158_1059 ();
 FILLCELL_X1 FILLER_158_1067 ();
 FILLCELL_X4 FILLER_158_1103 ();
 FILLCELL_X2 FILLER_158_1107 ();
 FILLCELL_X1 FILLER_158_1115 ();
 FILLCELL_X8 FILLER_158_1125 ();
 FILLCELL_X2 FILLER_158_1133 ();
 FILLCELL_X1 FILLER_158_1135 ();
 FILLCELL_X8 FILLER_158_1138 ();
 FILLCELL_X1 FILLER_158_1146 ();
 FILLCELL_X32 FILLER_158_1163 ();
 FILLCELL_X32 FILLER_158_1195 ();
 FILLCELL_X32 FILLER_158_1227 ();
 FILLCELL_X1 FILLER_158_1259 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X8 FILLER_159_193 ();
 FILLCELL_X2 FILLER_159_201 ();
 FILLCELL_X16 FILLER_159_223 ();
 FILLCELL_X8 FILLER_159_239 ();
 FILLCELL_X4 FILLER_159_247 ();
 FILLCELL_X8 FILLER_159_258 ();
 FILLCELL_X2 FILLER_159_266 ();
 FILLCELL_X8 FILLER_159_275 ();
 FILLCELL_X4 FILLER_159_283 ();
 FILLCELL_X1 FILLER_159_287 ();
 FILLCELL_X4 FILLER_159_318 ();
 FILLCELL_X2 FILLER_159_322 ();
 FILLCELL_X1 FILLER_159_331 ();
 FILLCELL_X1 FILLER_159_342 ();
 FILLCELL_X1 FILLER_159_350 ();
 FILLCELL_X1 FILLER_159_355 ();
 FILLCELL_X1 FILLER_159_399 ();
 FILLCELL_X4 FILLER_159_414 ();
 FILLCELL_X2 FILLER_159_418 ();
 FILLCELL_X1 FILLER_159_420 ();
 FILLCELL_X8 FILLER_159_449 ();
 FILLCELL_X4 FILLER_159_457 ();
 FILLCELL_X2 FILLER_159_461 ();
 FILLCELL_X1 FILLER_159_463 ();
 FILLCELL_X2 FILLER_159_518 ();
 FILLCELL_X1 FILLER_159_543 ();
 FILLCELL_X4 FILLER_159_576 ();
 FILLCELL_X1 FILLER_159_600 ();
 FILLCELL_X2 FILLER_159_618 ();
 FILLCELL_X1 FILLER_159_620 ();
 FILLCELL_X4 FILLER_159_628 ();
 FILLCELL_X2 FILLER_159_639 ();
 FILLCELL_X1 FILLER_159_641 ();
 FILLCELL_X1 FILLER_159_649 ();
 FILLCELL_X32 FILLER_159_670 ();
 FILLCELL_X32 FILLER_159_702 ();
 FILLCELL_X32 FILLER_159_734 ();
 FILLCELL_X8 FILLER_159_766 ();
 FILLCELL_X1 FILLER_159_780 ();
 FILLCELL_X4 FILLER_159_789 ();
 FILLCELL_X2 FILLER_159_793 ();
 FILLCELL_X1 FILLER_159_795 ();
 FILLCELL_X8 FILLER_159_798 ();
 FILLCELL_X4 FILLER_159_806 ();
 FILLCELL_X2 FILLER_159_810 ();
 FILLCELL_X1 FILLER_159_812 ();
 FILLCELL_X8 FILLER_159_831 ();
 FILLCELL_X1 FILLER_159_839 ();
 FILLCELL_X2 FILLER_159_846 ();
 FILLCELL_X1 FILLER_159_848 ();
 FILLCELL_X8 FILLER_159_852 ();
 FILLCELL_X1 FILLER_159_863 ();
 FILLCELL_X4 FILLER_159_868 ();
 FILLCELL_X2 FILLER_159_872 ();
 FILLCELL_X1 FILLER_159_922 ();
 FILLCELL_X1 FILLER_159_926 ();
 FILLCELL_X8 FILLER_159_945 ();
 FILLCELL_X2 FILLER_159_953 ();
 FILLCELL_X16 FILLER_159_971 ();
 FILLCELL_X1 FILLER_159_987 ();
 FILLCELL_X16 FILLER_159_993 ();
 FILLCELL_X8 FILLER_159_1009 ();
 FILLCELL_X1 FILLER_159_1017 ();
 FILLCELL_X2 FILLER_159_1021 ();
 FILLCELL_X2 FILLER_159_1101 ();
 FILLCELL_X4 FILLER_159_1135 ();
 FILLCELL_X32 FILLER_159_1155 ();
 FILLCELL_X32 FILLER_159_1187 ();
 FILLCELL_X32 FILLER_159_1219 ();
 FILLCELL_X8 FILLER_159_1251 ();
 FILLCELL_X1 FILLER_159_1259 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X16 FILLER_160_289 ();
 FILLCELL_X4 FILLER_160_305 ();
 FILLCELL_X2 FILLER_160_309 ();
 FILLCELL_X4 FILLER_160_363 ();
 FILLCELL_X2 FILLER_160_367 ();
 FILLCELL_X1 FILLER_160_369 ();
 FILLCELL_X4 FILLER_160_374 ();
 FILLCELL_X8 FILLER_160_381 ();
 FILLCELL_X2 FILLER_160_389 ();
 FILLCELL_X1 FILLER_160_395 ();
 FILLCELL_X4 FILLER_160_406 ();
 FILLCELL_X1 FILLER_160_417 ();
 FILLCELL_X2 FILLER_160_430 ();
 FILLCELL_X4 FILLER_160_439 ();
 FILLCELL_X1 FILLER_160_447 ();
 FILLCELL_X4 FILLER_160_451 ();
 FILLCELL_X2 FILLER_160_455 ();
 FILLCELL_X1 FILLER_160_457 ();
 FILLCELL_X2 FILLER_160_479 ();
 FILLCELL_X2 FILLER_160_508 ();
 FILLCELL_X2 FILLER_160_524 ();
 FILLCELL_X1 FILLER_160_526 ();
 FILLCELL_X8 FILLER_160_531 ();
 FILLCELL_X2 FILLER_160_539 ();
 FILLCELL_X1 FILLER_160_541 ();
 FILLCELL_X8 FILLER_160_596 ();
 FILLCELL_X4 FILLER_160_624 ();
 FILLCELL_X2 FILLER_160_628 ();
 FILLCELL_X1 FILLER_160_630 ();
 FILLCELL_X4 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_656 ();
 FILLCELL_X32 FILLER_160_688 ();
 FILLCELL_X32 FILLER_160_720 ();
 FILLCELL_X8 FILLER_160_752 ();
 FILLCELL_X4 FILLER_160_760 ();
 FILLCELL_X2 FILLER_160_764 ();
 FILLCELL_X1 FILLER_160_766 ();
 FILLCELL_X1 FILLER_160_789 ();
 FILLCELL_X2 FILLER_160_808 ();
 FILLCELL_X1 FILLER_160_812 ();
 FILLCELL_X4 FILLER_160_831 ();
 FILLCELL_X2 FILLER_160_851 ();
 FILLCELL_X2 FILLER_160_891 ();
 FILLCELL_X2 FILLER_160_895 ();
 FILLCELL_X1 FILLER_160_897 ();
 FILLCELL_X16 FILLER_160_925 ();
 FILLCELL_X2 FILLER_160_941 ();
 FILLCELL_X2 FILLER_160_946 ();
 FILLCELL_X1 FILLER_160_964 ();
 FILLCELL_X8 FILLER_160_989 ();
 FILLCELL_X1 FILLER_160_1015 ();
 FILLCELL_X16 FILLER_160_1048 ();
 FILLCELL_X4 FILLER_160_1064 ();
 FILLCELL_X2 FILLER_160_1116 ();
 FILLCELL_X1 FILLER_160_1118 ();
 FILLCELL_X32 FILLER_160_1140 ();
 FILLCELL_X32 FILLER_160_1172 ();
 FILLCELL_X32 FILLER_160_1204 ();
 FILLCELL_X16 FILLER_160_1236 ();
 FILLCELL_X8 FILLER_160_1252 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X8 FILLER_161_289 ();
 FILLCELL_X1 FILLER_161_297 ();
 FILLCELL_X4 FILLER_161_350 ();
 FILLCELL_X4 FILLER_161_361 ();
 FILLCELL_X1 FILLER_161_365 ();
 FILLCELL_X2 FILLER_161_406 ();
 FILLCELL_X1 FILLER_161_408 ();
 FILLCELL_X2 FILLER_161_416 ();
 FILLCELL_X1 FILLER_161_418 ();
 FILLCELL_X16 FILLER_161_478 ();
 FILLCELL_X4 FILLER_161_494 ();
 FILLCELL_X2 FILLER_161_498 ();
 FILLCELL_X1 FILLER_161_500 ();
 FILLCELL_X2 FILLER_161_519 ();
 FILLCELL_X1 FILLER_161_521 ();
 FILLCELL_X2 FILLER_161_526 ();
 FILLCELL_X1 FILLER_161_528 ();
 FILLCELL_X4 FILLER_161_532 ();
 FILLCELL_X1 FILLER_161_536 ();
 FILLCELL_X1 FILLER_161_548 ();
 FILLCELL_X16 FILLER_161_555 ();
 FILLCELL_X4 FILLER_161_571 ();
 FILLCELL_X8 FILLER_161_582 ();
 FILLCELL_X4 FILLER_161_590 ();
 FILLCELL_X2 FILLER_161_601 ();
 FILLCELL_X4 FILLER_161_633 ();
 FILLCELL_X2 FILLER_161_637 ();
 FILLCELL_X1 FILLER_161_639 ();
 FILLCELL_X2 FILLER_161_644 ();
 FILLCELL_X1 FILLER_161_646 ();
 FILLCELL_X32 FILLER_161_650 ();
 FILLCELL_X32 FILLER_161_682 ();
 FILLCELL_X32 FILLER_161_714 ();
 FILLCELL_X16 FILLER_161_746 ();
 FILLCELL_X8 FILLER_161_762 ();
 FILLCELL_X2 FILLER_161_770 ();
 FILLCELL_X1 FILLER_161_772 ();
 FILLCELL_X2 FILLER_161_779 ();
 FILLCELL_X1 FILLER_161_787 ();
 FILLCELL_X1 FILLER_161_796 ();
 FILLCELL_X4 FILLER_161_813 ();
 FILLCELL_X2 FILLER_161_819 ();
 FILLCELL_X1 FILLER_161_821 ();
 FILLCELL_X1 FILLER_161_824 ();
 FILLCELL_X1 FILLER_161_827 ();
 FILLCELL_X1 FILLER_161_830 ();
 FILLCELL_X1 FILLER_161_833 ();
 FILLCELL_X1 FILLER_161_840 ();
 FILLCELL_X4 FILLER_161_857 ();
 FILLCELL_X1 FILLER_161_861 ();
 FILLCELL_X8 FILLER_161_866 ();
 FILLCELL_X4 FILLER_161_874 ();
 FILLCELL_X1 FILLER_161_878 ();
 FILLCELL_X8 FILLER_161_882 ();
 FILLCELL_X2 FILLER_161_890 ();
 FILLCELL_X1 FILLER_161_892 ();
 FILLCELL_X2 FILLER_161_909 ();
 FILLCELL_X2 FILLER_161_917 ();
 FILLCELL_X2 FILLER_161_956 ();
 FILLCELL_X1 FILLER_161_1009 ();
 FILLCELL_X8 FILLER_161_1026 ();
 FILLCELL_X1 FILLER_161_1034 ();
 FILLCELL_X8 FILLER_161_1054 ();
 FILLCELL_X1 FILLER_161_1071 ();
 FILLCELL_X2 FILLER_161_1091 ();
 FILLCELL_X2 FILLER_161_1098 ();
 FILLCELL_X1 FILLER_161_1100 ();
 FILLCELL_X2 FILLER_161_1113 ();
 FILLCELL_X1 FILLER_161_1131 ();
 FILLCELL_X32 FILLER_161_1155 ();
 FILLCELL_X32 FILLER_161_1187 ();
 FILLCELL_X32 FILLER_161_1219 ();
 FILLCELL_X8 FILLER_161_1251 ();
 FILLCELL_X1 FILLER_161_1259 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X16 FILLER_162_257 ();
 FILLCELL_X8 FILLER_162_273 ();
 FILLCELL_X2 FILLER_162_281 ();
 FILLCELL_X8 FILLER_162_326 ();
 FILLCELL_X2 FILLER_162_334 ();
 FILLCELL_X1 FILLER_162_336 ();
 FILLCELL_X4 FILLER_162_347 ();
 FILLCELL_X2 FILLER_162_365 ();
 FILLCELL_X1 FILLER_162_367 ();
 FILLCELL_X16 FILLER_162_375 ();
 FILLCELL_X8 FILLER_162_391 ();
 FILLCELL_X4 FILLER_162_406 ();
 FILLCELL_X8 FILLER_162_417 ();
 FILLCELL_X4 FILLER_162_425 ();
 FILLCELL_X2 FILLER_162_429 ();
 FILLCELL_X1 FILLER_162_431 ();
 FILLCELL_X4 FILLER_162_445 ();
 FILLCELL_X2 FILLER_162_449 ();
 FILLCELL_X2 FILLER_162_455 ();
 FILLCELL_X1 FILLER_162_457 ();
 FILLCELL_X4 FILLER_162_465 ();
 FILLCELL_X2 FILLER_162_469 ();
 FILLCELL_X2 FILLER_162_514 ();
 FILLCELL_X1 FILLER_162_516 ();
 FILLCELL_X1 FILLER_162_557 ();
 FILLCELL_X8 FILLER_162_578 ();
 FILLCELL_X2 FILLER_162_586 ();
 FILLCELL_X16 FILLER_162_608 ();
 FILLCELL_X4 FILLER_162_624 ();
 FILLCELL_X2 FILLER_162_628 ();
 FILLCELL_X1 FILLER_162_630 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X4 FILLER_162_760 ();
 FILLCELL_X2 FILLER_162_764 ();
 FILLCELL_X1 FILLER_162_766 ();
 FILLCELL_X2 FILLER_162_783 ();
 FILLCELL_X2 FILLER_162_803 ();
 FILLCELL_X1 FILLER_162_805 ();
 FILLCELL_X16 FILLER_162_856 ();
 FILLCELL_X4 FILLER_162_872 ();
 FILLCELL_X2 FILLER_162_892 ();
 FILLCELL_X1 FILLER_162_894 ();
 FILLCELL_X4 FILLER_162_897 ();
 FILLCELL_X1 FILLER_162_901 ();
 FILLCELL_X4 FILLER_162_904 ();
 FILLCELL_X2 FILLER_162_908 ();
 FILLCELL_X2 FILLER_162_912 ();
 FILLCELL_X2 FILLER_162_933 ();
 FILLCELL_X1 FILLER_162_935 ();
 FILLCELL_X4 FILLER_162_941 ();
 FILLCELL_X8 FILLER_162_948 ();
 FILLCELL_X4 FILLER_162_960 ();
 FILLCELL_X1 FILLER_162_964 ();
 FILLCELL_X4 FILLER_162_971 ();
 FILLCELL_X4 FILLER_162_977 ();
 FILLCELL_X2 FILLER_162_981 ();
 FILLCELL_X1 FILLER_162_983 ();
 FILLCELL_X4 FILLER_162_987 ();
 FILLCELL_X2 FILLER_162_991 ();
 FILLCELL_X4 FILLER_162_1001 ();
 FILLCELL_X2 FILLER_162_1008 ();
 FILLCELL_X2 FILLER_162_1013 ();
 FILLCELL_X1 FILLER_162_1015 ();
 FILLCELL_X1 FILLER_162_1019 ();
 FILLCELL_X16 FILLER_162_1032 ();
 FILLCELL_X4 FILLER_162_1048 ();
 FILLCELL_X2 FILLER_162_1052 ();
 FILLCELL_X1 FILLER_162_1054 ();
 FILLCELL_X4 FILLER_162_1118 ();
 FILLCELL_X2 FILLER_162_1122 ();
 FILLCELL_X1 FILLER_162_1124 ();
 FILLCELL_X1 FILLER_162_1127 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X16 FILLER_162_1240 ();
 FILLCELL_X4 FILLER_162_1256 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X8 FILLER_163_289 ();
 FILLCELL_X4 FILLER_163_297 ();
 FILLCELL_X2 FILLER_163_301 ();
 FILLCELL_X4 FILLER_163_313 ();
 FILLCELL_X1 FILLER_163_317 ();
 FILLCELL_X1 FILLER_163_332 ();
 FILLCELL_X1 FILLER_163_368 ();
 FILLCELL_X4 FILLER_163_376 ();
 FILLCELL_X4 FILLER_163_387 ();
 FILLCELL_X2 FILLER_163_395 ();
 FILLCELL_X1 FILLER_163_400 ();
 FILLCELL_X4 FILLER_163_422 ();
 FILLCELL_X2 FILLER_163_470 ();
 FILLCELL_X4 FILLER_163_475 ();
 FILLCELL_X2 FILLER_163_479 ();
 FILLCELL_X2 FILLER_163_488 ();
 FILLCELL_X2 FILLER_163_499 ();
 FILLCELL_X1 FILLER_163_501 ();
 FILLCELL_X4 FILLER_163_520 ();
 FILLCELL_X2 FILLER_163_524 ();
 FILLCELL_X1 FILLER_163_526 ();
 FILLCELL_X8 FILLER_163_534 ();
 FILLCELL_X2 FILLER_163_542 ();
 FILLCELL_X1 FILLER_163_544 ();
 FILLCELL_X1 FILLER_163_572 ();
 FILLCELL_X1 FILLER_163_594 ();
 FILLCELL_X32 FILLER_163_598 ();
 FILLCELL_X32 FILLER_163_630 ();
 FILLCELL_X32 FILLER_163_662 ();
 FILLCELL_X32 FILLER_163_694 ();
 FILLCELL_X32 FILLER_163_726 ();
 FILLCELL_X32 FILLER_163_758 ();
 FILLCELL_X2 FILLER_163_790 ();
 FILLCELL_X32 FILLER_163_798 ();
 FILLCELL_X8 FILLER_163_830 ();
 FILLCELL_X4 FILLER_163_838 ();
 FILLCELL_X1 FILLER_163_842 ();
 FILLCELL_X32 FILLER_163_845 ();
 FILLCELL_X4 FILLER_163_877 ();
 FILLCELL_X2 FILLER_163_881 ();
 FILLCELL_X1 FILLER_163_883 ();
 FILLCELL_X1 FILLER_163_900 ();
 FILLCELL_X1 FILLER_163_903 ();
 FILLCELL_X1 FILLER_163_920 ();
 FILLCELL_X1 FILLER_163_923 ();
 FILLCELL_X8 FILLER_163_930 ();
 FILLCELL_X2 FILLER_163_938 ();
 FILLCELL_X1 FILLER_163_940 ();
 FILLCELL_X2 FILLER_163_944 ();
 FILLCELL_X2 FILLER_163_949 ();
 FILLCELL_X2 FILLER_163_954 ();
 FILLCELL_X1 FILLER_163_965 ();
 FILLCELL_X8 FILLER_163_1069 ();
 FILLCELL_X4 FILLER_163_1077 ();
 FILLCELL_X2 FILLER_163_1081 ();
 FILLCELL_X1 FILLER_163_1103 ();
 FILLCELL_X8 FILLER_163_1106 ();
 FILLCELL_X4 FILLER_163_1114 ();
 FILLCELL_X8 FILLER_163_1120 ();
 FILLCELL_X4 FILLER_163_1128 ();
 FILLCELL_X2 FILLER_163_1132 ();
 FILLCELL_X32 FILLER_163_1146 ();
 FILLCELL_X32 FILLER_163_1178 ();
 FILLCELL_X32 FILLER_163_1210 ();
 FILLCELL_X16 FILLER_163_1242 ();
 FILLCELL_X2 FILLER_163_1258 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X1 FILLER_164_289 ();
 FILLCELL_X2 FILLER_164_310 ();
 FILLCELL_X1 FILLER_164_326 ();
 FILLCELL_X2 FILLER_164_352 ();
 FILLCELL_X4 FILLER_164_382 ();
 FILLCELL_X8 FILLER_164_413 ();
 FILLCELL_X4 FILLER_164_441 ();
 FILLCELL_X2 FILLER_164_445 ();
 FILLCELL_X1 FILLER_164_447 ();
 FILLCELL_X8 FILLER_164_536 ();
 FILLCELL_X4 FILLER_164_544 ();
 FILLCELL_X4 FILLER_164_578 ();
 FILLCELL_X1 FILLER_164_582 ();
 FILLCELL_X16 FILLER_164_603 ();
 FILLCELL_X8 FILLER_164_619 ();
 FILLCELL_X4 FILLER_164_627 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X16 FILLER_164_856 ();
 FILLCELL_X8 FILLER_164_872 ();
 FILLCELL_X4 FILLER_164_880 ();
 FILLCELL_X2 FILLER_164_884 ();
 FILLCELL_X1 FILLER_164_886 ();
 FILLCELL_X8 FILLER_164_967 ();
 FILLCELL_X2 FILLER_164_975 ();
 FILLCELL_X1 FILLER_164_977 ();
 FILLCELL_X1 FILLER_164_994 ();
 FILLCELL_X8 FILLER_164_998 ();
 FILLCELL_X4 FILLER_164_1006 ();
 FILLCELL_X2 FILLER_164_1026 ();
 FILLCELL_X1 FILLER_164_1028 ();
 FILLCELL_X2 FILLER_164_1047 ();
 FILLCELL_X4 FILLER_164_1051 ();
 FILLCELL_X2 FILLER_164_1055 ();
 FILLCELL_X1 FILLER_164_1057 ();
 FILLCELL_X1 FILLER_164_1074 ();
 FILLCELL_X1 FILLER_164_1077 ();
 FILLCELL_X2 FILLER_164_1094 ();
 FILLCELL_X16 FILLER_164_1098 ();
 FILLCELL_X1 FILLER_164_1114 ();
 FILLCELL_X4 FILLER_164_1131 ();
 FILLCELL_X1 FILLER_164_1135 ();
 FILLCELL_X32 FILLER_164_1138 ();
 FILLCELL_X32 FILLER_164_1170 ();
 FILLCELL_X32 FILLER_164_1202 ();
 FILLCELL_X16 FILLER_164_1234 ();
 FILLCELL_X8 FILLER_164_1250 ();
 FILLCELL_X2 FILLER_164_1258 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X8 FILLER_165_289 ();
 FILLCELL_X4 FILLER_165_297 ();
 FILLCELL_X2 FILLER_165_301 ();
 FILLCELL_X1 FILLER_165_303 ();
 FILLCELL_X4 FILLER_165_331 ();
 FILLCELL_X1 FILLER_165_335 ();
 FILLCELL_X2 FILLER_165_340 ();
 FILLCELL_X2 FILLER_165_345 ();
 FILLCELL_X2 FILLER_165_370 ();
 FILLCELL_X8 FILLER_165_379 ();
 FILLCELL_X2 FILLER_165_387 ();
 FILLCELL_X2 FILLER_165_397 ();
 FILLCELL_X1 FILLER_165_403 ();
 FILLCELL_X1 FILLER_165_407 ();
 FILLCELL_X8 FILLER_165_415 ();
 FILLCELL_X1 FILLER_165_437 ();
 FILLCELL_X4 FILLER_165_445 ();
 FILLCELL_X8 FILLER_165_454 ();
 FILLCELL_X2 FILLER_165_462 ();
 FILLCELL_X1 FILLER_165_464 ();
 FILLCELL_X16 FILLER_165_469 ();
 FILLCELL_X8 FILLER_165_485 ();
 FILLCELL_X2 FILLER_165_493 ();
 FILLCELL_X1 FILLER_165_495 ();
 FILLCELL_X32 FILLER_165_506 ();
 FILLCELL_X8 FILLER_165_538 ();
 FILLCELL_X4 FILLER_165_546 ();
 FILLCELL_X2 FILLER_165_550 ();
 FILLCELL_X1 FILLER_165_552 ();
 FILLCELL_X16 FILLER_165_556 ();
 FILLCELL_X1 FILLER_165_572 ();
 FILLCELL_X32 FILLER_165_580 ();
 FILLCELL_X32 FILLER_165_612 ();
 FILLCELL_X32 FILLER_165_644 ();
 FILLCELL_X32 FILLER_165_676 ();
 FILLCELL_X32 FILLER_165_708 ();
 FILLCELL_X32 FILLER_165_740 ();
 FILLCELL_X32 FILLER_165_772 ();
 FILLCELL_X32 FILLER_165_804 ();
 FILLCELL_X32 FILLER_165_836 ();
 FILLCELL_X32 FILLER_165_868 ();
 FILLCELL_X8 FILLER_165_900 ();
 FILLCELL_X4 FILLER_165_910 ();
 FILLCELL_X4 FILLER_165_918 ();
 FILLCELL_X2 FILLER_165_922 ();
 FILLCELL_X8 FILLER_165_958 ();
 FILLCELL_X2 FILLER_165_966 ();
 FILLCELL_X1 FILLER_165_968 ();
 FILLCELL_X4 FILLER_165_985 ();
 FILLCELL_X8 FILLER_165_1005 ();
 FILLCELL_X2 FILLER_165_1013 ();
 FILLCELL_X1 FILLER_165_1015 ();
 FILLCELL_X2 FILLER_165_1026 ();
 FILLCELL_X4 FILLER_165_1030 ();
 FILLCELL_X2 FILLER_165_1034 ();
 FILLCELL_X1 FILLER_165_1036 ();
 FILLCELL_X2 FILLER_165_1071 ();
 FILLCELL_X4 FILLER_165_1091 ();
 FILLCELL_X2 FILLER_165_1095 ();
 FILLCELL_X16 FILLER_165_1115 ();
 FILLCELL_X32 FILLER_165_1147 ();
 FILLCELL_X32 FILLER_165_1179 ();
 FILLCELL_X32 FILLER_165_1211 ();
 FILLCELL_X16 FILLER_165_1243 ();
 FILLCELL_X1 FILLER_165_1259 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X8 FILLER_166_321 ();
 FILLCELL_X2 FILLER_166_329 ();
 FILLCELL_X2 FILLER_166_351 ();
 FILLCELL_X4 FILLER_166_381 ();
 FILLCELL_X2 FILLER_166_385 ();
 FILLCELL_X2 FILLER_166_415 ();
 FILLCELL_X8 FILLER_166_420 ();
 FILLCELL_X2 FILLER_166_428 ();
 FILLCELL_X2 FILLER_166_450 ();
 FILLCELL_X32 FILLER_166_475 ();
 FILLCELL_X32 FILLER_166_507 ();
 FILLCELL_X32 FILLER_166_539 ();
 FILLCELL_X32 FILLER_166_571 ();
 FILLCELL_X16 FILLER_166_603 ();
 FILLCELL_X8 FILLER_166_619 ();
 FILLCELL_X4 FILLER_166_627 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X8 FILLER_166_920 ();
 FILLCELL_X4 FILLER_166_928 ();
 FILLCELL_X1 FILLER_166_932 ();
 FILLCELL_X1 FILLER_166_981 ();
 FILLCELL_X2 FILLER_166_998 ();
 FILLCELL_X2 FILLER_166_1016 ();
 FILLCELL_X16 FILLER_166_1034 ();
 FILLCELL_X8 FILLER_166_1050 ();
 FILLCELL_X2 FILLER_166_1058 ();
 FILLCELL_X4 FILLER_166_1076 ();
 FILLCELL_X2 FILLER_166_1080 ();
 FILLCELL_X2 FILLER_166_1100 ();
 FILLCELL_X1 FILLER_166_1102 ();
 FILLCELL_X1 FILLER_166_1105 ();
 FILLCELL_X2 FILLER_166_1122 ();
 FILLCELL_X1 FILLER_166_1128 ();
 FILLCELL_X2 FILLER_166_1133 ();
 FILLCELL_X32 FILLER_166_1147 ();
 FILLCELL_X32 FILLER_166_1179 ();
 FILLCELL_X32 FILLER_166_1211 ();
 FILLCELL_X16 FILLER_166_1243 ();
 FILLCELL_X1 FILLER_166_1259 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X16 FILLER_167_353 ();
 FILLCELL_X4 FILLER_167_369 ();
 FILLCELL_X1 FILLER_167_373 ();
 FILLCELL_X2 FILLER_167_437 ();
 FILLCELL_X1 FILLER_167_439 ();
 FILLCELL_X32 FILLER_167_443 ();
 FILLCELL_X32 FILLER_167_475 ();
 FILLCELL_X32 FILLER_167_507 ();
 FILLCELL_X32 FILLER_167_539 ();
 FILLCELL_X32 FILLER_167_571 ();
 FILLCELL_X32 FILLER_167_603 ();
 FILLCELL_X32 FILLER_167_635 ();
 FILLCELL_X32 FILLER_167_667 ();
 FILLCELL_X32 FILLER_167_699 ();
 FILLCELL_X32 FILLER_167_731 ();
 FILLCELL_X32 FILLER_167_763 ();
 FILLCELL_X32 FILLER_167_795 ();
 FILLCELL_X32 FILLER_167_827 ();
 FILLCELL_X32 FILLER_167_859 ();
 FILLCELL_X32 FILLER_167_891 ();
 FILLCELL_X16 FILLER_167_923 ();
 FILLCELL_X8 FILLER_167_939 ();
 FILLCELL_X4 FILLER_167_947 ();
 FILLCELL_X2 FILLER_167_951 ();
 FILLCELL_X1 FILLER_167_953 ();
 FILLCELL_X8 FILLER_167_956 ();
 FILLCELL_X1 FILLER_167_964 ();
 FILLCELL_X2 FILLER_167_967 ();
 FILLCELL_X1 FILLER_167_969 ();
 FILLCELL_X4 FILLER_167_972 ();
 FILLCELL_X4 FILLER_167_994 ();
 FILLCELL_X2 FILLER_167_1010 ();
 FILLCELL_X1 FILLER_167_1012 ();
 FILLCELL_X8 FILLER_167_1029 ();
 FILLCELL_X4 FILLER_167_1039 ();
 FILLCELL_X2 FILLER_167_1043 ();
 FILLCELL_X1 FILLER_167_1061 ();
 FILLCELL_X8 FILLER_167_1064 ();
 FILLCELL_X2 FILLER_167_1072 ();
 FILLCELL_X4 FILLER_167_1097 ();
 FILLCELL_X1 FILLER_167_1101 ();
 FILLCELL_X1 FILLER_167_1116 ();
 FILLCELL_X1 FILLER_167_1120 ();
 FILLCELL_X1 FILLER_167_1127 ();
 FILLCELL_X32 FILLER_167_1155 ();
 FILLCELL_X32 FILLER_167_1187 ();
 FILLCELL_X32 FILLER_167_1219 ();
 FILLCELL_X8 FILLER_167_1251 ();
 FILLCELL_X1 FILLER_167_1259 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X8 FILLER_168_385 ();
 FILLCELL_X1 FILLER_168_393 ();
 FILLCELL_X32 FILLER_168_397 ();
 FILLCELL_X32 FILLER_168_429 ();
 FILLCELL_X32 FILLER_168_461 ();
 FILLCELL_X32 FILLER_168_493 ();
 FILLCELL_X32 FILLER_168_525 ();
 FILLCELL_X32 FILLER_168_557 ();
 FILLCELL_X32 FILLER_168_589 ();
 FILLCELL_X8 FILLER_168_621 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X8 FILLER_168_952 ();
 FILLCELL_X2 FILLER_168_960 ();
 FILLCELL_X4 FILLER_168_978 ();
 FILLCELL_X1 FILLER_168_982 ();
 FILLCELL_X4 FILLER_168_993 ();
 FILLCELL_X1 FILLER_168_997 ();
 FILLCELL_X8 FILLER_168_1016 ();
 FILLCELL_X4 FILLER_168_1026 ();
 FILLCELL_X1 FILLER_168_1030 ();
 FILLCELL_X2 FILLER_168_1047 ();
 FILLCELL_X1 FILLER_168_1049 ();
 FILLCELL_X4 FILLER_168_1052 ();
 FILLCELL_X2 FILLER_168_1056 ();
 FILLCELL_X4 FILLER_168_1068 ();
 FILLCELL_X2 FILLER_168_1072 ();
 FILLCELL_X4 FILLER_168_1112 ();
 FILLCELL_X2 FILLER_168_1116 ();
 FILLCELL_X1 FILLER_168_1118 ();
 FILLCELL_X8 FILLER_168_1126 ();
 FILLCELL_X32 FILLER_168_1138 ();
 FILLCELL_X32 FILLER_168_1170 ();
 FILLCELL_X32 FILLER_168_1202 ();
 FILLCELL_X16 FILLER_168_1234 ();
 FILLCELL_X8 FILLER_168_1250 ();
 FILLCELL_X2 FILLER_168_1258 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X16 FILLER_169_545 ();
 FILLCELL_X8 FILLER_169_561 ();
 FILLCELL_X2 FILLER_169_569 ();
 FILLCELL_X1 FILLER_169_575 ();
 FILLCELL_X8 FILLER_169_580 ();
 FILLCELL_X2 FILLER_169_588 ();
 FILLCELL_X1 FILLER_169_590 ();
 FILLCELL_X8 FILLER_169_595 ();
 FILLCELL_X2 FILLER_169_603 ();
 FILLCELL_X1 FILLER_169_605 ();
 FILLCELL_X4 FILLER_169_609 ();
 FILLCELL_X1 FILLER_169_613 ();
 FILLCELL_X2 FILLER_169_619 ();
 FILLCELL_X8 FILLER_169_624 ();
 FILLCELL_X1 FILLER_169_632 ();
 FILLCELL_X16 FILLER_169_636 ();
 FILLCELL_X2 FILLER_169_658 ();
 FILLCELL_X1 FILLER_169_660 ();
 FILLCELL_X8 FILLER_169_664 ();
 FILLCELL_X4 FILLER_169_672 ();
 FILLCELL_X2 FILLER_169_676 ();
 FILLCELL_X32 FILLER_169_681 ();
 FILLCELL_X32 FILLER_169_713 ();
 FILLCELL_X32 FILLER_169_745 ();
 FILLCELL_X4 FILLER_169_777 ();
 FILLCELL_X32 FILLER_169_784 ();
 FILLCELL_X32 FILLER_169_816 ();
 FILLCELL_X32 FILLER_169_848 ();
 FILLCELL_X32 FILLER_169_880 ();
 FILLCELL_X32 FILLER_169_912 ();
 FILLCELL_X32 FILLER_169_944 ();
 FILLCELL_X1 FILLER_169_976 ();
 FILLCELL_X4 FILLER_169_979 ();
 FILLCELL_X2 FILLER_169_983 ();
 FILLCELL_X1 FILLER_169_1003 ();
 FILLCELL_X2 FILLER_169_1020 ();
 FILLCELL_X4 FILLER_169_1049 ();
 FILLCELL_X2 FILLER_169_1063 ();
 FILLCELL_X2 FILLER_169_1067 ();
 FILLCELL_X4 FILLER_169_1071 ();
 FILLCELL_X2 FILLER_169_1075 ();
 FILLCELL_X32 FILLER_169_1095 ();
 FILLCELL_X32 FILLER_169_1127 ();
 FILLCELL_X32 FILLER_169_1159 ();
 FILLCELL_X32 FILLER_169_1191 ();
 FILLCELL_X32 FILLER_169_1223 ();
 FILLCELL_X4 FILLER_169_1255 ();
 FILLCELL_X1 FILLER_169_1259 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X4 FILLER_170_545 ();
 FILLCELL_X2 FILLER_170_549 ();
 FILLCELL_X1 FILLER_170_551 ();
 FILLCELL_X4 FILLER_170_556 ();
 FILLCELL_X2 FILLER_170_560 ();
 FILLCELL_X1 FILLER_170_566 ();
 FILLCELL_X4 FILLER_170_572 ();
 FILLCELL_X4 FILLER_170_583 ();
 FILLCELL_X1 FILLER_170_590 ();
 FILLCELL_X1 FILLER_170_595 ();
 FILLCELL_X1 FILLER_170_599 ();
 FILLCELL_X4 FILLER_170_617 ();
 FILLCELL_X1 FILLER_170_630 ();
 FILLCELL_X2 FILLER_170_641 ();
 FILLCELL_X1 FILLER_170_643 ();
 FILLCELL_X2 FILLER_170_650 ();
 FILLCELL_X1 FILLER_170_652 ();
 FILLCELL_X2 FILLER_170_663 ();
 FILLCELL_X4 FILLER_170_672 ();
 FILLCELL_X1 FILLER_170_676 ();
 FILLCELL_X32 FILLER_170_686 ();
 FILLCELL_X32 FILLER_170_718 ();
 FILLCELL_X32 FILLER_170_750 ();
 FILLCELL_X16 FILLER_170_782 ();
 FILLCELL_X2 FILLER_170_798 ();
 FILLCELL_X1 FILLER_170_800 ();
 FILLCELL_X8 FILLER_170_804 ();
 FILLCELL_X4 FILLER_170_812 ();
 FILLCELL_X2 FILLER_170_816 ();
 FILLCELL_X32 FILLER_170_821 ();
 FILLCELL_X32 FILLER_170_853 ();
 FILLCELL_X32 FILLER_170_885 ();
 FILLCELL_X32 FILLER_170_917 ();
 FILLCELL_X16 FILLER_170_949 ();
 FILLCELL_X4 FILLER_170_965 ();
 FILLCELL_X2 FILLER_170_969 ();
 FILLCELL_X4 FILLER_170_987 ();
 FILLCELL_X2 FILLER_170_991 ();
 FILLCELL_X1 FILLER_170_993 ();
 FILLCELL_X8 FILLER_170_1010 ();
 FILLCELL_X4 FILLER_170_1018 ();
 FILLCELL_X2 FILLER_170_1022 ();
 FILLCELL_X1 FILLER_170_1024 ();
 FILLCELL_X4 FILLER_170_1027 ();
 FILLCELL_X2 FILLER_170_1031 ();
 FILLCELL_X4 FILLER_170_1045 ();
 FILLCELL_X2 FILLER_170_1049 ();
 FILLCELL_X32 FILLER_170_1071 ();
 FILLCELL_X32 FILLER_170_1103 ();
 FILLCELL_X32 FILLER_170_1135 ();
 FILLCELL_X32 FILLER_170_1167 ();
 FILLCELL_X32 FILLER_170_1199 ();
 FILLCELL_X16 FILLER_170_1231 ();
 FILLCELL_X8 FILLER_170_1247 ();
 FILLCELL_X4 FILLER_170_1255 ();
 FILLCELL_X1 FILLER_170_1259 ();
endmodule
