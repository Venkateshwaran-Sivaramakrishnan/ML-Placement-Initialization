module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire net807;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire net928;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire net705;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire net834;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire net657;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire net765;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt_next[0] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net43;
 wire net44;
 wire net46;
 wire net48;
 wire net49;
 wire net50;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net65;
 wire net66;
 wire net67;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net12;
 wire net31;
 wire net42;
 wire net45;
 wire net47;
 wire net51;
 wire net64;
 wire net68;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net706;
 wire net707;
 wire net708;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net766;
 wire net767;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net927;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;

 INVx1_ASAP7_75t_R _16086_ (.A(_16081_),
    .Y(\u0.r0.rcnt[1] ));
 INVx2_ASAP7_75t_R _16087_ (.A(\u0.r0.rcnt_next[0] ),
    .Y(\u0.r0.rcnt[0] ));
 INVx4_ASAP7_75t_R _16088_ (.A(net195),
    .Y(_07939_));
 BUFx6f_ASAP7_75t_R _16089_ (.A(_07939_),
    .Y(_07940_));
 OR2x2_ASAP7_75t_R _16090_ (.A(net105),
    .B(net14),
    .Y(_07941_));
 BUFx4f_ASAP7_75t_R _16091_ (.A(_01005_),
    .Y(_07942_));
 XNOR2x2_ASAP7_75t_R _16092_ (.A(_07942_),
    .B(_01037_),
    .Y(_07943_));
 INVx1_ASAP7_75t_R _16093_ (.A(_07943_),
    .Y(_07944_));
 BUFx6f_ASAP7_75t_R _16094_ (.A(_01101_),
    .Y(_07945_));
 XOR2x2_ASAP7_75t_R _16095_ (.A(_01069_),
    .B(_07945_),
    .Y(_07946_));
 XNOR2x1_ASAP7_75t_R _16096_ (.B(_07946_),
    .Y(_07947_),
    .A(_00441_));
 NAND2x1_ASAP7_75t_R _16097_ (.A(_07944_),
    .B(_07947_),
    .Y(_07948_));
 XOR2x1_ASAP7_75t_R _16098_ (.A(_07946_),
    .Y(_07949_),
    .B(_00441_));
 NAND2x1_ASAP7_75t_R _16099_ (.A(_07943_),
    .B(_07949_),
    .Y(_07950_));
 BUFx12_ASAP7_75t_R _16100_ (.A(net195),
    .Y(_07951_));
 AO21x2_ASAP7_75t_R _16101_ (.A1(_07948_),
    .A2(_07950_),
    .B(_07951_),
    .Y(_07952_));
 NAND2x2_ASAP7_75t_R _16102_ (.A(_07941_),
    .B(_07952_),
    .Y(_07953_));
 CKINVDCx8_ASAP7_75t_R _16103_ (.A(_07953_),
    .Y(_07954_));
 BUFx6f_ASAP7_75t_R _16104_ (.A(_07954_),
    .Y(_07955_));
 BUFx6f_ASAP7_75t_R _16105_ (.A(_07955_),
    .Y(_00390_));
 BUFx12_ASAP7_75t_R _16106_ (.A(_07940_),
    .Y(_07956_));
 BUFx16f_ASAP7_75t_R _16107_ (.A(_07940_),
    .Y(_07957_));
 BUFx4f_ASAP7_75t_R _16108_ (.A(_01002_),
    .Y(_07958_));
 XNOR2x2_ASAP7_75t_R _16109_ (.A(_00439_),
    .B(_07958_),
    .Y(_07959_));
 BUFx6f_ASAP7_75t_R _16110_ (.A(_01034_),
    .Y(_07960_));
 BUFx6f_ASAP7_75t_R _16111_ (.A(_01066_),
    .Y(_07961_));
 XNOR2x1_ASAP7_75t_R _16112_ (.B(_07961_),
    .Y(_07962_),
    .A(_07960_));
 XOR2x2_ASAP7_75t_R _16113_ (.A(_07962_),
    .B(_07959_),
    .Y(_07963_));
 XOR2x1_ASAP7_75t_R _16114_ (.A(_07963_),
    .Y(_07964_),
    .B(_01098_));
 NAND2x1_ASAP7_75t_R _16115_ (.A(_07957_),
    .B(_07964_),
    .Y(_07965_));
 OAI21x1_ASAP7_75t_R _16116_ (.A1(net102),
    .A2(_07956_),
    .B(_07965_),
    .Y(_07966_));
 BUFx12_ASAP7_75t_R _16117_ (.A(net839),
    .Y(_15732_));
 BUFx12f_ASAP7_75t_R _16118_ (.A(_07951_),
    .Y(_07967_));
 INVx1_ASAP7_75t_R _16119_ (.A(net103),
    .Y(_07968_));
 BUFx4f_ASAP7_75t_R _16120_ (.A(_01003_),
    .Y(_07969_));
 BUFx3_ASAP7_75t_R _16121_ (.A(_01035_),
    .Y(_07970_));
 XOR2x2_ASAP7_75t_R _16122_ (.A(_07969_),
    .B(_07970_),
    .Y(_07971_));
 BUFx6f_ASAP7_75t_R _16123_ (.A(_01067_),
    .Y(_07972_));
 BUFx6f_ASAP7_75t_R _16124_ (.A(_01099_),
    .Y(_07973_));
 XOR2x1_ASAP7_75t_R _16125_ (.A(_07972_),
    .Y(_07974_),
    .B(_07973_));
 XOR2x1_ASAP7_75t_R _16126_ (.A(_07974_),
    .Y(_07975_),
    .B(_00440_));
 XNOR2x2_ASAP7_75t_R _16127_ (.A(_07971_),
    .B(_07975_),
    .Y(_07976_));
 NOR2x1_ASAP7_75t_R _16128_ (.A(_07967_),
    .B(_07976_),
    .Y(_07977_));
 AOI21x1_ASAP7_75t_R _16129_ (.A1(_07967_),
    .A2(_07968_),
    .B(_07977_),
    .Y(_07978_));
 BUFx16f_ASAP7_75t_R _16130_ (.A(_07978_),
    .Y(_15729_));
 CKINVDCx6p67_ASAP7_75t_R _16131_ (.A(_15729_),
    .Y(_15735_));
 BUFx6f_ASAP7_75t_R _16132_ (.A(_07957_),
    .Y(_07979_));
 BUFx6f_ASAP7_75t_R _16133_ (.A(_07979_),
    .Y(_07980_));
 XNOR2x1_ASAP7_75t_R _16134_ (.B(_01008_),
    .Y(_07981_),
    .A(_00443_));
 INVx1_ASAP7_75t_R _16135_ (.A(_01040_),
    .Y(_07982_));
 XOR2x2_ASAP7_75t_R _16136_ (.A(_07981_),
    .B(_07982_),
    .Y(_07983_));
 BUFx4f_ASAP7_75t_R _16137_ (.A(_01072_),
    .Y(_07984_));
 XOR2x2_ASAP7_75t_R _16138_ (.A(_07983_),
    .B(_07984_),
    .Y(_07985_));
 XOR2x1_ASAP7_75t_R _16139_ (.A(_07985_),
    .Y(_07986_),
    .B(_01104_));
 BUFx6f_ASAP7_75t_R _16140_ (.A(_07956_),
    .Y(_07987_));
 NOR2x1_ASAP7_75t_R _16141_ (.A(net108),
    .B(_07987_),
    .Y(_07988_));
 AOI21x1_ASAP7_75t_R _16142_ (.A1(_07980_),
    .A2(_07986_),
    .B(_07988_),
    .Y(_07989_));
 BUFx6f_ASAP7_75t_R _16143_ (.A(_07989_),
    .Y(_07990_));
 BUFx6f_ASAP7_75t_R _16144_ (.A(_07990_),
    .Y(_00392_));
 XNOR2x1_ASAP7_75t_R _16145_ (.B(_01007_),
    .Y(_07991_),
    .A(_00442_));
 INVx1_ASAP7_75t_R _16146_ (.A(_01039_),
    .Y(_07992_));
 XOR2x2_ASAP7_75t_R _16147_ (.A(_07991_),
    .B(_07992_),
    .Y(_07993_));
 BUFx4f_ASAP7_75t_R _16148_ (.A(_01071_),
    .Y(_07994_));
 XOR2x2_ASAP7_75t_R _16149_ (.A(_07993_),
    .B(_07994_),
    .Y(_07995_));
 BUFx4f_ASAP7_75t_R _16150_ (.A(_01103_),
    .Y(_07996_));
 XOR2x1_ASAP7_75t_R _16151_ (.A(_07995_),
    .Y(_07997_),
    .B(_07996_));
 NOR2x1_ASAP7_75t_R _16152_ (.A(net107),
    .B(_07956_),
    .Y(_07998_));
 AOI21x1_ASAP7_75t_R _16153_ (.A1(_07979_),
    .A2(_07997_),
    .B(_07998_),
    .Y(_07999_));
 BUFx6f_ASAP7_75t_R _16154_ (.A(_07999_),
    .Y(_08000_));
 BUFx6f_ASAP7_75t_R _16155_ (.A(_08000_),
    .Y(_08001_));
 BUFx6f_ASAP7_75t_R _16156_ (.A(_08001_),
    .Y(_00391_));
 BUFx4f_ASAP7_75t_R _16157_ (.A(_01004_),
    .Y(_08002_));
 XOR2x1_ASAP7_75t_R _16158_ (.A(_00416_),
    .Y(_08003_),
    .B(_08002_));
 BUFx4f_ASAP7_75t_R _16159_ (.A(_01036_),
    .Y(_08004_));
 XOR2x2_ASAP7_75t_R _16160_ (.A(_08003_),
    .B(_08004_),
    .Y(_08005_));
 NAND2x2_ASAP7_75t_R _16161_ (.A(_07940_),
    .B(_08005_),
    .Y(_08006_));
 BUFx6f_ASAP7_75t_R _16162_ (.A(_01068_),
    .Y(_08007_));
 BUFx6f_ASAP7_75t_R _16163_ (.A(_01100_),
    .Y(_08008_));
 XNOR2x2_ASAP7_75t_R _16164_ (.A(_08007_),
    .B(_08008_),
    .Y(_08009_));
 AND2x2_ASAP7_75t_R _16165_ (.A(_07951_),
    .B(net104),
    .Y(_08010_));
 AO21x1_ASAP7_75t_R _16166_ (.A1(_08009_),
    .A2(net14),
    .B(_08010_),
    .Y(_08011_));
 NAND2x1_ASAP7_75t_R _16167_ (.A(_08011_),
    .B(_08006_),
    .Y(_08012_));
 OAI21x1_ASAP7_75t_R _16168_ (.A1(_08006_),
    .A2(_08009_),
    .B(_08012_),
    .Y(_08013_));
 BUFx16f_ASAP7_75t_R _16169_ (.A(_08013_),
    .Y(_08014_));
 BUFx6f_ASAP7_75t_R _16170_ (.A(_08014_),
    .Y(_15742_));
 XNOR2x2_ASAP7_75t_R _16171_ (.A(_00425_),
    .B(_00995_),
    .Y(_08015_));
 BUFx6f_ASAP7_75t_R _16172_ (.A(_01027_),
    .Y(_08016_));
 XNOR2x1_ASAP7_75t_R _16173_ (.B(_01059_),
    .Y(_08017_),
    .A(_08016_));
 XOR2x2_ASAP7_75t_R _16174_ (.A(_08015_),
    .B(_08017_),
    .Y(_08018_));
 XOR2x1_ASAP7_75t_R _16175_ (.A(_08018_),
    .Y(_08019_),
    .B(_01091_));
 NAND2x1_ASAP7_75t_R _16176_ (.A(_08019_),
    .B(_07957_),
    .Y(_08020_));
 OAI21x1_ASAP7_75t_R _16177_ (.A1(_07957_),
    .A2(net12),
    .B(_08020_),
    .Y(_08021_));
 BUFx10_ASAP7_75t_R _16178_ (.A(_08021_),
    .Y(_15768_));
 NOR2x2_ASAP7_75t_R _16179_ (.A(net106),
    .B(_07957_),
    .Y(_08022_));
 BUFx6f_ASAP7_75t_R _16180_ (.A(_01006_),
    .Y(_08023_));
 BUFx6f_ASAP7_75t_R _16181_ (.A(_01038_),
    .Y(_08024_));
 XOR2x2_ASAP7_75t_R _16182_ (.A(_08023_),
    .B(_08024_),
    .Y(_08025_));
 BUFx6f_ASAP7_75t_R _16183_ (.A(_01070_),
    .Y(_08026_));
 XOR2x1_ASAP7_75t_R _16184_ (.A(_08026_),
    .Y(_08027_),
    .B(_01102_));
 XOR2x1_ASAP7_75t_R _16185_ (.A(_08027_),
    .Y(_08028_),
    .B(_00426_));
 XNOR2x1_ASAP7_75t_R _16186_ (.B(_08028_),
    .Y(_08029_),
    .A(_08025_));
 NOR2x2_ASAP7_75t_R _16187_ (.A(_07951_),
    .B(_08029_),
    .Y(_08030_));
 NOR2x2_ASAP7_75t_R _16188_ (.A(_08022_),
    .B(_08030_),
    .Y(_15765_));
 INVx5_ASAP7_75t_R _16189_ (.A(_15765_),
    .Y(_15771_));
 BUFx6f_ASAP7_75t_R _16190_ (.A(_01017_),
    .Y(_08031_));
 XOR2x1_ASAP7_75t_R _16191_ (.A(_00423_),
    .Y(_08032_),
    .B(_08031_));
 BUFx6f_ASAP7_75t_R _16192_ (.A(_01049_),
    .Y(_08033_));
 XOR2x2_ASAP7_75t_R _16193_ (.A(_08032_),
    .B(_08033_),
    .Y(_08034_));
 BUFx10_ASAP7_75t_R _16194_ (.A(_01081_),
    .Y(_08035_));
 XNOR2x1_ASAP7_75t_R _16195_ (.B(_01113_),
    .Y(_08036_),
    .A(_08035_));
 INVx1_ASAP7_75t_R _16196_ (.A(_08036_),
    .Y(_08037_));
 NAND3x2_ASAP7_75t_R _16197_ (.B(net14),
    .C(_08037_),
    .Y(_08038_),
    .A(_08034_));
 AND2x2_ASAP7_75t_R _16198_ (.A(net195),
    .B(net117),
    .Y(_08039_));
 AO21x1_ASAP7_75t_R _16199_ (.A1(_08036_),
    .A2(_07939_),
    .B(_08039_),
    .Y(_08040_));
 NAND2x2_ASAP7_75t_R _16200_ (.A(_07939_),
    .B(_08034_),
    .Y(_08041_));
 NAND2x2_ASAP7_75t_R _16201_ (.A(_08040_),
    .B(_08041_),
    .Y(_08042_));
 NAND2x2_ASAP7_75t_R _16202_ (.A(_08038_),
    .B(_08042_),
    .Y(_08043_));
 BUFx10_ASAP7_75t_R _16203_ (.A(_08043_),
    .Y(_15778_));
 OR2x2_ASAP7_75t_R _16204_ (.A(net128),
    .B(net14),
    .Y(_08044_));
 XNOR2x2_ASAP7_75t_R _16205_ (.A(_01020_),
    .B(_01052_),
    .Y(_08045_));
 INVx1_ASAP7_75t_R _16206_ (.A(_08045_),
    .Y(_08046_));
 BUFx6f_ASAP7_75t_R _16207_ (.A(_01084_),
    .Y(_08047_));
 XOR2x2_ASAP7_75t_R _16208_ (.A(_08047_),
    .B(_01116_),
    .Y(_08048_));
 XNOR2x1_ASAP7_75t_R _16209_ (.B(_08048_),
    .Y(_08049_),
    .A(_00427_));
 NAND2x1_ASAP7_75t_R _16210_ (.A(_08046_),
    .B(_08049_),
    .Y(_08050_));
 XOR2x1_ASAP7_75t_R _16211_ (.A(_08048_),
    .Y(_08051_),
    .B(_00427_));
 NAND2x1_ASAP7_75t_R _16212_ (.A(_08045_),
    .B(_08051_),
    .Y(_08052_));
 AO21x2_ASAP7_75t_R _16213_ (.A1(_08050_),
    .A2(_08052_),
    .B(_07951_),
    .Y(_08053_));
 NAND2x2_ASAP7_75t_R _16214_ (.A(_08044_),
    .B(_08053_),
    .Y(_08054_));
 INVx2_ASAP7_75t_R _16215_ (.A(_08054_),
    .Y(_08055_));
 BUFx6f_ASAP7_75t_R _16216_ (.A(_08055_),
    .Y(_08056_));
 BUFx6f_ASAP7_75t_R _16217_ (.A(_08056_),
    .Y(_00400_));
 XNOR2x1_ASAP7_75t_R _16218_ (.B(_01021_),
    .Y(_08057_),
    .A(_00428_));
 INVx2_ASAP7_75t_R _16219_ (.A(_01053_),
    .Y(_08058_));
 XOR2x2_ASAP7_75t_R _16220_ (.A(_08057_),
    .B(_08058_),
    .Y(_08059_));
 XOR2x2_ASAP7_75t_R _16221_ (.A(_08059_),
    .B(_01085_),
    .Y(_08060_));
 XOR2x1_ASAP7_75t_R _16222_ (.A(_08060_),
    .Y(_08061_),
    .B(_01117_));
 NOR2x1_ASAP7_75t_R _16223_ (.A(net139),
    .B(_07979_),
    .Y(_08062_));
 AOI21x1_ASAP7_75t_R _16224_ (.A1(_07980_),
    .A2(_08061_),
    .B(_08062_),
    .Y(_08063_));
 BUFx6f_ASAP7_75t_R _16225_ (.A(_08063_),
    .Y(_08064_));
 BUFx10_ASAP7_75t_R _16226_ (.A(_08064_),
    .Y(_00401_));
 XNOR2x1_ASAP7_75t_R _16227_ (.B(_01022_),
    .Y(_08065_),
    .A(_00429_));
 INVx2_ASAP7_75t_R _16228_ (.A(_01054_),
    .Y(_08066_));
 XOR2x2_ASAP7_75t_R _16229_ (.A(_08065_),
    .B(_08066_),
    .Y(_08067_));
 XOR2x2_ASAP7_75t_R _16230_ (.A(_08067_),
    .B(_01086_),
    .Y(_08068_));
 XOR2x1_ASAP7_75t_R _16231_ (.A(_08068_),
    .Y(_08069_),
    .B(_01118_));
 NOR2x1_ASAP7_75t_R _16232_ (.A(net150),
    .B(_07979_),
    .Y(_08070_));
 AOI21x1_ASAP7_75t_R _16233_ (.A1(_07987_),
    .A2(_08069_),
    .B(_08070_),
    .Y(_08071_));
 BUFx6f_ASAP7_75t_R _16234_ (.A(_08071_),
    .Y(_08072_));
 BUFx10_ASAP7_75t_R _16235_ (.A(_08072_),
    .Y(_00402_));
 XNOR2x2_ASAP7_75t_R _16236_ (.A(_00430_),
    .B(_01023_),
    .Y(_08073_));
 XNOR2x1_ASAP7_75t_R _16237_ (.B(_08073_),
    .Y(_08074_),
    .A(_01055_));
 XOR2x2_ASAP7_75t_R _16238_ (.A(_08074_),
    .B(_01087_),
    .Y(_08075_));
 XOR2x1_ASAP7_75t_R _16239_ (.A(_08075_),
    .Y(_08076_),
    .B(_01119_));
 NAND2x1_ASAP7_75t_R _16240_ (.A(_07980_),
    .B(_08076_),
    .Y(_08077_));
 OAI21x1_ASAP7_75t_R _16241_ (.A1(_07980_),
    .A2(net161),
    .B(_08077_),
    .Y(_08078_));
 CKINVDCx6p67_ASAP7_75t_R _16242_ (.A(_08078_),
    .Y(_08079_));
 BUFx10_ASAP7_75t_R _16243_ (.A(_08079_),
    .Y(_00403_));
 BUFx10_ASAP7_75t_R _16244_ (.A(_07987_),
    .Y(_08080_));
 XNOR2x1_ASAP7_75t_R _16245_ (.B(_01024_),
    .Y(_08081_),
    .A(_00431_));
 XNOR2x2_ASAP7_75t_R _16246_ (.A(_01056_),
    .B(_08081_),
    .Y(_08082_));
 XOR2x2_ASAP7_75t_R _16247_ (.A(_08082_),
    .B(_01088_),
    .Y(_08083_));
 XOR2x1_ASAP7_75t_R _16248_ (.A(_08083_),
    .Y(_08084_),
    .B(_01120_));
 NAND2x1_ASAP7_75t_R _16249_ (.A(_07980_),
    .B(_08084_),
    .Y(_08085_));
 OA21x2_ASAP7_75t_R _16250_ (.A1(_08080_),
    .A2(net172),
    .B(_08085_),
    .Y(_08086_));
 BUFx10_ASAP7_75t_R _16251_ (.A(_08086_),
    .Y(_00404_));
 INVx1_ASAP7_75t_R _16252_ (.A(net183),
    .Y(_08087_));
 XNOR2x1_ASAP7_75t_R _16253_ (.B(_01057_),
    .Y(_08088_),
    .A(_01025_));
 XOR2x2_ASAP7_75t_R _16254_ (.A(_01089_),
    .B(_01121_),
    .Y(_08089_));
 XOR2x1_ASAP7_75t_R _16255_ (.A(_08089_),
    .Y(_08090_),
    .B(_00432_));
 NAND2x1_ASAP7_75t_R _16256_ (.A(_08088_),
    .B(_08090_),
    .Y(_08091_));
 INVx1_ASAP7_75t_R _16257_ (.A(_08088_),
    .Y(_08092_));
 XNOR2x1_ASAP7_75t_R _16258_ (.B(_08089_),
    .Y(_08093_),
    .A(_00432_));
 NAND2x1_ASAP7_75t_R _16259_ (.A(_08092_),
    .B(_08093_),
    .Y(_08094_));
 AOI21x1_ASAP7_75t_R _16260_ (.A1(_08091_),
    .A2(_08094_),
    .B(_07951_),
    .Y(_08095_));
 AOI21x1_ASAP7_75t_R _16261_ (.A1(_07967_),
    .A2(_08087_),
    .B(_08095_),
    .Y(_08096_));
 BUFx16f_ASAP7_75t_R _16262_ (.A(_08096_),
    .Y(_15748_));
 INVx4_ASAP7_75t_R _16263_ (.A(_15748_),
    .Y(_15750_));
 BUFx2_ASAP7_75t_R rebuffer475 (.A(_01058_),
    .Y(net928));
 XOR2x2_ASAP7_75t_R _16265_ (.A(_01058_),
    .B(_00433_),
    .Y(_08098_));
 BUFx6f_ASAP7_75t_R _16266_ (.A(_01090_),
    .Y(_08099_));
 XOR2x1_ASAP7_75t_R _16267_ (.A(_08098_),
    .Y(_08100_),
    .B(_08099_));
 BUFx6f_ASAP7_75t_R _16268_ (.A(_01026_),
    .Y(_08101_));
 XOR2x1_ASAP7_75t_R _16269_ (.A(_00642_),
    .Y(_08102_),
    .B(_08101_));
 XOR2x1_ASAP7_75t_R _16270_ (.A(_08100_),
    .Y(_08103_),
    .B(_08102_));
 NAND2x1_ASAP7_75t_R _16271_ (.A(_07957_),
    .B(_08103_),
    .Y(_08104_));
 OAI21x1_ASAP7_75t_R _16272_ (.A1(_07956_),
    .A2(net194),
    .B(_08104_),
    .Y(_08105_));
 BUFx16f_ASAP7_75t_R _16273_ (.A(_08105_),
    .Y(_15753_));
 BUFx6f_ASAP7_75t_R _16274_ (.A(_00996_),
    .Y(_08106_));
 XOR2x1_ASAP7_75t_R _16275_ (.A(_00424_),
    .Y(_08107_),
    .B(_08106_));
 BUFx4f_ASAP7_75t_R _16276_ (.A(_01028_),
    .Y(_08108_));
 XOR2x2_ASAP7_75t_R _16277_ (.A(_08107_),
    .B(_08108_),
    .Y(_08109_));
 BUFx10_ASAP7_75t_R _16278_ (.A(_01060_),
    .Y(_08110_));
 BUFx6f_ASAP7_75t_R _16279_ (.A(_01092_),
    .Y(_08111_));
 XNOR2x1_ASAP7_75t_R _16280_ (.B(_08111_),
    .Y(_08112_),
    .A(_08110_));
 INVx1_ASAP7_75t_R _16281_ (.A(_08112_),
    .Y(_08113_));
 NAND3x2_ASAP7_75t_R _16282_ (.B(net14),
    .C(_08113_),
    .Y(_08114_),
    .A(_08109_));
 AND2x2_ASAP7_75t_R _16283_ (.A(net195),
    .B(net78),
    .Y(_08115_));
 AO21x1_ASAP7_75t_R _16284_ (.A1(_08112_),
    .A2(_07939_),
    .B(_08115_),
    .Y(_08116_));
 NAND2x2_ASAP7_75t_R _16285_ (.A(_07939_),
    .B(_08109_),
    .Y(_08117_));
 NAND2x2_ASAP7_75t_R _16286_ (.A(_08116_),
    .B(_08117_),
    .Y(_08118_));
 NAND2x2_ASAP7_75t_R _16287_ (.A(_08114_),
    .B(_08118_),
    .Y(_08119_));
 BUFx12_ASAP7_75t_R _16288_ (.A(_08119_),
    .Y(_15760_));
 XNOR2x1_ASAP7_75t_R _16289_ (.B(_00997_),
    .Y(_08120_),
    .A(_00434_));
 INVx1_ASAP7_75t_R _16290_ (.A(_01029_),
    .Y(_08121_));
 XOR2x2_ASAP7_75t_R _16291_ (.A(_08120_),
    .B(_08121_),
    .Y(_08122_));
 XOR2x2_ASAP7_75t_R _16292_ (.A(_08122_),
    .B(_01061_),
    .Y(_08123_));
 BUFx3_ASAP7_75t_R _16293_ (.A(_01093_),
    .Y(_08124_));
 XOR2x2_ASAP7_75t_R _16294_ (.A(_08123_),
    .B(_08124_),
    .Y(_08125_));
 NOR2x2_ASAP7_75t_R _16295_ (.A(net89),
    .B(_07957_),
    .Y(_08126_));
 AOI21x1_ASAP7_75t_R _16296_ (.A1(_07979_),
    .A2(_08125_),
    .B(_08126_),
    .Y(_08127_));
 BUFx6f_ASAP7_75t_R _16297_ (.A(_08127_),
    .Y(_08128_));
 BUFx6f_ASAP7_75t_R _16298_ (.A(_08128_),
    .Y(_00385_));
 XNOR2x2_ASAP7_75t_R _16299_ (.A(_00435_),
    .B(_00998_),
    .Y(_08129_));
 INVx1_ASAP7_75t_R _16300_ (.A(_01030_),
    .Y(_08130_));
 XOR2x1_ASAP7_75t_R _16301_ (.A(_08129_),
    .Y(_08131_),
    .B(_08130_));
 XOR2x2_ASAP7_75t_R _16302_ (.A(_08131_),
    .B(_01062_),
    .Y(_08132_));
 BUFx4f_ASAP7_75t_R _16303_ (.A(_01094_),
    .Y(_08133_));
 XOR2x1_ASAP7_75t_R _16304_ (.A(_08132_),
    .Y(_08134_),
    .B(_08133_));
 NOR2x1_ASAP7_75t_R _16305_ (.A(net98),
    .B(_07956_),
    .Y(_08135_));
 AOI21x1_ASAP7_75t_R _16306_ (.A1(_07956_),
    .A2(_08134_),
    .B(_08135_),
    .Y(_08136_));
 BUFx6f_ASAP7_75t_R _16307_ (.A(_08136_),
    .Y(_08137_));
 BUFx6f_ASAP7_75t_R _16308_ (.A(_08137_),
    .Y(_00386_));
 XNOR2x2_ASAP7_75t_R _16309_ (.A(_00436_),
    .B(_00999_),
    .Y(_08138_));
 INVx2_ASAP7_75t_R _16310_ (.A(_01031_),
    .Y(_08139_));
 XOR2x1_ASAP7_75t_R _16311_ (.A(_08138_),
    .Y(_08140_),
    .B(_08139_));
 XOR2x2_ASAP7_75t_R _16312_ (.A(_08140_),
    .B(_01063_),
    .Y(_08141_));
 XOR2x2_ASAP7_75t_R _16313_ (.A(_08141_),
    .B(_01095_),
    .Y(_08142_));
 NAND2x1_ASAP7_75t_R _16314_ (.A(_07987_),
    .B(_08142_),
    .Y(_08143_));
 OAI21x1_ASAP7_75t_R _16315_ (.A1(_07987_),
    .A2(net99),
    .B(_08143_),
    .Y(_08144_));
 INVx5_ASAP7_75t_R _16316_ (.A(_08144_),
    .Y(_08145_));
 BUFx10_ASAP7_75t_R _16317_ (.A(_08145_),
    .Y(_00387_));
 XNOR2x2_ASAP7_75t_R _16318_ (.A(_00437_),
    .B(_01000_),
    .Y(_08146_));
 INVx1_ASAP7_75t_R _16319_ (.A(_01032_),
    .Y(_08147_));
 XOR2x1_ASAP7_75t_R _16320_ (.A(_08146_),
    .Y(_08148_),
    .B(_08147_));
 XOR2x2_ASAP7_75t_R _16321_ (.A(_08148_),
    .B(_01064_),
    .Y(_08149_));
 XOR2x2_ASAP7_75t_R _16322_ (.A(_08149_),
    .B(_01096_),
    .Y(_08150_));
 NAND2x1_ASAP7_75t_R _16323_ (.A(_07979_),
    .B(_08150_),
    .Y(_08151_));
 OA21x2_ASAP7_75t_R _16324_ (.A1(_07987_),
    .A2(net100),
    .B(_08151_),
    .Y(_08152_));
 BUFx10_ASAP7_75t_R _16325_ (.A(_08152_),
    .Y(_08153_));
 BUFx6f_ASAP7_75t_R _16326_ (.A(_08153_),
    .Y(_00388_));
 XNOR2x2_ASAP7_75t_R _16327_ (.A(_00438_),
    .B(_01001_),
    .Y(_08154_));
 XNOR2x1_ASAP7_75t_R _16328_ (.B(_08154_),
    .Y(_08155_),
    .A(_01033_));
 XOR2x2_ASAP7_75t_R _16329_ (.A(_08155_),
    .B(_01065_),
    .Y(_08156_));
 XOR2x1_ASAP7_75t_R _16330_ (.A(_08156_),
    .Y(_08157_),
    .B(_01097_));
 NAND2x1_ASAP7_75t_R _16331_ (.A(_07980_),
    .B(_08157_),
    .Y(_08158_));
 OA21x2_ASAP7_75t_R _16332_ (.A1(_08080_),
    .A2(net101),
    .B(_08158_),
    .Y(_08159_));
 BUFx12f_ASAP7_75t_R _16333_ (.A(_08159_),
    .Y(_00389_));
 XNOR2x2_ASAP7_75t_R _16334_ (.A(_00444_),
    .B(_01009_),
    .Y(_08160_));
 XNOR2x1_ASAP7_75t_R _16335_ (.B(_08160_),
    .Y(_08161_),
    .A(_01041_));
 XOR2x2_ASAP7_75t_R _16336_ (.A(_08161_),
    .B(_01073_),
    .Y(_08162_));
 XOR2x1_ASAP7_75t_R _16337_ (.A(_08162_),
    .Y(_08163_),
    .B(_01105_));
 NAND2x1_ASAP7_75t_R _16338_ (.A(_07979_),
    .B(_08163_),
    .Y(_08164_));
 OA21x2_ASAP7_75t_R _16339_ (.A1(_07987_),
    .A2(net109),
    .B(_08164_),
    .Y(_08165_));
 BUFx4f_ASAP7_75t_R _16340_ (.A(_08165_),
    .Y(_08166_));
 BUFx6f_ASAP7_75t_R _16341_ (.A(_08166_),
    .Y(_00393_));
 XNOR2x2_ASAP7_75t_R _16342_ (.A(_00445_),
    .B(_01010_),
    .Y(_08167_));
 XNOR2x2_ASAP7_75t_R _16343_ (.A(_01042_),
    .B(_08167_),
    .Y(_08168_));
 XOR2x2_ASAP7_75t_R _16344_ (.A(_08168_),
    .B(_01074_),
    .Y(_08169_));
 XOR2x1_ASAP7_75t_R _16345_ (.A(_08169_),
    .Y(_08170_),
    .B(_01106_));
 NAND2x1_ASAP7_75t_R _16346_ (.A(_07987_),
    .B(_08170_),
    .Y(_08171_));
 OA21x2_ASAP7_75t_R _16347_ (.A1(_07980_),
    .A2(net110),
    .B(_08171_),
    .Y(_08172_));
 BUFx10_ASAP7_75t_R _16348_ (.A(_08172_),
    .Y(_00394_));
 XNOR2x2_ASAP7_75t_R _16349_ (.A(_01011_),
    .B(_01043_),
    .Y(_08173_));
 XOR2x2_ASAP7_75t_R _16350_ (.A(_00446_),
    .B(_00987_),
    .Y(_08174_));
 XOR2x1_ASAP7_75t_R _16351_ (.A(_08173_),
    .Y(_08175_),
    .B(_08174_));
 NAND2x2_ASAP7_75t_R _16352_ (.A(_07940_),
    .B(_08175_),
    .Y(_08176_));
 BUFx12_ASAP7_75t_R _16353_ (.A(_01075_),
    .Y(_08177_));
 XNOR2x1_ASAP7_75t_R _16354_ (.B(_01107_),
    .Y(_08178_),
    .A(_08177_));
 AND2x2_ASAP7_75t_R _16355_ (.A(_07951_),
    .B(net111),
    .Y(_08179_));
 AO21x1_ASAP7_75t_R _16356_ (.A1(_08178_),
    .A2(_07940_),
    .B(_08179_),
    .Y(_08180_));
 NAND2x1_ASAP7_75t_R _16357_ (.A(_08180_),
    .B(_08176_),
    .Y(_08181_));
 OAI21x1_ASAP7_75t_R _16358_ (.A1(_08176_),
    .A2(_08178_),
    .B(_08181_),
    .Y(_15784_));
 INVx6_ASAP7_75t_R _16359_ (.A(net822),
    .Y(_15786_));
 NOR2x2_ASAP7_75t_R _16360_ (.A(net112),
    .B(_07957_),
    .Y(_08182_));
 INVx4_ASAP7_75t_R _16361_ (.A(_08182_),
    .Y(_08183_));
 XOR2x2_ASAP7_75t_R _16362_ (.A(_00447_),
    .B(_00988_),
    .Y(_08184_));
 BUFx4f_ASAP7_75t_R _16363_ (.A(_01012_),
    .Y(_08185_));
 BUFx6f_ASAP7_75t_R _16364_ (.A(_01044_),
    .Y(_08186_));
 XNOR2x2_ASAP7_75t_R _16365_ (.A(_08185_),
    .B(_08186_),
    .Y(_08187_));
 OR2x2_ASAP7_75t_R _16366_ (.A(_08184_),
    .B(_08187_),
    .Y(_08188_));
 NAND2x2_ASAP7_75t_R _16367_ (.A(_08184_),
    .B(_08187_),
    .Y(_08189_));
 BUFx6f_ASAP7_75t_R _16368_ (.A(_01076_),
    .Y(_08190_));
 BUFx4f_ASAP7_75t_R _16369_ (.A(_01108_),
    .Y(_08191_));
 XNOR2x2_ASAP7_75t_R _16370_ (.A(_08190_),
    .B(_08191_),
    .Y(_08192_));
 AO21x1_ASAP7_75t_R _16371_ (.A1(_08188_),
    .A2(_08189_),
    .B(_08192_),
    .Y(_08193_));
 INVx1_ASAP7_75t_R _16372_ (.A(_08193_),
    .Y(_08194_));
 AND3x1_ASAP7_75t_R _16373_ (.A(_08188_),
    .B(_08192_),
    .C(_08189_),
    .Y(_08195_));
 OAI21x1_ASAP7_75t_R _16374_ (.A1(_08195_),
    .A2(_08194_),
    .B(_07957_),
    .Y(_08196_));
 NAND2x2_ASAP7_75t_R _16375_ (.A(_08183_),
    .B(_08196_),
    .Y(_15789_));
 BUFx10_ASAP7_75t_R _16376_ (.A(_01077_),
    .Y(_08197_));
 BUFx6f_ASAP7_75t_R _16377_ (.A(_01109_),
    .Y(_08198_));
 XOR2x2_ASAP7_75t_R _16378_ (.A(_08197_),
    .B(_08198_),
    .Y(_08199_));
 XOR2x2_ASAP7_75t_R _16379_ (.A(_01013_),
    .B(_01045_),
    .Y(_08200_));
 XOR2x2_ASAP7_75t_R _16380_ (.A(_00448_),
    .B(_00989_),
    .Y(_08201_));
 XOR2x1_ASAP7_75t_R _16381_ (.A(_08200_),
    .Y(_08202_),
    .B(_08201_));
 NOR2x2_ASAP7_75t_R _16382_ (.A(_07951_),
    .B(_08202_),
    .Y(_08203_));
 NAND2x2_ASAP7_75t_R _16383_ (.A(_08199_),
    .B(_08203_),
    .Y(_08204_));
 NAND2x1_ASAP7_75t_R _16384_ (.A(_07951_),
    .B(net113),
    .Y(_08205_));
 OA21x2_ASAP7_75t_R _16385_ (.A1(_08199_),
    .A2(_07951_),
    .B(_08205_),
    .Y(_08206_));
 OR2x4_ASAP7_75t_R _16386_ (.A(_08206_),
    .B(_08203_),
    .Y(_08207_));
 NAND2x2_ASAP7_75t_R _16387_ (.A(_08204_),
    .B(_08207_),
    .Y(_08208_));
 CKINVDCx12_ASAP7_75t_R _16388_ (.A(_08208_),
    .Y(_15796_));
 XOR2x1_ASAP7_75t_R _16389_ (.A(_00990_),
    .Y(_08209_),
    .B(_01014_));
 XOR2x2_ASAP7_75t_R _16390_ (.A(_08209_),
    .B(_00449_),
    .Y(_08210_));
 BUFx6f_ASAP7_75t_R _16391_ (.A(_01078_),
    .Y(_08211_));
 XOR2x1_ASAP7_75t_R _16392_ (.A(_01046_),
    .Y(_08212_),
    .B(_08211_));
 XOR2x2_ASAP7_75t_R _16393_ (.A(_08210_),
    .B(_08212_),
    .Y(_08213_));
 XOR2x2_ASAP7_75t_R _16394_ (.A(_08213_),
    .B(_01110_),
    .Y(_08214_));
 AND2x6_ASAP7_75t_R _16395_ (.A(_07967_),
    .B(net114),
    .Y(_08215_));
 AO21x2_ASAP7_75t_R _16396_ (.A1(_08214_),
    .A2(_07979_),
    .B(_08215_),
    .Y(_08216_));
 BUFx6f_ASAP7_75t_R _16397_ (.A(_08216_),
    .Y(_08217_));
 BUFx6f_ASAP7_75t_R _16398_ (.A(_08217_),
    .Y(_00395_));
 XOR2x1_ASAP7_75t_R _16399_ (.A(_00991_),
    .Y(_08218_),
    .B(_01015_));
 XOR2x2_ASAP7_75t_R _16400_ (.A(_08218_),
    .B(_00450_),
    .Y(_08219_));
 BUFx3_ASAP7_75t_R _16401_ (.A(_01047_),
    .Y(_08220_));
 XOR2x2_ASAP7_75t_R _16402_ (.A(_08219_),
    .B(_08220_),
    .Y(_08221_));
 XNOR2x1_ASAP7_75t_R _16403_ (.B(_01111_),
    .Y(_08222_),
    .A(_01079_));
 XOR2x2_ASAP7_75t_R _16404_ (.A(_08221_),
    .B(_08222_),
    .Y(_08223_));
 NOR2x1_ASAP7_75t_R _16405_ (.A(net115),
    .B(_07957_),
    .Y(_08224_));
 AOI21x1_ASAP7_75t_R _16406_ (.A1(_07956_),
    .A2(_08223_),
    .B(_08224_),
    .Y(_08225_));
 BUFx6f_ASAP7_75t_R _16407_ (.A(_08225_),
    .Y(_08226_));
 BUFx6f_ASAP7_75t_R _16408_ (.A(_08226_),
    .Y(_00396_));
 XOR2x1_ASAP7_75t_R _16409_ (.A(_00992_),
    .Y(_08227_),
    .B(_01016_));
 XOR2x2_ASAP7_75t_R _16410_ (.A(_08227_),
    .B(_00451_),
    .Y(_08228_));
 XOR2x2_ASAP7_75t_R _16411_ (.A(_08228_),
    .B(_01048_),
    .Y(_08229_));
 XNOR2x1_ASAP7_75t_R _16412_ (.B(_01112_),
    .Y(_08230_),
    .A(_01080_));
 XOR2x1_ASAP7_75t_R _16413_ (.A(_08229_),
    .Y(_08231_),
    .B(_08230_));
 NOR2x1_ASAP7_75t_R _16414_ (.A(net116),
    .B(_07956_),
    .Y(_08232_));
 AO21x1_ASAP7_75t_R _16415_ (.A1(_08231_),
    .A2(_07979_),
    .B(_08232_),
    .Y(_08233_));
 BUFx10_ASAP7_75t_R _16416_ (.A(_08233_),
    .Y(_08234_));
 CKINVDCx5p33_ASAP7_75t_R _16417_ (.A(_08234_),
    .Y(_08235_));
 BUFx6f_ASAP7_75t_R _16418_ (.A(_08235_),
    .Y(_00397_));
 XOR2x1_ASAP7_75t_R _16419_ (.A(_00993_),
    .Y(_08236_),
    .B(_01018_));
 XOR2x2_ASAP7_75t_R _16420_ (.A(_08236_),
    .B(_00452_),
    .Y(_08237_));
 XOR2x1_ASAP7_75t_R _16421_ (.A(_08237_),
    .Y(_08238_),
    .B(_01050_));
 XOR2x2_ASAP7_75t_R _16422_ (.A(_08238_),
    .B(_01082_),
    .Y(_08239_));
 XNOR2x1_ASAP7_75t_R _16423_ (.B(_08239_),
    .Y(_08240_),
    .A(_01114_));
 NOR2x1_ASAP7_75t_R _16424_ (.A(net118),
    .B(_07987_),
    .Y(_08241_));
 AOI21x1_ASAP7_75t_R _16425_ (.A1(_07980_),
    .A2(_08240_),
    .B(_08241_),
    .Y(_08242_));
 BUFx10_ASAP7_75t_R _16426_ (.A(_08242_),
    .Y(_08243_));
 BUFx10_ASAP7_75t_R _16427_ (.A(_08243_),
    .Y(_00398_));
 XOR2x1_ASAP7_75t_R _16428_ (.A(_00994_),
    .Y(_08244_),
    .B(_01019_));
 XOR2x2_ASAP7_75t_R _16429_ (.A(_08244_),
    .B(_00453_),
    .Y(_08245_));
 XOR2x2_ASAP7_75t_R _16430_ (.A(_08245_),
    .B(_01051_),
    .Y(_08246_));
 XOR2x2_ASAP7_75t_R _16431_ (.A(_08246_),
    .B(_01083_),
    .Y(_08247_));
 XNOR2x1_ASAP7_75t_R _16432_ (.B(_08247_),
    .Y(_08248_),
    .A(_01115_));
 NOR2x1_ASAP7_75t_R _16433_ (.A(net119),
    .B(_07987_),
    .Y(_08249_));
 AOI21x1_ASAP7_75t_R _16434_ (.A1(_07980_),
    .A2(_08248_),
    .B(_08249_),
    .Y(_08250_));
 BUFx6f_ASAP7_75t_R _16435_ (.A(_08250_),
    .Y(_00399_));
 BUFx6f_ASAP7_75t_R _16436_ (.A(_08080_),
    .Y(_08251_));
 BUFx6f_ASAP7_75t_R _16437_ (.A(_07967_),
    .Y(_08252_));
 BUFx6f_ASAP7_75t_R _16438_ (.A(_08252_),
    .Y(_08253_));
 AND2x2_ASAP7_75t_R _16439_ (.A(_08253_),
    .B(net120),
    .Y(_08254_));
 AO21x1_ASAP7_75t_R _16440_ (.A1(_08018_),
    .A2(_08251_),
    .B(_08254_),
    .Y(_00353_));
 XOR2x2_ASAP7_75t_R _16441_ (.A(_08025_),
    .B(_00426_),
    .Y(_08255_));
 XOR2x1_ASAP7_75t_R _16442_ (.A(_08255_),
    .Y(_08256_),
    .B(_08026_));
 AND2x2_ASAP7_75t_R _16443_ (.A(_08253_),
    .B(net121),
    .Y(_08257_));
 AO21x1_ASAP7_75t_R _16444_ (.A1(_08256_),
    .A2(_08251_),
    .B(_08257_),
    .Y(_00364_));
 INVx4_ASAP7_75t_R _16445_ (.A(_08035_),
    .Y(_08258_));
 AO21x1_ASAP7_75t_R _16446_ (.A1(_08034_),
    .A2(_08258_),
    .B(_08253_),
    .Y(_08259_));
 NOR2x1_ASAP7_75t_R _16447_ (.A(_08258_),
    .B(_08034_),
    .Y(_08260_));
 OA22x2_ASAP7_75t_R _16448_ (.A1(_08251_),
    .A2(net122),
    .B1(_08259_),
    .B2(_08260_),
    .Y(_00375_));
 XNOR2x1_ASAP7_75t_R _16449_ (.B(_01020_),
    .Y(_08261_),
    .A(_00427_));
 INVx1_ASAP7_75t_R _16450_ (.A(_01052_),
    .Y(_08262_));
 XOR2x2_ASAP7_75t_R _16451_ (.A(_08261_),
    .B(_08262_),
    .Y(_08263_));
 XOR2x1_ASAP7_75t_R _16452_ (.A(_08263_),
    .Y(_08264_),
    .B(_08047_));
 BUFx4f_ASAP7_75t_R _16453_ (.A(_08080_),
    .Y(_08265_));
 AND2x2_ASAP7_75t_R _16454_ (.A(_08253_),
    .B(net123),
    .Y(_08266_));
 AO21x1_ASAP7_75t_R _16455_ (.A1(_08264_),
    .A2(_08265_),
    .B(_08266_),
    .Y(_00378_));
 BUFx4f_ASAP7_75t_R _16456_ (.A(_08252_),
    .Y(_08267_));
 AND2x2_ASAP7_75t_R _16457_ (.A(_08267_),
    .B(net124),
    .Y(_08268_));
 AO21x1_ASAP7_75t_R _16458_ (.A1(_08060_),
    .A2(_08265_),
    .B(_08268_),
    .Y(_00379_));
 AND2x2_ASAP7_75t_R _16459_ (.A(_08267_),
    .B(net125),
    .Y(_08269_));
 AO21x1_ASAP7_75t_R _16460_ (.A1(_08068_),
    .A2(_08265_),
    .B(_08269_),
    .Y(_00380_));
 AND2x2_ASAP7_75t_R _16461_ (.A(_08267_),
    .B(net126),
    .Y(_08270_));
 AO21x1_ASAP7_75t_R _16462_ (.A1(_08075_),
    .A2(_08265_),
    .B(_08270_),
    .Y(_00381_));
 AND2x2_ASAP7_75t_R _16463_ (.A(_08267_),
    .B(net127),
    .Y(_08271_));
 AO21x1_ASAP7_75t_R _16464_ (.A1(_08083_),
    .A2(_08265_),
    .B(_08271_),
    .Y(_00382_));
 XNOR2x1_ASAP7_75t_R _16465_ (.B(_01025_),
    .Y(_08272_),
    .A(_00432_));
 XNOR2x2_ASAP7_75t_R _16466_ (.A(_01057_),
    .B(_08272_),
    .Y(_08273_));
 XOR2x1_ASAP7_75t_R _16467_ (.A(_08273_),
    .Y(_08274_),
    .B(_01089_));
 AND2x2_ASAP7_75t_R _16468_ (.A(_08267_),
    .B(net129),
    .Y(_08275_));
 AO21x1_ASAP7_75t_R _16469_ (.A1(_08274_),
    .A2(_08265_),
    .B(_08275_),
    .Y(_00383_));
 XOR2x2_ASAP7_75t_R _16470_ (.A(_08098_),
    .B(_08101_),
    .Y(_08276_));
 XOR2x1_ASAP7_75t_R _16471_ (.A(_08276_),
    .Y(_08277_),
    .B(_08099_));
 AND2x2_ASAP7_75t_R _16472_ (.A(_08267_),
    .B(net130),
    .Y(_08278_));
 AO21x1_ASAP7_75t_R _16473_ (.A1(_08277_),
    .A2(_08265_),
    .B(_08278_),
    .Y(_00384_));
 INVx5_ASAP7_75t_R _16474_ (.A(_08110_),
    .Y(_08279_));
 AO21x1_ASAP7_75t_R _16475_ (.A1(_08109_),
    .A2(_08279_),
    .B(_08253_),
    .Y(_08280_));
 NOR2x1_ASAP7_75t_R _16476_ (.A(_08279_),
    .B(_08109_),
    .Y(_08281_));
 OA22x2_ASAP7_75t_R _16477_ (.A1(_08251_),
    .A2(net131),
    .B1(_08280_),
    .B2(_08281_),
    .Y(_00354_));
 AND2x2_ASAP7_75t_R _16478_ (.A(_08267_),
    .B(net132),
    .Y(_08282_));
 AO21x1_ASAP7_75t_R _16479_ (.A1(_08123_),
    .A2(_08265_),
    .B(_08282_),
    .Y(_00355_));
 AND2x2_ASAP7_75t_R _16480_ (.A(_08267_),
    .B(net133),
    .Y(_08283_));
 AO21x1_ASAP7_75t_R _16481_ (.A1(_08132_),
    .A2(_08265_),
    .B(_08283_),
    .Y(_00356_));
 AND2x2_ASAP7_75t_R _16482_ (.A(_08267_),
    .B(net134),
    .Y(_08284_));
 AO21x1_ASAP7_75t_R _16483_ (.A1(_08141_),
    .A2(_08265_),
    .B(_08284_),
    .Y(_00357_));
 BUFx4f_ASAP7_75t_R _16484_ (.A(_08080_),
    .Y(_08285_));
 AND2x2_ASAP7_75t_R _16485_ (.A(_08267_),
    .B(net135),
    .Y(_08286_));
 AO21x1_ASAP7_75t_R _16486_ (.A1(_08149_),
    .A2(_08285_),
    .B(_08286_),
    .Y(_00358_));
 BUFx3_ASAP7_75t_R _16487_ (.A(_08252_),
    .Y(_08287_));
 AND2x2_ASAP7_75t_R _16488_ (.A(_08287_),
    .B(net136),
    .Y(_08288_));
 AO21x1_ASAP7_75t_R _16489_ (.A1(_08156_),
    .A2(_08285_),
    .B(_08288_),
    .Y(_00359_));
 AND2x2_ASAP7_75t_R _16490_ (.A(_08287_),
    .B(net137),
    .Y(_08289_));
 AO21x1_ASAP7_75t_R _16491_ (.A1(_07963_),
    .A2(_08285_),
    .B(_08289_),
    .Y(_00360_));
 XOR2x2_ASAP7_75t_R _16492_ (.A(_07971_),
    .B(_00440_),
    .Y(_08290_));
 XOR2x1_ASAP7_75t_R _16493_ (.A(_08290_),
    .Y(_08291_),
    .B(_07972_));
 AND2x2_ASAP7_75t_R _16494_ (.A(_08287_),
    .B(net138),
    .Y(_08292_));
 AO21x1_ASAP7_75t_R _16495_ (.A1(_08291_),
    .A2(_08285_),
    .B(_08292_),
    .Y(_00361_));
 INVx4_ASAP7_75t_R _16496_ (.A(_08007_),
    .Y(_08293_));
 AO21x1_ASAP7_75t_R _16497_ (.A1(_08005_),
    .A2(_08293_),
    .B(_08253_),
    .Y(_08294_));
 NOR2x1_ASAP7_75t_R _16498_ (.A(_08293_),
    .B(_08005_),
    .Y(_08295_));
 OA22x2_ASAP7_75t_R _16499_ (.A1(_08251_),
    .A2(net140),
    .B1(_08294_),
    .B2(_08295_),
    .Y(_00362_));
 XNOR2x1_ASAP7_75t_R _16500_ (.B(_07942_),
    .Y(_08296_),
    .A(_00441_));
 INVx2_ASAP7_75t_R _16501_ (.A(_01037_),
    .Y(_08297_));
 XOR2x2_ASAP7_75t_R _16502_ (.A(_08296_),
    .B(_08297_),
    .Y(_08298_));
 XOR2x1_ASAP7_75t_R _16503_ (.A(_08298_),
    .Y(_08299_),
    .B(_01069_));
 AND2x2_ASAP7_75t_R _16504_ (.A(_08287_),
    .B(net141),
    .Y(_08300_));
 AO21x1_ASAP7_75t_R _16505_ (.A1(_08299_),
    .A2(_08285_),
    .B(_08300_),
    .Y(_00363_));
 AND2x2_ASAP7_75t_R _16506_ (.A(_08287_),
    .B(net142),
    .Y(_08301_));
 AO21x1_ASAP7_75t_R _16507_ (.A1(_07995_),
    .A2(_08285_),
    .B(_08301_),
    .Y(_00365_));
 AND2x2_ASAP7_75t_R _16508_ (.A(_08287_),
    .B(net143),
    .Y(_08302_));
 AO21x1_ASAP7_75t_R _16509_ (.A1(_07985_),
    .A2(_08285_),
    .B(_08302_),
    .Y(_00366_));
 AND2x2_ASAP7_75t_R _16510_ (.A(_08287_),
    .B(net144),
    .Y(_08303_));
 AO21x1_ASAP7_75t_R _16511_ (.A1(_08162_),
    .A2(_08285_),
    .B(_08303_),
    .Y(_00367_));
 AND2x2_ASAP7_75t_R _16512_ (.A(_08287_),
    .B(net145),
    .Y(_08304_));
 AO21x1_ASAP7_75t_R _16513_ (.A1(_08169_),
    .A2(_08285_),
    .B(_08304_),
    .Y(_00368_));
 XOR2x1_ASAP7_75t_R _16514_ (.A(_08173_),
    .Y(_08305_),
    .B(_08177_));
 XOR2x1_ASAP7_75t_R _16515_ (.A(_08305_),
    .Y(_08306_),
    .B(_08174_));
 AND2x2_ASAP7_75t_R _16516_ (.A(_08287_),
    .B(net146),
    .Y(_08307_));
 AO21x1_ASAP7_75t_R _16517_ (.A1(_08306_),
    .A2(_08285_),
    .B(_08307_),
    .Y(_00369_));
 XOR2x1_ASAP7_75t_R _16518_ (.A(_08186_),
    .Y(_08308_),
    .B(_08190_));
 XOR2x1_ASAP7_75t_R _16519_ (.A(_00988_),
    .Y(_08309_),
    .B(_08185_));
 XOR2x2_ASAP7_75t_R _16520_ (.A(_08309_),
    .B(_00447_),
    .Y(_08310_));
 XNOR2x1_ASAP7_75t_R _16521_ (.B(_08310_),
    .Y(_08311_),
    .A(_08308_));
 BUFx6f_ASAP7_75t_R _16522_ (.A(_08080_),
    .Y(_08312_));
 AND2x2_ASAP7_75t_R _16523_ (.A(_08287_),
    .B(net147),
    .Y(_08313_));
 AO21x1_ASAP7_75t_R _16524_ (.A1(_08311_),
    .A2(_08312_),
    .B(_08313_),
    .Y(_00370_));
 INVx6_ASAP7_75t_R _16525_ (.A(_08197_),
    .Y(_08314_));
 XOR2x1_ASAP7_75t_R _16526_ (.A(_08200_),
    .Y(_08315_),
    .B(_08314_));
 XOR2x1_ASAP7_75t_R _16527_ (.A(_08315_),
    .Y(_08316_),
    .B(_08201_));
 BUFx6f_ASAP7_75t_R _16528_ (.A(_08252_),
    .Y(_08317_));
 AND2x2_ASAP7_75t_R _16529_ (.A(_08317_),
    .B(net148),
    .Y(_08318_));
 AO21x1_ASAP7_75t_R _16530_ (.A1(_08316_),
    .A2(_08312_),
    .B(_08318_),
    .Y(_00371_));
 BUFx10_ASAP7_75t_R _16531_ (.A(_08252_),
    .Y(_08319_));
 BUFx6f_ASAP7_75t_R _16532_ (.A(_08319_),
    .Y(_08320_));
 BUFx6f_ASAP7_75t_R _16533_ (.A(_08252_),
    .Y(_08321_));
 NOR2x1_ASAP7_75t_R _16534_ (.A(_08321_),
    .B(_08213_),
    .Y(_08322_));
 AO21x1_ASAP7_75t_R _16535_ (.A1(_08320_),
    .A2(net149),
    .B(_08322_),
    .Y(_00372_));
 INVx2_ASAP7_75t_R _16536_ (.A(_01079_),
    .Y(_08323_));
 XOR2x1_ASAP7_75t_R _16537_ (.A(_08221_),
    .Y(_08324_),
    .B(_08323_));
 AND2x2_ASAP7_75t_R _16538_ (.A(_08317_),
    .B(net151),
    .Y(_08325_));
 AO21x1_ASAP7_75t_R _16539_ (.A1(_08324_),
    .A2(_08312_),
    .B(_08325_),
    .Y(_00373_));
 INVx1_ASAP7_75t_R _16540_ (.A(_01080_),
    .Y(_08326_));
 XOR2x1_ASAP7_75t_R _16541_ (.A(_08229_),
    .Y(_08327_),
    .B(_08326_));
 AND2x2_ASAP7_75t_R _16542_ (.A(_08317_),
    .B(net152),
    .Y(_08328_));
 AO21x1_ASAP7_75t_R _16543_ (.A1(_08327_),
    .A2(_08312_),
    .B(_08328_),
    .Y(_00374_));
 NOR2x1_ASAP7_75t_R _16544_ (.A(_08321_),
    .B(_08239_),
    .Y(_08329_));
 AO21x1_ASAP7_75t_R _16545_ (.A1(_08320_),
    .A2(net153),
    .B(_08329_),
    .Y(_00376_));
 BUFx10_ASAP7_75t_R _16546_ (.A(_08319_),
    .Y(_08330_));
 NOR2x1_ASAP7_75t_R _16547_ (.A(_08330_),
    .B(_08247_),
    .Y(_08331_));
 AO21x1_ASAP7_75t_R _16548_ (.A1(_08320_),
    .A2(net154),
    .B(_08331_),
    .Y(_00377_));
 XOR2x1_ASAP7_75t_R _16549_ (.A(net861),
    .Y(_08332_),
    .B(_08016_));
 AND2x2_ASAP7_75t_R _16550_ (.A(_08317_),
    .B(net155),
    .Y(_08333_));
 AO21x1_ASAP7_75t_R _16551_ (.A1(_08332_),
    .A2(_08312_),
    .B(_08333_),
    .Y(_00321_));
 NOR2x1_ASAP7_75t_R _16552_ (.A(_08330_),
    .B(_08255_),
    .Y(_08334_));
 AO21x1_ASAP7_75t_R _16553_ (.A1(_08320_),
    .A2(net156),
    .B(_08334_),
    .Y(_00332_));
 OA21x2_ASAP7_75t_R _16554_ (.A1(_08251_),
    .A2(net157),
    .B(_08041_),
    .Y(_00343_));
 NOR2x1_ASAP7_75t_R _16555_ (.A(_08330_),
    .B(_08263_),
    .Y(_08335_));
 AO21x1_ASAP7_75t_R _16556_ (.A1(_08320_),
    .A2(net158),
    .B(_08335_),
    .Y(_00346_));
 NOR2x1_ASAP7_75t_R _16557_ (.A(_08330_),
    .B(_08059_),
    .Y(_08336_));
 AO21x1_ASAP7_75t_R _16558_ (.A1(_08320_),
    .A2(net159),
    .B(_08336_),
    .Y(_00347_));
 NOR2x1_ASAP7_75t_R _16559_ (.A(_08330_),
    .B(_08067_),
    .Y(_08337_));
 AO21x1_ASAP7_75t_R _16560_ (.A1(_08320_),
    .A2(net160),
    .B(_08337_),
    .Y(_00348_));
 NOR2x1_ASAP7_75t_R _16561_ (.A(_08330_),
    .B(_08074_),
    .Y(_08338_));
 AO21x1_ASAP7_75t_R _16562_ (.A1(_08320_),
    .A2(net162),
    .B(_08338_),
    .Y(_00349_));
 NOR2x1_ASAP7_75t_R _16563_ (.A(_08330_),
    .B(_08082_),
    .Y(_08339_));
 AO21x1_ASAP7_75t_R _16564_ (.A1(_08320_),
    .A2(net163),
    .B(_08339_),
    .Y(_00350_));
 BUFx6f_ASAP7_75t_R _16565_ (.A(_08252_),
    .Y(_08340_));
 BUFx6f_ASAP7_75t_R _16566_ (.A(_08340_),
    .Y(_08341_));
 NOR2x1_ASAP7_75t_R _16567_ (.A(_08330_),
    .B(_08273_),
    .Y(_08342_));
 AO21x1_ASAP7_75t_R _16568_ (.A1(_08341_),
    .A2(net164),
    .B(_08342_),
    .Y(_00351_));
 NOR2x1_ASAP7_75t_R _16569_ (.A(_08330_),
    .B(_08276_),
    .Y(_08343_));
 AO21x1_ASAP7_75t_R _16570_ (.A1(_08341_),
    .A2(net165),
    .B(_08343_),
    .Y(_00352_));
 OA21x2_ASAP7_75t_R _16571_ (.A1(_08251_),
    .A2(net166),
    .B(_08117_),
    .Y(_00322_));
 NOR2x1_ASAP7_75t_R _16572_ (.A(_08330_),
    .B(_08122_),
    .Y(_08344_));
 AO21x1_ASAP7_75t_R _16573_ (.A1(_08341_),
    .A2(net167),
    .B(_08344_),
    .Y(_00323_));
 BUFx6f_ASAP7_75t_R _16574_ (.A(_08319_),
    .Y(_08345_));
 NOR2x1_ASAP7_75t_R _16575_ (.A(_08345_),
    .B(_08131_),
    .Y(_08346_));
 AO21x1_ASAP7_75t_R _16576_ (.A1(_08341_),
    .A2(net168),
    .B(_08346_),
    .Y(_00324_));
 NOR2x1_ASAP7_75t_R _16577_ (.A(_08345_),
    .B(_08140_),
    .Y(_08347_));
 AO21x1_ASAP7_75t_R _16578_ (.A1(_08341_),
    .A2(net169),
    .B(_08347_),
    .Y(_00325_));
 NOR2x1_ASAP7_75t_R _16579_ (.A(_08345_),
    .B(_08148_),
    .Y(_08348_));
 AO21x1_ASAP7_75t_R _16580_ (.A1(_08341_),
    .A2(net170),
    .B(_08348_),
    .Y(_00326_));
 NOR2x1_ASAP7_75t_R _16581_ (.A(_08345_),
    .B(_08155_),
    .Y(_08349_));
 AO21x1_ASAP7_75t_R _16582_ (.A1(_08341_),
    .A2(net171),
    .B(_08349_),
    .Y(_00327_));
 XOR2x1_ASAP7_75t_R _16583_ (.A(_07959_),
    .Y(_08350_),
    .B(_07960_));
 AND2x2_ASAP7_75t_R _16584_ (.A(_08317_),
    .B(net173),
    .Y(_08351_));
 AO21x1_ASAP7_75t_R _16585_ (.A1(_08350_),
    .A2(_08312_),
    .B(_08351_),
    .Y(_00328_));
 NOR2x1_ASAP7_75t_R _16586_ (.A(_08345_),
    .B(_08290_),
    .Y(_08352_));
 AO21x1_ASAP7_75t_R _16587_ (.A1(_08341_),
    .A2(net174),
    .B(_08352_),
    .Y(_00329_));
 OA21x2_ASAP7_75t_R _16588_ (.A1(_08251_),
    .A2(net175),
    .B(_08006_),
    .Y(_00330_));
 NOR2x1_ASAP7_75t_R _16589_ (.A(_08345_),
    .B(_08298_),
    .Y(_08353_));
 AO21x1_ASAP7_75t_R _16590_ (.A1(_08341_),
    .A2(net176),
    .B(_08353_),
    .Y(_00331_));
 NOR2x1_ASAP7_75t_R _16591_ (.A(_08345_),
    .B(_07993_),
    .Y(_08354_));
 AO21x1_ASAP7_75t_R _16592_ (.A1(_08341_),
    .A2(net177),
    .B(_08354_),
    .Y(_00333_));
 BUFx10_ASAP7_75t_R _16593_ (.A(_08340_),
    .Y(_08355_));
 NOR2x1_ASAP7_75t_R _16594_ (.A(_08345_),
    .B(_07983_),
    .Y(_08356_));
 AO21x1_ASAP7_75t_R _16595_ (.A1(_08355_),
    .A2(net178),
    .B(_08356_),
    .Y(_00334_));
 NOR2x1_ASAP7_75t_R _16596_ (.A(_08345_),
    .B(_08161_),
    .Y(_08357_));
 AO21x1_ASAP7_75t_R _16597_ (.A1(_08355_),
    .A2(net179),
    .B(_08357_),
    .Y(_00335_));
 NOR2x1_ASAP7_75t_R _16598_ (.A(_08345_),
    .B(_08168_),
    .Y(_08358_));
 AO21x1_ASAP7_75t_R _16599_ (.A1(_08355_),
    .A2(net180),
    .B(_08358_),
    .Y(_00336_));
 OA21x2_ASAP7_75t_R _16600_ (.A1(_08251_),
    .A2(net181),
    .B(_08176_),
    .Y(_00337_));
 AOI21x1_ASAP7_75t_R _16601_ (.A1(_08189_),
    .A2(_08188_),
    .B(_08321_),
    .Y(_08359_));
 AO21x1_ASAP7_75t_R _16602_ (.A1(_08355_),
    .A2(net182),
    .B(_08359_),
    .Y(_00338_));
 BUFx6f_ASAP7_75t_R _16603_ (.A(_08253_),
    .Y(_08360_));
 INVx2_ASAP7_75t_R _16604_ (.A(net184),
    .Y(_08361_));
 AOI21x1_ASAP7_75t_R _16605_ (.A1(_08360_),
    .A2(_08361_),
    .B(_08203_),
    .Y(_00339_));
 XOR2x1_ASAP7_75t_R _16606_ (.A(_08210_),
    .Y(_08362_),
    .B(_01046_));
 AND2x2_ASAP7_75t_R _16607_ (.A(_08317_),
    .B(net185),
    .Y(_08363_));
 AO21x1_ASAP7_75t_R _16608_ (.A1(_08362_),
    .A2(_08312_),
    .B(_08363_),
    .Y(_00340_));
 AND2x2_ASAP7_75t_R _16609_ (.A(_08317_),
    .B(net186),
    .Y(_08364_));
 AO21x1_ASAP7_75t_R _16610_ (.A1(_08221_),
    .A2(_08312_),
    .B(_08364_),
    .Y(_00341_));
 AND2x2_ASAP7_75t_R _16611_ (.A(_08317_),
    .B(net187),
    .Y(_08365_));
 AO21x1_ASAP7_75t_R _16612_ (.A1(_08229_),
    .A2(_08312_),
    .B(_08365_),
    .Y(_00342_));
 AND2x2_ASAP7_75t_R _16613_ (.A(_08317_),
    .B(net188),
    .Y(_08366_));
 AO21x1_ASAP7_75t_R _16614_ (.A1(_08238_),
    .A2(_08312_),
    .B(_08366_),
    .Y(_00344_));
 BUFx6f_ASAP7_75t_R _16615_ (.A(_08080_),
    .Y(_08367_));
 AND2x2_ASAP7_75t_R _16616_ (.A(_08317_),
    .B(net189),
    .Y(_08368_));
 AO21x1_ASAP7_75t_R _16617_ (.A1(_08246_),
    .A2(_08367_),
    .B(_08368_),
    .Y(_00345_));
 BUFx10_ASAP7_75t_R _16618_ (.A(_08319_),
    .Y(_08369_));
 NOR2x1_ASAP7_75t_R _16619_ (.A(_08369_),
    .B(net862),
    .Y(_08370_));
 AO21x1_ASAP7_75t_R _16620_ (.A1(_08355_),
    .A2(net190),
    .B(_08370_),
    .Y(_00289_));
 XOR2x1_ASAP7_75t_R _16621_ (.A(_00426_),
    .Y(_08371_),
    .B(_08023_));
 AND2x2_ASAP7_75t_R _16622_ (.A(_08340_),
    .B(net191),
    .Y(_08372_));
 AO21x1_ASAP7_75t_R _16623_ (.A1(_08371_),
    .A2(_08367_),
    .B(_08372_),
    .Y(_00300_));
 AND2x2_ASAP7_75t_R _16624_ (.A(_08340_),
    .B(net192),
    .Y(_08373_));
 AO21x1_ASAP7_75t_R _16625_ (.A1(_08032_),
    .A2(_08367_),
    .B(_08373_),
    .Y(_00311_));
 NOR2x1_ASAP7_75t_R _16626_ (.A(_08369_),
    .B(_08261_),
    .Y(_08374_));
 AO21x1_ASAP7_75t_R _16627_ (.A1(_08355_),
    .A2(net193),
    .B(_08374_),
    .Y(_00314_));
 NOR2x1_ASAP7_75t_R _16628_ (.A(_08369_),
    .B(_08057_),
    .Y(_08375_));
 AO21x1_ASAP7_75t_R _16629_ (.A1(_08355_),
    .A2(net31),
    .B(_08375_),
    .Y(_00315_));
 NOR2x1_ASAP7_75t_R _16630_ (.A(_08369_),
    .B(_08065_),
    .Y(_08376_));
 AO21x1_ASAP7_75t_R _16631_ (.A1(_08355_),
    .A2(net42),
    .B(_08376_),
    .Y(_00316_));
 NOR2x1_ASAP7_75t_R _16632_ (.A(_08369_),
    .B(_08073_),
    .Y(_08377_));
 AO21x1_ASAP7_75t_R _16633_ (.A1(_08355_),
    .A2(net45),
    .B(_08377_),
    .Y(_00317_));
 NOR2x1_ASAP7_75t_R _16634_ (.A(_08369_),
    .B(_08081_),
    .Y(_08378_));
 AO21x1_ASAP7_75t_R _16635_ (.A1(_08355_),
    .A2(net47),
    .B(_08378_),
    .Y(_00318_));
 BUFx10_ASAP7_75t_R _16636_ (.A(_08252_),
    .Y(_08379_));
 BUFx4f_ASAP7_75t_R _16637_ (.A(_08379_),
    .Y(_08380_));
 NOR2x1_ASAP7_75t_R _16638_ (.A(_08369_),
    .B(_08272_),
    .Y(_08381_));
 AO21x1_ASAP7_75t_R _16639_ (.A1(_08380_),
    .A2(net51),
    .B(_08381_),
    .Y(_00319_));
 XOR2x1_ASAP7_75t_R _16640_ (.A(_00433_),
    .Y(_08382_),
    .B(_08101_));
 AND2x2_ASAP7_75t_R _16641_ (.A(_08340_),
    .B(net64),
    .Y(_08383_));
 AO21x1_ASAP7_75t_R _16642_ (.A1(_08382_),
    .A2(_08367_),
    .B(_08383_),
    .Y(_00320_));
 AND2x2_ASAP7_75t_R _16643_ (.A(_08340_),
    .B(net68),
    .Y(_08384_));
 AO21x1_ASAP7_75t_R _16644_ (.A1(_08107_),
    .A2(_08367_),
    .B(_08384_),
    .Y(_00290_));
 NOR2x1_ASAP7_75t_R _16645_ (.A(_08369_),
    .B(_08120_),
    .Y(_08385_));
 AO21x1_ASAP7_75t_R _16646_ (.A1(_08380_),
    .A2(net75),
    .B(_08385_),
    .Y(_00291_));
 NOR2x1_ASAP7_75t_R _16647_ (.A(_08369_),
    .B(_08129_),
    .Y(_08386_));
 AO21x1_ASAP7_75t_R _16648_ (.A1(_08380_),
    .A2(net76),
    .B(_08386_),
    .Y(_00292_));
 NOR2x1_ASAP7_75t_R _16649_ (.A(_08369_),
    .B(_08138_),
    .Y(_08387_));
 AO21x1_ASAP7_75t_R _16650_ (.A1(_08380_),
    .A2(net77),
    .B(_08387_),
    .Y(_00293_));
 BUFx6f_ASAP7_75t_R _16651_ (.A(_08319_),
    .Y(_08388_));
 NOR2x1_ASAP7_75t_R _16652_ (.A(_08388_),
    .B(_08146_),
    .Y(_08389_));
 AO21x1_ASAP7_75t_R _16653_ (.A1(_08380_),
    .A2(net79),
    .B(_08389_),
    .Y(_00294_));
 NOR2x1_ASAP7_75t_R _16654_ (.A(_08388_),
    .B(_08154_),
    .Y(_08390_));
 AO21x1_ASAP7_75t_R _16655_ (.A1(_08380_),
    .A2(net80),
    .B(_08390_),
    .Y(_00295_));
 NOR2x1_ASAP7_75t_R _16656_ (.A(_08388_),
    .B(_07959_),
    .Y(_08391_));
 AO21x1_ASAP7_75t_R _16657_ (.A1(_08380_),
    .A2(net81),
    .B(_08391_),
    .Y(_00296_));
 XOR2x1_ASAP7_75t_R _16658_ (.A(_00440_),
    .Y(_08392_),
    .B(_07969_));
 AND2x2_ASAP7_75t_R _16659_ (.A(_08340_),
    .B(net82),
    .Y(_08393_));
 AO21x1_ASAP7_75t_R _16660_ (.A1(_08392_),
    .A2(_08367_),
    .B(_08393_),
    .Y(_00297_));
 AND2x2_ASAP7_75t_R _16661_ (.A(_08340_),
    .B(net83),
    .Y(_08394_));
 AO21x1_ASAP7_75t_R _16662_ (.A1(_08003_),
    .A2(_08367_),
    .B(_08394_),
    .Y(_00298_));
 NOR2x1_ASAP7_75t_R _16663_ (.A(_08388_),
    .B(_08296_),
    .Y(_08395_));
 AO21x1_ASAP7_75t_R _16664_ (.A1(_08380_),
    .A2(net84),
    .B(_08395_),
    .Y(_00299_));
 NOR2x1_ASAP7_75t_R _16665_ (.A(_08388_),
    .B(_07991_),
    .Y(_08396_));
 AO21x1_ASAP7_75t_R _16666_ (.A1(_08380_),
    .A2(net85),
    .B(_08396_),
    .Y(_00301_));
 NOR2x1_ASAP7_75t_R _16667_ (.A(_08388_),
    .B(_07981_),
    .Y(_08397_));
 AO21x1_ASAP7_75t_R _16668_ (.A1(_08380_),
    .A2(net86),
    .B(_08397_),
    .Y(_00302_));
 BUFx4f_ASAP7_75t_R _16669_ (.A(_08379_),
    .Y(_08398_));
 NOR2x1_ASAP7_75t_R _16670_ (.A(_08388_),
    .B(_08160_),
    .Y(_08399_));
 AO21x1_ASAP7_75t_R _16671_ (.A1(_08398_),
    .A2(net87),
    .B(_08399_),
    .Y(_00303_));
 NOR2x1_ASAP7_75t_R _16672_ (.A(_08388_),
    .B(_08167_),
    .Y(_08400_));
 AO21x1_ASAP7_75t_R _16673_ (.A1(_08398_),
    .A2(net88),
    .B(_08400_),
    .Y(_00304_));
 INVx3_ASAP7_75t_R _16674_ (.A(_01011_),
    .Y(_08401_));
 XOR2x1_ASAP7_75t_R _16675_ (.A(_08174_),
    .Y(_08402_),
    .B(_08401_));
 AND2x2_ASAP7_75t_R _16676_ (.A(_08340_),
    .B(net90),
    .Y(_08403_));
 AO21x1_ASAP7_75t_R _16677_ (.A1(_08402_),
    .A2(_08367_),
    .B(_08403_),
    .Y(_00305_));
 NOR2x1_ASAP7_75t_R _16678_ (.A(_08388_),
    .B(_08310_),
    .Y(_08404_));
 AO21x1_ASAP7_75t_R _16679_ (.A1(_08398_),
    .A2(net91),
    .B(_08404_),
    .Y(_00306_));
 INVx4_ASAP7_75t_R _16680_ (.A(_01013_),
    .Y(_08405_));
 XOR2x1_ASAP7_75t_R _16681_ (.A(_08201_),
    .Y(_08406_),
    .B(_08405_));
 AND2x2_ASAP7_75t_R _16682_ (.A(_08340_),
    .B(net92),
    .Y(_08407_));
 AO21x1_ASAP7_75t_R _16683_ (.A1(_08406_),
    .A2(_08367_),
    .B(_08407_),
    .Y(_00307_));
 NOR2x1_ASAP7_75t_R _16684_ (.A(_08388_),
    .B(_08210_),
    .Y(_08408_));
 AO21x1_ASAP7_75t_R _16685_ (.A1(_08398_),
    .A2(net93),
    .B(_08408_),
    .Y(_00308_));
 BUFx6f_ASAP7_75t_R _16686_ (.A(_08319_),
    .Y(_08409_));
 NOR2x1_ASAP7_75t_R _16687_ (.A(_08409_),
    .B(_08219_),
    .Y(_08410_));
 AO21x1_ASAP7_75t_R _16688_ (.A1(_08398_),
    .A2(net94),
    .B(_08410_),
    .Y(_00309_));
 NOR2x1_ASAP7_75t_R _16689_ (.A(_08409_),
    .B(_08228_),
    .Y(_08411_));
 AO21x1_ASAP7_75t_R _16690_ (.A1(_08398_),
    .A2(net95),
    .B(_08411_),
    .Y(_00310_));
 NOR2x1_ASAP7_75t_R _16691_ (.A(_08409_),
    .B(_08237_),
    .Y(_08412_));
 AO21x1_ASAP7_75t_R _16692_ (.A1(_08398_),
    .A2(net96),
    .B(_08412_),
    .Y(_00312_));
 NOR2x1_ASAP7_75t_R _16693_ (.A(_08409_),
    .B(_08245_),
    .Y(_08413_));
 AO21x1_ASAP7_75t_R _16694_ (.A1(_08398_),
    .A2(net97),
    .B(_08413_),
    .Y(_00313_));
 NOR2x1_ASAP7_75t_R _16695_ (.A(_08009_),
    .B(_08006_),
    .Y(_08414_));
 AOI21x1_ASAP7_75t_R _16696_ (.A1(_08006_),
    .A2(_08011_),
    .B(_08414_),
    .Y(_08415_));
 BUFx10_ASAP7_75t_R _16697_ (.A(_08415_),
    .Y(_15740_));
 INVx6_ASAP7_75t_R _16698_ (.A(net838),
    .Y(_15730_));
 INVx2_ASAP7_75t_R _16699_ (.A(_07999_),
    .Y(_08416_));
 BUFx6f_ASAP7_75t_R _16700_ (.A(_08416_),
    .Y(_08417_));
 BUFx6f_ASAP7_75t_R _16701_ (.A(_08417_),
    .Y(_08418_));
 NOR2x2_ASAP7_75t_R _16702_ (.A(_08014_),
    .B(net802),
    .Y(_08419_));
 INVx4_ASAP7_75t_R _16703_ (.A(_08419_),
    .Y(_08420_));
 BUFx4f_ASAP7_75t_R _16704_ (.A(_07954_),
    .Y(_08421_));
 NAND2x2_ASAP7_75t_R _16705_ (.A(net803),
    .B(_15729_),
    .Y(_08422_));
 AND3x1_ASAP7_75t_R _16706_ (.A(_08420_),
    .B(_08421_),
    .C(_08422_),
    .Y(_08423_));
 NOR2x1_ASAP7_75t_R _16707_ (.A(_08418_),
    .B(_08423_),
    .Y(_08424_));
 NAND2x2_ASAP7_75t_R _16708_ (.A(net803),
    .B(_15735_),
    .Y(_08425_));
 NOR2x2_ASAP7_75t_R _16709_ (.A(_08415_),
    .B(net839),
    .Y(_08426_));
 NOR2x2_ASAP7_75t_R _16710_ (.A(_07955_),
    .B(_08426_),
    .Y(_08427_));
 NAND2x1_ASAP7_75t_R _16711_ (.A(_08425_),
    .B(_08427_),
    .Y(_08428_));
 BUFx6f_ASAP7_75t_R _16712_ (.A(_00457_),
    .Y(_08429_));
 BUFx12f_ASAP7_75t_R _16713_ (.A(_08013_),
    .Y(_08430_));
 NOR2x2_ASAP7_75t_R _16714_ (.A(_08429_),
    .B(_08430_),
    .Y(_08431_));
 INVx2_ASAP7_75t_R _16715_ (.A(_08431_),
    .Y(_08432_));
 NAND2x2_ASAP7_75t_R _16716_ (.A(_08013_),
    .B(net480),
    .Y(_08433_));
 INVx4_ASAP7_75t_R _16717_ (.A(_08433_),
    .Y(_08434_));
 NOR2x2_ASAP7_75t_R _16718_ (.A(_07955_),
    .B(_08434_),
    .Y(_08435_));
 INVx1_ASAP7_75t_R _16719_ (.A(_00454_),
    .Y(_08436_));
 NOR2x2_ASAP7_75t_R _16720_ (.A(_08436_),
    .B(_15740_),
    .Y(_08437_));
 INVx1_ASAP7_75t_R _16721_ (.A(_00455_),
    .Y(_08438_));
 NOR2x2_ASAP7_75t_R _16722_ (.A(_08438_),
    .B(_08430_),
    .Y(_08439_));
 BUFx10_ASAP7_75t_R _16723_ (.A(_07954_),
    .Y(_08440_));
 BUFx4f_ASAP7_75t_R _16724_ (.A(_08440_),
    .Y(_08441_));
 OA21x2_ASAP7_75t_R _16725_ (.A1(_08437_),
    .A2(_08439_),
    .B(_08441_),
    .Y(_08442_));
 BUFx6f_ASAP7_75t_R _16726_ (.A(_08000_),
    .Y(_08443_));
 AOI211x1_ASAP7_75t_R _16727_ (.A1(_08432_),
    .A2(_08435_),
    .B(_08442_),
    .C(_08443_),
    .Y(_08444_));
 BUFx6f_ASAP7_75t_R _16728_ (.A(_08166_),
    .Y(_08445_));
 AOI211x1_ASAP7_75t_R _16729_ (.A1(_08424_),
    .A2(_08428_),
    .B(_08444_),
    .C(_08445_),
    .Y(_08446_));
 INVx5_ASAP7_75t_R _16730_ (.A(_08166_),
    .Y(_08447_));
 BUFx10_ASAP7_75t_R _16731_ (.A(_08447_),
    .Y(_08448_));
 BUFx10_ASAP7_75t_R _16732_ (.A(_07953_),
    .Y(_08449_));
 INVx3_ASAP7_75t_R _16733_ (.A(_01122_),
    .Y(_08450_));
 NOR2x2_ASAP7_75t_R _16734_ (.A(_08450_),
    .B(_08013_),
    .Y(_08451_));
 NOR2x2_ASAP7_75t_R _16735_ (.A(_08449_),
    .B(_08451_),
    .Y(_08452_));
 BUFx6f_ASAP7_75t_R _16736_ (.A(_08449_),
    .Y(_08453_));
 INVx3_ASAP7_75t_R _16737_ (.A(_00458_),
    .Y(_08454_));
 NAND2x2_ASAP7_75t_R _16738_ (.A(_08454_),
    .B(_08415_),
    .Y(_08455_));
 NAND2x2_ASAP7_75t_R _16739_ (.A(_08453_),
    .B(_08455_),
    .Y(_08456_));
 NAND2x2_ASAP7_75t_R _16740_ (.A(_08430_),
    .B(_15732_),
    .Y(_08457_));
 INVx1_ASAP7_75t_R _16741_ (.A(_08457_),
    .Y(_08458_));
 NOR2x1_ASAP7_75t_R _16742_ (.A(_08456_),
    .B(_08458_),
    .Y(_08459_));
 AO21x1_ASAP7_75t_R _16743_ (.A1(_08433_),
    .A2(_08452_),
    .B(_08459_),
    .Y(_08460_));
 NAND2x2_ASAP7_75t_R _16744_ (.A(_08415_),
    .B(_15732_),
    .Y(_08461_));
 AND2x2_ASAP7_75t_R _16745_ (.A(_08461_),
    .B(_08453_),
    .Y(_08462_));
 NAND2x2_ASAP7_75t_R _16746_ (.A(_08014_),
    .B(_01123_),
    .Y(_08463_));
 AND3x1_ASAP7_75t_R _16747_ (.A(_08455_),
    .B(_07955_),
    .C(_08463_),
    .Y(_08464_));
 BUFx6f_ASAP7_75t_R _16748_ (.A(_08416_),
    .Y(_08465_));
 BUFx6f_ASAP7_75t_R _16749_ (.A(_08465_),
    .Y(_08466_));
 OA21x2_ASAP7_75t_R _16750_ (.A1(_08462_),
    .A2(_08464_),
    .B(_08466_),
    .Y(_08467_));
 AOI21x1_ASAP7_75t_R _16751_ (.A1(_00391_),
    .A2(_08460_),
    .B(_08467_),
    .Y(_08468_));
 OAI21x1_ASAP7_75t_R _16752_ (.A1(_08448_),
    .A2(_08468_),
    .B(_00392_),
    .Y(_08469_));
 NOR2x1_ASAP7_75t_R _16753_ (.A(_08446_),
    .B(_08469_),
    .Y(_08470_));
 NOR2x2_ASAP7_75t_R _16754_ (.A(_08449_),
    .B(_08434_),
    .Y(_08471_));
 NOR2x1_ASAP7_75t_R _16755_ (.A(_00455_),
    .B(_08430_),
    .Y(_08472_));
 INVx1_ASAP7_75t_R _16756_ (.A(_08472_),
    .Y(_08473_));
 BUFx6f_ASAP7_75t_R _16757_ (.A(_08453_),
    .Y(_08474_));
 NAND2x2_ASAP7_75t_R _16758_ (.A(_00454_),
    .B(_08415_),
    .Y(_08475_));
 INVx1_ASAP7_75t_R _16759_ (.A(_08475_),
    .Y(_08476_));
 AOI22x1_ASAP7_75t_R _16760_ (.A1(_08471_),
    .A2(_08473_),
    .B1(_08474_),
    .B2(_08476_),
    .Y(_08477_));
 BUFx6f_ASAP7_75t_R _16761_ (.A(_08000_),
    .Y(_08478_));
 NAND2x2_ASAP7_75t_R _16762_ (.A(_08014_),
    .B(_00455_),
    .Y(_08479_));
 NOR2x2_ASAP7_75t_R _16763_ (.A(_08440_),
    .B(_08479_),
    .Y(_08480_));
 NOR2x2_ASAP7_75t_R _16764_ (.A(_08478_),
    .B(_08480_),
    .Y(_08481_));
 BUFx4f_ASAP7_75t_R _16765_ (.A(_08453_),
    .Y(_08482_));
 INVx2_ASAP7_75t_R _16766_ (.A(net480),
    .Y(_08483_));
 NOR2x2_ASAP7_75t_R _16767_ (.A(_08483_),
    .B(_08013_),
    .Y(_08484_));
 NOR2x2_ASAP7_75t_R _16768_ (.A(_08449_),
    .B(_08484_),
    .Y(_08485_));
 AO21x1_ASAP7_75t_R _16769_ (.A1(_08482_),
    .A2(_08434_),
    .B(_08485_),
    .Y(_08486_));
 NOR2x1_ASAP7_75t_R _16770_ (.A(_07954_),
    .B(_15729_),
    .Y(_08487_));
 AND2x2_ASAP7_75t_R _16771_ (.A(_08487_),
    .B(_15740_),
    .Y(_08488_));
 OA21x2_ASAP7_75t_R _16772_ (.A1(_08486_),
    .A2(_08488_),
    .B(_08443_),
    .Y(_08489_));
 AOI211x1_ASAP7_75t_R _16773_ (.A1(_08477_),
    .A2(_08481_),
    .B(_08489_),
    .C(_00393_),
    .Y(_08490_));
 AO21x2_ASAP7_75t_R _16774_ (.A1(_15732_),
    .A2(_08415_),
    .B(_08449_),
    .Y(_08491_));
 INVx1_ASAP7_75t_R _16775_ (.A(_08491_),
    .Y(_08492_));
 INVx2_ASAP7_75t_R _16776_ (.A(_08429_),
    .Y(_08493_));
 NAND2x2_ASAP7_75t_R _16777_ (.A(_08493_),
    .B(_08430_),
    .Y(_08494_));
 AO21x1_ASAP7_75t_R _16778_ (.A1(_08487_),
    .A2(_15740_),
    .B(_08478_),
    .Y(_08495_));
 INVx3_ASAP7_75t_R _16779_ (.A(_01125_),
    .Y(_08496_));
 NAND2x2_ASAP7_75t_R _16780_ (.A(_08496_),
    .B(_08014_),
    .Y(_08497_));
 NOR2x2_ASAP7_75t_R _16781_ (.A(_08440_),
    .B(_08497_),
    .Y(_08498_));
 AOI211x1_ASAP7_75t_R _16782_ (.A1(_08492_),
    .A2(_08494_),
    .B(_08495_),
    .C(_08498_),
    .Y(_08499_));
 NOR2x2_ASAP7_75t_R _16783_ (.A(_08450_),
    .B(_15740_),
    .Y(_08500_));
 OA21x2_ASAP7_75t_R _16784_ (.A1(_08491_),
    .A2(_08500_),
    .B(_08001_),
    .Y(_08501_));
 NAND2x2_ASAP7_75t_R _16785_ (.A(_08430_),
    .B(net805),
    .Y(_08502_));
 NOR2x2_ASAP7_75t_R _16786_ (.A(_08454_),
    .B(_08014_),
    .Y(_08503_));
 INVx2_ASAP7_75t_R _16787_ (.A(_08503_),
    .Y(_08504_));
 AO21x1_ASAP7_75t_R _16788_ (.A1(_08502_),
    .A2(_08504_),
    .B(_08441_),
    .Y(_08505_));
 AO21x1_ASAP7_75t_R _16789_ (.A1(_08501_),
    .A2(_08505_),
    .B(_08447_),
    .Y(_08506_));
 INVx2_ASAP7_75t_R _16790_ (.A(_07989_),
    .Y(_08507_));
 BUFx6f_ASAP7_75t_R _16791_ (.A(_08507_),
    .Y(_08508_));
 OAI21x1_ASAP7_75t_R _16792_ (.A1(_08499_),
    .A2(_08506_),
    .B(_08508_),
    .Y(_08509_));
 INVx1_ASAP7_75t_R _16793_ (.A(_00394_),
    .Y(_08510_));
 BUFx10_ASAP7_75t_R _16794_ (.A(_08510_),
    .Y(_08511_));
 OAI21x1_ASAP7_75t_R _16795_ (.A1(_08490_),
    .A2(_08509_),
    .B(_08511_),
    .Y(_08512_));
 NAND2x2_ASAP7_75t_R _16796_ (.A(net837),
    .B(_08430_),
    .Y(_08513_));
 AO21x1_ASAP7_75t_R _16797_ (.A1(_08475_),
    .A2(_08513_),
    .B(_08421_),
    .Y(_08514_));
 BUFx6f_ASAP7_75t_R _16798_ (.A(_08449_),
    .Y(_08515_));
 OA21x2_ASAP7_75t_R _16799_ (.A1(_08515_),
    .A2(_08497_),
    .B(_08000_),
    .Y(_08516_));
 AOI21x1_ASAP7_75t_R _16800_ (.A1(_08514_),
    .A2(_08516_),
    .B(_08166_),
    .Y(_08517_));
 NAND2x2_ASAP7_75t_R _16801_ (.A(_08454_),
    .B(_08014_),
    .Y(_08518_));
 NAND2x2_ASAP7_75t_R _16802_ (.A(_07954_),
    .B(_08518_),
    .Y(_08519_));
 INVx3_ASAP7_75t_R _16803_ (.A(_01124_),
    .Y(_08520_));
 NOR2x2_ASAP7_75t_R _16804_ (.A(_08520_),
    .B(_08430_),
    .Y(_08521_));
 OA21x2_ASAP7_75t_R _16805_ (.A1(_08519_),
    .A2(_08521_),
    .B(_08465_),
    .Y(_08522_));
 OAI21x1_ASAP7_75t_R _16806_ (.A1(_00390_),
    .A2(_08497_),
    .B(_08522_),
    .Y(_08523_));
 AOI21x1_ASAP7_75t_R _16807_ (.A1(_08517_),
    .A2(_08523_),
    .B(_08508_),
    .Y(_08524_));
 NAND2x2_ASAP7_75t_R _16808_ (.A(_07954_),
    .B(_08463_),
    .Y(_08525_));
 INVx1_ASAP7_75t_R _16809_ (.A(_08439_),
    .Y(_08526_));
 AO21x1_ASAP7_75t_R _16810_ (.A1(_08526_),
    .A2(_08497_),
    .B(_08421_),
    .Y(_08527_));
 BUFx6f_ASAP7_75t_R _16811_ (.A(_08465_),
    .Y(_08528_));
 AOI21x1_ASAP7_75t_R _16812_ (.A1(_08525_),
    .A2(_08527_),
    .B(_08528_),
    .Y(_08529_));
 NOR2x2_ASAP7_75t_R _16813_ (.A(net481),
    .B(_08014_),
    .Y(_08530_));
 NOR2x2_ASAP7_75t_R _16814_ (.A(_08440_),
    .B(_08530_),
    .Y(_08531_));
 NAND2x1_ASAP7_75t_R _16815_ (.A(_08531_),
    .B(_08502_),
    .Y(_08532_));
 INVx3_ASAP7_75t_R _16816_ (.A(_08426_),
    .Y(_08533_));
 AO21x1_ASAP7_75t_R _16817_ (.A1(_08533_),
    .A2(_08475_),
    .B(_08482_),
    .Y(_08534_));
 BUFx6f_ASAP7_75t_R _16818_ (.A(_08000_),
    .Y(_08535_));
 AOI21x1_ASAP7_75t_R _16819_ (.A1(_08532_),
    .A2(_08534_),
    .B(_08535_),
    .Y(_08536_));
 OAI21x1_ASAP7_75t_R _16820_ (.A1(_08529_),
    .A2(_08536_),
    .B(_08445_),
    .Y(_08537_));
 AOI21x1_ASAP7_75t_R _16821_ (.A1(_08524_),
    .A2(_08537_),
    .B(_08511_),
    .Y(_08538_));
 INVx1_ASAP7_75t_R _16822_ (.A(_08494_),
    .Y(_08539_));
 OAI21x1_ASAP7_75t_R _16823_ (.A1(_08539_),
    .A2(_08491_),
    .B(_08466_),
    .Y(_08540_));
 INVx1_ASAP7_75t_R _16824_ (.A(_08471_),
    .Y(_08541_));
 NAND2x2_ASAP7_75t_R _16825_ (.A(_08520_),
    .B(_08013_),
    .Y(_08542_));
 INVx2_ASAP7_75t_R _16826_ (.A(_08542_),
    .Y(_08543_));
 AO21x1_ASAP7_75t_R _16827_ (.A1(_08453_),
    .A2(_08543_),
    .B(_08416_),
    .Y(_08544_));
 INVx1_ASAP7_75t_R _16828_ (.A(_08544_),
    .Y(_08545_));
 NAND2x1_ASAP7_75t_R _16829_ (.A(_08541_),
    .B(_08545_),
    .Y(_08546_));
 BUFx6f_ASAP7_75t_R _16830_ (.A(_07954_),
    .Y(_08547_));
 NOR2x2_ASAP7_75t_R _16831_ (.A(_01123_),
    .B(_08013_),
    .Y(_08548_));
 INVx4_ASAP7_75t_R _16832_ (.A(_08548_),
    .Y(_08549_));
 NOR2x1_ASAP7_75t_R _16833_ (.A(_08547_),
    .B(_08549_),
    .Y(_08550_));
 AOI21x1_ASAP7_75t_R _16834_ (.A1(_08540_),
    .A2(_08546_),
    .B(_08550_),
    .Y(_08551_));
 BUFx4f_ASAP7_75t_R _16835_ (.A(_08440_),
    .Y(_08552_));
 AO21x1_ASAP7_75t_R _16836_ (.A1(_01127_),
    .A2(_08552_),
    .B(_08531_),
    .Y(_08553_));
 AOI21x1_ASAP7_75t_R _16837_ (.A1(_08443_),
    .A2(_08553_),
    .B(_08445_),
    .Y(_08554_));
 AO21x1_ASAP7_75t_R _16838_ (.A1(_08461_),
    .A2(_08513_),
    .B(_08552_),
    .Y(_08555_));
 NOR2x1_ASAP7_75t_R _16839_ (.A(_00455_),
    .B(_15740_),
    .Y(_08556_));
 OA21x2_ASAP7_75t_R _16840_ (.A1(_08491_),
    .A2(_08556_),
    .B(_08417_),
    .Y(_08557_));
 NAND2x1_ASAP7_75t_R _16841_ (.A(_08555_),
    .B(_08557_),
    .Y(_08558_));
 AOI21x1_ASAP7_75t_R _16842_ (.A1(_08554_),
    .A2(_08558_),
    .B(_00392_),
    .Y(_08559_));
 OAI21x1_ASAP7_75t_R _16843_ (.A1(_08448_),
    .A2(_08551_),
    .B(_08559_),
    .Y(_08560_));
 NAND2x1_ASAP7_75t_R _16844_ (.A(_08538_),
    .B(_08560_),
    .Y(_08561_));
 OAI21x1_ASAP7_75t_R _16845_ (.A1(_08470_),
    .A2(_08512_),
    .B(_08561_),
    .Y(_00000_));
 AO21x1_ASAP7_75t_R _16846_ (.A1(_08420_),
    .A2(_08479_),
    .B(_08421_),
    .Y(_08562_));
 BUFx4f_ASAP7_75t_R _16847_ (.A(_08449_),
    .Y(_08563_));
 AO21x1_ASAP7_75t_R _16848_ (.A1(_08549_),
    .A2(_08433_),
    .B(_08563_),
    .Y(_08564_));
 AND3x1_ASAP7_75t_R _16849_ (.A(_08562_),
    .B(_08535_),
    .C(_08564_),
    .Y(_08565_));
 AO21x1_ASAP7_75t_R _16850_ (.A1(net803),
    .A2(_15742_),
    .B(_08440_),
    .Y(_08566_));
 NAND2x2_ASAP7_75t_R _16851_ (.A(_15729_),
    .B(_15730_),
    .Y(_08567_));
 AO21x1_ASAP7_75t_R _16852_ (.A1(_08567_),
    .A2(_08457_),
    .B(_08515_),
    .Y(_08568_));
 OAI21x1_ASAP7_75t_R _16853_ (.A1(_08530_),
    .A2(_08566_),
    .B(_08568_),
    .Y(_08569_));
 BUFx6f_ASAP7_75t_R _16854_ (.A(_08507_),
    .Y(_08570_));
 OAI21x1_ASAP7_75t_R _16855_ (.A1(_08443_),
    .A2(_08569_),
    .B(_08570_),
    .Y(_08571_));
 NAND2x2_ASAP7_75t_R _16856_ (.A(_08429_),
    .B(_08415_),
    .Y(_08572_));
 BUFx4f_ASAP7_75t_R _16857_ (.A(_08449_),
    .Y(_08573_));
 AO21x1_ASAP7_75t_R _16858_ (.A1(_08572_),
    .A2(_08433_),
    .B(_08573_),
    .Y(_08574_));
 INVx1_ASAP7_75t_R _16859_ (.A(_01123_),
    .Y(_08575_));
 NAND2x1_ASAP7_75t_R _16860_ (.A(_08575_),
    .B(_15742_),
    .Y(_08576_));
 OA21x2_ASAP7_75t_R _16861_ (.A1(_08547_),
    .A2(_08576_),
    .B(_08465_),
    .Y(_08577_));
 BUFx6f_ASAP7_75t_R _16862_ (.A(_08507_),
    .Y(_08578_));
 AOI21x1_ASAP7_75t_R _16863_ (.A1(_08574_),
    .A2(_08577_),
    .B(_08578_),
    .Y(_08579_));
 NAND2x2_ASAP7_75t_R _16864_ (.A(_08429_),
    .B(_08013_),
    .Y(_08580_));
 INVx1_ASAP7_75t_R _16865_ (.A(_08452_),
    .Y(_08581_));
 NOR2x2_ASAP7_75t_R _16866_ (.A(_08415_),
    .B(net805),
    .Y(_08582_));
 OA21x2_ASAP7_75t_R _16867_ (.A1(_08581_),
    .A2(_08582_),
    .B(_08000_),
    .Y(_08583_));
 OAI21x1_ASAP7_75t_R _16868_ (.A1(_00390_),
    .A2(_08580_),
    .B(_08583_),
    .Y(_08584_));
 AOI21x1_ASAP7_75t_R _16869_ (.A1(_08579_),
    .A2(_08584_),
    .B(_08448_),
    .Y(_08585_));
 OAI21x1_ASAP7_75t_R _16870_ (.A1(_08565_),
    .A2(_08571_),
    .B(_08585_),
    .Y(_08586_));
 INVx1_ASAP7_75t_R _16871_ (.A(_08530_),
    .Y(_08587_));
 NAND2x2_ASAP7_75t_R _16872_ (.A(_08450_),
    .B(_08430_),
    .Y(_08588_));
 AO21x1_ASAP7_75t_R _16873_ (.A1(_08587_),
    .A2(_08588_),
    .B(_08573_),
    .Y(_08589_));
 AO21x1_ASAP7_75t_R _16874_ (.A1(_08549_),
    .A2(_08513_),
    .B(_08547_),
    .Y(_08590_));
 NAND3x1_ASAP7_75t_R _16875_ (.A(_08589_),
    .B(_08590_),
    .C(_08466_),
    .Y(_08591_));
 AOI21x1_ASAP7_75t_R _16876_ (.A1(_00460_),
    .A2(_08552_),
    .B(_08417_),
    .Y(_08592_));
 INVx2_ASAP7_75t_R _16877_ (.A(_08582_),
    .Y(_08593_));
 AO21x1_ASAP7_75t_R _16878_ (.A1(_08593_),
    .A2(_08549_),
    .B(_08421_),
    .Y(_08594_));
 AOI21x1_ASAP7_75t_R _16879_ (.A1(_08592_),
    .A2(_08594_),
    .B(_07990_),
    .Y(_08595_));
 AOI21x1_ASAP7_75t_R _16880_ (.A1(_08591_),
    .A2(_08595_),
    .B(_08445_),
    .Y(_08596_));
 OA21x2_ASAP7_75t_R _16881_ (.A1(_08515_),
    .A2(_08504_),
    .B(_08465_),
    .Y(_08597_));
 NAND3x2_ASAP7_75t_R _16882_ (.B(_08515_),
    .C(_08502_),
    .Y(_08598_),
    .A(_08425_));
 AOI21x1_ASAP7_75t_R _16883_ (.A1(_08597_),
    .A2(_08598_),
    .B(_08578_),
    .Y(_08599_));
 AND2x2_ASAP7_75t_R _16884_ (.A(_08463_),
    .B(_08453_),
    .Y(_08600_));
 AO221x1_ASAP7_75t_R _16885_ (.A1(_08461_),
    .A2(_08471_),
    .B1(_08600_),
    .B2(_08420_),
    .C(_08417_),
    .Y(_08601_));
 NAND2x1_ASAP7_75t_R _16886_ (.A(_08599_),
    .B(_08601_),
    .Y(_08602_));
 AOI21x1_ASAP7_75t_R _16887_ (.A1(_08596_),
    .A2(_08602_),
    .B(_08510_),
    .Y(_08603_));
 NAND2x1_ASAP7_75t_R _16888_ (.A(_08586_),
    .B(_08603_),
    .Y(_08604_));
 NAND2x2_ASAP7_75t_R _16889_ (.A(_08496_),
    .B(_08415_),
    .Y(_08605_));
 AO21x1_ASAP7_75t_R _16890_ (.A1(_08605_),
    .A2(_08588_),
    .B(_08421_),
    .Y(_08606_));
 AOI21x1_ASAP7_75t_R _16891_ (.A1(_08574_),
    .A2(_08606_),
    .B(_08466_),
    .Y(_08607_));
 AND3x1_ASAP7_75t_R _16892_ (.A(_08461_),
    .B(_08453_),
    .C(_08494_),
    .Y(_08608_));
 OA21x2_ASAP7_75t_R _16893_ (.A1(_08608_),
    .A2(_08471_),
    .B(_08417_),
    .Y(_08609_));
 OAI21x1_ASAP7_75t_R _16894_ (.A1(_08607_),
    .A2(_08609_),
    .B(_08570_),
    .Y(_08610_));
 NOR2x2_ASAP7_75t_R _16895_ (.A(_08014_),
    .B(net805),
    .Y(_08611_));
 NOR2x2_ASAP7_75t_R _16896_ (.A(_08525_),
    .B(_08611_),
    .Y(_08612_));
 AO211x2_ASAP7_75t_R _16897_ (.A1(_08473_),
    .A2(_08427_),
    .B(_08478_),
    .C(_08612_),
    .Y(_08613_));
 OA21x2_ASAP7_75t_R _16898_ (.A1(_08420_),
    .A2(_08547_),
    .B(_08000_),
    .Y(_08614_));
 OA21x2_ASAP7_75t_R _16899_ (.A1(_00455_),
    .A2(_15740_),
    .B(_08485_),
    .Y(_08615_));
 NOR2x1_ASAP7_75t_R _16900_ (.A(_08498_),
    .B(_08615_),
    .Y(_08616_));
 AOI21x1_ASAP7_75t_R _16901_ (.A1(_08614_),
    .A2(_08616_),
    .B(_08578_),
    .Y(_08617_));
 AOI21x1_ASAP7_75t_R _16902_ (.A1(_08613_),
    .A2(_08617_),
    .B(_08447_),
    .Y(_08618_));
 NAND2x1_ASAP7_75t_R _16903_ (.A(_08610_),
    .B(_08618_),
    .Y(_08619_));
 NAND2x1_ASAP7_75t_R _16904_ (.A(_00459_),
    .B(_07955_),
    .Y(_08620_));
 AO21x1_ASAP7_75t_R _16905_ (.A1(_08475_),
    .A2(_08580_),
    .B(_07954_),
    .Y(_08621_));
 OA21x2_ASAP7_75t_R _16906_ (.A1(_07989_),
    .A2(_08620_),
    .B(_08621_),
    .Y(_08622_));
 OA21x2_ASAP7_75t_R _16907_ (.A1(_08622_),
    .A2(_08535_),
    .B(_08447_),
    .Y(_08623_));
 BUFx6f_ASAP7_75t_R _16908_ (.A(_07990_),
    .Y(_08624_));
 NAND2x2_ASAP7_75t_R _16909_ (.A(_15740_),
    .B(_15729_),
    .Y(_08625_));
 AO21x1_ASAP7_75t_R _16910_ (.A1(_08427_),
    .A2(_08625_),
    .B(_08612_),
    .Y(_08626_));
 AO21x1_ASAP7_75t_R _16911_ (.A1(_08504_),
    .A2(_08580_),
    .B(_08563_),
    .Y(_08627_));
 OA21x2_ASAP7_75t_R _16912_ (.A1(_08566_),
    .A2(_08472_),
    .B(_07990_),
    .Y(_08628_));
 AOI21x1_ASAP7_75t_R _16913_ (.A1(_08627_),
    .A2(_08628_),
    .B(_08466_),
    .Y(_08629_));
 OAI21x1_ASAP7_75t_R _16914_ (.A1(_08624_),
    .A2(_08626_),
    .B(_08629_),
    .Y(_08630_));
 AOI21x1_ASAP7_75t_R _16915_ (.A1(_08623_),
    .A2(_08630_),
    .B(_00394_),
    .Y(_08631_));
 NAND2x1_ASAP7_75t_R _16916_ (.A(_08619_),
    .B(_08631_),
    .Y(_08632_));
 NAND2x1_ASAP7_75t_R _16917_ (.A(_08604_),
    .B(_08632_),
    .Y(_00001_));
 NAND2x1_ASAP7_75t_R _16918_ (.A(_08456_),
    .B(_08465_),
    .Y(_08633_));
 AND3x1_ASAP7_75t_R _16919_ (.A(_07952_),
    .B(_00461_),
    .C(_07941_),
    .Y(_08634_));
 OA21x2_ASAP7_75t_R _16920_ (.A1(_08633_),
    .A2(_08634_),
    .B(_08447_),
    .Y(_08635_));
 OA21x2_ASAP7_75t_R _16921_ (.A1(_01126_),
    .A2(_08421_),
    .B(_08478_),
    .Y(_08636_));
 NAND2x2_ASAP7_75t_R _16922_ (.A(_07954_),
    .B(_08455_),
    .Y(_08637_));
 AO21x1_ASAP7_75t_R _16923_ (.A1(_15729_),
    .A2(_15742_),
    .B(_08637_),
    .Y(_08638_));
 NAND2x1_ASAP7_75t_R _16924_ (.A(_08636_),
    .B(_08638_),
    .Y(_08639_));
 AO21x1_ASAP7_75t_R _16925_ (.A1(_08635_),
    .A2(_08639_),
    .B(_00392_),
    .Y(_08640_));
 AO21x1_ASAP7_75t_R _16926_ (.A1(_08502_),
    .A2(_08526_),
    .B(_08547_),
    .Y(_08641_));
 OR3x1_ASAP7_75t_R _16927_ (.A(_08573_),
    .B(_08436_),
    .C(_15740_),
    .Y(_08642_));
 NAND2x2_ASAP7_75t_R _16928_ (.A(_08440_),
    .B(_08530_),
    .Y(_08643_));
 AND4x1_ASAP7_75t_R _16929_ (.A(_08641_),
    .B(_08001_),
    .C(_08642_),
    .D(_08643_),
    .Y(_08644_));
 NOR2x1_ASAP7_75t_R _16930_ (.A(_15729_),
    .B(_15730_),
    .Y(_08645_));
 AO21x2_ASAP7_75t_R _16931_ (.A1(_15729_),
    .A2(_08430_),
    .B(_08449_),
    .Y(_08646_));
 OAI21x1_ASAP7_75t_R _16932_ (.A1(_08645_),
    .A2(_08646_),
    .B(_08465_),
    .Y(_08647_));
 AO21x1_ASAP7_75t_R _16933_ (.A1(_00459_),
    .A2(_08474_),
    .B(_08647_),
    .Y(_08648_));
 NAND2x1_ASAP7_75t_R _16934_ (.A(_08445_),
    .B(_08648_),
    .Y(_08649_));
 NOR2x1_ASAP7_75t_R _16935_ (.A(_08644_),
    .B(_08649_),
    .Y(_08650_));
 NOR2x1_ASAP7_75t_R _16936_ (.A(_01127_),
    .B(_08440_),
    .Y(_08651_));
 AO21x1_ASAP7_75t_R _16937_ (.A1(_08485_),
    .A2(_08518_),
    .B(_08651_),
    .Y(_08652_));
 AND2x2_ASAP7_75t_R _16938_ (.A(_08652_),
    .B(_08417_),
    .Y(_08653_));
 AO21x1_ASAP7_75t_R _16939_ (.A1(_08533_),
    .A2(_01126_),
    .B(_08515_),
    .Y(_08654_));
 AOI21x1_ASAP7_75t_R _16940_ (.A1(_08532_),
    .A2(_08654_),
    .B(_08466_),
    .Y(_08655_));
 OAI21x1_ASAP7_75t_R _16941_ (.A1(_08653_),
    .A2(_08655_),
    .B(_08445_),
    .Y(_08656_));
 NAND2x2_ASAP7_75t_R _16942_ (.A(_08483_),
    .B(_08013_),
    .Y(_08657_));
 AO21x1_ASAP7_75t_R _16943_ (.A1(_08549_),
    .A2(_08657_),
    .B(_08563_),
    .Y(_08658_));
 AOI21x1_ASAP7_75t_R _16944_ (.A1(_08481_),
    .A2(_08658_),
    .B(_08166_),
    .Y(_08659_));
 AO21x2_ASAP7_75t_R _16945_ (.A1(_15730_),
    .A2(_15742_),
    .B(_08453_),
    .Y(_08660_));
 AND2x2_ASAP7_75t_R _16946_ (.A(_08621_),
    .B(_08000_),
    .Y(_08661_));
 OAI21x1_ASAP7_75t_R _16947_ (.A1(_08431_),
    .A2(_08660_),
    .B(_08661_),
    .Y(_08662_));
 AOI21x1_ASAP7_75t_R _16948_ (.A1(_08659_),
    .A2(_08662_),
    .B(_08570_),
    .Y(_08663_));
 AOI21x1_ASAP7_75t_R _16949_ (.A1(_08656_),
    .A2(_08663_),
    .B(_08511_),
    .Y(_08664_));
 OAI21x1_ASAP7_75t_R _16950_ (.A1(_08640_),
    .A2(_08650_),
    .B(_08664_),
    .Y(_08665_));
 NOR2x2_ASAP7_75t_R _16951_ (.A(_01122_),
    .B(_08014_),
    .Y(_08666_));
 INVx2_ASAP7_75t_R _16952_ (.A(_08666_),
    .Y(_08667_));
 AO21x1_ASAP7_75t_R _16953_ (.A1(_08667_),
    .A2(_08576_),
    .B(_08547_),
    .Y(_08668_));
 AOI21x1_ASAP7_75t_R _16954_ (.A1(_08668_),
    .A2(_08638_),
    .B(_08466_),
    .Y(_08669_));
 NOR2x1_ASAP7_75t_R _16955_ (.A(_08453_),
    .B(_08548_),
    .Y(_08670_));
 AO21x1_ASAP7_75t_R _16956_ (.A1(_08670_),
    .A2(_08513_),
    .B(_08000_),
    .Y(_08671_));
 AOI21x1_ASAP7_75t_R _16957_ (.A1(_08502_),
    .A2(_08531_),
    .B(_08671_),
    .Y(_08672_));
 OAI21x1_ASAP7_75t_R _16958_ (.A1(_08669_),
    .A2(_08672_),
    .B(_08447_),
    .Y(_08673_));
 AO21x1_ASAP7_75t_R _16959_ (.A1(_08502_),
    .A2(_08549_),
    .B(_08573_),
    .Y(_08674_));
 AO21x1_ASAP7_75t_R _16960_ (.A1(_08549_),
    .A2(_08542_),
    .B(_07955_),
    .Y(_08675_));
 NAND3x1_ASAP7_75t_R _16961_ (.A(_08674_),
    .B(_08466_),
    .C(_08675_),
    .Y(_08676_));
 NOR2x1_ASAP7_75t_R _16962_ (.A(_08440_),
    .B(_08666_),
    .Y(_08677_));
 AO21x1_ASAP7_75t_R _16963_ (.A1(_08533_),
    .A2(_08670_),
    .B(_08677_),
    .Y(_08678_));
 AOI21x1_ASAP7_75t_R _16964_ (.A1(_08678_),
    .A2(_08545_),
    .B(_08447_),
    .Y(_08679_));
 AOI21x1_ASAP7_75t_R _16965_ (.A1(_08676_),
    .A2(_08679_),
    .B(_08624_),
    .Y(_08680_));
 NAND2x1_ASAP7_75t_R _16966_ (.A(_08673_),
    .B(_08680_),
    .Y(_08681_));
 INVx2_ASAP7_75t_R _16967_ (.A(_08484_),
    .Y(_08682_));
 AO21x1_ASAP7_75t_R _16968_ (.A1(_08682_),
    .A2(_08657_),
    .B(_08515_),
    .Y(_08683_));
 NAND2x2_ASAP7_75t_R _16969_ (.A(_08520_),
    .B(_08415_),
    .Y(_08684_));
 AO21x1_ASAP7_75t_R _16970_ (.A1(_08533_),
    .A2(_08684_),
    .B(_08547_),
    .Y(_08685_));
 AOI21x1_ASAP7_75t_R _16971_ (.A1(_08683_),
    .A2(_08685_),
    .B(_08535_),
    .Y(_08686_));
 AO21x1_ASAP7_75t_R _16972_ (.A1(_15730_),
    .A2(_15742_),
    .B(_07955_),
    .Y(_08687_));
 OAI21x1_ASAP7_75t_R _16973_ (.A1(_08666_),
    .A2(_08687_),
    .B(_08478_),
    .Y(_08688_));
 INVx2_ASAP7_75t_R _16974_ (.A(_08611_),
    .Y(_08689_));
 AND3x1_ASAP7_75t_R _16975_ (.A(_08689_),
    .B(_08547_),
    .C(_08542_),
    .Y(_08690_));
 NOR2x1_ASAP7_75t_R _16976_ (.A(_08688_),
    .B(_08690_),
    .Y(_08691_));
 OAI21x1_ASAP7_75t_R _16977_ (.A1(_08686_),
    .A2(_08691_),
    .B(_08445_),
    .Y(_08692_));
 AOI21x1_ASAP7_75t_R _16978_ (.A1(_08588_),
    .A2(_08572_),
    .B(_08515_),
    .Y(_08693_));
 OA21x2_ASAP7_75t_R _16979_ (.A1(_08633_),
    .A2(_08693_),
    .B(_08447_),
    .Y(_08694_));
 INVx1_ASAP7_75t_R _16980_ (.A(_08605_),
    .Y(_08695_));
 NAND2x2_ASAP7_75t_R _16981_ (.A(_08657_),
    .B(_08449_),
    .Y(_08696_));
 AO21x1_ASAP7_75t_R _16982_ (.A1(_15735_),
    .A2(_15740_),
    .B(_08696_),
    .Y(_08697_));
 OAI21x1_ASAP7_75t_R _16983_ (.A1(_08695_),
    .A2(_08660_),
    .B(_08697_),
    .Y(_08698_));
 NAND2x1_ASAP7_75t_R _16984_ (.A(_08535_),
    .B(_08698_),
    .Y(_08699_));
 AOI21x1_ASAP7_75t_R _16985_ (.A1(_08694_),
    .A2(_08699_),
    .B(_08570_),
    .Y(_08700_));
 AOI21x1_ASAP7_75t_R _16986_ (.A1(_08692_),
    .A2(_08700_),
    .B(_00394_),
    .Y(_08701_));
 NAND2x1_ASAP7_75t_R _16987_ (.A(_08681_),
    .B(_08701_),
    .Y(_08702_));
 NAND2x1_ASAP7_75t_R _16988_ (.A(_08665_),
    .B(_08702_),
    .Y(_00002_));
 NAND2x1_ASAP7_75t_R _16989_ (.A(_08422_),
    .B(_08533_),
    .Y(_08703_));
 NOR2x1_ASAP7_75t_R _16990_ (.A(_00390_),
    .B(_08703_),
    .Y(_08704_));
 NAND2x1_ASAP7_75t_R _16991_ (.A(_08637_),
    .B(_08528_),
    .Y(_08705_));
 OA21x2_ASAP7_75t_R _16992_ (.A1(_08704_),
    .A2(_08705_),
    .B(_08508_),
    .Y(_08706_));
 OAI21x1_ASAP7_75t_R _16993_ (.A1(_08521_),
    .A2(_08696_),
    .B(_08583_),
    .Y(_08707_));
 NAND2x2_ASAP7_75t_R _16994_ (.A(_08515_),
    .B(_08494_),
    .Y(_08708_));
 NOR2x1_ASAP7_75t_R _16995_ (.A(_08484_),
    .B(_08708_),
    .Y(_08709_));
 OA21x2_ASAP7_75t_R _16996_ (.A1(_08437_),
    .A2(_08503_),
    .B(_08441_),
    .Y(_08710_));
 OAI21x1_ASAP7_75t_R _16997_ (.A1(_08709_),
    .A2(_08710_),
    .B(_08418_),
    .Y(_08711_));
 OA21x2_ASAP7_75t_R _16998_ (.A1(_08476_),
    .A2(_08434_),
    .B(_08474_),
    .Y(_08712_));
 AOI21x1_ASAP7_75t_R _16999_ (.A1(_08422_),
    .A2(_08420_),
    .B(_08474_),
    .Y(_08713_));
 OAI21x1_ASAP7_75t_R _17000_ (.A1(_08712_),
    .A2(_08713_),
    .B(_00391_),
    .Y(_08714_));
 AOI21x1_ASAP7_75t_R _17001_ (.A1(_08711_),
    .A2(_08714_),
    .B(_08508_),
    .Y(_08715_));
 AOI211x1_ASAP7_75t_R _17002_ (.A1(_08706_),
    .A2(_08707_),
    .B(_08715_),
    .C(_08448_),
    .Y(_08716_));
 OAI22x1_ASAP7_75t_R _17003_ (.A1(_08703_),
    .A2(_00390_),
    .B1(_08541_),
    .B2(_08611_),
    .Y(_08717_));
 AND2x2_ASAP7_75t_R _17004_ (.A(_08533_),
    .B(_01126_),
    .Y(_08718_));
 NAND2x2_ASAP7_75t_R _17005_ (.A(_07955_),
    .B(_08484_),
    .Y(_08719_));
 NAND2x1_ASAP7_75t_R _17006_ (.A(_08719_),
    .B(_08001_),
    .Y(_08720_));
 AOI21x1_ASAP7_75t_R _17007_ (.A1(_08474_),
    .A2(_08718_),
    .B(_08720_),
    .Y(_08721_));
 AOI21x1_ASAP7_75t_R _17008_ (.A1(_08418_),
    .A2(_08717_),
    .B(_08721_),
    .Y(_08722_));
 AO21x1_ASAP7_75t_R _17009_ (.A1(_08682_),
    .A2(_08479_),
    .B(_08563_),
    .Y(_08723_));
 OAI21x1_ASAP7_75t_R _17010_ (.A1(_08437_),
    .A2(_08419_),
    .B(_08474_),
    .Y(_08724_));
 AOI21x1_ASAP7_75t_R _17011_ (.A1(_08723_),
    .A2(_08724_),
    .B(_08528_),
    .Y(_08725_));
 AO21x1_ASAP7_75t_R _17012_ (.A1(_08549_),
    .A2(_08588_),
    .B(_08482_),
    .Y(_08726_));
 AOI21x1_ASAP7_75t_R _17013_ (.A1(_08726_),
    .A2(_08697_),
    .B(_08443_),
    .Y(_08727_));
 OAI21x1_ASAP7_75t_R _17014_ (.A1(_08725_),
    .A2(_08727_),
    .B(_00392_),
    .Y(_08728_));
 OAI21x1_ASAP7_75t_R _17015_ (.A1(_00392_),
    .A2(_08722_),
    .B(_08728_),
    .Y(_08729_));
 OAI21x1_ASAP7_75t_R _17016_ (.A1(_00393_),
    .A2(_08729_),
    .B(_00394_),
    .Y(_08730_));
 OA21x2_ASAP7_75t_R _17017_ (.A1(_00454_),
    .A2(_15742_),
    .B(_08573_),
    .Y(_08731_));
 NAND2x1_ASAP7_75t_R _17018_ (.A(_08502_),
    .B(_08731_),
    .Y(_08732_));
 AOI21x1_ASAP7_75t_R _17019_ (.A1(_08719_),
    .A2(_08732_),
    .B(_07990_),
    .Y(_08733_));
 NAND2x1_ASAP7_75t_R _17020_ (.A(_08482_),
    .B(_08434_),
    .Y(_08734_));
 OAI21x1_ASAP7_75t_R _17021_ (.A1(_08578_),
    .A2(_08734_),
    .B(_08516_),
    .Y(_08735_));
 OAI21x1_ASAP7_75t_R _17022_ (.A1(_08733_),
    .A2(_08735_),
    .B(_08448_),
    .Y(_08736_));
 AOI21x1_ASAP7_75t_R _17023_ (.A1(_08461_),
    .A2(_08435_),
    .B(_07990_),
    .Y(_08737_));
 OAI21x1_ASAP7_75t_R _17024_ (.A1(_08426_),
    .A2(_08581_),
    .B(_08737_),
    .Y(_08738_));
 NAND2x2_ASAP7_75t_R _17025_ (.A(_08440_),
    .B(_08543_),
    .Y(_08739_));
 AND2x2_ASAP7_75t_R _17026_ (.A(_08739_),
    .B(_07989_),
    .Y(_08740_));
 NAND2x1_ASAP7_75t_R _17027_ (.A(_08740_),
    .B(_08685_),
    .Y(_08741_));
 AOI21x1_ASAP7_75t_R _17028_ (.A1(_08738_),
    .A2(_08741_),
    .B(_00391_),
    .Y(_08742_));
 NOR2x1_ASAP7_75t_R _17029_ (.A(_08736_),
    .B(_08742_),
    .Y(_08743_));
 AO21x2_ASAP7_75t_R _17030_ (.A1(_08457_),
    .A2(_08684_),
    .B(_08515_),
    .Y(_08744_));
 AOI21x1_ASAP7_75t_R _17031_ (.A1(_08621_),
    .A2(_08744_),
    .B(_08535_),
    .Y(_08745_));
 NAND2x1_ASAP7_75t_R _17032_ (.A(_08578_),
    .B(_08688_),
    .Y(_08746_));
 OAI21x1_ASAP7_75t_R _17033_ (.A1(_08745_),
    .A2(_08746_),
    .B(_08445_),
    .Y(_08747_));
 AO21x1_ASAP7_75t_R _17034_ (.A1(_08667_),
    .A2(_08657_),
    .B(_08552_),
    .Y(_08748_));
 AOI21x1_ASAP7_75t_R _17035_ (.A1(_08542_),
    .A2(_08461_),
    .B(_08573_),
    .Y(_08749_));
 NOR2x1_ASAP7_75t_R _17036_ (.A(_08417_),
    .B(_08749_),
    .Y(_08750_));
 NAND2x1_ASAP7_75t_R _17037_ (.A(_08748_),
    .B(_08750_),
    .Y(_08751_));
 NAND2x1_ASAP7_75t_R _17038_ (.A(_08598_),
    .B(_08557_),
    .Y(_08752_));
 AOI21x1_ASAP7_75t_R _17039_ (.A1(_08751_),
    .A2(_08752_),
    .B(_08508_),
    .Y(_08753_));
 NOR2x1_ASAP7_75t_R _17040_ (.A(_08747_),
    .B(_08753_),
    .Y(_08754_));
 OAI21x1_ASAP7_75t_R _17041_ (.A1(_08743_),
    .A2(_08754_),
    .B(_08511_),
    .Y(_08755_));
 OAI21x1_ASAP7_75t_R _17042_ (.A1(_08716_),
    .A2(_08730_),
    .B(_08755_),
    .Y(_00003_));
 OAI21x1_ASAP7_75t_R _17043_ (.A1(_08429_),
    .A2(_00390_),
    .B(_08643_),
    .Y(_08756_));
 AO21x1_ASAP7_75t_R _17044_ (.A1(_08756_),
    .A2(_08528_),
    .B(_08570_),
    .Y(_08757_));
 NOR2x2_ASAP7_75t_R _17045_ (.A(_08573_),
    .B(_08521_),
    .Y(_08758_));
 INVx1_ASAP7_75t_R _17046_ (.A(_08758_),
    .Y(_08759_));
 OA21x2_ASAP7_75t_R _17047_ (.A1(_08552_),
    .A2(_08513_),
    .B(_08478_),
    .Y(_08760_));
 OA21x2_ASAP7_75t_R _17048_ (.A1(_08582_),
    .A2(_08759_),
    .B(_08760_),
    .Y(_08761_));
 OAI21x1_ASAP7_75t_R _17049_ (.A1(_08757_),
    .A2(_08761_),
    .B(_08511_),
    .Y(_08762_));
 AOI21x1_ASAP7_75t_R _17050_ (.A1(_08567_),
    .A2(_08593_),
    .B(_00390_),
    .Y(_08763_));
 INVx1_ASAP7_75t_R _17051_ (.A(_08744_),
    .Y(_08764_));
 OAI21x1_ASAP7_75t_R _17052_ (.A1(_08763_),
    .A2(_08764_),
    .B(_00391_),
    .Y(_08765_));
 INVx1_ASAP7_75t_R _17053_ (.A(_08527_),
    .Y(_08766_));
 OAI21x1_ASAP7_75t_R _17054_ (.A1(_08766_),
    .A2(_08423_),
    .B(_08418_),
    .Y(_08767_));
 AOI21x1_ASAP7_75t_R _17055_ (.A1(_08765_),
    .A2(_08767_),
    .B(_00392_),
    .Y(_08768_));
 OAI21x1_ASAP7_75t_R _17056_ (.A1(_08762_),
    .A2(_08768_),
    .B(_08448_),
    .Y(_08769_));
 INVx2_ASAP7_75t_R _17057_ (.A(_08519_),
    .Y(_08770_));
 NAND2x1_ASAP7_75t_R _17058_ (.A(_08770_),
    .B(_08689_),
    .Y(_08771_));
 AO21x1_ASAP7_75t_R _17059_ (.A1(_08771_),
    .A2(_08668_),
    .B(_08528_),
    .Y(_08772_));
 AO21x1_ASAP7_75t_R _17060_ (.A1(_08625_),
    .A2(_08479_),
    .B(_08482_),
    .Y(_08773_));
 AO21x1_ASAP7_75t_R _17061_ (.A1(_08773_),
    .A2(_08590_),
    .B(_08443_),
    .Y(_08774_));
 AOI21x1_ASAP7_75t_R _17062_ (.A1(_08772_),
    .A2(_08774_),
    .B(_00392_),
    .Y(_08775_));
 AO21x1_ASAP7_75t_R _17063_ (.A1(_08587_),
    .A2(_08588_),
    .B(_08552_),
    .Y(_08776_));
 AO21x1_ASAP7_75t_R _17064_ (.A1(_08522_),
    .A2(_08776_),
    .B(_08578_),
    .Y(_08777_));
 AND4x1_ASAP7_75t_R _17065_ (.A(_08675_),
    .B(_08001_),
    .C(_08643_),
    .D(_08739_),
    .Y(_08778_));
 OAI21x1_ASAP7_75t_R _17066_ (.A1(_08777_),
    .A2(_08778_),
    .B(_00394_),
    .Y(_08779_));
 NOR2x1_ASAP7_75t_R _17067_ (.A(_08775_),
    .B(_08779_),
    .Y(_08780_));
 OAI21x1_ASAP7_75t_R _17068_ (.A1(_08439_),
    .A2(_08646_),
    .B(_00391_),
    .Y(_08781_));
 NOR2x1_ASAP7_75t_R _17069_ (.A(_08645_),
    .B(_08646_),
    .Y(_08782_));
 AND2x2_ASAP7_75t_R _17070_ (.A(_08427_),
    .B(_08625_),
    .Y(_08783_));
 OAI21x1_ASAP7_75t_R _17071_ (.A1(_08782_),
    .A2(_08783_),
    .B(_08418_),
    .Y(_08784_));
 OAI21x1_ASAP7_75t_R _17072_ (.A1(_08763_),
    .A2(_08781_),
    .B(_08784_),
    .Y(_08785_));
 OAI21x1_ASAP7_75t_R _17073_ (.A1(_01128_),
    .A2(_08515_),
    .B(_08465_),
    .Y(_08786_));
 AO22x1_ASAP7_75t_R _17074_ (.A1(_08482_),
    .A2(_08439_),
    .B1(_15730_),
    .B2(_15742_),
    .Y(_08787_));
 NOR2x1_ASAP7_75t_R _17075_ (.A(_08786_),
    .B(_08787_),
    .Y(_08788_));
 NOR2x1_ASAP7_75t_R _17076_ (.A(_08758_),
    .B(_08498_),
    .Y(_08789_));
 AO21x1_ASAP7_75t_R _17077_ (.A1(_08789_),
    .A2(_08443_),
    .B(_08570_),
    .Y(_08790_));
 OAI21x1_ASAP7_75t_R _17078_ (.A1(_08788_),
    .A2(_08790_),
    .B(_00394_),
    .Y(_08791_));
 AOI21x1_ASAP7_75t_R _17079_ (.A1(_08508_),
    .A2(_08785_),
    .B(_08791_),
    .Y(_08792_));
 OA21x2_ASAP7_75t_R _17080_ (.A1(_08496_),
    .A2(_15742_),
    .B(_08573_),
    .Y(_08793_));
 AO21x1_ASAP7_75t_R _17081_ (.A1(_08441_),
    .A2(_08432_),
    .B(_08793_),
    .Y(_08794_));
 OAI21x1_ASAP7_75t_R _17082_ (.A1(_08418_),
    .A2(_08794_),
    .B(_00392_),
    .Y(_08795_));
 AOI21x1_ASAP7_75t_R _17083_ (.A1(_08587_),
    .A2(_08600_),
    .B(_08540_),
    .Y(_08796_));
 OAI21x1_ASAP7_75t_R _17084_ (.A1(_08795_),
    .A2(_08796_),
    .B(_08511_),
    .Y(_08797_));
 NOR2x1_ASAP7_75t_R _17085_ (.A(_08480_),
    .B(_08465_),
    .Y(_08798_));
 NOR2x1_ASAP7_75t_R _17086_ (.A(_08612_),
    .B(_08488_),
    .Y(_08799_));
 AO21x1_ASAP7_75t_R _17087_ (.A1(_08457_),
    .A2(_08667_),
    .B(_08441_),
    .Y(_08800_));
 NOR2x2_ASAP7_75t_R _17088_ (.A(_15742_),
    .B(_08453_),
    .Y(_08801_));
 NOR2x1_ASAP7_75t_R _17089_ (.A(_08801_),
    .B(_08001_),
    .Y(_08802_));
 AO21x1_ASAP7_75t_R _17090_ (.A1(_08800_),
    .A2(_08802_),
    .B(_08624_),
    .Y(_08803_));
 AOI21x1_ASAP7_75t_R _17091_ (.A1(_08798_),
    .A2(_08799_),
    .B(_08803_),
    .Y(_08804_));
 OAI21x1_ASAP7_75t_R _17092_ (.A1(_08797_),
    .A2(_08804_),
    .B(_00393_),
    .Y(_08805_));
 OAI22x1_ASAP7_75t_R _17093_ (.A1(_08769_),
    .A2(_08780_),
    .B1(_08792_),
    .B2(_08805_),
    .Y(_00004_));
 OA21x2_ASAP7_75t_R _17094_ (.A1(_08600_),
    .A2(_08503_),
    .B(_08001_),
    .Y(_08806_));
 OA21x2_ASAP7_75t_R _17095_ (.A1(_08749_),
    .A2(_08435_),
    .B(_08417_),
    .Y(_08807_));
 OAI21x1_ASAP7_75t_R _17096_ (.A1(_08806_),
    .A2(_08807_),
    .B(_08570_),
    .Y(_08808_));
 NAND2x1_ASAP7_75t_R _17097_ (.A(_08445_),
    .B(_08808_),
    .Y(_08809_));
 AO21x1_ASAP7_75t_R _17098_ (.A1(_08457_),
    .A2(_08549_),
    .B(_08482_),
    .Y(_08810_));
 AO21x1_ASAP7_75t_R _17099_ (.A1(_08684_),
    .A2(_08513_),
    .B(_08552_),
    .Y(_08811_));
 AO21x1_ASAP7_75t_R _17100_ (.A1(_08810_),
    .A2(_08811_),
    .B(_08528_),
    .Y(_08812_));
 AO21x1_ASAP7_75t_R _17101_ (.A1(_08689_),
    .A2(_08497_),
    .B(_08441_),
    .Y(_08813_));
 NAND2x1_ASAP7_75t_R _17102_ (.A(_08463_),
    .B(_08452_),
    .Y(_08814_));
 AO21x1_ASAP7_75t_R _17103_ (.A1(_08813_),
    .A2(_08814_),
    .B(_08443_),
    .Y(_08815_));
 AOI21x1_ASAP7_75t_R _17104_ (.A1(_08812_),
    .A2(_08815_),
    .B(_08508_),
    .Y(_08816_));
 NOR2x1_ASAP7_75t_R _17105_ (.A(_08809_),
    .B(_08816_),
    .Y(_08817_));
 OA21x2_ASAP7_75t_R _17106_ (.A1(net803),
    .A2(_08441_),
    .B(_15729_),
    .Y(_08818_));
 OAI21x1_ASAP7_75t_R _17107_ (.A1(_08818_),
    .A2(_08495_),
    .B(_08624_),
    .Y(_08819_));
 NAND3x1_ASAP7_75t_R _17108_ (.A(_08475_),
    .B(_08580_),
    .C(_00390_),
    .Y(_08820_));
 NAND2x1_ASAP7_75t_R _17109_ (.A(_08567_),
    .B(_08462_),
    .Y(_08821_));
 AOI21x1_ASAP7_75t_R _17110_ (.A1(_08820_),
    .A2(_08821_),
    .B(_08418_),
    .Y(_08822_));
 NOR2x1_ASAP7_75t_R _17111_ (.A(_08819_),
    .B(_08822_),
    .Y(_08823_));
 AO21x1_ASAP7_75t_R _17112_ (.A1(_08471_),
    .A2(_08526_),
    .B(_08677_),
    .Y(_08824_));
 AND2x2_ASAP7_75t_R _17113_ (.A(_08824_),
    .B(_08528_),
    .Y(_08825_));
 NAND2x1_ASAP7_75t_R _17114_ (.A(_08643_),
    .B(_08478_),
    .Y(_08826_));
 AO21x1_ASAP7_75t_R _17115_ (.A1(_08502_),
    .A2(_08793_),
    .B(_08826_),
    .Y(_08827_));
 NAND2x1_ASAP7_75t_R _17116_ (.A(_08570_),
    .B(_08827_),
    .Y(_08828_));
 OAI21x1_ASAP7_75t_R _17117_ (.A1(_08825_),
    .A2(_08828_),
    .B(_08448_),
    .Y(_08829_));
 OAI21x1_ASAP7_75t_R _17118_ (.A1(_08823_),
    .A2(_08829_),
    .B(_00394_),
    .Y(_08830_));
 OA21x2_ASAP7_75t_R _17119_ (.A1(_08426_),
    .A2(_08548_),
    .B(_08474_),
    .Y(_08831_));
 NOR2x1_ASAP7_75t_R _17120_ (.A(_08831_),
    .B(_08540_),
    .Y(_08832_));
 OAI22x1_ASAP7_75t_R _17121_ (.A1(_08708_),
    .A2(_08451_),
    .B1(_08474_),
    .B2(_08475_),
    .Y(_08833_));
 OAI21x1_ASAP7_75t_R _17122_ (.A1(_08418_),
    .A2(_08833_),
    .B(_08508_),
    .Y(_08834_));
 OAI21x1_ASAP7_75t_R _17123_ (.A1(_08832_),
    .A2(_08834_),
    .B(_00393_),
    .Y(_08835_));
 OA21x2_ASAP7_75t_R _17124_ (.A1(_08563_),
    .A2(net803),
    .B(_08417_),
    .Y(_08836_));
 AO21x1_ASAP7_75t_R _17125_ (.A1(_08836_),
    .A2(_08428_),
    .B(_08578_),
    .Y(_08837_));
 INVx1_ASAP7_75t_R _17126_ (.A(_08521_),
    .Y(_08838_));
 NOR2x2_ASAP7_75t_R _17127_ (.A(_08547_),
    .B(_08582_),
    .Y(_08839_));
 AOI221x1_ASAP7_75t_R _17128_ (.A1(_08455_),
    .A2(_08471_),
    .B1(_08838_),
    .B2(_08839_),
    .C(_08418_),
    .Y(_08840_));
 NOR2x1_ASAP7_75t_R _17129_ (.A(_08837_),
    .B(_08840_),
    .Y(_08841_));
 OAI21x1_ASAP7_75t_R _17130_ (.A1(_08835_),
    .A2(_08841_),
    .B(_08511_),
    .Y(_08842_));
 AO21x1_ASAP7_75t_R _17131_ (.A1(_08475_),
    .A2(_08657_),
    .B(_08563_),
    .Y(_08843_));
 AO21x1_ASAP7_75t_R _17132_ (.A1(_08667_),
    .A2(_08433_),
    .B(_08552_),
    .Y(_08844_));
 AOI21x1_ASAP7_75t_R _17133_ (.A1(_08843_),
    .A2(_08844_),
    .B(_08528_),
    .Y(_08845_));
 NAND2x1_ASAP7_75t_R _17134_ (.A(_00454_),
    .B(_08441_),
    .Y(_08846_));
 AOI21x1_ASAP7_75t_R _17135_ (.A1(_08846_),
    .A2(_08708_),
    .B(_08535_),
    .Y(_08847_));
 OR3x1_ASAP7_75t_R _17136_ (.A(_08845_),
    .B(_08624_),
    .C(_08847_),
    .Y(_08848_));
 AO21x1_ASAP7_75t_R _17137_ (.A1(_08504_),
    .A2(_08580_),
    .B(_08552_),
    .Y(_08849_));
 AOI21x1_ASAP7_75t_R _17138_ (.A1(_08660_),
    .A2(_08849_),
    .B(_08535_),
    .Y(_08850_));
 OA21x2_ASAP7_75t_R _17139_ (.A1(_08550_),
    .A2(_08452_),
    .B(_08001_),
    .Y(_08851_));
 OR3x1_ASAP7_75t_R _17140_ (.A(_08850_),
    .B(_08570_),
    .C(_08851_),
    .Y(_08852_));
 AOI21x1_ASAP7_75t_R _17141_ (.A1(_08848_),
    .A2(_08852_),
    .B(_00393_),
    .Y(_08853_));
 OAI22x1_ASAP7_75t_R _17142_ (.A1(_08817_),
    .A2(_08830_),
    .B1(_08842_),
    .B2(_08853_),
    .Y(_00005_));
 AO21x1_ASAP7_75t_R _17143_ (.A1(_08533_),
    .A2(_08422_),
    .B(_08563_),
    .Y(_08854_));
 NAND2x1_ASAP7_75t_R _17144_ (.A(_08504_),
    .B(_08839_),
    .Y(_08855_));
 AOI21x1_ASAP7_75t_R _17145_ (.A1(_08854_),
    .A2(_08855_),
    .B(_08443_),
    .Y(_08856_));
 NOR2x2_ASAP7_75t_R _17146_ (.A(_08547_),
    .B(_08500_),
    .Y(_08857_));
 AOI21x1_ASAP7_75t_R _17147_ (.A1(_08420_),
    .A2(_08857_),
    .B(_08417_),
    .Y(_08858_));
 AO21x1_ASAP7_75t_R _17148_ (.A1(_08854_),
    .A2(_08858_),
    .B(_08570_),
    .Y(_08859_));
 NOR2x1_ASAP7_75t_R _17149_ (.A(_08856_),
    .B(_08859_),
    .Y(_08860_));
 INVx1_ASAP7_75t_R _17150_ (.A(_08459_),
    .Y(_08861_));
 AO21x1_ASAP7_75t_R _17151_ (.A1(_08592_),
    .A2(_08861_),
    .B(_08624_),
    .Y(_08862_));
 INVx1_ASAP7_75t_R _17152_ (.A(_08749_),
    .Y(_08863_));
 AO21x1_ASAP7_75t_R _17153_ (.A1(_07941_),
    .A2(_07952_),
    .B(_08657_),
    .Y(_08864_));
 AND3x1_ASAP7_75t_R _17154_ (.A(_08863_),
    .B(_08864_),
    .C(_08528_),
    .Y(_08865_));
 OAI21x1_ASAP7_75t_R _17155_ (.A1(_08862_),
    .A2(_08865_),
    .B(_00393_),
    .Y(_08866_));
 OAI21x1_ASAP7_75t_R _17156_ (.A1(_08860_),
    .A2(_08866_),
    .B(_08511_),
    .Y(_08867_));
 AO21x1_ASAP7_75t_R _17157_ (.A1(_08593_),
    .A2(_08758_),
    .B(_08731_),
    .Y(_08868_));
 NAND2x1_ASAP7_75t_R _17158_ (.A(_08578_),
    .B(_08671_),
    .Y(_08869_));
 AO21x1_ASAP7_75t_R _17159_ (.A1(_00391_),
    .A2(_08868_),
    .B(_08869_),
    .Y(_08870_));
 AO21x1_ASAP7_75t_R _17160_ (.A1(_00462_),
    .A2(_08441_),
    .B(_08001_),
    .Y(_08871_));
 AOI21x1_ASAP7_75t_R _17161_ (.A1(_08839_),
    .A2(_08838_),
    .B(_08871_),
    .Y(_08872_));
 NAND2x1_ASAP7_75t_R _17162_ (.A(_08657_),
    .B(_08452_),
    .Y(_08873_));
 AND2x2_ASAP7_75t_R _17163_ (.A(_08614_),
    .B(_08873_),
    .Y(_08874_));
 OAI21x1_ASAP7_75t_R _17164_ (.A1(_08872_),
    .A2(_08874_),
    .B(_00392_),
    .Y(_08875_));
 AOI21x1_ASAP7_75t_R _17165_ (.A1(_08870_),
    .A2(_08875_),
    .B(_00393_),
    .Y(_08876_));
 NAND2x1_ASAP7_75t_R _17166_ (.A(_08496_),
    .B(_08801_),
    .Y(_08877_));
 AND3x1_ASAP7_75t_R _17167_ (.A(_08798_),
    .B(_08739_),
    .C(_08877_),
    .Y(_08878_));
 AO21x1_ASAP7_75t_R _17168_ (.A1(_08593_),
    .A2(_08567_),
    .B(_08563_),
    .Y(_08879_));
 NOR2x1_ASAP7_75t_R _17169_ (.A(_08478_),
    .B(_08487_),
    .Y(_08880_));
 AO21x1_ASAP7_75t_R _17170_ (.A1(_08879_),
    .A2(_08880_),
    .B(_08578_),
    .Y(_08881_));
 NOR2x1_ASAP7_75t_R _17171_ (.A(_08878_),
    .B(_08881_),
    .Y(_08882_));
 AO21x1_ASAP7_75t_R _17172_ (.A1(_08684_),
    .A2(_08588_),
    .B(_08421_),
    .Y(_08883_));
 AO21x1_ASAP7_75t_R _17173_ (.A1(_08572_),
    .A2(_08497_),
    .B(_08563_),
    .Y(_08884_));
 AND3x1_ASAP7_75t_R _17174_ (.A(_08883_),
    .B(_08884_),
    .C(_08466_),
    .Y(_08885_));
 NAND2x1_ASAP7_75t_R _17175_ (.A(_08531_),
    .B(_08533_),
    .Y(_08886_));
 AO21x1_ASAP7_75t_R _17176_ (.A1(_08750_),
    .A2(_08886_),
    .B(_08624_),
    .Y(_08887_));
 OAI21x1_ASAP7_75t_R _17177_ (.A1(_08885_),
    .A2(_08887_),
    .B(_00393_),
    .Y(_08888_));
 NOR2x1_ASAP7_75t_R _17178_ (.A(_08882_),
    .B(_08888_),
    .Y(_08889_));
 OA21x2_ASAP7_75t_R _17179_ (.A1(_08552_),
    .A2(_08475_),
    .B(_08478_),
    .Y(_08890_));
 NAND2x1_ASAP7_75t_R _17180_ (.A(_08625_),
    .B(_08770_),
    .Y(_08891_));
 AO21x1_ASAP7_75t_R _17181_ (.A1(_08890_),
    .A2(_08891_),
    .B(_08624_),
    .Y(_08892_));
 NAND2x1_ASAP7_75t_R _17182_ (.A(_08420_),
    .B(_08770_),
    .Y(_08893_));
 AND3x1_ASAP7_75t_R _17183_ (.A(_08893_),
    .B(_08886_),
    .C(_08466_),
    .Y(_08894_));
 OAI21x1_ASAP7_75t_R _17184_ (.A1(_08892_),
    .A2(_08894_),
    .B(_08448_),
    .Y(_08895_));
 INVx1_ASAP7_75t_R _17185_ (.A(_08456_),
    .Y(_08896_));
 AOI21x1_ASAP7_75t_R _17186_ (.A1(_08433_),
    .A2(_08896_),
    .B(_08634_),
    .Y(_08897_));
 AO21x1_ASAP7_75t_R _17187_ (.A1(_08605_),
    .A2(_08433_),
    .B(_00390_),
    .Y(_08898_));
 OA21x2_ASAP7_75t_R _17188_ (.A1(_08582_),
    .A2(_08637_),
    .B(_08528_),
    .Y(_08899_));
 AOI221x1_ASAP7_75t_R _17189_ (.A1(_00391_),
    .A2(_08897_),
    .B1(_08898_),
    .B2(_08899_),
    .C(_08508_),
    .Y(_08900_));
 OAI21x1_ASAP7_75t_R _17190_ (.A1(_08895_),
    .A2(_08900_),
    .B(_00394_),
    .Y(_08901_));
 OAI22x1_ASAP7_75t_R _17191_ (.A1(_08867_),
    .A2(_08876_),
    .B1(_08889_),
    .B2(_08901_),
    .Y(_00006_));
 AO21x1_ASAP7_75t_R _17192_ (.A1(_08593_),
    .A2(_08758_),
    .B(_08857_),
    .Y(_08902_));
 NAND2x1_ASAP7_75t_R _17193_ (.A(_08624_),
    .B(_08902_),
    .Y(_08903_));
 OA21x2_ASAP7_75t_R _17194_ (.A1(_08654_),
    .A2(_07990_),
    .B(_08883_),
    .Y(_08904_));
 AOI21x1_ASAP7_75t_R _17195_ (.A1(_08903_),
    .A2(_08904_),
    .B(_00391_),
    .Y(_08905_));
 AND2x2_ASAP7_75t_R _17196_ (.A(_08737_),
    .B(_08589_),
    .Y(_08906_));
 AND3x1_ASAP7_75t_R _17197_ (.A(_08461_),
    .B(_08482_),
    .C(_08518_),
    .Y(_08907_));
 OAI21x1_ASAP7_75t_R _17198_ (.A1(_08482_),
    .A2(_08479_),
    .B(_07990_),
    .Y(_08908_));
 AO21x1_ASAP7_75t_R _17199_ (.A1(_08429_),
    .A2(_08801_),
    .B(_08908_),
    .Y(_08909_));
 OAI21x1_ASAP7_75t_R _17200_ (.A1(_08907_),
    .A2(_08909_),
    .B(_00391_),
    .Y(_08910_));
 OAI21x1_ASAP7_75t_R _17201_ (.A1(_08906_),
    .A2(_08910_),
    .B(_00393_),
    .Y(_08911_));
 NOR2x1_ASAP7_75t_R _17202_ (.A(_08905_),
    .B(_08911_),
    .Y(_08912_));
 OA211x2_ASAP7_75t_R _17203_ (.A1(_08431_),
    .A2(_08696_),
    .B(_08535_),
    .C(_08519_),
    .Y(_08913_));
 AO21x1_ASAP7_75t_R _17204_ (.A1(_08441_),
    .A2(_08580_),
    .B(_08435_),
    .Y(_08914_));
 AO21x1_ASAP7_75t_R _17205_ (.A1(_08914_),
    .A2(_08418_),
    .B(_08624_),
    .Y(_08915_));
 OAI21x1_ASAP7_75t_R _17206_ (.A1(_08913_),
    .A2(_08915_),
    .B(_08448_),
    .Y(_08916_));
 AO21x1_ASAP7_75t_R _17207_ (.A1(_08625_),
    .A2(_08457_),
    .B(_08474_),
    .Y(_08917_));
 OA21x2_ASAP7_75t_R _17208_ (.A1(_00390_),
    .A2(net803),
    .B(_08443_),
    .Y(_08918_));
 AOI21x1_ASAP7_75t_R _17209_ (.A1(_08432_),
    .A2(_08839_),
    .B(_08647_),
    .Y(_08919_));
 AOI211x1_ASAP7_75t_R _17210_ (.A1(_08917_),
    .A2(_08918_),
    .B(_08919_),
    .C(_08508_),
    .Y(_08920_));
 OAI21x1_ASAP7_75t_R _17211_ (.A1(_08916_),
    .A2(_08920_),
    .B(_08511_),
    .Y(_08921_));
 NOR2x1_ASAP7_75t_R _17212_ (.A(_08493_),
    .B(_08563_),
    .Y(_08922_));
 AO21x1_ASAP7_75t_R _17213_ (.A1(_08573_),
    .A2(_08695_),
    .B(_08000_),
    .Y(_08923_));
 OAI21x1_ASAP7_75t_R _17214_ (.A1(_08922_),
    .A2(_08923_),
    .B(_07990_),
    .Y(_08924_));
 AO21x1_ASAP7_75t_R _17215_ (.A1(_08799_),
    .A2(_08760_),
    .B(_08924_),
    .Y(_08925_));
 OA21x2_ASAP7_75t_R _17216_ (.A1(_08543_),
    .A2(_08484_),
    .B(_08573_),
    .Y(_08926_));
 OA21x2_ASAP7_75t_R _17217_ (.A1(_08786_),
    .A2(_08926_),
    .B(_08507_),
    .Y(_08927_));
 AND3x1_ASAP7_75t_R _17218_ (.A(_08682_),
    .B(_07955_),
    .C(_08657_),
    .Y(_08928_));
 NOR2x1_ASAP7_75t_R _17219_ (.A(_08651_),
    .B(_08928_),
    .Y(_08929_));
 NAND2x1_ASAP7_75t_R _17220_ (.A(_08614_),
    .B(_08929_),
    .Y(_08930_));
 AOI21x1_ASAP7_75t_R _17221_ (.A1(_08927_),
    .A2(_08930_),
    .B(_08445_),
    .Y(_08931_));
 NAND2x1_ASAP7_75t_R _17222_ (.A(_08925_),
    .B(_08931_),
    .Y(_08932_));
 OA21x2_ASAP7_75t_R _17223_ (.A1(_08605_),
    .A2(_08421_),
    .B(_08479_),
    .Y(_08933_));
 AOI21x1_ASAP7_75t_R _17224_ (.A1(_15735_),
    .A2(_08801_),
    .B(_08001_),
    .Y(_08934_));
 AOI21x1_ASAP7_75t_R _17225_ (.A1(_08933_),
    .A2(_08934_),
    .B(_07990_),
    .Y(_08935_));
 OA21x2_ASAP7_75t_R _17226_ (.A1(_01123_),
    .A2(_08421_),
    .B(_08478_),
    .Y(_08936_));
 NAND2x1_ASAP7_75t_R _17227_ (.A(_08936_),
    .B(_08879_),
    .Y(_08937_));
 AOI21x1_ASAP7_75t_R _17228_ (.A1(_08935_),
    .A2(_08937_),
    .B(_08448_),
    .Y(_08938_));
 AND3x1_ASAP7_75t_R _17229_ (.A(_08502_),
    .B(_08474_),
    .C(_08432_),
    .Y(_08939_));
 NAND2x1_ASAP7_75t_R _17230_ (.A(_08535_),
    .B(_08744_),
    .Y(_08940_));
 AO21x1_ASAP7_75t_R _17231_ (.A1(_08475_),
    .A2(_08433_),
    .B(_08482_),
    .Y(_08941_));
 AO21x1_ASAP7_75t_R _17232_ (.A1(_08572_),
    .A2(_08479_),
    .B(_07955_),
    .Y(_08942_));
 AND2x2_ASAP7_75t_R _17233_ (.A(_08942_),
    .B(_08465_),
    .Y(_08943_));
 AOI21x1_ASAP7_75t_R _17234_ (.A1(_08941_),
    .A2(_08943_),
    .B(_08578_),
    .Y(_08944_));
 OAI21x1_ASAP7_75t_R _17235_ (.A1(_08939_),
    .A2(_08940_),
    .B(_08944_),
    .Y(_08945_));
 AOI21x1_ASAP7_75t_R _17236_ (.A1(_08938_),
    .A2(_08945_),
    .B(_08511_),
    .Y(_08946_));
 NAND2x1_ASAP7_75t_R _17237_ (.A(_08932_),
    .B(_08946_),
    .Y(_08947_));
 OAI21x1_ASAP7_75t_R _17238_ (.A1(_08912_),
    .A2(_08921_),
    .B(_08947_),
    .Y(_00007_));
 INVx8_ASAP7_75t_R _17239_ (.A(_15753_),
    .Y(_15747_));
 CKINVDCx6p67_ASAP7_75t_R _17240_ (.A(_08119_),
    .Y(_08948_));
 BUFx12f_ASAP7_75t_R _17241_ (.A(_08948_),
    .Y(_15758_));
 BUFx12f_ASAP7_75t_R _17242_ (.A(_08119_),
    .Y(_08949_));
 NOR2x2_ASAP7_75t_R _17243_ (.A(_01129_),
    .B(_08949_),
    .Y(_08950_));
 INVx3_ASAP7_75t_R _17244_ (.A(_08950_),
    .Y(_08951_));
 NOR2x2_ASAP7_75t_R _17245_ (.A(net554),
    .B(_08948_),
    .Y(_08952_));
 INVx3_ASAP7_75t_R _17246_ (.A(_08952_),
    .Y(_08953_));
 INVx4_ASAP7_75t_R _17247_ (.A(_08126_),
    .Y(_08954_));
 INVx3_ASAP7_75t_R _17248_ (.A(_01061_),
    .Y(_08955_));
 XOR2x1_ASAP7_75t_R _17249_ (.A(_08122_),
    .Y(_08956_),
    .B(_08955_));
 NOR2x1_ASAP7_75t_R _17250_ (.A(_08124_),
    .B(_08956_),
    .Y(_08957_));
 INVx1_ASAP7_75t_R _17251_ (.A(_08124_),
    .Y(_08958_));
 NOR2x1_ASAP7_75t_R _17252_ (.A(_08958_),
    .B(_08123_),
    .Y(_08959_));
 OAI21x1_ASAP7_75t_R _17253_ (.A1(_08957_),
    .A2(_08959_),
    .B(_07956_),
    .Y(_08960_));
 NAND2x2_ASAP7_75t_R _17254_ (.A(_08954_),
    .B(_08960_),
    .Y(_08961_));
 BUFx4f_ASAP7_75t_R _17255_ (.A(_08961_),
    .Y(_08962_));
 AO21x1_ASAP7_75t_R _17256_ (.A1(_08951_),
    .A2(_08953_),
    .B(_08962_),
    .Y(_08963_));
 NAND2x2_ASAP7_75t_R _17257_ (.A(net944),
    .B(_15758_),
    .Y(_08964_));
 NAND2x2_ASAP7_75t_R _17258_ (.A(_08949_),
    .B(_15748_),
    .Y(_08965_));
 BUFx4f_ASAP7_75t_R _17259_ (.A(_08965_),
    .Y(_08966_));
 BUFx4f_ASAP7_75t_R _17260_ (.A(_08128_),
    .Y(_08967_));
 AO21x1_ASAP7_75t_R _17261_ (.A1(_08964_),
    .A2(_08966_),
    .B(_08967_),
    .Y(_08968_));
 INVx4_ASAP7_75t_R _17262_ (.A(_08136_),
    .Y(_08969_));
 BUFx4f_ASAP7_75t_R _17263_ (.A(_08969_),
    .Y(_08970_));
 AO21x1_ASAP7_75t_R _17264_ (.A1(_08963_),
    .A2(_08968_),
    .B(_08970_),
    .Y(_08971_));
 AO21x2_ASAP7_75t_R _17265_ (.A1(_08118_),
    .A2(_08114_),
    .B(_01130_),
    .Y(_08972_));
 AO21x1_ASAP7_75t_R _17266_ (.A1(_08964_),
    .A2(_08972_),
    .B(_08962_),
    .Y(_08973_));
 NOR2x2_ASAP7_75t_R _17267_ (.A(_08949_),
    .B(_15748_),
    .Y(_08974_));
 INVx1_ASAP7_75t_R _17268_ (.A(_08974_),
    .Y(_08975_));
 BUFx4f_ASAP7_75t_R _17269_ (.A(_08961_),
    .Y(_08976_));
 NAND2x1_ASAP7_75t_R _17270_ (.A(_08975_),
    .B(_08976_),
    .Y(_08977_));
 BUFx4f_ASAP7_75t_R _17271_ (.A(_08136_),
    .Y(_08978_));
 AO21x1_ASAP7_75t_R _17272_ (.A1(_08973_),
    .A2(_08977_),
    .B(_08978_),
    .Y(_08979_));
 BUFx10_ASAP7_75t_R _17273_ (.A(_08144_),
    .Y(_08980_));
 AOI21x1_ASAP7_75t_R _17274_ (.A1(_08971_),
    .A2(_08979_),
    .B(_08980_),
    .Y(_08981_));
 NAND2x2_ASAP7_75t_R _17275_ (.A(_08948_),
    .B(_15748_),
    .Y(_08982_));
 INVx4_ASAP7_75t_R _17276_ (.A(_00466_),
    .Y(_08983_));
 AO21x2_ASAP7_75t_R _17277_ (.A1(_08118_),
    .A2(_08114_),
    .B(_08983_),
    .Y(_08984_));
 BUFx10_ASAP7_75t_R _17278_ (.A(_08961_),
    .Y(_08985_));
 AO21x2_ASAP7_75t_R _17279_ (.A1(_08982_),
    .A2(_08984_),
    .B(_08985_),
    .Y(_08986_));
 AO21x2_ASAP7_75t_R _17280_ (.A1(_08118_),
    .A2(_08114_),
    .B(_01132_),
    .Y(_08987_));
 NAND2x2_ASAP7_75t_R _17281_ (.A(_08948_),
    .B(_15753_),
    .Y(_08988_));
 BUFx4f_ASAP7_75t_R _17282_ (.A(_08988_),
    .Y(_08989_));
 BUFx6f_ASAP7_75t_R _17283_ (.A(_08128_),
    .Y(_08990_));
 AO21x1_ASAP7_75t_R _17284_ (.A1(_08987_),
    .A2(_08989_),
    .B(_08990_),
    .Y(_08991_));
 AO21x1_ASAP7_75t_R _17285_ (.A1(_08986_),
    .A2(_08991_),
    .B(_08978_),
    .Y(_08992_));
 NOR2x2_ASAP7_75t_R _17286_ (.A(_08948_),
    .B(_15753_),
    .Y(_08993_));
 INVx4_ASAP7_75t_R _17287_ (.A(_08993_),
    .Y(_08994_));
 BUFx6f_ASAP7_75t_R _17288_ (.A(_08128_),
    .Y(_08995_));
 AO21x1_ASAP7_75t_R _17289_ (.A1(_08994_),
    .A2(_08964_),
    .B(_08995_),
    .Y(_08996_));
 BUFx4f_ASAP7_75t_R _17290_ (.A(_08982_),
    .Y(_08997_));
 AO21x2_ASAP7_75t_R _17291_ (.A1(_08118_),
    .A2(_08114_),
    .B(_01129_),
    .Y(_08998_));
 BUFx4f_ASAP7_75t_R _17292_ (.A(_08961_),
    .Y(_08999_));
 AO21x1_ASAP7_75t_R _17293_ (.A1(_08997_),
    .A2(_08998_),
    .B(_08999_),
    .Y(_09000_));
 AO21x1_ASAP7_75t_R _17294_ (.A1(_08996_),
    .A2(_09000_),
    .B(_08970_),
    .Y(_09001_));
 AOI21x1_ASAP7_75t_R _17295_ (.A1(_08992_),
    .A2(_09001_),
    .B(_00387_),
    .Y(_09002_));
 OAI21x1_ASAP7_75t_R _17296_ (.A1(_08981_),
    .A2(_09002_),
    .B(_00388_),
    .Y(_09003_));
 INVx1_ASAP7_75t_R _17297_ (.A(_00463_),
    .Y(_09004_));
 AO21x2_ASAP7_75t_R _17298_ (.A1(_08118_),
    .A2(_08114_),
    .B(_09004_),
    .Y(_09005_));
 NAND2x2_ASAP7_75t_R _17299_ (.A(_00464_),
    .B(_15758_),
    .Y(_09006_));
 BUFx4f_ASAP7_75t_R _17300_ (.A(_08961_),
    .Y(_09007_));
 AO21x1_ASAP7_75t_R _17301_ (.A1(_09005_),
    .A2(_09006_),
    .B(_09007_),
    .Y(_09008_));
 NOR2x1_ASAP7_75t_R _17302_ (.A(_08983_),
    .B(_08949_),
    .Y(_09009_));
 INVx2_ASAP7_75t_R _17303_ (.A(_09009_),
    .Y(_09010_));
 BUFx4f_ASAP7_75t_R _17304_ (.A(_08128_),
    .Y(_09011_));
 AO21x1_ASAP7_75t_R _17305_ (.A1(_08953_),
    .A2(_09010_),
    .B(_09011_),
    .Y(_09012_));
 AO21x1_ASAP7_75t_R _17306_ (.A1(_09008_),
    .A2(_09012_),
    .B(_08978_),
    .Y(_09013_));
 NAND2x2_ASAP7_75t_R _17307_ (.A(_15750_),
    .B(net927),
    .Y(_09014_));
 INVx3_ASAP7_75t_R _17308_ (.A(_09014_),
    .Y(_09015_));
 NAND2x2_ASAP7_75t_R _17309_ (.A(_08966_),
    .B(_08985_),
    .Y(_09016_));
 NOR2x2_ASAP7_75t_R _17310_ (.A(_09015_),
    .B(_09016_),
    .Y(_09017_));
 INVx3_ASAP7_75t_R _17311_ (.A(_08965_),
    .Y(_09018_));
 BUFx4f_ASAP7_75t_R _17312_ (.A(_08128_),
    .Y(_09019_));
 OA21x2_ASAP7_75t_R _17313_ (.A1(_09015_),
    .A2(_09018_),
    .B(_09019_),
    .Y(_09020_));
 OAI21x1_ASAP7_75t_R _17314_ (.A1(_09017_),
    .A2(_09020_),
    .B(_00386_),
    .Y(_09021_));
 BUFx10_ASAP7_75t_R _17315_ (.A(_08145_),
    .Y(_09022_));
 NAND3x1_ASAP7_75t_R _17316_ (.A(_09013_),
    .B(_09021_),
    .C(_09022_),
    .Y(_09023_));
 BUFx4f_ASAP7_75t_R _17317_ (.A(_08961_),
    .Y(_09024_));
 OAI21x1_ASAP7_75t_R _17318_ (.A1(_15760_),
    .A2(net927),
    .B(_08953_),
    .Y(_09025_));
 NAND2x1_ASAP7_75t_R _17319_ (.A(_09024_),
    .B(_09025_),
    .Y(_09026_));
 INVx1_ASAP7_75t_R _17320_ (.A(_00465_),
    .Y(_09027_));
 NOR2x2_ASAP7_75t_R _17321_ (.A(_09027_),
    .B(_08949_),
    .Y(_09028_));
 INVx3_ASAP7_75t_R _17322_ (.A(_09028_),
    .Y(_09029_));
 NOR2x1_ASAP7_75t_R _17323_ (.A(_09029_),
    .B(_08985_),
    .Y(_09030_));
 INVx1_ASAP7_75t_R _17324_ (.A(_09030_),
    .Y(_09031_));
 AO21x1_ASAP7_75t_R _17325_ (.A1(_09026_),
    .A2(_09031_),
    .B(_08970_),
    .Y(_09032_));
 BUFx4f_ASAP7_75t_R _17326_ (.A(_08969_),
    .Y(_09033_));
 BUFx10_ASAP7_75t_R _17327_ (.A(_09033_),
    .Y(_09034_));
 AO21x2_ASAP7_75t_R _17328_ (.A1(_08118_),
    .A2(_08114_),
    .B(_09027_),
    .Y(_09035_));
 INVx2_ASAP7_75t_R _17329_ (.A(_09035_),
    .Y(_09036_));
 NOR2x2_ASAP7_75t_R _17330_ (.A(_09036_),
    .B(_08961_),
    .Y(_09037_));
 INVx1_ASAP7_75t_R _17331_ (.A(_09037_),
    .Y(_09038_));
 NOR2x2_ASAP7_75t_R _17332_ (.A(_00464_),
    .B(_15760_),
    .Y(_09039_));
 NOR2x2_ASAP7_75t_R _17333_ (.A(_09004_),
    .B(_08949_),
    .Y(_09040_));
 INVx4_ASAP7_75t_R _17334_ (.A(_09040_),
    .Y(_09041_));
 NAND2x2_ASAP7_75t_R _17335_ (.A(_00464_),
    .B(_08949_),
    .Y(_09042_));
 AO21x1_ASAP7_75t_R _17336_ (.A1(_09041_),
    .A2(_09042_),
    .B(_09011_),
    .Y(_09043_));
 OAI21x1_ASAP7_75t_R _17337_ (.A1(_09038_),
    .A2(_09039_),
    .B(_09043_),
    .Y(_09044_));
 AOI21x1_ASAP7_75t_R _17338_ (.A1(_09034_),
    .A2(_09044_),
    .B(_09022_),
    .Y(_09045_));
 AOI21x1_ASAP7_75t_R _17339_ (.A1(_09032_),
    .A2(_09045_),
    .B(_00388_),
    .Y(_09046_));
 AOI21x1_ASAP7_75t_R _17340_ (.A1(_09023_),
    .A2(_09046_),
    .B(_00389_),
    .Y(_09047_));
 NAND2x2_ASAP7_75t_R _17341_ (.A(_08119_),
    .B(net944),
    .Y(_09048_));
 INVx1_ASAP7_75t_R _17342_ (.A(_09048_),
    .Y(_09049_));
 OA21x2_ASAP7_75t_R _17343_ (.A1(_08974_),
    .A2(_09049_),
    .B(_08999_),
    .Y(_09050_));
 NAND2x1_ASAP7_75t_R _17344_ (.A(_09042_),
    .B(_08982_),
    .Y(_09051_));
 AO21x1_ASAP7_75t_R _17345_ (.A1(_09051_),
    .A2(_08995_),
    .B(_08137_),
    .Y(_09052_));
 NOR2x1_ASAP7_75t_R _17346_ (.A(_09050_),
    .B(_09052_),
    .Y(_09053_));
 INVx1_ASAP7_75t_R _17347_ (.A(_01134_),
    .Y(_09054_));
 NOR2x2_ASAP7_75t_R _17348_ (.A(net553),
    .B(_08119_),
    .Y(_09055_));
 AO21x2_ASAP7_75t_R _17349_ (.A1(_08960_),
    .A2(_08954_),
    .B(_09055_),
    .Y(_09056_));
 OAI21x1_ASAP7_75t_R _17350_ (.A1(_09054_),
    .A2(_09024_),
    .B(_09056_),
    .Y(_09057_));
 BUFx6f_ASAP7_75t_R _17351_ (.A(_08145_),
    .Y(_09058_));
 AO21x1_ASAP7_75t_R _17352_ (.A1(_09057_),
    .A2(_08978_),
    .B(_09058_),
    .Y(_09059_));
 OR2x4_ASAP7_75t_R _17353_ (.A(_01131_),
    .B(_08949_),
    .Y(_09060_));
 NAND2x2_ASAP7_75t_R _17354_ (.A(_09048_),
    .B(_09060_),
    .Y(_09061_));
 NAND2x2_ASAP7_75t_R _17355_ (.A(_08990_),
    .B(_09061_),
    .Y(_09062_));
 INVx2_ASAP7_75t_R _17356_ (.A(_08987_),
    .Y(_09063_));
 AOI21x1_ASAP7_75t_R _17357_ (.A1(_09063_),
    .A2(_08999_),
    .B(_08137_),
    .Y(_09064_));
 BUFx6f_ASAP7_75t_R _17358_ (.A(_08144_),
    .Y(_09065_));
 AOI21x1_ASAP7_75t_R _17359_ (.A1(_09062_),
    .A2(_09064_),
    .B(_09065_),
    .Y(_09066_));
 OAI21x1_ASAP7_75t_R _17360_ (.A1(_09040_),
    .A2(_09049_),
    .B(_08962_),
    .Y(_09067_));
 BUFx6f_ASAP7_75t_R _17361_ (.A(_08136_),
    .Y(_09068_));
 BUFx4f_ASAP7_75t_R _17362_ (.A(_08128_),
    .Y(_09069_));
 NAND2x1_ASAP7_75t_R _17363_ (.A(_09063_),
    .B(_09069_),
    .Y(_09070_));
 NAND3x1_ASAP7_75t_R _17364_ (.A(_09067_),
    .B(_09068_),
    .C(_09070_),
    .Y(_09071_));
 BUFx10_ASAP7_75t_R _17365_ (.A(_08153_),
    .Y(_09072_));
 AOI21x1_ASAP7_75t_R _17366_ (.A1(_09066_),
    .A2(_09071_),
    .B(_09072_),
    .Y(_09073_));
 OAI21x1_ASAP7_75t_R _17367_ (.A1(_09053_),
    .A2(_09059_),
    .B(_09073_),
    .Y(_09074_));
 AO21x1_ASAP7_75t_R _17368_ (.A1(_08966_),
    .A2(_09041_),
    .B(_08976_),
    .Y(_09075_));
 BUFx4f_ASAP7_75t_R _17369_ (.A(_08961_),
    .Y(_09076_));
 AO21x1_ASAP7_75t_R _17370_ (.A1(net927),
    .A2(_15760_),
    .B(_09028_),
    .Y(_09077_));
 BUFx4f_ASAP7_75t_R _17371_ (.A(_08136_),
    .Y(_09078_));
 AOI21x1_ASAP7_75t_R _17372_ (.A1(_09076_),
    .A2(_09077_),
    .B(_09078_),
    .Y(_09079_));
 NAND2x1_ASAP7_75t_R _17373_ (.A(_09075_),
    .B(_09079_),
    .Y(_09080_));
 AO21x1_ASAP7_75t_R _17374_ (.A1(_08987_),
    .A2(_09006_),
    .B(_09019_),
    .Y(_09081_));
 INVx1_ASAP7_75t_R _17375_ (.A(_01130_),
    .Y(_09082_));
 NOR2x2_ASAP7_75t_R _17376_ (.A(_09082_),
    .B(_15758_),
    .Y(_09083_));
 OA21x2_ASAP7_75t_R _17377_ (.A1(_08976_),
    .A2(_09083_),
    .B(_09078_),
    .Y(_09084_));
 AOI21x1_ASAP7_75t_R _17378_ (.A1(_09081_),
    .A2(_09084_),
    .B(_09065_),
    .Y(_09085_));
 CKINVDCx5p33_ASAP7_75t_R _17379_ (.A(_08153_),
    .Y(_09086_));
 AOI21x1_ASAP7_75t_R _17380_ (.A1(_09080_),
    .A2(_09085_),
    .B(_09086_),
    .Y(_09087_));
 NOR2x2_ASAP7_75t_R _17381_ (.A(_01130_),
    .B(_08119_),
    .Y(_09088_));
 INVx4_ASAP7_75t_R _17382_ (.A(_09088_),
    .Y(_09089_));
 OAI21x1_ASAP7_75t_R _17383_ (.A1(_00385_),
    .A2(_09089_),
    .B(_08986_),
    .Y(_09090_));
 AO21x2_ASAP7_75t_R _17384_ (.A1(_08118_),
    .A2(_08114_),
    .B(_01131_),
    .Y(_09091_));
 AO21x2_ASAP7_75t_R _17385_ (.A1(_09089_),
    .A2(_09091_),
    .B(_08128_),
    .Y(_09092_));
 BUFx6f_ASAP7_75t_R _17386_ (.A(_08969_),
    .Y(_09093_));
 NOR2x1_ASAP7_75t_R _17387_ (.A(_09093_),
    .B(_09037_),
    .Y(_09094_));
 AOI21x1_ASAP7_75t_R _17388_ (.A1(_09092_),
    .A2(_09094_),
    .B(_08145_),
    .Y(_09095_));
 OAI21x1_ASAP7_75t_R _17389_ (.A1(_00386_),
    .A2(_09090_),
    .B(_09095_),
    .Y(_09096_));
 NAND2x1_ASAP7_75t_R _17390_ (.A(_09087_),
    .B(_09096_),
    .Y(_09097_));
 INVx8_ASAP7_75t_R _17391_ (.A(_00389_),
    .Y(_09098_));
 AOI21x1_ASAP7_75t_R _17392_ (.A1(_09074_),
    .A2(_09097_),
    .B(_09098_),
    .Y(_09099_));
 AOI21x1_ASAP7_75t_R _17393_ (.A1(_09003_),
    .A2(_09047_),
    .B(_09099_),
    .Y(_00008_));
 BUFx4f_ASAP7_75t_R _17394_ (.A(_09035_),
    .Y(_09100_));
 AO21x1_ASAP7_75t_R _17395_ (.A1(_09100_),
    .A2(_09089_),
    .B(_09007_),
    .Y(_09101_));
 NAND2x1_ASAP7_75t_R _17396_ (.A(_08999_),
    .B(_09051_),
    .Y(_09102_));
 BUFx6f_ASAP7_75t_R _17397_ (.A(_08969_),
    .Y(_09103_));
 AO21x1_ASAP7_75t_R _17398_ (.A1(_09101_),
    .A2(_09102_),
    .B(_09103_),
    .Y(_09104_));
 NAND2x2_ASAP7_75t_R _17399_ (.A(_15748_),
    .B(_15747_),
    .Y(_09105_));
 NAND2x2_ASAP7_75t_R _17400_ (.A(_08949_),
    .B(_15750_),
    .Y(_09106_));
 AO21x1_ASAP7_75t_R _17401_ (.A1(_09105_),
    .A2(_09106_),
    .B(_09007_),
    .Y(_09107_));
 AO21x1_ASAP7_75t_R _17402_ (.A1(_08966_),
    .A2(_09029_),
    .B(_08995_),
    .Y(_09108_));
 AO21x1_ASAP7_75t_R _17403_ (.A1(_09107_),
    .A2(_09108_),
    .B(_08978_),
    .Y(_09109_));
 AOI21x1_ASAP7_75t_R _17404_ (.A1(_09104_),
    .A2(_09109_),
    .B(_09022_),
    .Y(_09110_));
 NAND2x2_ASAP7_75t_R _17405_ (.A(_08949_),
    .B(_15753_),
    .Y(_09111_));
 INVx1_ASAP7_75t_R _17406_ (.A(_01129_),
    .Y(_09112_));
 NOR2x2_ASAP7_75t_R _17407_ (.A(_09112_),
    .B(_15760_),
    .Y(_09113_));
 NOR2x2_ASAP7_75t_R _17408_ (.A(_09113_),
    .B(_08985_),
    .Y(_09114_));
 AOI21x1_ASAP7_75t_R _17409_ (.A1(_09111_),
    .A2(_09114_),
    .B(_09093_),
    .Y(_09115_));
 OA21x2_ASAP7_75t_R _17410_ (.A1(_00385_),
    .A2(_08984_),
    .B(_09115_),
    .Y(_09116_));
 AO21x1_ASAP7_75t_R _17411_ (.A1(_09035_),
    .A2(_09010_),
    .B(_08985_),
    .Y(_09117_));
 OAI21x1_ASAP7_75t_R _17412_ (.A1(_00385_),
    .A2(_08972_),
    .B(_09117_),
    .Y(_09118_));
 OAI21x1_ASAP7_75t_R _17413_ (.A1(_00386_),
    .A2(_09118_),
    .B(_09022_),
    .Y(_09119_));
 OAI21x1_ASAP7_75t_R _17414_ (.A1(_09116_),
    .A2(_09119_),
    .B(_00388_),
    .Y(_09120_));
 NOR2x1_ASAP7_75t_R _17415_ (.A(_09110_),
    .B(_09120_),
    .Y(_09121_));
 BUFx6f_ASAP7_75t_R _17416_ (.A(_08985_),
    .Y(_09122_));
 INVx2_ASAP7_75t_R _17417_ (.A(_09111_),
    .Y(_09123_));
 AND3x2_ASAP7_75t_R _17418_ (.A(_08960_),
    .B(_00469_),
    .C(_08954_),
    .Y(_09124_));
 AO21x1_ASAP7_75t_R _17419_ (.A1(_08962_),
    .A2(_09088_),
    .B(_09093_),
    .Y(_09125_));
 AOI211x1_ASAP7_75t_R _17420_ (.A1(_09122_),
    .A2(_09123_),
    .B(_09124_),
    .C(_09125_),
    .Y(_09126_));
 NAND2x2_ASAP7_75t_R _17421_ (.A(_09048_),
    .B(_09089_),
    .Y(_09127_));
 NAND2x1_ASAP7_75t_R _17422_ (.A(_09127_),
    .B(_08985_),
    .Y(_09128_));
 AND2x2_ASAP7_75t_R _17423_ (.A(_09128_),
    .B(_09093_),
    .Y(_09129_));
 INVx3_ASAP7_75t_R _17424_ (.A(_09055_),
    .Y(_09130_));
 NAND2x1_ASAP7_75t_R _17425_ (.A(_08998_),
    .B(_09130_),
    .Y(_09131_));
 NAND2x1_ASAP7_75t_R _17426_ (.A(_08995_),
    .B(_09131_),
    .Y(_09132_));
 AO21x1_ASAP7_75t_R _17427_ (.A1(_09129_),
    .A2(_09132_),
    .B(_09058_),
    .Y(_09133_));
 BUFx6f_ASAP7_75t_R _17428_ (.A(_09086_),
    .Y(_09134_));
 OAI21x1_ASAP7_75t_R _17429_ (.A1(_09126_),
    .A2(_09133_),
    .B(_09134_),
    .Y(_09135_));
 OA21x2_ASAP7_75t_R _17430_ (.A1(_08976_),
    .A2(_08964_),
    .B(_08969_),
    .Y(_09136_));
 OR3x1_ASAP7_75t_R _17431_ (.A(_09015_),
    .B(_09069_),
    .C(_08993_),
    .Y(_09137_));
 AO21x1_ASAP7_75t_R _17432_ (.A1(_08997_),
    .A2(_08953_),
    .B(_09122_),
    .Y(_09138_));
 AO21x1_ASAP7_75t_R _17433_ (.A1(_08960_),
    .A2(_08954_),
    .B(_09083_),
    .Y(_09139_));
 INVx1_ASAP7_75t_R _17434_ (.A(_08997_),
    .Y(_09140_));
 BUFx6f_ASAP7_75t_R _17435_ (.A(_08136_),
    .Y(_09141_));
 OA21x2_ASAP7_75t_R _17436_ (.A1(_09139_),
    .A2(_09140_),
    .B(_09141_),
    .Y(_09142_));
 AOI221x1_ASAP7_75t_R _17437_ (.A1(_09136_),
    .A2(_09137_),
    .B1(_09138_),
    .B2(_09142_),
    .C(_08980_),
    .Y(_09143_));
 OAI21x1_ASAP7_75t_R _17438_ (.A1(_09135_),
    .A2(_09143_),
    .B(_00389_),
    .Y(_09144_));
 AO21x1_ASAP7_75t_R _17439_ (.A1(_08997_),
    .A2(_08987_),
    .B(_09069_),
    .Y(_09145_));
 AO21x1_ASAP7_75t_R _17440_ (.A1(_09042_),
    .A2(_09130_),
    .B(_09076_),
    .Y(_09146_));
 AOI21x1_ASAP7_75t_R _17441_ (.A1(_09145_),
    .A2(_09146_),
    .B(_09103_),
    .Y(_09147_));
 AO21x1_ASAP7_75t_R _17442_ (.A1(_09106_),
    .A2(_09006_),
    .B(_09069_),
    .Y(_09148_));
 NOR2x2_ASAP7_75t_R _17443_ (.A(_09083_),
    .B(_08961_),
    .Y(_09149_));
 NAND2x1_ASAP7_75t_R _17444_ (.A(_08989_),
    .B(_09149_),
    .Y(_09150_));
 AOI21x1_ASAP7_75t_R _17445_ (.A1(_09148_),
    .A2(_09150_),
    .B(_09141_),
    .Y(_09151_));
 OAI21x1_ASAP7_75t_R _17446_ (.A1(_09147_),
    .A2(_09151_),
    .B(_09058_),
    .Y(_09152_));
 AO21x1_ASAP7_75t_R _17447_ (.A1(_08997_),
    .A2(_08984_),
    .B(_08967_),
    .Y(_09153_));
 NOR2x1_ASAP7_75t_R _17448_ (.A(_09078_),
    .B(_09037_),
    .Y(_09154_));
 AOI21x1_ASAP7_75t_R _17449_ (.A1(_09153_),
    .A2(_09154_),
    .B(_08145_),
    .Y(_09155_));
 INVx1_ASAP7_75t_R _17450_ (.A(_01132_),
    .Y(_09156_));
 NAND2x2_ASAP7_75t_R _17451_ (.A(_09156_),
    .B(_08948_),
    .Y(_09157_));
 AO21x1_ASAP7_75t_R _17452_ (.A1(_08998_),
    .A2(_09157_),
    .B(_09019_),
    .Y(_09158_));
 NAND3x1_ASAP7_75t_R _17453_ (.A(_09117_),
    .B(_09158_),
    .C(_09068_),
    .Y(_09159_));
 AOI21x1_ASAP7_75t_R _17454_ (.A1(_09155_),
    .A2(_09159_),
    .B(_09086_),
    .Y(_09160_));
 NAND2x1_ASAP7_75t_R _17455_ (.A(_09152_),
    .B(_09160_),
    .Y(_09161_));
 AOI21x1_ASAP7_75t_R _17456_ (.A1(_08988_),
    .A2(_09106_),
    .B(_08967_),
    .Y(_09162_));
 AO21x1_ASAP7_75t_R _17457_ (.A1(_08989_),
    .A2(_09149_),
    .B(_09162_),
    .Y(_09163_));
 AO21x1_ASAP7_75t_R _17458_ (.A1(_08966_),
    .A2(_09006_),
    .B(_09019_),
    .Y(_09164_));
 BUFx6f_ASAP7_75t_R _17459_ (.A(_08128_),
    .Y(_09165_));
 NAND2x1_ASAP7_75t_R _17460_ (.A(_08984_),
    .B(_08964_),
    .Y(_09166_));
 AOI21x1_ASAP7_75t_R _17461_ (.A1(_09165_),
    .A2(_09166_),
    .B(_08144_),
    .Y(_09167_));
 AOI21x1_ASAP7_75t_R _17462_ (.A1(_09164_),
    .A2(_09167_),
    .B(_09103_),
    .Y(_09168_));
 OAI21x1_ASAP7_75t_R _17463_ (.A1(_09022_),
    .A2(_09163_),
    .B(_09168_),
    .Y(_09169_));
 INVx1_ASAP7_75t_R _17464_ (.A(_00468_),
    .Y(_09170_));
 BUFx4f_ASAP7_75t_R _17465_ (.A(_08961_),
    .Y(_09171_));
 NOR2x1_ASAP7_75t_R _17466_ (.A(_09170_),
    .B(_09171_),
    .Y(_09172_));
 INVx1_ASAP7_75t_R _17467_ (.A(_08984_),
    .Y(_09173_));
 OA21x2_ASAP7_75t_R _17468_ (.A1(_09173_),
    .A2(_09040_),
    .B(_08985_),
    .Y(_09174_));
 AO21x1_ASAP7_75t_R _17469_ (.A1(_08144_),
    .A2(_09172_),
    .B(_09174_),
    .Y(_09175_));
 AOI21x1_ASAP7_75t_R _17470_ (.A1(_09034_),
    .A2(_09175_),
    .B(_09072_),
    .Y(_09176_));
 AOI21x1_ASAP7_75t_R _17471_ (.A1(_09169_),
    .A2(_09176_),
    .B(_00389_),
    .Y(_09177_));
 NAND2x2_ASAP7_75t_R _17472_ (.A(_09161_),
    .B(_09177_),
    .Y(_09178_));
 OAI21x1_ASAP7_75t_R _17473_ (.A1(_09121_),
    .A2(_09144_),
    .B(_09178_),
    .Y(_00009_));
 AO21x1_ASAP7_75t_R _17474_ (.A1(_09111_),
    .A2(_08964_),
    .B(_09076_),
    .Y(_09179_));
 AO21x1_ASAP7_75t_R _17475_ (.A1(_08951_),
    .A2(_08972_),
    .B(_08967_),
    .Y(_09180_));
 AO21x1_ASAP7_75t_R _17476_ (.A1(_09179_),
    .A2(_09180_),
    .B(_09103_),
    .Y(_09181_));
 OAI21x1_ASAP7_75t_R _17477_ (.A1(_09122_),
    .A2(_09127_),
    .B(_09079_),
    .Y(_09182_));
 NAND3x1_ASAP7_75t_R _17478_ (.A(_09181_),
    .B(_09182_),
    .C(_09134_),
    .Y(_09183_));
 INVx2_ASAP7_75t_R _17479_ (.A(_09091_),
    .Y(_09184_));
 AO21x1_ASAP7_75t_R _17480_ (.A1(_08999_),
    .A2(_08950_),
    .B(_09033_),
    .Y(_09185_));
 NAND2x1_ASAP7_75t_R _17481_ (.A(_01130_),
    .B(_15758_),
    .Y(_09186_));
 AND3x1_ASAP7_75t_R _17482_ (.A(_08995_),
    .B(_09106_),
    .C(_09186_),
    .Y(_09187_));
 AOI211x1_ASAP7_75t_R _17483_ (.A1(_09122_),
    .A2(_09184_),
    .B(_09185_),
    .C(_09187_),
    .Y(_09188_));
 AO21x1_ASAP7_75t_R _17484_ (.A1(_08994_),
    .A2(_09089_),
    .B(_09007_),
    .Y(_09189_));
 AND3x1_ASAP7_75t_R _17485_ (.A(_09189_),
    .B(_09103_),
    .C(_09092_),
    .Y(_09190_));
 OAI21x1_ASAP7_75t_R _17486_ (.A1(_09188_),
    .A2(_09190_),
    .B(_00388_),
    .Y(_09191_));
 AOI21x1_ASAP7_75t_R _17487_ (.A1(_09183_),
    .A2(_09191_),
    .B(_00387_),
    .Y(_09192_));
 AO21x1_ASAP7_75t_R _17488_ (.A1(net927),
    .A2(_15758_),
    .B(_08952_),
    .Y(_09193_));
 INVx1_ASAP7_75t_R _17489_ (.A(_09157_),
    .Y(_09194_));
 OA21x2_ASAP7_75t_R _17490_ (.A1(_09018_),
    .A2(_09194_),
    .B(_09165_),
    .Y(_09195_));
 AOI211x1_ASAP7_75t_R _17491_ (.A1(_09122_),
    .A2(_09193_),
    .B(_09195_),
    .C(_08970_),
    .Y(_09196_));
 NOR2x2_ASAP7_75t_R _17492_ (.A(net945),
    .B(_15760_),
    .Y(_09197_));
 NOR2x1_ASAP7_75t_R _17493_ (.A(_09197_),
    .B(_08128_),
    .Y(_09198_));
 NOR2x1_ASAP7_75t_R _17494_ (.A(_09068_),
    .B(_09198_),
    .Y(_09199_));
 AO21x1_ASAP7_75t_R _17495_ (.A1(_08998_),
    .A2(_09010_),
    .B(_08999_),
    .Y(_09200_));
 AO21x1_ASAP7_75t_R _17496_ (.A1(_09199_),
    .A2(_09200_),
    .B(_08153_),
    .Y(_09201_));
 OAI21x1_ASAP7_75t_R _17497_ (.A1(_09196_),
    .A2(_09201_),
    .B(_00387_),
    .Y(_09202_));
 AND3x1_ASAP7_75t_R _17498_ (.A(_09165_),
    .B(_09100_),
    .C(_09130_),
    .Y(_09203_));
 NAND2x2_ASAP7_75t_R _17499_ (.A(_01131_),
    .B(_15758_),
    .Y(_09204_));
 AND3x1_ASAP7_75t_R _17500_ (.A(_09007_),
    .B(_09106_),
    .C(_09204_),
    .Y(_09205_));
 OAI21x1_ASAP7_75t_R _17501_ (.A1(_09203_),
    .A2(_09205_),
    .B(_09034_),
    .Y(_09206_));
 NOR2x1_ASAP7_75t_R _17502_ (.A(_09184_),
    .B(_09024_),
    .Y(_09207_));
 OAI21x1_ASAP7_75t_R _17503_ (.A1(_08950_),
    .A2(_09016_),
    .B(_09068_),
    .Y(_09208_));
 AO21x1_ASAP7_75t_R _17504_ (.A1(_08989_),
    .A2(_09207_),
    .B(_09208_),
    .Y(_09209_));
 AOI21x1_ASAP7_75t_R _17505_ (.A1(_09206_),
    .A2(_09209_),
    .B(_09134_),
    .Y(_09210_));
 OAI21x1_ASAP7_75t_R _17506_ (.A1(_09202_),
    .A2(_09210_),
    .B(_09098_),
    .Y(_09211_));
 AO21x1_ASAP7_75t_R _17507_ (.A1(_08994_),
    .A2(_09006_),
    .B(_09011_),
    .Y(_09212_));
 AO21x1_ASAP7_75t_R _17508_ (.A1(_09005_),
    .A2(_09130_),
    .B(_09171_),
    .Y(_09213_));
 AND3x1_ASAP7_75t_R _17509_ (.A(_09212_),
    .B(_09141_),
    .C(_09213_),
    .Y(_09214_));
 NOR2x1_ASAP7_75t_R _17510_ (.A(_09170_),
    .B(_00385_),
    .Y(_09215_));
 NAND2x1_ASAP7_75t_R _17511_ (.A(_09019_),
    .B(_08994_),
    .Y(_09216_));
 OAI21x1_ASAP7_75t_R _17512_ (.A1(_09015_),
    .A2(_09216_),
    .B(_09033_),
    .Y(_09217_));
 OAI21x1_ASAP7_75t_R _17513_ (.A1(_09215_),
    .A2(_09217_),
    .B(_09072_),
    .Y(_09218_));
 OA21x2_ASAP7_75t_R _17514_ (.A1(_09069_),
    .A2(_01133_),
    .B(_09078_),
    .Y(_09219_));
 AOI21x1_ASAP7_75t_R _17515_ (.A1(_09219_),
    .A2(_09179_),
    .B(_08153_),
    .Y(_09220_));
 INVx1_ASAP7_75t_R _17516_ (.A(_00470_),
    .Y(_09221_));
 NOR2x1_ASAP7_75t_R _17517_ (.A(_09221_),
    .B(_08985_),
    .Y(_09222_));
 OR3x1_ASAP7_75t_R _17518_ (.A(_09222_),
    .B(_08137_),
    .C(_09198_),
    .Y(_09223_));
 AOI21x1_ASAP7_75t_R _17519_ (.A1(_09220_),
    .A2(_09223_),
    .B(_09022_),
    .Y(_09224_));
 OAI21x1_ASAP7_75t_R _17520_ (.A1(_09214_),
    .A2(_09218_),
    .B(_09224_),
    .Y(_09225_));
 AO21x1_ASAP7_75t_R _17521_ (.A1(_01133_),
    .A2(_08966_),
    .B(_09076_),
    .Y(_09226_));
 OAI21x1_ASAP7_75t_R _17522_ (.A1(_08993_),
    .A2(_09056_),
    .B(_09226_),
    .Y(_09227_));
 AO21x1_ASAP7_75t_R _17523_ (.A1(_09130_),
    .A2(_09048_),
    .B(_09171_),
    .Y(_09228_));
 AO21x1_ASAP7_75t_R _17524_ (.A1(_08960_),
    .A2(_08954_),
    .B(_01134_),
    .Y(_09229_));
 AND2x2_ASAP7_75t_R _17525_ (.A(_09229_),
    .B(_08969_),
    .Y(_09230_));
 AOI21x1_ASAP7_75t_R _17526_ (.A1(_09228_),
    .A2(_09230_),
    .B(_09086_),
    .Y(_09231_));
 OAI21x1_ASAP7_75t_R _17527_ (.A1(_09034_),
    .A2(_09227_),
    .B(_09231_),
    .Y(_09232_));
 AO21x1_ASAP7_75t_R _17528_ (.A1(_08953_),
    .A2(_09089_),
    .B(_09171_),
    .Y(_09233_));
 OA21x2_ASAP7_75t_R _17529_ (.A1(_08967_),
    .A2(_09042_),
    .B(_09093_),
    .Y(_09234_));
 AOI21x1_ASAP7_75t_R _17530_ (.A1(_09233_),
    .A2(_09234_),
    .B(_08153_),
    .Y(_09235_));
 AO21x1_ASAP7_75t_R _17531_ (.A1(_09106_),
    .A2(_09010_),
    .B(_09076_),
    .Y(_09236_));
 AO21x1_ASAP7_75t_R _17532_ (.A1(_08984_),
    .A2(_09041_),
    .B(_09069_),
    .Y(_09237_));
 NAND3x1_ASAP7_75t_R _17533_ (.A(_09236_),
    .B(_09237_),
    .C(_09068_),
    .Y(_09238_));
 AOI21x1_ASAP7_75t_R _17534_ (.A1(_09235_),
    .A2(_09238_),
    .B(_08980_),
    .Y(_09239_));
 AOI21x1_ASAP7_75t_R _17535_ (.A1(_09232_),
    .A2(_09239_),
    .B(_09098_),
    .Y(_09240_));
 NAND2x1_ASAP7_75t_R _17536_ (.A(_09225_),
    .B(_09240_),
    .Y(_09241_));
 OAI21x1_ASAP7_75t_R _17537_ (.A1(_09192_),
    .A2(_09211_),
    .B(_09241_),
    .Y(_00010_));
 AO21x1_ASAP7_75t_R _17538_ (.A1(_09111_),
    .A2(_09041_),
    .B(_09011_),
    .Y(_09242_));
 AO21x1_ASAP7_75t_R _17539_ (.A1(_09242_),
    .A2(_09031_),
    .B(_09058_),
    .Y(_09243_));
 AO21x1_ASAP7_75t_R _17540_ (.A1(_08960_),
    .A2(_08954_),
    .B(_09035_),
    .Y(_09244_));
 OA211x2_ASAP7_75t_R _17541_ (.A1(_09065_),
    .A2(_09244_),
    .B(_09070_),
    .C(_09068_),
    .Y(_09245_));
 NAND2x1_ASAP7_75t_R _17542_ (.A(_09243_),
    .B(_09245_),
    .Y(_09246_));
 AO21x1_ASAP7_75t_R _17543_ (.A1(_09106_),
    .A2(_08951_),
    .B(_09007_),
    .Y(_09247_));
 AO21x1_ASAP7_75t_R _17544_ (.A1(_08997_),
    .A2(_08953_),
    .B(_08990_),
    .Y(_09248_));
 AND3x1_ASAP7_75t_R _17545_ (.A(_09247_),
    .B(_09065_),
    .C(_09248_),
    .Y(_09249_));
 AOI211x1_ASAP7_75t_R _17546_ (.A1(_00385_),
    .A2(_09184_),
    .B(_09205_),
    .C(_09065_),
    .Y(_09250_));
 OAI21x1_ASAP7_75t_R _17547_ (.A1(_09249_),
    .A2(_09250_),
    .B(_09034_),
    .Y(_09251_));
 AOI21x1_ASAP7_75t_R _17548_ (.A1(_09246_),
    .A2(_09251_),
    .B(_00388_),
    .Y(_09252_));
 AND3x1_ASAP7_75t_R _17549_ (.A(_08990_),
    .B(_08966_),
    .C(_09204_),
    .Y(_09253_));
 OAI21x1_ASAP7_75t_R _17550_ (.A1(_09174_),
    .A2(_09253_),
    .B(_09034_),
    .Y(_09254_));
 AOI21x1_ASAP7_75t_R _17551_ (.A1(_09208_),
    .A2(_09254_),
    .B(_00387_),
    .Y(_09255_));
 INVx1_ASAP7_75t_R _17552_ (.A(_09113_),
    .Y(_09256_));
 NOR2x2_ASAP7_75t_R _17553_ (.A(_09036_),
    .B(_08990_),
    .Y(_09257_));
 OA21x2_ASAP7_75t_R _17554_ (.A1(_08974_),
    .A2(_09184_),
    .B(_09019_),
    .Y(_09258_));
 AOI211x1_ASAP7_75t_R _17555_ (.A1(_09256_),
    .A2(_09257_),
    .B(_09258_),
    .C(_09034_),
    .Y(_09259_));
 INVx1_ASAP7_75t_R _17556_ (.A(_09137_),
    .Y(_09260_));
 OAI21x1_ASAP7_75t_R _17557_ (.A1(_09052_),
    .A2(_09260_),
    .B(_09022_),
    .Y(_09261_));
 OAI21x1_ASAP7_75t_R _17558_ (.A1(_09259_),
    .A2(_09261_),
    .B(_00388_),
    .Y(_09262_));
 OAI21x1_ASAP7_75t_R _17559_ (.A1(_09255_),
    .A2(_09262_),
    .B(_09098_),
    .Y(_09263_));
 AO21x1_ASAP7_75t_R _17560_ (.A1(_09029_),
    .A2(_09042_),
    .B(_09171_),
    .Y(_09264_));
 AO21x1_ASAP7_75t_R _17561_ (.A1(_08997_),
    .A2(_09005_),
    .B(_08990_),
    .Y(_09265_));
 AND3x1_ASAP7_75t_R _17562_ (.A(_09264_),
    .B(_09141_),
    .C(_09265_),
    .Y(_09266_));
 OA21x2_ASAP7_75t_R _17563_ (.A1(_09193_),
    .A2(_09011_),
    .B(_09093_),
    .Y(_09267_));
 AO21x1_ASAP7_75t_R _17564_ (.A1(_08998_),
    .A2(_09089_),
    .B(_08962_),
    .Y(_09268_));
 AO21x1_ASAP7_75t_R _17565_ (.A1(_09267_),
    .A2(_09268_),
    .B(_09065_),
    .Y(_09269_));
 AO21x1_ASAP7_75t_R _17566_ (.A1(_09014_),
    .A2(_08997_),
    .B(_09069_),
    .Y(_09270_));
 AOI21x1_ASAP7_75t_R _17567_ (.A1(_08995_),
    .A2(_09025_),
    .B(_08137_),
    .Y(_09271_));
 AOI21x1_ASAP7_75t_R _17568_ (.A1(_09270_),
    .A2(_09271_),
    .B(_08145_),
    .Y(_09272_));
 AND3x1_ASAP7_75t_R _17569_ (.A(_08976_),
    .B(_01133_),
    .C(_08966_),
    .Y(_09273_));
 OAI21x1_ASAP7_75t_R _17570_ (.A1(_09030_),
    .A2(_09273_),
    .B(_08978_),
    .Y(_09274_));
 AOI21x1_ASAP7_75t_R _17571_ (.A1(_09272_),
    .A2(_09274_),
    .B(_09072_),
    .Y(_09275_));
 OAI21x1_ASAP7_75t_R _17572_ (.A1(_09266_),
    .A2(_09269_),
    .B(_09275_),
    .Y(_09276_));
 OA21x2_ASAP7_75t_R _17573_ (.A1(_08976_),
    .A2(_09197_),
    .B(_08969_),
    .Y(_09277_));
 AOI21x1_ASAP7_75t_R _17574_ (.A1(_09270_),
    .A2(_09277_),
    .B(_08145_),
    .Y(_09278_));
 AO21x1_ASAP7_75t_R _17575_ (.A1(_09100_),
    .A2(_09060_),
    .B(_08967_),
    .Y(_09279_));
 NAND2x1_ASAP7_75t_R _17576_ (.A(_09279_),
    .B(_09115_),
    .Y(_09280_));
 AOI21x1_ASAP7_75t_R _17577_ (.A1(_09278_),
    .A2(_09280_),
    .B(_09134_),
    .Y(_09281_));
 OA21x2_ASAP7_75t_R _17578_ (.A1(_09069_),
    .A2(_09041_),
    .B(_09078_),
    .Y(_09282_));
 OAI21x1_ASAP7_75t_R _17579_ (.A1(_09257_),
    .A2(_09020_),
    .B(_09282_),
    .Y(_09283_));
 AOI22x1_ASAP7_75t_R _17580_ (.A1(_08960_),
    .A2(_08954_),
    .B1(_08983_),
    .B2(_15760_),
    .Y(_09284_));
 NOR2x1_ASAP7_75t_R _17581_ (.A(_09005_),
    .B(_08976_),
    .Y(_09285_));
 AOI21x1_ASAP7_75t_R _17582_ (.A1(_09029_),
    .A2(_09284_),
    .B(_09285_),
    .Y(_09286_));
 AOI21x1_ASAP7_75t_R _17583_ (.A1(_09136_),
    .A2(_09286_),
    .B(_09065_),
    .Y(_09287_));
 NAND2x1_ASAP7_75t_R _17584_ (.A(_09283_),
    .B(_09287_),
    .Y(_09288_));
 AOI21x1_ASAP7_75t_R _17585_ (.A1(_09281_),
    .A2(_09288_),
    .B(_09098_),
    .Y(_09289_));
 NAND2x1_ASAP7_75t_R _17586_ (.A(_09276_),
    .B(_09289_),
    .Y(_09290_));
 OAI21x1_ASAP7_75t_R _17587_ (.A1(_09252_),
    .A2(_09263_),
    .B(_09290_),
    .Y(_00011_));
 NAND2x1_ASAP7_75t_R _17588_ (.A(_09131_),
    .B(_08962_),
    .Y(_09291_));
 AND3x1_ASAP7_75t_R _17589_ (.A(_09062_),
    .B(_09033_),
    .C(_09291_),
    .Y(_09292_));
 OA21x2_ASAP7_75t_R _17590_ (.A1(_08976_),
    .A2(_09091_),
    .B(_08136_),
    .Y(_09293_));
 INVx1_ASAP7_75t_R _17591_ (.A(_09293_),
    .Y(_09294_));
 NAND2x2_ASAP7_75t_R _17592_ (.A(_09055_),
    .B(_09069_),
    .Y(_09295_));
 NAND2x1_ASAP7_75t_R _17593_ (.A(_09295_),
    .B(_09092_),
    .Y(_09296_));
 OAI21x1_ASAP7_75t_R _17594_ (.A1(_09294_),
    .A2(_09296_),
    .B(_09086_),
    .Y(_09297_));
 NOR2x1_ASAP7_75t_R _17595_ (.A(_09292_),
    .B(_09297_),
    .Y(_09298_));
 NOR2x1_ASAP7_75t_R _17596_ (.A(_09063_),
    .B(_09033_),
    .Y(_09299_));
 NAND2x2_ASAP7_75t_R _17597_ (.A(_09204_),
    .B(_09019_),
    .Y(_09300_));
 AO21x1_ASAP7_75t_R _17598_ (.A1(_09299_),
    .A2(_09300_),
    .B(_09086_),
    .Y(_09301_));
 AO21x1_ASAP7_75t_R _17599_ (.A1(_01135_),
    .A2(_08966_),
    .B(_08976_),
    .Y(_09302_));
 NAND2x1_ASAP7_75t_R _17600_ (.A(_09164_),
    .B(_09302_),
    .Y(_09303_));
 NOR2x1_ASAP7_75t_R _17601_ (.A(_08978_),
    .B(_09303_),
    .Y(_09304_));
 OAI21x1_ASAP7_75t_R _17602_ (.A1(_09301_),
    .A2(_09304_),
    .B(_00387_),
    .Y(_09305_));
 OAI21x1_ASAP7_75t_R _17603_ (.A1(_09298_),
    .A2(_09305_),
    .B(_00389_),
    .Y(_09306_));
 OA21x2_ASAP7_75t_R _17604_ (.A1(net944),
    .A2(_15758_),
    .B(_08995_),
    .Y(_09307_));
 NAND2x1_ASAP7_75t_R _17605_ (.A(_09141_),
    .B(_09180_),
    .Y(_09308_));
 AO21x1_ASAP7_75t_R _17606_ (.A1(_08989_),
    .A2(_09307_),
    .B(_09308_),
    .Y(_09309_));
 NAND2x1_ASAP7_75t_R _17607_ (.A(_15747_),
    .B(_09011_),
    .Y(_09310_));
 OAI21x1_ASAP7_75t_R _17608_ (.A1(_15760_),
    .A2(_09310_),
    .B(_09128_),
    .Y(_09311_));
 INVx1_ASAP7_75t_R _17609_ (.A(_09042_),
    .Y(_09312_));
 AO21x1_ASAP7_75t_R _17610_ (.A1(_00385_),
    .A2(_09312_),
    .B(_09068_),
    .Y(_09313_));
 OA21x2_ASAP7_75t_R _17611_ (.A1(_09311_),
    .A2(_09313_),
    .B(_09134_),
    .Y(_09314_));
 NOR2x1_ASAP7_75t_R _17612_ (.A(_09162_),
    .B(_09217_),
    .Y(_09315_));
 NAND2x2_ASAP7_75t_R _17613_ (.A(_09111_),
    .B(_09105_),
    .Y(_09316_));
 NOR2x2_ASAP7_75t_R _17614_ (.A(_09165_),
    .B(_09316_),
    .Y(_09317_));
 NAND2x1_ASAP7_75t_R _17615_ (.A(_09111_),
    .B(_08995_),
    .Y(_09318_));
 OAI21x1_ASAP7_75t_R _17616_ (.A1(_09039_),
    .A2(_09318_),
    .B(_09141_),
    .Y(_09319_));
 OAI21x1_ASAP7_75t_R _17617_ (.A1(_09317_),
    .A2(_09319_),
    .B(_09072_),
    .Y(_09320_));
 OAI21x1_ASAP7_75t_R _17618_ (.A1(_09315_),
    .A2(_09320_),
    .B(_08980_),
    .Y(_09321_));
 AOI21x1_ASAP7_75t_R _17619_ (.A1(_09309_),
    .A2(_09314_),
    .B(_09321_),
    .Y(_09322_));
 AO21x1_ASAP7_75t_R _17620_ (.A1(_09106_),
    .A2(_08951_),
    .B(_09011_),
    .Y(_09323_));
 NAND2x1_ASAP7_75t_R _17621_ (.A(_15758_),
    .B(_08995_),
    .Y(_09324_));
 AO21x1_ASAP7_75t_R _17622_ (.A1(_09323_),
    .A2(_09324_),
    .B(_09141_),
    .Y(_09325_));
 AO21x1_ASAP7_75t_R _17623_ (.A1(_08989_),
    .A2(_09042_),
    .B(_09011_),
    .Y(_09326_));
 AO21x1_ASAP7_75t_R _17624_ (.A1(_09150_),
    .A2(_09326_),
    .B(_08970_),
    .Y(_09327_));
 AOI21x1_ASAP7_75t_R _17625_ (.A1(_09325_),
    .A2(_09327_),
    .B(_09134_),
    .Y(_09328_));
 AND2x2_ASAP7_75t_R _17626_ (.A(_09316_),
    .B(_09007_),
    .Y(_09329_));
 NOR2x2_ASAP7_75t_R _17627_ (.A(_09018_),
    .B(_08985_),
    .Y(_09330_));
 AO21x1_ASAP7_75t_R _17628_ (.A1(_09330_),
    .A2(_09204_),
    .B(_09033_),
    .Y(_09331_));
 NOR2x1_ASAP7_75t_R _17629_ (.A(_09329_),
    .B(_09331_),
    .Y(_09332_));
 NAND2x1_ASAP7_75t_R _17630_ (.A(_09103_),
    .B(_09081_),
    .Y(_09333_));
 OAI21x1_ASAP7_75t_R _17631_ (.A1(_09020_),
    .A2(_09333_),
    .B(_09134_),
    .Y(_09334_));
 OAI21x1_ASAP7_75t_R _17632_ (.A1(_09332_),
    .A2(_09334_),
    .B(_08980_),
    .Y(_09335_));
 NOR2x1_ASAP7_75t_R _17633_ (.A(_09328_),
    .B(_09335_),
    .Y(_09336_));
 AO21x1_ASAP7_75t_R _17634_ (.A1(_08999_),
    .A2(_00466_),
    .B(_08137_),
    .Y(_09337_));
 AOI21x1_ASAP7_75t_R _17635_ (.A1(_00385_),
    .A2(_09130_),
    .B(_09337_),
    .Y(_09338_));
 NOR2x1_ASAP7_75t_R _17636_ (.A(_09123_),
    .B(_09300_),
    .Y(_09339_));
 AO21x1_ASAP7_75t_R _17637_ (.A1(_09024_),
    .A2(_09049_),
    .B(_09033_),
    .Y(_09340_));
 OAI21x1_ASAP7_75t_R _17638_ (.A1(_09339_),
    .A2(_09340_),
    .B(_09086_),
    .Y(_09341_));
 OAI21x1_ASAP7_75t_R _17639_ (.A1(_09338_),
    .A2(_09341_),
    .B(_00387_),
    .Y(_09342_));
 OA21x2_ASAP7_75t_R _17640_ (.A1(_09139_),
    .A2(_09055_),
    .B(_08986_),
    .Y(_09343_));
 OA21x2_ASAP7_75t_R _17641_ (.A1(_09156_),
    .A2(_15760_),
    .B(_08999_),
    .Y(_09344_));
 NAND2x2_ASAP7_75t_R _17642_ (.A(_08983_),
    .B(_15758_),
    .Y(_09345_));
 AO21x1_ASAP7_75t_R _17643_ (.A1(_09165_),
    .A2(_09345_),
    .B(_09033_),
    .Y(_09346_));
 OAI21x1_ASAP7_75t_R _17644_ (.A1(_09344_),
    .A2(_09346_),
    .B(_09072_),
    .Y(_09347_));
 AOI21x1_ASAP7_75t_R _17645_ (.A1(_09034_),
    .A2(_09343_),
    .B(_09347_),
    .Y(_09348_));
 OAI21x1_ASAP7_75t_R _17646_ (.A1(_09342_),
    .A2(_09348_),
    .B(_09098_),
    .Y(_09349_));
 OAI22x1_ASAP7_75t_R _17647_ (.A1(_09306_),
    .A2(_09322_),
    .B1(_09336_),
    .B2(_09349_),
    .Y(_00012_));
 AO21x1_ASAP7_75t_R _17648_ (.A1(_08994_),
    .A2(_09060_),
    .B(_08967_),
    .Y(_09350_));
 OA21x2_ASAP7_75t_R _17649_ (.A1(_09197_),
    .A2(_09038_),
    .B(_09350_),
    .Y(_09351_));
 AO21x1_ASAP7_75t_R _17650_ (.A1(_08995_),
    .A2(_15748_),
    .B(_08137_),
    .Y(_09352_));
 OAI21x1_ASAP7_75t_R _17651_ (.A1(_09352_),
    .A2(_09017_),
    .B(_09058_),
    .Y(_09353_));
 AOI21x1_ASAP7_75t_R _17652_ (.A1(_00386_),
    .A2(_09351_),
    .B(_09353_),
    .Y(_09354_));
 OA21x2_ASAP7_75t_R _17653_ (.A1(_09076_),
    .A2(_09041_),
    .B(_09078_),
    .Y(_09355_));
 AO21x1_ASAP7_75t_R _17654_ (.A1(_08984_),
    .A2(_08951_),
    .B(_09011_),
    .Y(_09356_));
 AO21x1_ASAP7_75t_R _17655_ (.A1(_09355_),
    .A2(_09356_),
    .B(_09058_),
    .Y(_09357_));
 AO21x1_ASAP7_75t_R _17656_ (.A1(_08966_),
    .A2(_09089_),
    .B(_08990_),
    .Y(_09358_));
 AND3x1_ASAP7_75t_R _17657_ (.A(_08986_),
    .B(_09103_),
    .C(_09358_),
    .Y(_09359_));
 OAI21x1_ASAP7_75t_R _17658_ (.A1(_09357_),
    .A2(_09359_),
    .B(_09098_),
    .Y(_09360_));
 NOR2x1_ASAP7_75t_R _17659_ (.A(_09354_),
    .B(_09360_),
    .Y(_09361_));
 AO21x1_ASAP7_75t_R _17660_ (.A1(_08976_),
    .A2(_09100_),
    .B(_09078_),
    .Y(_09362_));
 NOR2x1_ASAP7_75t_R _17661_ (.A(_09258_),
    .B(_09362_),
    .Y(_09363_));
 AND2x2_ASAP7_75t_R _17662_ (.A(_09078_),
    .B(_08964_),
    .Y(_09364_));
 AO21x1_ASAP7_75t_R _17663_ (.A1(_09364_),
    .A2(_09139_),
    .B(_09058_),
    .Y(_09365_));
 OAI21x1_ASAP7_75t_R _17664_ (.A1(_09363_),
    .A2(_09365_),
    .B(_00389_),
    .Y(_09366_));
 AO21x1_ASAP7_75t_R _17665_ (.A1(_08951_),
    .A2(_08972_),
    .B(_09007_),
    .Y(_09367_));
 AO21x1_ASAP7_75t_R _17666_ (.A1(_09367_),
    .A2(_08991_),
    .B(_08978_),
    .Y(_09368_));
 AO21x1_ASAP7_75t_R _17667_ (.A1(_09106_),
    .A2(_09089_),
    .B(_08962_),
    .Y(_09369_));
 NAND2x1_ASAP7_75t_R _17668_ (.A(_09024_),
    .B(_09061_),
    .Y(_09370_));
 AO21x1_ASAP7_75t_R _17669_ (.A1(_09369_),
    .A2(_09370_),
    .B(_08970_),
    .Y(_09371_));
 AOI21x1_ASAP7_75t_R _17670_ (.A1(_09368_),
    .A2(_09371_),
    .B(_08980_),
    .Y(_09372_));
 OAI21x1_ASAP7_75t_R _17671_ (.A1(_09366_),
    .A2(_09372_),
    .B(_00388_),
    .Y(_09373_));
 NAND2x1_ASAP7_75t_R _17672_ (.A(_09068_),
    .B(_09295_),
    .Y(_09374_));
 AOI21x1_ASAP7_75t_R _17673_ (.A1(_08994_),
    .A2(_09344_),
    .B(_09374_),
    .Y(_09375_));
 OA21x2_ASAP7_75t_R _17674_ (.A1(_08967_),
    .A2(_08951_),
    .B(_09093_),
    .Y(_09376_));
 AO21x1_ASAP7_75t_R _17675_ (.A1(_09100_),
    .A2(_09006_),
    .B(_09171_),
    .Y(_09377_));
 AND2x2_ASAP7_75t_R _17676_ (.A(_09376_),
    .B(_09377_),
    .Y(_09378_));
 OAI21x1_ASAP7_75t_R _17677_ (.A1(_09375_),
    .A2(_09378_),
    .B(_08980_),
    .Y(_09379_));
 INVx1_ASAP7_75t_R _17678_ (.A(_09310_),
    .Y(_09380_));
 OAI21x1_ASAP7_75t_R _17679_ (.A1(_09380_),
    .A2(_09317_),
    .B(_09034_),
    .Y(_09381_));
 NOR2x1_ASAP7_75t_R _17680_ (.A(_09173_),
    .B(_09171_),
    .Y(_09382_));
 AOI21x1_ASAP7_75t_R _17681_ (.A1(_09041_),
    .A2(_09382_),
    .B(_09103_),
    .Y(_09383_));
 AO21x1_ASAP7_75t_R _17682_ (.A1(_15748_),
    .A2(_15747_),
    .B(_08977_),
    .Y(_09384_));
 AOI21x1_ASAP7_75t_R _17683_ (.A1(_09383_),
    .A2(_09384_),
    .B(_09065_),
    .Y(_09385_));
 NAND2x1_ASAP7_75t_R _17684_ (.A(_09381_),
    .B(_09385_),
    .Y(_09386_));
 AOI21x1_ASAP7_75t_R _17685_ (.A1(_09379_),
    .A2(_09386_),
    .B(_09098_),
    .Y(_09387_));
 AOI211x1_ASAP7_75t_R _17686_ (.A1(_09122_),
    .A2(_09166_),
    .B(_09330_),
    .C(_08978_),
    .Y(_09388_));
 OAI21x1_ASAP7_75t_R _17687_ (.A1(_09114_),
    .A2(_09125_),
    .B(_09058_),
    .Y(_09389_));
 NOR2x1_ASAP7_75t_R _17688_ (.A(_09388_),
    .B(_09389_),
    .Y(_09390_));
 AO21x1_ASAP7_75t_R _17689_ (.A1(_09165_),
    .A2(_00463_),
    .B(_09068_),
    .Y(_09391_));
 OAI21x1_ASAP7_75t_R _17690_ (.A1(_09284_),
    .A2(_09391_),
    .B(_09065_),
    .Y(_09392_));
 OA21x2_ASAP7_75t_R _17691_ (.A1(_08952_),
    .A2(_09040_),
    .B(_09165_),
    .Y(_09393_));
 OAI21x1_ASAP7_75t_R _17692_ (.A1(_09100_),
    .A2(_00385_),
    .B(_09141_),
    .Y(_09394_));
 AOI211x1_ASAP7_75t_R _17693_ (.A1(_09122_),
    .A2(_08950_),
    .B(_09393_),
    .C(_09394_),
    .Y(_09395_));
 OAI21x1_ASAP7_75t_R _17694_ (.A1(_09392_),
    .A2(_09395_),
    .B(_09098_),
    .Y(_09396_));
 OAI21x1_ASAP7_75t_R _17695_ (.A1(_09390_),
    .A2(_09396_),
    .B(_09134_),
    .Y(_09397_));
 OAI22x1_ASAP7_75t_R _17696_ (.A1(_09361_),
    .A2(_09373_),
    .B1(_09387_),
    .B2(_09397_),
    .Y(_00013_));
 AO21x1_ASAP7_75t_R _17697_ (.A1(_08989_),
    .A2(_09048_),
    .B(_08962_),
    .Y(_09398_));
 AO21x1_ASAP7_75t_R _17698_ (.A1(_09398_),
    .A2(_09282_),
    .B(_08153_),
    .Y(_09399_));
 NOR2x2_ASAP7_75t_R _17699_ (.A(_09018_),
    .B(_09056_),
    .Y(_09400_));
 AOI211x1_ASAP7_75t_R _17700_ (.A1(_09307_),
    .A2(_08997_),
    .B(_09400_),
    .C(_00386_),
    .Y(_09401_));
 OAI21x1_ASAP7_75t_R _17701_ (.A1(_09399_),
    .A2(_09401_),
    .B(_08980_),
    .Y(_09402_));
 AO21x1_ASAP7_75t_R _17702_ (.A1(_08987_),
    .A2(_09010_),
    .B(_09076_),
    .Y(_09403_));
 AO21x1_ASAP7_75t_R _17703_ (.A1(_08998_),
    .A2(_09060_),
    .B(_09069_),
    .Y(_09404_));
 AND3x1_ASAP7_75t_R _17704_ (.A(_09403_),
    .B(_09103_),
    .C(_09404_),
    .Y(_09405_));
 OAI21x1_ASAP7_75t_R _17705_ (.A1(_15748_),
    .A2(_09324_),
    .B(_09293_),
    .Y(_09406_));
 OAI21x1_ASAP7_75t_R _17706_ (.A1(_09400_),
    .A2(_09406_),
    .B(_09072_),
    .Y(_09407_));
 NOR2x1_ASAP7_75t_R _17707_ (.A(_09405_),
    .B(_09407_),
    .Y(_09408_));
 OAI21x1_ASAP7_75t_R _17708_ (.A1(_09402_),
    .A2(_09408_),
    .B(_00389_),
    .Y(_09409_));
 OA211x2_ASAP7_75t_R _17709_ (.A1(_09222_),
    .A2(_09198_),
    .B(_09244_),
    .C(_09078_),
    .Y(_09410_));
 AO21x1_ASAP7_75t_R _17710_ (.A1(_09100_),
    .A2(_09157_),
    .B(_08990_),
    .Y(_09411_));
 AO21x1_ASAP7_75t_R _17711_ (.A1(_08994_),
    .A2(_08964_),
    .B(_09171_),
    .Y(_09412_));
 AOI21x1_ASAP7_75t_R _17712_ (.A1(_09411_),
    .A2(_09412_),
    .B(_09141_),
    .Y(_09413_));
 OA21x2_ASAP7_75t_R _17713_ (.A1(_09410_),
    .A2(_09413_),
    .B(_09134_),
    .Y(_09414_));
 AND2x2_ASAP7_75t_R _17714_ (.A(_09316_),
    .B(_08990_),
    .Y(_09415_));
 AOI211x1_ASAP7_75t_R _17715_ (.A1(net927),
    .A2(_09122_),
    .B(_09415_),
    .C(_00386_),
    .Y(_09416_));
 OA21x2_ASAP7_75t_R _17716_ (.A1(_09184_),
    .A2(_09194_),
    .B(_09019_),
    .Y(_09417_));
 AO21x1_ASAP7_75t_R _17717_ (.A1(_09024_),
    .A2(_09312_),
    .B(_09417_),
    .Y(_09418_));
 OAI21x1_ASAP7_75t_R _17718_ (.A1(_09034_),
    .A2(_09418_),
    .B(_09072_),
    .Y(_09419_));
 OAI21x1_ASAP7_75t_R _17719_ (.A1(_09416_),
    .A2(_09419_),
    .B(_00387_),
    .Y(_09420_));
 NOR2x1_ASAP7_75t_R _17720_ (.A(_09414_),
    .B(_09420_),
    .Y(_09421_));
 AND3x1_ASAP7_75t_R _17721_ (.A(_09076_),
    .B(_09111_),
    .C(_08964_),
    .Y(_09422_));
 AND3x1_ASAP7_75t_R _17722_ (.A(_09019_),
    .B(_09014_),
    .C(_08982_),
    .Y(_09423_));
 OA21x2_ASAP7_75t_R _17723_ (.A1(_09422_),
    .A2(_09423_),
    .B(_08970_),
    .Y(_09424_));
 NAND2x1_ASAP7_75t_R _17724_ (.A(_08998_),
    .B(_08975_),
    .Y(_09425_));
 AO21x1_ASAP7_75t_R _17725_ (.A1(_09425_),
    .A2(_09024_),
    .B(_09033_),
    .Y(_09426_));
 OAI21x1_ASAP7_75t_R _17726_ (.A1(_09423_),
    .A2(_09426_),
    .B(_09072_),
    .Y(_09427_));
 OA21x2_ASAP7_75t_R _17727_ (.A1(_09019_),
    .A2(_08982_),
    .B(_08136_),
    .Y(_09428_));
 AO21x1_ASAP7_75t_R _17728_ (.A1(_09100_),
    .A2(_08951_),
    .B(_09076_),
    .Y(_09429_));
 NAND2x1_ASAP7_75t_R _17729_ (.A(_09428_),
    .B(_09429_),
    .Y(_09430_));
 AOI21x1_ASAP7_75t_R _17730_ (.A1(_00471_),
    .A2(_09165_),
    .B(_08137_),
    .Y(_09431_));
 AOI21x1_ASAP7_75t_R _17731_ (.A1(_09431_),
    .A2(_09350_),
    .B(_08153_),
    .Y(_09432_));
 AOI21x1_ASAP7_75t_R _17732_ (.A1(_09430_),
    .A2(_09432_),
    .B(_08980_),
    .Y(_09433_));
 OAI21x1_ASAP7_75t_R _17733_ (.A1(_09424_),
    .A2(_09427_),
    .B(_09433_),
    .Y(_09434_));
 NOR2x1_ASAP7_75t_R _17734_ (.A(_09127_),
    .B(_08999_),
    .Y(_09435_));
 AOI21x1_ASAP7_75t_R _17735_ (.A1(_09103_),
    .A2(_09435_),
    .B(_08153_),
    .Y(_09436_));
 NOR2x1_ASAP7_75t_R _17736_ (.A(_00463_),
    .B(_15760_),
    .Y(_09437_));
 OA21x2_ASAP7_75t_R _17737_ (.A1(_08967_),
    .A2(_09437_),
    .B(_09078_),
    .Y(_09438_));
 OAI21x1_ASAP7_75t_R _17738_ (.A1(_09123_),
    .A2(_09300_),
    .B(_09438_),
    .Y(_09439_));
 AOI21x1_ASAP7_75t_R _17739_ (.A1(_09436_),
    .A2(_09439_),
    .B(_09022_),
    .Y(_09440_));
 AO21x1_ASAP7_75t_R _17740_ (.A1(_09024_),
    .A2(_08952_),
    .B(_09258_),
    .Y(_09441_));
 NOR2x1_ASAP7_75t_R _17741_ (.A(_09093_),
    .B(_09124_),
    .Y(_09442_));
 AOI21x1_ASAP7_75t_R _17742_ (.A1(_08968_),
    .A2(_09442_),
    .B(_09086_),
    .Y(_09443_));
 OAI21x1_ASAP7_75t_R _17743_ (.A1(_00386_),
    .A2(_09441_),
    .B(_09443_),
    .Y(_09444_));
 AOI21x1_ASAP7_75t_R _17744_ (.A1(_09440_),
    .A2(_09444_),
    .B(_00389_),
    .Y(_09445_));
 NAND2x1_ASAP7_75t_R _17745_ (.A(_09434_),
    .B(_09445_),
    .Y(_09446_));
 OAI21x1_ASAP7_75t_R _17746_ (.A1(_09409_),
    .A2(_09421_),
    .B(_09446_),
    .Y(_00014_));
 NOR2x1_ASAP7_75t_R _17747_ (.A(_08983_),
    .B(_09122_),
    .Y(_09447_));
 AO21x1_ASAP7_75t_R _17748_ (.A1(_09024_),
    .A2(_09194_),
    .B(_08137_),
    .Y(_09448_));
 OAI21x1_ASAP7_75t_R _17749_ (.A1(_09447_),
    .A2(_09448_),
    .B(_09022_),
    .Y(_09449_));
 AOI21x1_ASAP7_75t_R _17750_ (.A1(_08989_),
    .A2(_09048_),
    .B(_00385_),
    .Y(_09450_));
 AOI211x1_ASAP7_75t_R _17751_ (.A1(_09149_),
    .A2(_08989_),
    .B(_09450_),
    .C(_08970_),
    .Y(_09451_));
 OAI21x1_ASAP7_75t_R _17752_ (.A1(_09449_),
    .A2(_09451_),
    .B(_09134_),
    .Y(_09452_));
 AO21x1_ASAP7_75t_R _17753_ (.A1(_09029_),
    .A2(_09091_),
    .B(_09011_),
    .Y(_09453_));
 INVx1_ASAP7_75t_R _17754_ (.A(_01135_),
    .Y(_09454_));
 AOI21x1_ASAP7_75t_R _17755_ (.A1(_09454_),
    .A2(_09165_),
    .B(_08137_),
    .Y(_09455_));
 AO21x1_ASAP7_75t_R _17756_ (.A1(_09453_),
    .A2(_09455_),
    .B(_09058_),
    .Y(_09456_));
 AO21x1_ASAP7_75t_R _17757_ (.A1(_09100_),
    .A2(_09130_),
    .B(_09171_),
    .Y(_09457_));
 AND3x1_ASAP7_75t_R _17758_ (.A(_09457_),
    .B(_09428_),
    .C(_09229_),
    .Y(_09458_));
 NOR2x1_ASAP7_75t_R _17759_ (.A(_09456_),
    .B(_09458_),
    .Y(_09459_));
 OAI21x1_ASAP7_75t_R _17760_ (.A1(_09452_),
    .A2(_09459_),
    .B(_00389_),
    .Y(_09460_));
 AO21x1_ASAP7_75t_R _17761_ (.A1(_09100_),
    .A2(_09041_),
    .B(_09171_),
    .Y(_09461_));
 AO21x1_ASAP7_75t_R _17762_ (.A1(_09010_),
    .A2(_09042_),
    .B(_08990_),
    .Y(_09462_));
 AO21x1_ASAP7_75t_R _17763_ (.A1(_09461_),
    .A2(_09462_),
    .B(_09141_),
    .Y(_09463_));
 AND3x1_ASAP7_75t_R _17764_ (.A(_08994_),
    .B(_09007_),
    .C(_09345_),
    .Y(_09464_));
 OAI21x1_ASAP7_75t_R _17765_ (.A1(_09253_),
    .A2(_09464_),
    .B(_00386_),
    .Y(_09465_));
 AOI21x1_ASAP7_75t_R _17766_ (.A1(_09463_),
    .A2(_09465_),
    .B(_08980_),
    .Y(_09466_));
 AO21x1_ASAP7_75t_R _17767_ (.A1(_09082_),
    .A2(_08962_),
    .B(_09093_),
    .Y(_09467_));
 NOR2x1_ASAP7_75t_R _17768_ (.A(_09467_),
    .B(_09415_),
    .Y(_09468_));
 OA21x2_ASAP7_75t_R _17769_ (.A1(_09076_),
    .A2(_08988_),
    .B(_09093_),
    .Y(_09469_));
 OA21x2_ASAP7_75t_R _17770_ (.A1(_08967_),
    .A2(_09157_),
    .B(_09042_),
    .Y(_09470_));
 AO21x1_ASAP7_75t_R _17771_ (.A1(_09469_),
    .A2(_09470_),
    .B(_09058_),
    .Y(_09471_));
 OAI21x1_ASAP7_75t_R _17772_ (.A1(_09468_),
    .A2(_09471_),
    .B(_09072_),
    .Y(_09472_));
 NOR2x1_ASAP7_75t_R _17773_ (.A(_09466_),
    .B(_09472_),
    .Y(_09473_));
 AO21x1_ASAP7_75t_R _17774_ (.A1(_09248_),
    .A2(_09132_),
    .B(_08970_),
    .Y(_09474_));
 AO21x1_ASAP7_75t_R _17775_ (.A1(_09226_),
    .A2(_09404_),
    .B(_08978_),
    .Y(_09475_));
 AOI21x1_ASAP7_75t_R _17776_ (.A1(_09474_),
    .A2(_09475_),
    .B(_00387_),
    .Y(_09476_));
 AO21x1_ASAP7_75t_R _17777_ (.A1(_08118_),
    .A2(_08114_),
    .B(_09112_),
    .Y(_09477_));
 AO21x1_ASAP7_75t_R _17778_ (.A1(_09024_),
    .A2(_09477_),
    .B(_09068_),
    .Y(_09478_));
 OAI21x1_ASAP7_75t_R _17779_ (.A1(_09478_),
    .A2(_09339_),
    .B(_09022_),
    .Y(_09479_));
 NAND2x1_ASAP7_75t_R _17780_ (.A(_09048_),
    .B(_08997_),
    .Y(_09480_));
 OA21x2_ASAP7_75t_R _17781_ (.A1(_09009_),
    .A2(_09312_),
    .B(_09165_),
    .Y(_09481_));
 AOI211x1_ASAP7_75t_R _17782_ (.A1(_09122_),
    .A2(_09480_),
    .B(_09481_),
    .C(_08970_),
    .Y(_09482_));
 OAI21x1_ASAP7_75t_R _17783_ (.A1(_09479_),
    .A2(_09482_),
    .B(_00388_),
    .Y(_09483_));
 OAI21x1_ASAP7_75t_R _17784_ (.A1(_09476_),
    .A2(_09483_),
    .B(_09098_),
    .Y(_09484_));
 AND3x1_ASAP7_75t_R _17785_ (.A(_09007_),
    .B(_08953_),
    .C(_09345_),
    .Y(_09485_));
 OAI21x1_ASAP7_75t_R _17786_ (.A1(_09307_),
    .A2(_09485_),
    .B(_00386_),
    .Y(_09486_));
 OA21x2_ASAP7_75t_R _17787_ (.A1(_09362_),
    .A2(_09382_),
    .B(_09065_),
    .Y(_09487_));
 NAND2x1_ASAP7_75t_R _17788_ (.A(_09486_),
    .B(_09487_),
    .Y(_09488_));
 AO21x1_ASAP7_75t_R _17789_ (.A1(_15748_),
    .A2(_08999_),
    .B(_09033_),
    .Y(_09489_));
 AOI21x1_ASAP7_75t_R _17790_ (.A1(_08989_),
    .A2(_09330_),
    .B(_09489_),
    .Y(_09490_));
 AND3x1_ASAP7_75t_R _17791_ (.A(_08962_),
    .B(_09111_),
    .C(_09345_),
    .Y(_09491_));
 NOR2x1_ASAP7_75t_R _17792_ (.A(_09491_),
    .B(_09217_),
    .Y(_09492_));
 OAI21x1_ASAP7_75t_R _17793_ (.A1(_09490_),
    .A2(_09492_),
    .B(_00387_),
    .Y(_09493_));
 AOI21x1_ASAP7_75t_R _17794_ (.A1(_09488_),
    .A2(_09493_),
    .B(_00388_),
    .Y(_09494_));
 OAI22x1_ASAP7_75t_R _17795_ (.A1(_09460_),
    .A2(_09473_),
    .B1(_09484_),
    .B2(_09494_),
    .Y(_00015_));
 INVx6_ASAP7_75t_R _17796_ (.A(_08043_),
    .Y(_09495_));
 BUFx12f_ASAP7_75t_R _17797_ (.A(_09495_),
    .Y(_15776_));
 INVx6_ASAP7_75t_R _17798_ (.A(_15768_),
    .Y(_15766_));
 NAND2x2_ASAP7_75t_R _17799_ (.A(_09495_),
    .B(net17),
    .Y(_09496_));
 BUFx3_ASAP7_75t_R _17800_ (.A(_08042_),
    .Y(_09497_));
 BUFx3_ASAP7_75t_R _17801_ (.A(_08038_),
    .Y(_09498_));
 AO21x2_ASAP7_75t_R _17802_ (.A1(_09497_),
    .A2(_09498_),
    .B(_00474_),
    .Y(_09499_));
 BUFx10_ASAP7_75t_R _17803_ (.A(_08055_),
    .Y(_09500_));
 BUFx4f_ASAP7_75t_R _17804_ (.A(_09500_),
    .Y(_09501_));
 AO21x1_ASAP7_75t_R _17805_ (.A1(_09496_),
    .A2(_09499_),
    .B(_09501_),
    .Y(_09502_));
 INVx1_ASAP7_75t_R _17806_ (.A(_00474_),
    .Y(_09503_));
 BUFx12_ASAP7_75t_R _17807_ (.A(_08043_),
    .Y(_09504_));
 NOR2x2_ASAP7_75t_R _17808_ (.A(net857),
    .B(_09504_),
    .Y(_09505_));
 NAND2x1_ASAP7_75t_R _17809_ (.A(_09505_),
    .B(_08056_),
    .Y(_09506_));
 INVx2_ASAP7_75t_R _17810_ (.A(_01117_),
    .Y(_09507_));
 XOR2x1_ASAP7_75t_R _17811_ (.A(_08060_),
    .Y(_09508_),
    .B(_09507_));
 INVx1_ASAP7_75t_R _17812_ (.A(_08062_),
    .Y(_09509_));
 OAI21x1_ASAP7_75t_R _17813_ (.A1(_07967_),
    .A2(_09508_),
    .B(_09509_),
    .Y(_09510_));
 BUFx6f_ASAP7_75t_R _17814_ (.A(_09510_),
    .Y(_09511_));
 AO21x1_ASAP7_75t_R _17815_ (.A1(_09502_),
    .A2(_09506_),
    .B(_09511_),
    .Y(_09512_));
 INVx2_ASAP7_75t_R _17816_ (.A(_00473_),
    .Y(_09513_));
 AO21x2_ASAP7_75t_R _17817_ (.A1(_09497_),
    .A2(_09498_),
    .B(_09513_),
    .Y(_09514_));
 NOR2x2_ASAP7_75t_R _17818_ (.A(_09514_),
    .B(_09500_),
    .Y(_09515_));
 AO21x1_ASAP7_75t_R _17819_ (.A1(_08042_),
    .A2(_08038_),
    .B(_09503_),
    .Y(_09516_));
 BUFx3_ASAP7_75t_R _17820_ (.A(_09516_),
    .Y(_09517_));
 INVx4_ASAP7_75t_R _17821_ (.A(_09517_),
    .Y(_09518_));
 NOR2x2_ASAP7_75t_R _17822_ (.A(_08054_),
    .B(_09518_),
    .Y(_09519_));
 NAND2x2_ASAP7_75t_R _17823_ (.A(_09513_),
    .B(_15776_),
    .Y(_09520_));
 BUFx10_ASAP7_75t_R _17824_ (.A(_08055_),
    .Y(_09521_));
 NAND2x2_ASAP7_75t_R _17825_ (.A(_00472_),
    .B(_15776_),
    .Y(_09522_));
 NOR2x2_ASAP7_75t_R _17826_ (.A(_09521_),
    .B(_09522_),
    .Y(_09523_));
 AO21x1_ASAP7_75t_R _17827_ (.A1(_09519_),
    .A2(_09520_),
    .B(_09523_),
    .Y(_09524_));
 BUFx6f_ASAP7_75t_R _17828_ (.A(_09510_),
    .Y(_09525_));
 BUFx6f_ASAP7_75t_R _17829_ (.A(_09525_),
    .Y(_09526_));
 OAI21x1_ASAP7_75t_R _17830_ (.A1(_09515_),
    .A2(_09524_),
    .B(_09526_),
    .Y(_09527_));
 INVx4_ASAP7_75t_R _17831_ (.A(_08071_),
    .Y(_09528_));
 BUFx10_ASAP7_75t_R _17832_ (.A(_09528_),
    .Y(_09529_));
 NAND3x1_ASAP7_75t_R _17833_ (.A(_09512_),
    .B(_09527_),
    .C(_09529_),
    .Y(_09530_));
 AND2x2_ASAP7_75t_R _17834_ (.A(_09504_),
    .B(_00472_),
    .Y(_09531_));
 INVx1_ASAP7_75t_R _17835_ (.A(_09531_),
    .Y(_09532_));
 NOR2x2_ASAP7_75t_R _17836_ (.A(_09513_),
    .B(_08043_),
    .Y(_09533_));
 INVx2_ASAP7_75t_R _17837_ (.A(_09533_),
    .Y(_09534_));
 BUFx6f_ASAP7_75t_R _17838_ (.A(_08054_),
    .Y(_09535_));
 BUFx4f_ASAP7_75t_R _17839_ (.A(_09535_),
    .Y(_09536_));
 AO21x1_ASAP7_75t_R _17840_ (.A1(_09532_),
    .A2(_09534_),
    .B(_09536_),
    .Y(_09537_));
 NAND2x2_ASAP7_75t_R _17841_ (.A(net527),
    .B(_15776_),
    .Y(_09538_));
 AO21x1_ASAP7_75t_R _17842_ (.A1(_09538_),
    .A2(_09499_),
    .B(_09501_),
    .Y(_09539_));
 AND3x1_ASAP7_75t_R _17843_ (.A(_09537_),
    .B(_09511_),
    .C(_09539_),
    .Y(_09540_));
 NOR2x1_ASAP7_75t_R _17844_ (.A(net2),
    .B(_15766_),
    .Y(_09541_));
 INVx1_ASAP7_75t_R _17845_ (.A(_09541_),
    .Y(_09542_));
 NOR2x2_ASAP7_75t_R _17846_ (.A(_09495_),
    .B(_15768_),
    .Y(_09543_));
 NOR2x1_ASAP7_75t_R _17847_ (.A(_09500_),
    .B(_09543_),
    .Y(_09544_));
 NAND2x1_ASAP7_75t_R _17848_ (.A(_09542_),
    .B(_09544_),
    .Y(_09545_));
 BUFx6f_ASAP7_75t_R _17849_ (.A(_08063_),
    .Y(_09546_));
 BUFx4f_ASAP7_75t_R _17850_ (.A(_09500_),
    .Y(_09547_));
 OAI21x1_ASAP7_75t_R _17851_ (.A1(_09543_),
    .A2(_09541_),
    .B(_09547_),
    .Y(_09548_));
 AND3x1_ASAP7_75t_R _17852_ (.A(_09545_),
    .B(_09546_),
    .C(_09548_),
    .Y(_09549_));
 OAI21x1_ASAP7_75t_R _17853_ (.A1(_09540_),
    .A2(_09549_),
    .B(_00402_),
    .Y(_09550_));
 AOI21x1_ASAP7_75t_R _17854_ (.A1(_09530_),
    .A2(_09550_),
    .B(_00403_),
    .Y(_09551_));
 INVx1_ASAP7_75t_R _17855_ (.A(_01136_),
    .Y(_09552_));
 NOR2x2_ASAP7_75t_R _17856_ (.A(_09552_),
    .B(_09504_),
    .Y(_09553_));
 INVx2_ASAP7_75t_R _17857_ (.A(_09553_),
    .Y(_09554_));
 NAND2x2_ASAP7_75t_R _17858_ (.A(_08056_),
    .B(_09554_),
    .Y(_09555_));
 NOR2x1_ASAP7_75t_R _17859_ (.A(_09518_),
    .B(_09555_),
    .Y(_09556_));
 INVx1_ASAP7_75t_R _17860_ (.A(_00476_),
    .Y(_09557_));
 NAND2x2_ASAP7_75t_R _17861_ (.A(_09557_),
    .B(_09495_),
    .Y(_09558_));
 AND2x2_ASAP7_75t_R _17862_ (.A(_09558_),
    .B(_09535_),
    .Y(_09559_));
 NAND2x2_ASAP7_75t_R _17863_ (.A(_15778_),
    .B(net13),
    .Y(_09560_));
 AND2x2_ASAP7_75t_R _17864_ (.A(_09559_),
    .B(_09560_),
    .Y(_09561_));
 OAI21x1_ASAP7_75t_R _17865_ (.A1(_09556_),
    .A2(_09561_),
    .B(_00401_),
    .Y(_09562_));
 BUFx6f_ASAP7_75t_R _17866_ (.A(_09510_),
    .Y(_09563_));
 BUFx6f_ASAP7_75t_R _17867_ (.A(_09563_),
    .Y(_09564_));
 INVx1_ASAP7_75t_R _17868_ (.A(_01137_),
    .Y(_09565_));
 OA21x2_ASAP7_75t_R _17869_ (.A1(_09565_),
    .A2(_15776_),
    .B(_09500_),
    .Y(_09566_));
 NAND2x2_ASAP7_75t_R _17870_ (.A(_09495_),
    .B(_15768_),
    .Y(_09567_));
 INVx3_ASAP7_75t_R _17871_ (.A(_09567_),
    .Y(_09568_));
 NOR2x2_ASAP7_75t_R _17872_ (.A(_08056_),
    .B(_09568_),
    .Y(_09569_));
 AO21x1_ASAP7_75t_R _17873_ (.A1(_09558_),
    .A2(_09566_),
    .B(_09569_),
    .Y(_09570_));
 NAND2x1_ASAP7_75t_R _17874_ (.A(_09564_),
    .B(_09570_),
    .Y(_09571_));
 AOI21x1_ASAP7_75t_R _17875_ (.A1(_09562_),
    .A2(_09571_),
    .B(_09529_),
    .Y(_09572_));
 NOR2x2_ASAP7_75t_R _17876_ (.A(_09504_),
    .B(net17),
    .Y(_09573_));
 NAND2x1_ASAP7_75t_R _17877_ (.A(_09535_),
    .B(_09573_),
    .Y(_09574_));
 AND2x2_ASAP7_75t_R _17878_ (.A(_09574_),
    .B(_09525_),
    .Y(_09575_));
 BUFx6f_ASAP7_75t_R _17879_ (.A(_09521_),
    .Y(_09576_));
 INVx2_ASAP7_75t_R _17880_ (.A(_00475_),
    .Y(_09577_));
 NOR2x1_ASAP7_75t_R _17881_ (.A(_09577_),
    .B(_15776_),
    .Y(_09578_));
 AO21x1_ASAP7_75t_R _17882_ (.A1(_15766_),
    .A2(_15776_),
    .B(_09578_),
    .Y(_09579_));
 NAND2x1_ASAP7_75t_R _17883_ (.A(_09576_),
    .B(_09579_),
    .Y(_09580_));
 BUFx6f_ASAP7_75t_R _17884_ (.A(_08054_),
    .Y(_09581_));
 AO21x2_ASAP7_75t_R _17885_ (.A1(_09497_),
    .A2(_09498_),
    .B(_01139_),
    .Y(_09582_));
 INVx2_ASAP7_75t_R _17886_ (.A(_09582_),
    .Y(_09583_));
 NAND2x2_ASAP7_75t_R _17887_ (.A(_09581_),
    .B(_09583_),
    .Y(_09584_));
 AND3x1_ASAP7_75t_R _17888_ (.A(_09575_),
    .B(_09580_),
    .C(_09584_),
    .Y(_09585_));
 AO21x2_ASAP7_75t_R _17889_ (.A1(_09497_),
    .A2(_09498_),
    .B(_09552_),
    .Y(_09586_));
 NOR2x1_ASAP7_75t_R _17890_ (.A(_09581_),
    .B(_09568_),
    .Y(_09587_));
 BUFx6f_ASAP7_75t_R _17891_ (.A(_09510_),
    .Y(_09588_));
 AOI21x1_ASAP7_75t_R _17892_ (.A1(_09586_),
    .A2(_09587_),
    .B(_09588_),
    .Y(_09589_));
 BUFx6f_ASAP7_75t_R _17893_ (.A(_08054_),
    .Y(_09590_));
 OAI21x1_ASAP7_75t_R _17894_ (.A1(_08022_),
    .A2(_08030_),
    .B(_09504_),
    .Y(_09591_));
 NAND2x1_ASAP7_75t_R _17895_ (.A(_09590_),
    .B(_09591_),
    .Y(_09592_));
 INVx2_ASAP7_75t_R _17896_ (.A(_09592_),
    .Y(_09593_));
 NAND2x1_ASAP7_75t_R _17897_ (.A(_09558_),
    .B(_09593_),
    .Y(_09594_));
 BUFx6f_ASAP7_75t_R _17898_ (.A(_08071_),
    .Y(_09595_));
 AO21x1_ASAP7_75t_R _17899_ (.A1(_09589_),
    .A2(_09594_),
    .B(_09595_),
    .Y(_09596_));
 OAI21x1_ASAP7_75t_R _17900_ (.A1(_09585_),
    .A2(_09596_),
    .B(_00403_),
    .Y(_09597_));
 INVx2_ASAP7_75t_R _17901_ (.A(_08086_),
    .Y(_09598_));
 BUFx10_ASAP7_75t_R _17902_ (.A(_09598_),
    .Y(_09599_));
 OAI21x1_ASAP7_75t_R _17903_ (.A1(_09572_),
    .A2(_09597_),
    .B(_09599_),
    .Y(_09600_));
 AO21x1_ASAP7_75t_R _17904_ (.A1(_09497_),
    .A2(_09498_),
    .B(_09557_),
    .Y(_09601_));
 BUFx4f_ASAP7_75t_R _17905_ (.A(_09500_),
    .Y(_09602_));
 AO21x1_ASAP7_75t_R _17906_ (.A1(_09567_),
    .A2(_09601_),
    .B(_09602_),
    .Y(_09603_));
 OAI21x1_ASAP7_75t_R _17907_ (.A1(_15778_),
    .A2(net13),
    .B(_09514_),
    .Y(_09604_));
 AOI21x1_ASAP7_75t_R _17908_ (.A1(_09501_),
    .A2(_09604_),
    .B(_08064_),
    .Y(_09605_));
 NOR2x2_ASAP7_75t_R _17909_ (.A(net499),
    .B(_08043_),
    .Y(_09606_));
 INVx4_ASAP7_75t_R _17910_ (.A(_09606_),
    .Y(_09607_));
 NAND2x1_ASAP7_75t_R _17911_ (.A(_09535_),
    .B(_09607_),
    .Y(_09608_));
 NAND2x1_ASAP7_75t_R _17912_ (.A(_01141_),
    .B(_09521_),
    .Y(_09609_));
 AO21x1_ASAP7_75t_R _17913_ (.A1(_09608_),
    .A2(_09609_),
    .B(_09525_),
    .Y(_09610_));
 NAND2x1_ASAP7_75t_R _17914_ (.A(_09528_),
    .B(_09610_),
    .Y(_09611_));
 AO21x1_ASAP7_75t_R _17915_ (.A1(_09603_),
    .A2(_09605_),
    .B(_09611_),
    .Y(_09612_));
 AO21x2_ASAP7_75t_R _17916_ (.A1(_09497_),
    .A2(_09498_),
    .B(_00476_),
    .Y(_09613_));
 NAND2x2_ASAP7_75t_R _17917_ (.A(_09613_),
    .B(_09521_),
    .Y(_09614_));
 INVx1_ASAP7_75t_R _17918_ (.A(_01138_),
    .Y(_09615_));
 NOR2x2_ASAP7_75t_R _17919_ (.A(_09615_),
    .B(_09504_),
    .Y(_09616_));
 OA21x2_ASAP7_75t_R _17920_ (.A1(_09614_),
    .A2(_09616_),
    .B(_09525_),
    .Y(_09617_));
 BUFx6f_ASAP7_75t_R _17921_ (.A(_09528_),
    .Y(_09618_));
 AOI21x1_ASAP7_75t_R _17922_ (.A1(_09584_),
    .A2(_09617_),
    .B(_09618_),
    .Y(_09619_));
 INVx1_ASAP7_75t_R _17923_ (.A(_09601_),
    .Y(_09620_));
 NAND2x2_ASAP7_75t_R _17924_ (.A(_09535_),
    .B(_09620_),
    .Y(_09621_));
 NAND2x1_ASAP7_75t_R _17925_ (.A(_09583_),
    .B(_09521_),
    .Y(_09622_));
 NAND2x1_ASAP7_75t_R _17926_ (.A(_09621_),
    .B(_09622_),
    .Y(_09623_));
 OR3x1_ASAP7_75t_R _17927_ (.A(_09623_),
    .B(_09563_),
    .C(_09523_),
    .Y(_09624_));
 AOI21x1_ASAP7_75t_R _17928_ (.A1(_09619_),
    .A2(_09624_),
    .B(_08079_),
    .Y(_09625_));
 AOI21x1_ASAP7_75t_R _17929_ (.A1(_09612_),
    .A2(_09625_),
    .B(_09599_),
    .Y(_09626_));
 NOR2x2_ASAP7_75t_R _17930_ (.A(_01137_),
    .B(_08043_),
    .Y(_09627_));
 INVx3_ASAP7_75t_R _17931_ (.A(_09627_),
    .Y(_09628_));
 AO21x2_ASAP7_75t_R _17932_ (.A1(_08042_),
    .A2(_08038_),
    .B(_01138_),
    .Y(_09629_));
 AO21x2_ASAP7_75t_R _17933_ (.A1(_09628_),
    .A2(_09629_),
    .B(_08056_),
    .Y(_09630_));
 BUFx6f_ASAP7_75t_R _17934_ (.A(_08063_),
    .Y(_09631_));
 INVx3_ASAP7_75t_R _17935_ (.A(_09519_),
    .Y(_09632_));
 NAND3x1_ASAP7_75t_R _17936_ (.A(_09630_),
    .B(_09631_),
    .C(_09632_),
    .Y(_09633_));
 NOR2x1_ASAP7_75t_R _17937_ (.A(_09500_),
    .B(_09628_),
    .Y(_09634_));
 INVx2_ASAP7_75t_R _17938_ (.A(_09634_),
    .Y(_09635_));
 AOI21x1_ASAP7_75t_R _17939_ (.A1(_09602_),
    .A2(_09579_),
    .B(_08064_),
    .Y(_09636_));
 NAND2x1_ASAP7_75t_R _17940_ (.A(_09635_),
    .B(_09636_),
    .Y(_09637_));
 AOI21x1_ASAP7_75t_R _17941_ (.A1(_09633_),
    .A2(_09637_),
    .B(_09595_),
    .Y(_09638_));
 NOR2x1_ASAP7_75t_R _17942_ (.A(_09505_),
    .B(_09592_),
    .Y(_09639_));
 AND3x1_ASAP7_75t_R _17943_ (.A(_09497_),
    .B(_00472_),
    .C(_09498_),
    .Y(_09640_));
 AO21x1_ASAP7_75t_R _17944_ (.A1(net16),
    .A2(_15778_),
    .B(_09590_),
    .Y(_09641_));
 OAI21x1_ASAP7_75t_R _17945_ (.A1(_09640_),
    .A2(_09641_),
    .B(_09563_),
    .Y(_09642_));
 OAI21x1_ASAP7_75t_R _17946_ (.A1(_09639_),
    .A2(_09642_),
    .B(_08072_),
    .Y(_09643_));
 BUFx4f_ASAP7_75t_R _17947_ (.A(_08054_),
    .Y(_09644_));
 NAND2x1_ASAP7_75t_R _17948_ (.A(_09582_),
    .B(_09534_),
    .Y(_09645_));
 AO21x1_ASAP7_75t_R _17949_ (.A1(_09644_),
    .A2(_09645_),
    .B(_09566_),
    .Y(_09646_));
 BUFx6f_ASAP7_75t_R _17950_ (.A(_08063_),
    .Y(_09647_));
 AND2x2_ASAP7_75t_R _17951_ (.A(_09646_),
    .B(_09647_),
    .Y(_09648_));
 NOR2x1_ASAP7_75t_R _17952_ (.A(_09643_),
    .B(_09648_),
    .Y(_09649_));
 OAI21x1_ASAP7_75t_R _17953_ (.A1(_09638_),
    .A2(_09649_),
    .B(_00403_),
    .Y(_09650_));
 NAND2x1_ASAP7_75t_R _17954_ (.A(_09626_),
    .B(_09650_),
    .Y(_09651_));
 OAI21x1_ASAP7_75t_R _17955_ (.A1(_09551_),
    .A2(_09600_),
    .B(_09651_),
    .Y(_00016_));
 INVx2_ASAP7_75t_R _17956_ (.A(_09591_),
    .Y(_09652_));
 NOR2x1_ASAP7_75t_R _17957_ (.A(_09652_),
    .B(_09555_),
    .Y(_09653_));
 INVx2_ASAP7_75t_R _17958_ (.A(_09578_),
    .Y(_09654_));
 NOR2x1_ASAP7_75t_R _17959_ (.A(_00400_),
    .B(_09654_),
    .Y(_09655_));
 OR3x1_ASAP7_75t_R _17960_ (.A(_09653_),
    .B(_09526_),
    .C(_09655_),
    .Y(_09656_));
 AO21x2_ASAP7_75t_R _17961_ (.A1(_09497_),
    .A2(_09498_),
    .B(_01137_),
    .Y(_09657_));
 AO21x1_ASAP7_75t_R _17962_ (.A1(_09538_),
    .A2(_09517_),
    .B(_09644_),
    .Y(_09658_));
 OA21x2_ASAP7_75t_R _17963_ (.A1(_00400_),
    .A2(_09657_),
    .B(_09658_),
    .Y(_09659_));
 AOI21x1_ASAP7_75t_R _17964_ (.A1(_09564_),
    .A2(_09659_),
    .B(_09529_),
    .Y(_09660_));
 BUFx6f_ASAP7_75t_R _17965_ (.A(_09590_),
    .Y(_09661_));
 NAND2x1_ASAP7_75t_R _17966_ (.A(_09661_),
    .B(_09604_),
    .Y(_09662_));
 BUFx6f_ASAP7_75t_R _17967_ (.A(_09535_),
    .Y(_09663_));
 AO21x1_ASAP7_75t_R _17968_ (.A1(_09628_),
    .A2(net15),
    .B(_09663_),
    .Y(_09664_));
 AO21x1_ASAP7_75t_R _17969_ (.A1(_09662_),
    .A2(_09664_),
    .B(_09526_),
    .Y(_09665_));
 NAND2x2_ASAP7_75t_R _17970_ (.A(net2),
    .B(_15766_),
    .Y(_09666_));
 AOI21x1_ASAP7_75t_R _17971_ (.A1(_09560_),
    .A2(_09666_),
    .B(_09661_),
    .Y(_09667_));
 AND3x1_ASAP7_75t_R _17972_ (.A(_09560_),
    .B(_09663_),
    .C(_09607_),
    .Y(_09668_));
 OAI21x1_ASAP7_75t_R _17973_ (.A1(_09667_),
    .A2(_09668_),
    .B(_09564_),
    .Y(_09669_));
 AOI21x1_ASAP7_75t_R _17974_ (.A1(_09665_),
    .A2(_09669_),
    .B(_00402_),
    .Y(_09670_));
 BUFx10_ASAP7_75t_R _17975_ (.A(_08078_),
    .Y(_09671_));
 AOI211x1_ASAP7_75t_R _17976_ (.A1(_09656_),
    .A2(_09660_),
    .B(_09670_),
    .C(_09671_),
    .Y(_09672_));
 NAND2x2_ASAP7_75t_R _17977_ (.A(_00476_),
    .B(_15776_),
    .Y(_09673_));
 OA21x2_ASAP7_75t_R _17978_ (.A1(_09536_),
    .A2(_09673_),
    .B(_09563_),
    .Y(_09674_));
 NOR2x2_ASAP7_75t_R _17979_ (.A(net2),
    .B(net13),
    .Y(_09675_));
 INVx1_ASAP7_75t_R _17980_ (.A(_09496_),
    .Y(_09676_));
 OAI21x1_ASAP7_75t_R _17981_ (.A1(_09675_),
    .A2(_09676_),
    .B(_09663_),
    .Y(_09677_));
 BUFx6f_ASAP7_75t_R _17982_ (.A(_09528_),
    .Y(_09678_));
 AO21x1_ASAP7_75t_R _17983_ (.A1(_09674_),
    .A2(_09677_),
    .B(_09678_),
    .Y(_09679_));
 AO21x2_ASAP7_75t_R _17984_ (.A1(_01137_),
    .A2(_15778_),
    .B(_09500_),
    .Y(_09680_));
 NOR2x2_ASAP7_75t_R _17985_ (.A(_15778_),
    .B(net13),
    .Y(_09681_));
 OA21x2_ASAP7_75t_R _17986_ (.A1(_09680_),
    .A2(_09681_),
    .B(_08064_),
    .Y(_09682_));
 OA21x2_ASAP7_75t_R _17987_ (.A1(_09632_),
    .A2(_09568_),
    .B(_09682_),
    .Y(_09683_));
 OAI21x1_ASAP7_75t_R _17988_ (.A1(_09679_),
    .A2(_09683_),
    .B(_09671_),
    .Y(_09684_));
 OA21x2_ASAP7_75t_R _17989_ (.A1(_09652_),
    .A2(_09627_),
    .B(_09581_),
    .Y(_09685_));
 AO21x1_ASAP7_75t_R _17990_ (.A1(_00478_),
    .A2(_00400_),
    .B(_09685_),
    .Y(_09686_));
 NAND3x2_ASAP7_75t_R _17991_ (.B(_09525_),
    .C(_09621_),
    .Y(_09687_),
    .A(_09635_));
 AO21x2_ASAP7_75t_R _17992_ (.A1(_09497_),
    .A2(_09498_),
    .B(_01136_),
    .Y(_09688_));
 AO21x1_ASAP7_75t_R _17993_ (.A1(_09607_),
    .A2(_09688_),
    .B(_09590_),
    .Y(_09689_));
 INVx1_ASAP7_75t_R _17994_ (.A(_09689_),
    .Y(_09690_));
 OA21x2_ASAP7_75t_R _17995_ (.A1(_09687_),
    .A2(_09690_),
    .B(_09618_),
    .Y(_09691_));
 OA21x2_ASAP7_75t_R _17996_ (.A1(_09564_),
    .A2(_09686_),
    .B(_09691_),
    .Y(_09692_));
 OAI21x1_ASAP7_75t_R _17997_ (.A1(_09684_),
    .A2(_09692_),
    .B(_00404_),
    .Y(_09693_));
 AND3x1_ASAP7_75t_R _17998_ (.A(_09560_),
    .B(_09663_),
    .C(_09520_),
    .Y(_09694_));
 NAND2x2_ASAP7_75t_R _17999_ (.A(_09500_),
    .B(_09558_),
    .Y(_09695_));
 INVx1_ASAP7_75t_R _18000_ (.A(_09695_),
    .Y(_09696_));
 AO21x2_ASAP7_75t_R _18001_ (.A1(_09497_),
    .A2(_09498_),
    .B(_00475_),
    .Y(_09697_));
 AO21x1_ASAP7_75t_R _18002_ (.A1(_09696_),
    .A2(_09697_),
    .B(_09528_),
    .Y(_09698_));
 OAI21x1_ASAP7_75t_R _18003_ (.A1(_09694_),
    .A2(_09698_),
    .B(_00401_),
    .Y(_09699_));
 INVx2_ASAP7_75t_R _18004_ (.A(_09573_),
    .Y(_09700_));
 AND2x2_ASAP7_75t_R _18005_ (.A(_09544_),
    .B(_09496_),
    .Y(_09701_));
 AOI211x1_ASAP7_75t_R _18006_ (.A1(_09700_),
    .A2(_09566_),
    .B(_09701_),
    .C(_09595_),
    .Y(_09702_));
 NAND2x1_ASAP7_75t_R _18007_ (.A(_00477_),
    .B(_08056_),
    .Y(_09703_));
 OA21x2_ASAP7_75t_R _18008_ (.A1(_00472_),
    .A2(_09504_),
    .B(_08054_),
    .Y(_09704_));
 NAND2x2_ASAP7_75t_R _18009_ (.A(_09697_),
    .B(_09704_),
    .Y(_09705_));
 OA21x2_ASAP7_75t_R _18010_ (.A1(_08071_),
    .A2(_09703_),
    .B(_09705_),
    .Y(_09706_));
 OA21x2_ASAP7_75t_R _18011_ (.A1(_09706_),
    .A2(_09546_),
    .B(_08078_),
    .Y(_09707_));
 OAI21x1_ASAP7_75t_R _18012_ (.A1(_09699_),
    .A2(_09702_),
    .B(_09707_),
    .Y(_09708_));
 NOR2x2_ASAP7_75t_R _18013_ (.A(_01139_),
    .B(_09504_),
    .Y(_09709_));
 INVx2_ASAP7_75t_R _18014_ (.A(_09709_),
    .Y(_09710_));
 AO21x1_ASAP7_75t_R _18015_ (.A1(_09710_),
    .A2(_09688_),
    .B(_09547_),
    .Y(_09711_));
 NAND3x1_ASAP7_75t_R _18016_ (.A(_09711_),
    .B(_09658_),
    .C(_09647_),
    .Y(_09712_));
 NAND2x2_ASAP7_75t_R _18017_ (.A(_09697_),
    .B(_09590_),
    .Y(_09713_));
 NOR2x1_ASAP7_75t_R _18018_ (.A(_09713_),
    .B(_09568_),
    .Y(_09714_));
 NAND2x1_ASAP7_75t_R _18019_ (.A(_09525_),
    .B(_09632_),
    .Y(_09715_));
 OA21x2_ASAP7_75t_R _18020_ (.A1(_09714_),
    .A2(_09715_),
    .B(_09528_),
    .Y(_09716_));
 AOI21x1_ASAP7_75t_R _18021_ (.A1(_09712_),
    .A2(_09716_),
    .B(_09671_),
    .Y(_09717_));
 AO21x2_ASAP7_75t_R _18022_ (.A1(_09496_),
    .A2(_09657_),
    .B(_09644_),
    .Y(_09718_));
 AO21x1_ASAP7_75t_R _18023_ (.A1(_09560_),
    .A2(_09534_),
    .B(_09501_),
    .Y(_09719_));
 AOI21x1_ASAP7_75t_R _18024_ (.A1(_09718_),
    .A2(_09719_),
    .B(_09631_),
    .Y(_09720_));
 AO21x1_ASAP7_75t_R _18025_ (.A1(_09607_),
    .A2(_09514_),
    .B(_09536_),
    .Y(_09721_));
 INVx1_ASAP7_75t_R _18026_ (.A(_09681_),
    .Y(_09722_));
 AO21x1_ASAP7_75t_R _18027_ (.A1(_09722_),
    .A2(_09582_),
    .B(_09501_),
    .Y(_09723_));
 AOI21x1_ASAP7_75t_R _18028_ (.A1(_09721_),
    .A2(_09723_),
    .B(_09511_),
    .Y(_09724_));
 OAI21x1_ASAP7_75t_R _18029_ (.A1(_09720_),
    .A2(_09724_),
    .B(_00402_),
    .Y(_09725_));
 AOI21x1_ASAP7_75t_R _18030_ (.A1(_09725_),
    .A2(_09717_),
    .B(_00404_),
    .Y(_09726_));
 NAND2x1_ASAP7_75t_R _18031_ (.A(_09708_),
    .B(_09726_),
    .Y(_09727_));
 OAI21x1_ASAP7_75t_R _18032_ (.A1(_09672_),
    .A2(_09693_),
    .B(_09727_),
    .Y(_00017_));
 NOR2x2_ASAP7_75t_R _18033_ (.A(_09535_),
    .B(_09543_),
    .Y(_09728_));
 NAND2x1_ASAP7_75t_R _18034_ (.A(_09499_),
    .B(_09590_),
    .Y(_09729_));
 INVx1_ASAP7_75t_R _18035_ (.A(_09729_),
    .Y(_09730_));
 AOI22x1_ASAP7_75t_R _18036_ (.A1(_09728_),
    .A2(_09710_),
    .B1(_09700_),
    .B2(_09730_),
    .Y(_09731_));
 AO21x1_ASAP7_75t_R _18037_ (.A1(_09538_),
    .A2(_09688_),
    .B(_09644_),
    .Y(_09732_));
 NOR2x1_ASAP7_75t_R _18038_ (.A(_08064_),
    .B(_09559_),
    .Y(_09733_));
 AOI21x1_ASAP7_75t_R _18039_ (.A1(_09732_),
    .A2(_09733_),
    .B(_09618_),
    .Y(_09734_));
 OAI21x1_ASAP7_75t_R _18040_ (.A1(_09526_),
    .A2(_09731_),
    .B(_09734_),
    .Y(_09735_));
 AO21x1_ASAP7_75t_R _18041_ (.A1(_09591_),
    .A2(_09673_),
    .B(_09590_),
    .Y(_09736_));
 NOR2x2_ASAP7_75t_R _18042_ (.A(_01136_),
    .B(_09504_),
    .Y(_09737_));
 INVx2_ASAP7_75t_R _18043_ (.A(_09737_),
    .Y(_09738_));
 AO21x1_ASAP7_75t_R _18044_ (.A1(_09738_),
    .A2(_09657_),
    .B(_09547_),
    .Y(_09739_));
 AOI21x1_ASAP7_75t_R _18045_ (.A1(_09736_),
    .A2(_09739_),
    .B(_09588_),
    .Y(_09740_));
 NOR2x1_ASAP7_75t_R _18046_ (.A(_09535_),
    .B(_09627_),
    .Y(_09741_));
 AO21x1_ASAP7_75t_R _18047_ (.A1(_09601_),
    .A2(_09741_),
    .B(_08063_),
    .Y(_09742_));
 NAND2x1_ASAP7_75t_R _18048_ (.A(_09504_),
    .B(net2),
    .Y(_09743_));
 AND3x1_ASAP7_75t_R _18049_ (.A(_09743_),
    .B(_09535_),
    .C(_09607_),
    .Y(_09744_));
 NOR2x1_ASAP7_75t_R _18050_ (.A(_09742_),
    .B(_09744_),
    .Y(_09745_));
 OAI21x1_ASAP7_75t_R _18051_ (.A1(_09740_),
    .A2(_09745_),
    .B(_09678_),
    .Y(_09746_));
 AOI21x1_ASAP7_75t_R _18052_ (.A1(_09735_),
    .A2(_09746_),
    .B(_08079_),
    .Y(_09747_));
 AO21x1_ASAP7_75t_R _18053_ (.A1(_09738_),
    .A2(_09629_),
    .B(_09547_),
    .Y(_09748_));
 OAI21x1_ASAP7_75t_R _18054_ (.A1(_09627_),
    .A2(_09543_),
    .B(_09576_),
    .Y(_09749_));
 AOI21x1_ASAP7_75t_R _18055_ (.A1(_09748_),
    .A2(_09749_),
    .B(_09588_),
    .Y(_09750_));
 AO21x1_ASAP7_75t_R _18056_ (.A1(_09743_),
    .A2(_09628_),
    .B(_09581_),
    .Y(_09751_));
 AOI21x1_ASAP7_75t_R _18057_ (.A1(_09630_),
    .A2(_09751_),
    .B(_09631_),
    .Y(_09752_));
 OAI21x1_ASAP7_75t_R _18058_ (.A1(_09750_),
    .A2(_09752_),
    .B(_09678_),
    .Y(_09753_));
 NAND2x1_ASAP7_75t_R _18059_ (.A(_09607_),
    .B(_09519_),
    .Y(_09754_));
 INVx5_ASAP7_75t_R _18060_ (.A(_09616_),
    .Y(_09755_));
 NAND3x2_ASAP7_75t_R _18061_ (.B(_09644_),
    .C(_09755_),
    .Y(_09756_),
    .A(_09560_));
 AOI21x1_ASAP7_75t_R _18062_ (.A1(_09754_),
    .A2(_09756_),
    .B(_09631_),
    .Y(_09757_));
 OAI21x1_ASAP7_75t_R _18063_ (.A1(_09737_),
    .A2(_09543_),
    .B(_09663_),
    .Y(_09758_));
 AO21x1_ASAP7_75t_R _18064_ (.A1(_09700_),
    .A2(_09629_),
    .B(_09581_),
    .Y(_09759_));
 AOI21x1_ASAP7_75t_R _18065_ (.A1(_09758_),
    .A2(_09759_),
    .B(_09511_),
    .Y(_09760_));
 OAI21x1_ASAP7_75t_R _18066_ (.A1(_09757_),
    .A2(_09760_),
    .B(_09595_),
    .Y(_09761_));
 AOI21x1_ASAP7_75t_R _18067_ (.A1(_09753_),
    .A2(_09761_),
    .B(_09671_),
    .Y(_09762_));
 OAI21x1_ASAP7_75t_R _18068_ (.A1(_09747_),
    .A2(_09762_),
    .B(_09599_),
    .Y(_09763_));
 AO21x1_ASAP7_75t_R _18069_ (.A1(_09560_),
    .A2(_09538_),
    .B(_09644_),
    .Y(_09764_));
 AOI21x1_ASAP7_75t_R _18070_ (.A1(_09705_),
    .A2(_09764_),
    .B(_09588_),
    .Y(_09765_));
 NOR2x1_ASAP7_75t_R _18071_ (.A(_09565_),
    .B(_15778_),
    .Y(_09766_));
 INVx1_ASAP7_75t_R _18072_ (.A(_09766_),
    .Y(_09767_));
 AO21x1_ASAP7_75t_R _18073_ (.A1(_09519_),
    .A2(_09767_),
    .B(_09515_),
    .Y(_09768_));
 AND2x2_ASAP7_75t_R _18074_ (.A(_09768_),
    .B(_09563_),
    .Y(_09769_));
 OAI21x1_ASAP7_75t_R _18075_ (.A1(_09765_),
    .A2(_09769_),
    .B(_09595_),
    .Y(_09770_));
 AO21x1_ASAP7_75t_R _18076_ (.A1(_08053_),
    .A2(_08044_),
    .B(_01140_),
    .Y(_09771_));
 AO21x1_ASAP7_75t_R _18077_ (.A1(_09736_),
    .A2(_09771_),
    .B(_09525_),
    .Y(_09772_));
 AND3x1_ASAP7_75t_R _18078_ (.A(_08053_),
    .B(_00479_),
    .C(_08044_),
    .Y(_09773_));
 OAI21x1_ASAP7_75t_R _18079_ (.A1(_09773_),
    .A2(_09559_),
    .B(_09588_),
    .Y(_09774_));
 AO21x1_ASAP7_75t_R _18080_ (.A1(_09772_),
    .A2(_09774_),
    .B(_08072_),
    .Y(_09775_));
 AOI21x1_ASAP7_75t_R _18081_ (.A1(_09770_),
    .A2(_09775_),
    .B(_08079_),
    .Y(_09776_));
 NAND2x1_ASAP7_75t_R _18082_ (.A(_00477_),
    .B(_09663_),
    .Y(_09777_));
 OAI21x1_ASAP7_75t_R _18083_ (.A1(_09675_),
    .A2(_09676_),
    .B(_09521_),
    .Y(_09778_));
 AOI21x1_ASAP7_75t_R _18084_ (.A1(_09777_),
    .A2(_09778_),
    .B(_09631_),
    .Y(_09779_));
 AO21x1_ASAP7_75t_R _18085_ (.A1(_09591_),
    .A2(_09520_),
    .B(_08056_),
    .Y(_09780_));
 NOR2x1_ASAP7_75t_R _18086_ (.A(_09535_),
    .B(_09606_),
    .Y(_09781_));
 NAND2x1_ASAP7_75t_R _18087_ (.A(_09532_),
    .B(_09781_),
    .Y(_09782_));
 AND3x1_ASAP7_75t_R _18088_ (.A(_09780_),
    .B(_08064_),
    .C(_09782_),
    .Y(_09783_));
 OAI21x1_ASAP7_75t_R _18089_ (.A1(_09779_),
    .A2(_09783_),
    .B(_09678_),
    .Y(_09784_));
 INVx1_ASAP7_75t_R _18090_ (.A(_01140_),
    .Y(_09785_));
 OA21x2_ASAP7_75t_R _18091_ (.A1(_09543_),
    .A2(_09785_),
    .B(_09521_),
    .Y(_09786_));
 OR2x2_ASAP7_75t_R _18092_ (.A(_09786_),
    .B(_09744_),
    .Y(_09787_));
 NOR2x2_ASAP7_75t_R _18093_ (.A(_01141_),
    .B(_09521_),
    .Y(_09788_));
 INVx1_ASAP7_75t_R _18094_ (.A(_09505_),
    .Y(_09789_));
 AND3x1_ASAP7_75t_R _18095_ (.A(_09789_),
    .B(_09521_),
    .C(_09613_),
    .Y(_09790_));
 NOR2x1_ASAP7_75t_R _18096_ (.A(_09788_),
    .B(_09790_),
    .Y(_09791_));
 AOI21x1_ASAP7_75t_R _18097_ (.A1(_09511_),
    .A2(_09791_),
    .B(_09618_),
    .Y(_09792_));
 OAI21x1_ASAP7_75t_R _18098_ (.A1(_09564_),
    .A2(_09787_),
    .B(_09792_),
    .Y(_09793_));
 AOI21x1_ASAP7_75t_R _18099_ (.A1(_09784_),
    .A2(_09793_),
    .B(_09671_),
    .Y(_09794_));
 OAI21x1_ASAP7_75t_R _18100_ (.A1(_09776_),
    .A2(_09794_),
    .B(_00404_),
    .Y(_09795_));
 NAND2x1_ASAP7_75t_R _18101_ (.A(_09763_),
    .B(_09795_),
    .Y(_00018_));
 AO21x1_ASAP7_75t_R _18102_ (.A1(_09532_),
    .A2(_09673_),
    .B(_09663_),
    .Y(_09796_));
 AO21x1_ASAP7_75t_R _18103_ (.A1(_09654_),
    .A2(_09607_),
    .B(_09602_),
    .Y(_09797_));
 AO21x1_ASAP7_75t_R _18104_ (.A1(_09796_),
    .A2(_09797_),
    .B(_09546_),
    .Y(_09798_));
 AND2x2_ASAP7_75t_R _18105_ (.A(_08054_),
    .B(_09517_),
    .Y(_09799_));
 NAND2x1_ASAP7_75t_R _18106_ (.A(_09647_),
    .B(_09548_),
    .Y(_09800_));
 AO21x1_ASAP7_75t_R _18107_ (.A1(_09522_),
    .A2(_09799_),
    .B(_09800_),
    .Y(_09801_));
 NAND2x1_ASAP7_75t_R _18108_ (.A(_09798_),
    .B(_09801_),
    .Y(_09802_));
 AND3x1_ASAP7_75t_R _18109_ (.A(_09755_),
    .B(_09536_),
    .C(_09499_),
    .Y(_09803_));
 NOR3x1_ASAP7_75t_R _18110_ (.A(_09803_),
    .B(_09653_),
    .C(_09526_),
    .Y(_09804_));
 NAND2x1_ASAP7_75t_R _18111_ (.A(_09588_),
    .B(_09695_),
    .Y(_09805_));
 INVx1_ASAP7_75t_R _18112_ (.A(_09543_),
    .Y(_09806_));
 NAND2x2_ASAP7_75t_R _18113_ (.A(net2),
    .B(net13),
    .Y(_09807_));
 AND3x1_ASAP7_75t_R _18114_ (.A(_09806_),
    .B(_09663_),
    .C(_09807_),
    .Y(_09808_));
 OAI21x1_ASAP7_75t_R _18115_ (.A1(_09805_),
    .A2(_09808_),
    .B(_09529_),
    .Y(_09809_));
 OAI21x1_ASAP7_75t_R _18116_ (.A1(_09804_),
    .A2(_09809_),
    .B(_00403_),
    .Y(_09810_));
 AOI21x1_ASAP7_75t_R _18117_ (.A1(_00402_),
    .A2(_09802_),
    .B(_09810_),
    .Y(_09811_));
 NOR2x1_ASAP7_75t_R _18118_ (.A(_09573_),
    .B(_09632_),
    .Y(_09812_));
 OAI21x1_ASAP7_75t_R _18119_ (.A1(_09812_),
    .A2(_09808_),
    .B(_09564_),
    .Y(_09813_));
 AND2x2_ASAP7_75t_R _18120_ (.A(_09647_),
    .B(_09506_),
    .Y(_09814_));
 OR3x1_ASAP7_75t_R _18121_ (.A(_09543_),
    .B(_09785_),
    .C(_09602_),
    .Y(_09815_));
 AOI21x1_ASAP7_75t_R _18122_ (.A1(_09814_),
    .A2(_09815_),
    .B(_09595_),
    .Y(_09816_));
 INVx2_ASAP7_75t_R _18123_ (.A(_09514_),
    .Y(_09817_));
 OA21x2_ASAP7_75t_R _18124_ (.A1(_09817_),
    .A2(_09505_),
    .B(_00400_),
    .Y(_09818_));
 OA21x2_ASAP7_75t_R _18125_ (.A1(_09681_),
    .A2(_09531_),
    .B(_09661_),
    .Y(_09819_));
 OAI21x1_ASAP7_75t_R _18126_ (.A1(_09818_),
    .A2(_09819_),
    .B(_00401_),
    .Y(_09820_));
 AO21x1_ASAP7_75t_R _18127_ (.A1(_09628_),
    .A2(_09688_),
    .B(_09581_),
    .Y(_09821_));
 OAI21x1_ASAP7_75t_R _18128_ (.A1(_09573_),
    .A2(_09729_),
    .B(_09821_),
    .Y(_09822_));
 AOI21x1_ASAP7_75t_R _18129_ (.A1(_09564_),
    .A2(_09822_),
    .B(_09678_),
    .Y(_09823_));
 AOI22x1_ASAP7_75t_R _18130_ (.A1(_09813_),
    .A2(_09816_),
    .B1(_09820_),
    .B2(_09823_),
    .Y(_09824_));
 OAI21x1_ASAP7_75t_R _18131_ (.A1(_00403_),
    .A2(_09824_),
    .B(_00404_),
    .Y(_09825_));
 NAND2x1_ASAP7_75t_R _18132_ (.A(_09677_),
    .B(_09605_),
    .Y(_09826_));
 INVx1_ASAP7_75t_R _18133_ (.A(_09799_),
    .Y(_09827_));
 NOR2x2_ASAP7_75t_R _18134_ (.A(_09590_),
    .B(_09567_),
    .Y(_09828_));
 OR2x4_ASAP7_75t_R _18135_ (.A(_09629_),
    .B(_08054_),
    .Y(_09829_));
 NAND2x2_ASAP7_75t_R _18136_ (.A(_08063_),
    .B(_09829_),
    .Y(_09830_));
 NOR2x1_ASAP7_75t_R _18137_ (.A(_09828_),
    .B(_09830_),
    .Y(_09831_));
 OAI21x1_ASAP7_75t_R _18138_ (.A1(_09827_),
    .A2(_09553_),
    .B(_09831_),
    .Y(_09832_));
 AOI21x1_ASAP7_75t_R _18139_ (.A1(_09826_),
    .A2(_09832_),
    .B(_09678_),
    .Y(_09833_));
 NAND2x1_ASAP7_75t_R _18140_ (.A(_09755_),
    .B(_09728_),
    .Y(_09834_));
 AOI21x1_ASAP7_75t_R _18141_ (.A1(_09705_),
    .A2(_09834_),
    .B(_09631_),
    .Y(_09835_));
 AO21x1_ASAP7_75t_R _18142_ (.A1(net16),
    .A2(_15778_),
    .B(_09737_),
    .Y(_09836_));
 OAI21x1_ASAP7_75t_R _18143_ (.A1(_09576_),
    .A2(_09836_),
    .B(_09647_),
    .Y(_09837_));
 NAND2x1_ASAP7_75t_R _18144_ (.A(_09618_),
    .B(_09837_),
    .Y(_09838_));
 OAI21x1_ASAP7_75t_R _18145_ (.A1(_09835_),
    .A2(_09838_),
    .B(_08079_),
    .Y(_09839_));
 NOR2x1_ASAP7_75t_R _18146_ (.A(_09833_),
    .B(_09839_),
    .Y(_09840_));
 NOR2x1_ASAP7_75t_R _18147_ (.A(_09517_),
    .B(_09547_),
    .Y(_09841_));
 AOI221x1_ASAP7_75t_R _18148_ (.A1(_09576_),
    .A2(_09583_),
    .B1(_09841_),
    .B2(_08072_),
    .C(_09588_),
    .Y(_09842_));
 AO21x1_ASAP7_75t_R _18149_ (.A1(_09591_),
    .A2(_09522_),
    .B(_08056_),
    .Y(_09843_));
 AO21x1_ASAP7_75t_R _18150_ (.A1(_09843_),
    .A2(_09506_),
    .B(_08071_),
    .Y(_09844_));
 AO21x1_ASAP7_75t_R _18151_ (.A1(_09842_),
    .A2(_09844_),
    .B(_08079_),
    .Y(_09845_));
 NAND3x1_ASAP7_75t_R _18152_ (.A(_09756_),
    .B(_08072_),
    .C(_09829_),
    .Y(_09846_));
 AO21x1_ASAP7_75t_R _18153_ (.A1(_09799_),
    .A2(_09567_),
    .B(_08071_),
    .Y(_09847_));
 AO21x1_ASAP7_75t_R _18154_ (.A1(_09554_),
    .A2(_09728_),
    .B(_09847_),
    .Y(_09848_));
 AOI21x1_ASAP7_75t_R _18155_ (.A1(_09846_),
    .A2(_09848_),
    .B(_00401_),
    .Y(_09849_));
 NOR2x1_ASAP7_75t_R _18156_ (.A(_09845_),
    .B(_09849_),
    .Y(_09850_));
 OAI21x1_ASAP7_75t_R _18157_ (.A1(_09840_),
    .A2(_09850_),
    .B(_09599_),
    .Y(_09851_));
 OAI21x1_ASAP7_75t_R _18158_ (.A1(_09811_),
    .A2(_09825_),
    .B(_09851_),
    .Y(_00019_));
 OA21x2_ASAP7_75t_R _18159_ (.A1(_09676_),
    .A2(_09817_),
    .B(_00400_),
    .Y(_09852_));
 OAI21x1_ASAP7_75t_R _18160_ (.A1(_09852_),
    .A2(_09687_),
    .B(_09671_),
    .Y(_09853_));
 OA211x2_ASAP7_75t_R _18161_ (.A1(_09573_),
    .A2(_09614_),
    .B(_09739_),
    .C(_09647_),
    .Y(_09854_));
 OAI21x1_ASAP7_75t_R _18162_ (.A1(_09853_),
    .A2(_09854_),
    .B(_09529_),
    .Y(_09855_));
 NAND2x1_ASAP7_75t_R _18163_ (.A(_09525_),
    .B(_09778_),
    .Y(_09856_));
 OA21x2_ASAP7_75t_R _18164_ (.A1(_09856_),
    .A2(_09701_),
    .B(_08079_),
    .Y(_09857_));
 AO21x1_ASAP7_75t_R _18165_ (.A1(_09666_),
    .A2(_09591_),
    .B(_09547_),
    .Y(_09858_));
 AO21x1_ASAP7_75t_R _18166_ (.A1(_09591_),
    .A2(_09520_),
    .B(_09581_),
    .Y(_09859_));
 AO21x1_ASAP7_75t_R _18167_ (.A1(_09858_),
    .A2(_09859_),
    .B(_09511_),
    .Y(_09860_));
 AND2x2_ASAP7_75t_R _18168_ (.A(_09857_),
    .B(_09860_),
    .Y(_09861_));
 NAND2x1_ASAP7_75t_R _18169_ (.A(_09606_),
    .B(_09521_),
    .Y(_09862_));
 AND4x1_ASAP7_75t_R _18170_ (.A(_09630_),
    .B(_09631_),
    .C(_09862_),
    .D(_09829_),
    .Y(_09863_));
 AO21x1_ASAP7_75t_R _18171_ (.A1(_09607_),
    .A2(_09688_),
    .B(_09576_),
    .Y(_09864_));
 AO21x1_ASAP7_75t_R _18172_ (.A1(_09617_),
    .A2(_09864_),
    .B(_08079_),
    .Y(_09865_));
 AOI22x1_ASAP7_75t_R _18173_ (.A1(net16),
    .A2(_15778_),
    .B1(_09663_),
    .B2(_09533_),
    .Y(_09866_));
 OA21x2_ASAP7_75t_R _18174_ (.A1(_01142_),
    .A2(_09644_),
    .B(_09525_),
    .Y(_09867_));
 NAND2x1_ASAP7_75t_R _18175_ (.A(_09866_),
    .B(_09867_),
    .Y(_09868_));
 NAND2x2_ASAP7_75t_R _18176_ (.A(_09500_),
    .B(_09755_),
    .Y(_09869_));
 AND3x1_ASAP7_75t_R _18177_ (.A(_09869_),
    .B(_08063_),
    .C(_09582_),
    .Y(_09870_));
 NOR2x1_ASAP7_75t_R _18178_ (.A(_08078_),
    .B(_09870_),
    .Y(_09871_));
 AOI21x1_ASAP7_75t_R _18179_ (.A1(_09868_),
    .A2(_09871_),
    .B(_09529_),
    .Y(_09872_));
 OAI21x1_ASAP7_75t_R _18180_ (.A1(_09863_),
    .A2(_09865_),
    .B(_09872_),
    .Y(_09873_));
 OAI21x1_ASAP7_75t_R _18181_ (.A1(_09855_),
    .A2(_09861_),
    .B(_09873_),
    .Y(_09874_));
 INVx1_ASAP7_75t_R _18182_ (.A(_09858_),
    .Y(_09875_));
 AO21x1_ASAP7_75t_R _18183_ (.A1(_09728_),
    .A2(_09755_),
    .B(_09563_),
    .Y(_09876_));
 AOI21x1_ASAP7_75t_R _18184_ (.A1(_09661_),
    .A2(_09645_),
    .B(_09647_),
    .Y(_09877_));
 AOI21x1_ASAP7_75t_R _18185_ (.A1(_09877_),
    .A2(_09548_),
    .B(_08072_),
    .Y(_09878_));
 OAI21x1_ASAP7_75t_R _18186_ (.A1(_09875_),
    .A2(_09876_),
    .B(_09878_),
    .Y(_09879_));
 AO21x1_ASAP7_75t_R _18187_ (.A1(net528),
    .A2(_09661_),
    .B(_09781_),
    .Y(_09880_));
 NOR2x1_ASAP7_75t_R _18188_ (.A(_09652_),
    .B(_09869_),
    .Y(_09881_));
 NAND2x1_ASAP7_75t_R _18189_ (.A(_09621_),
    .B(_08064_),
    .Y(_09882_));
 OA21x2_ASAP7_75t_R _18190_ (.A1(_09881_),
    .A2(_09882_),
    .B(_08072_),
    .Y(_09883_));
 OAI21x1_ASAP7_75t_R _18191_ (.A1(_00401_),
    .A2(_09880_),
    .B(_09883_),
    .Y(_09884_));
 AOI21x1_ASAP7_75t_R _18192_ (.A1(_09879_),
    .A2(_09884_),
    .B(_00403_),
    .Y(_09885_));
 NOR2x1_ASAP7_75t_R _18193_ (.A(_09606_),
    .B(_09680_),
    .Y(_09886_));
 INVx1_ASAP7_75t_R _18194_ (.A(_09636_),
    .Y(_09887_));
 AO21x1_ASAP7_75t_R _18195_ (.A1(_01139_),
    .A2(_15776_),
    .B(_09501_),
    .Y(_09888_));
 NAND2x2_ASAP7_75t_R _18196_ (.A(_09577_),
    .B(_15776_),
    .Y(_09889_));
 AOI21x1_ASAP7_75t_R _18197_ (.A1(_00400_),
    .A2(_09889_),
    .B(_09588_),
    .Y(_09890_));
 AOI21x1_ASAP7_75t_R _18198_ (.A1(_09888_),
    .A2(_09890_),
    .B(_09618_),
    .Y(_09891_));
 OAI21x1_ASAP7_75t_R _18199_ (.A1(_09886_),
    .A2(_09887_),
    .B(_09891_),
    .Y(_09892_));
 OAI21x1_ASAP7_75t_R _18200_ (.A1(_09817_),
    .A2(_09573_),
    .B(_09661_),
    .Y(_09893_));
 AOI21x1_ASAP7_75t_R _18201_ (.A1(_09893_),
    .A2(_09718_),
    .B(_09526_),
    .Y(_09894_));
 NOR2x1_ASAP7_75t_R _18202_ (.A(_15778_),
    .B(_09581_),
    .Y(_09895_));
 INVx1_ASAP7_75t_R _18203_ (.A(_09895_),
    .Y(_09896_));
 AO21x1_ASAP7_75t_R _18204_ (.A1(_09560_),
    .A2(_09738_),
    .B(_09602_),
    .Y(_09897_));
 AOI21x1_ASAP7_75t_R _18205_ (.A1(_09896_),
    .A2(_09897_),
    .B(_09546_),
    .Y(_09898_));
 OAI21x1_ASAP7_75t_R _18206_ (.A1(_09894_),
    .A2(_09898_),
    .B(_09529_),
    .Y(_09899_));
 AOI21x1_ASAP7_75t_R _18207_ (.A1(_09892_),
    .A2(_09899_),
    .B(_09671_),
    .Y(_09900_));
 OAI21x1_ASAP7_75t_R _18208_ (.A1(_09885_),
    .A2(_09900_),
    .B(_09599_),
    .Y(_09901_));
 OAI21x1_ASAP7_75t_R _18209_ (.A1(_09599_),
    .A2(_09874_),
    .B(_09901_),
    .Y(_00020_));
 AND3x1_ASAP7_75t_R _18210_ (.A(_09755_),
    .B(_09591_),
    .C(_09536_),
    .Y(_09902_));
 NOR2x1_ASAP7_75t_R _18211_ (.A(_09518_),
    .B(_09695_),
    .Y(_09903_));
 OR3x1_ASAP7_75t_R _18212_ (.A(_09902_),
    .B(_09526_),
    .C(_09903_),
    .Y(_09904_));
 NAND2x1_ASAP7_75t_R _18213_ (.A(_09576_),
    .B(net16),
    .Y(_09905_));
 AND3x1_ASAP7_75t_R _18214_ (.A(_09545_),
    .B(_09511_),
    .C(_09905_),
    .Y(_09906_));
 NOR2x1_ASAP7_75t_R _18215_ (.A(_09529_),
    .B(_09906_),
    .Y(_09907_));
 OA21x2_ASAP7_75t_R _18216_ (.A1(_09536_),
    .A2(_09522_),
    .B(_08064_),
    .Y(_09908_));
 OA21x2_ASAP7_75t_R _18217_ (.A1(_09553_),
    .A2(_09713_),
    .B(_09908_),
    .Y(_09909_));
 AO21x1_ASAP7_75t_R _18218_ (.A1(_09806_),
    .A2(_09628_),
    .B(_09602_),
    .Y(_09910_));
 AO21x1_ASAP7_75t_R _18219_ (.A1(_09636_),
    .A2(_09910_),
    .B(_09595_),
    .Y(_09911_));
 OAI21x1_ASAP7_75t_R _18220_ (.A1(_09909_),
    .A2(_09911_),
    .B(_08079_),
    .Y(_09912_));
 AOI21x1_ASAP7_75t_R _18221_ (.A1(_09904_),
    .A2(_09907_),
    .B(_09912_),
    .Y(_09913_));
 AND3x1_ASAP7_75t_R _18222_ (.A(_09635_),
    .B(_09546_),
    .C(_09555_),
    .Y(_09914_));
 NOR2x1_ASAP7_75t_R _18223_ (.A(_09647_),
    .B(_09728_),
    .Y(_09915_));
 AO21x1_ASAP7_75t_R _18224_ (.A1(_09654_),
    .A2(_09673_),
    .B(_09576_),
    .Y(_09916_));
 AO21x1_ASAP7_75t_R _18225_ (.A1(_09915_),
    .A2(_09916_),
    .B(_09678_),
    .Y(_09917_));
 AO21x1_ASAP7_75t_R _18226_ (.A1(_09738_),
    .A2(_09517_),
    .B(_08056_),
    .Y(_09918_));
 AO21x1_ASAP7_75t_R _18227_ (.A1(_09522_),
    .A2(_09499_),
    .B(_09590_),
    .Y(_09919_));
 AO21x1_ASAP7_75t_R _18228_ (.A1(_09918_),
    .A2(_09919_),
    .B(_09563_),
    .Y(_09920_));
 NAND2x1_ASAP7_75t_R _18229_ (.A(_00472_),
    .B(_09547_),
    .Y(_09921_));
 AO21x1_ASAP7_75t_R _18230_ (.A1(_09921_),
    .A2(_09713_),
    .B(_09647_),
    .Y(_09922_));
 AO21x1_ASAP7_75t_R _18231_ (.A1(_09920_),
    .A2(_09922_),
    .B(_09595_),
    .Y(_09923_));
 OAI21x1_ASAP7_75t_R _18232_ (.A1(_09914_),
    .A2(_09917_),
    .B(_09923_),
    .Y(_09924_));
 OAI21x1_ASAP7_75t_R _18233_ (.A1(_00403_),
    .A2(_09924_),
    .B(_09599_),
    .Y(_09925_));
 AND3x1_ASAP7_75t_R _18234_ (.A(_09654_),
    .B(_09547_),
    .C(_09522_),
    .Y(_09926_));
 AOI21x1_ASAP7_75t_R _18235_ (.A1(_09666_),
    .A2(_09569_),
    .B(_09926_),
    .Y(_09927_));
 AO21x1_ASAP7_75t_R _18236_ (.A1(net16),
    .A2(_09581_),
    .B(_15771_),
    .Y(_09928_));
 AOI21x1_ASAP7_75t_R _18237_ (.A1(_09928_),
    .A2(_09575_),
    .B(_09618_),
    .Y(_09929_));
 OAI21x1_ASAP7_75t_R _18238_ (.A1(_09564_),
    .A2(_09927_),
    .B(_09929_),
    .Y(_09930_));
 OA21x2_ASAP7_75t_R _18239_ (.A1(_09652_),
    .A2(_09709_),
    .B(_09644_),
    .Y(_09931_));
 NAND2x1_ASAP7_75t_R _18240_ (.A(_09862_),
    .B(_08064_),
    .Y(_09932_));
 OA21x2_ASAP7_75t_R _18241_ (.A1(_09931_),
    .A2(_09932_),
    .B(_09528_),
    .Y(_09933_));
 AO22x1_ASAP7_75t_R _18242_ (.A1(_09644_),
    .A2(_09738_),
    .B1(_09519_),
    .B2(_09534_),
    .Y(_09934_));
 NAND2x1_ASAP7_75t_R _18243_ (.A(_09511_),
    .B(_09934_),
    .Y(_09935_));
 AOI21x1_ASAP7_75t_R _18244_ (.A1(_09933_),
    .A2(_09935_),
    .B(_08079_),
    .Y(_09936_));
 AOI21x1_ASAP7_75t_R _18245_ (.A1(_09930_),
    .A2(_09936_),
    .B(_09599_),
    .Y(_09937_));
 AND3x1_ASAP7_75t_R _18246_ (.A(_09755_),
    .B(_09661_),
    .C(_09613_),
    .Y(_09938_));
 AO21x1_ASAP7_75t_R _18247_ (.A1(_09728_),
    .A2(_09767_),
    .B(_09588_),
    .Y(_09939_));
 OAI21x1_ASAP7_75t_R _18248_ (.A1(_09938_),
    .A2(_09939_),
    .B(_00402_),
    .Y(_09940_));
 AO21x1_ASAP7_75t_R _18249_ (.A1(_09738_),
    .A2(_09657_),
    .B(_09536_),
    .Y(_09941_));
 AND3x1_ASAP7_75t_R _18250_ (.A(_09575_),
    .B(_09584_),
    .C(_09941_),
    .Y(_09942_));
 NAND2x1_ASAP7_75t_R _18251_ (.A(_09673_),
    .B(_09680_),
    .Y(_09943_));
 OA21x2_ASAP7_75t_R _18252_ (.A1(_09943_),
    .A2(_09588_),
    .B(_09618_),
    .Y(_09944_));
 NAND2x1_ASAP7_75t_R _18253_ (.A(_09525_),
    .B(_09829_),
    .Y(_09945_));
 OR3x1_ASAP7_75t_R _18254_ (.A(_09945_),
    .B(_09828_),
    .C(_09799_),
    .Y(_09946_));
 AOI21x1_ASAP7_75t_R _18255_ (.A1(_09944_),
    .A2(_09946_),
    .B(_09671_),
    .Y(_09947_));
 OAI21x1_ASAP7_75t_R _18256_ (.A1(_09940_),
    .A2(_09942_),
    .B(_09947_),
    .Y(_09948_));
 NAND2x1_ASAP7_75t_R _18257_ (.A(_09937_),
    .B(_09948_),
    .Y(_09949_));
 OAI21x1_ASAP7_75t_R _18258_ (.A1(_09913_),
    .A2(_09925_),
    .B(_09949_),
    .Y(_00021_));
 AND3x1_ASAP7_75t_R _18259_ (.A(_09755_),
    .B(_09536_),
    .C(_09586_),
    .Y(_09950_));
 NOR2x1_ASAP7_75t_R _18260_ (.A(_09661_),
    .B(_09538_),
    .Y(_09951_));
 NAND2x1_ASAP7_75t_R _18261_ (.A(_09622_),
    .B(_09511_),
    .Y(_09952_));
 OR3x1_ASAP7_75t_R _18262_ (.A(_09950_),
    .B(_09951_),
    .C(_09952_),
    .Y(_09953_));
 NOR2x1_ASAP7_75t_R _18263_ (.A(_09543_),
    .B(_09608_),
    .Y(_09954_));
 OR3x1_ASAP7_75t_R _18264_ (.A(_09830_),
    .B(_09954_),
    .C(_09828_),
    .Y(_09955_));
 AND2x2_ASAP7_75t_R _18265_ (.A(_09955_),
    .B(_09678_),
    .Y(_09956_));
 AO21x1_ASAP7_75t_R _18266_ (.A1(_09576_),
    .A2(_09709_),
    .B(_09515_),
    .Y(_09957_));
 OAI21x1_ASAP7_75t_R _18267_ (.A1(_09830_),
    .A2(_09957_),
    .B(_09595_),
    .Y(_09958_));
 AO21x1_ASAP7_75t_R _18268_ (.A1(_15771_),
    .A2(_09661_),
    .B(_09647_),
    .Y(_09959_));
 AND3x1_ASAP7_75t_R _18269_ (.A(_09700_),
    .B(_09547_),
    .C(_09807_),
    .Y(_09960_));
 NOR2x1_ASAP7_75t_R _18270_ (.A(_09959_),
    .B(_09960_),
    .Y(_09961_));
 OAI21x1_ASAP7_75t_R _18271_ (.A1(_09958_),
    .A2(_09961_),
    .B(_00404_),
    .Y(_09962_));
 AOI21x1_ASAP7_75t_R _18272_ (.A1(_09953_),
    .A2(_09956_),
    .B(_09962_),
    .Y(_09963_));
 INVx1_ASAP7_75t_R _18273_ (.A(_09499_),
    .Y(_09964_));
 AOI211x1_ASAP7_75t_R _18274_ (.A1(_09661_),
    .A2(_09964_),
    .B(_09945_),
    .C(_09828_),
    .Y(_09965_));
 AO21x1_ASAP7_75t_R _18275_ (.A1(_00478_),
    .A2(_09576_),
    .B(_09563_),
    .Y(_09966_));
 OAI21x1_ASAP7_75t_R _18276_ (.A1(_09966_),
    .A2(_09561_),
    .B(_09678_),
    .Y(_09967_));
 OAI21x1_ASAP7_75t_R _18277_ (.A1(_09965_),
    .A2(_09967_),
    .B(_09598_),
    .Y(_09968_));
 NAND2x1_ASAP7_75t_R _18278_ (.A(_09673_),
    .B(_09593_),
    .Y(_09969_));
 AO21x1_ASAP7_75t_R _18279_ (.A1(_09806_),
    .A2(_09807_),
    .B(_09581_),
    .Y(_09970_));
 AOI21x1_ASAP7_75t_R _18280_ (.A1(_09969_),
    .A2(_09970_),
    .B(_09546_),
    .Y(_09971_));
 NAND2x1_ASAP7_75t_R _18281_ (.A(_09586_),
    .B(_09590_),
    .Y(_09972_));
 OA21x2_ASAP7_75t_R _18282_ (.A1(_09681_),
    .A2(_09972_),
    .B(_08064_),
    .Y(_09973_));
 AO21x1_ASAP7_75t_R _18283_ (.A1(_09970_),
    .A2(_09973_),
    .B(_09618_),
    .Y(_09974_));
 NOR2x1_ASAP7_75t_R _18284_ (.A(_09971_),
    .B(_09974_),
    .Y(_09975_));
 OAI21x1_ASAP7_75t_R _18285_ (.A1(_09968_),
    .A2(_09975_),
    .B(_00403_),
    .Y(_09976_));
 OAI21x1_ASAP7_75t_R _18286_ (.A1(_09704_),
    .A2(_09881_),
    .B(_00401_),
    .Y(_09977_));
 NAND3x1_ASAP7_75t_R _18287_ (.A(_09977_),
    .B(_09529_),
    .C(_09742_),
    .Y(_09978_));
 AND3x1_ASAP7_75t_R _18288_ (.A(_09554_),
    .B(_09602_),
    .C(_09499_),
    .Y(_09979_));
 AO21x2_ASAP7_75t_R _18289_ (.A1(_09681_),
    .A2(_09663_),
    .B(_09563_),
    .Y(_09980_));
 NOR2x1_ASAP7_75t_R _18290_ (.A(_09979_),
    .B(_09980_),
    .Y(_09981_));
 AOI211x1_ASAP7_75t_R _18291_ (.A1(_00480_),
    .A2(_00400_),
    .B(_09902_),
    .C(_00401_),
    .Y(_09982_));
 OAI21x1_ASAP7_75t_R _18292_ (.A1(_09981_),
    .A2(_09982_),
    .B(_00402_),
    .Y(_09983_));
 AOI21x1_ASAP7_75t_R _18293_ (.A1(_09978_),
    .A2(_09983_),
    .B(_00404_),
    .Y(_09984_));
 NAND2x1_ASAP7_75t_R _18294_ (.A(_09591_),
    .B(_09696_),
    .Y(_09985_));
 AO21x1_ASAP7_75t_R _18295_ (.A1(_09710_),
    .A2(net15),
    .B(_09602_),
    .Y(_09986_));
 AO21x1_ASAP7_75t_R _18296_ (.A1(_09985_),
    .A2(_09986_),
    .B(_09546_),
    .Y(_09987_));
 AO21x1_ASAP7_75t_R _18297_ (.A1(_09559_),
    .A2(net15),
    .B(_09773_),
    .Y(_09988_));
 NAND2x1_ASAP7_75t_R _18298_ (.A(_09546_),
    .B(_09988_),
    .Y(_09989_));
 AOI21x1_ASAP7_75t_R _18299_ (.A1(_09987_),
    .A2(_09989_),
    .B(_09529_),
    .Y(_09990_));
 INVx1_ASAP7_75t_R _18300_ (.A(_09614_),
    .Y(_09991_));
 AOI211x1_ASAP7_75t_R _18301_ (.A1(_09722_),
    .A2(_09991_),
    .B(_09954_),
    .C(_00401_),
    .Y(_09992_));
 AOI21x1_ASAP7_75t_R _18302_ (.A1(_09496_),
    .A2(_09991_),
    .B(_09523_),
    .Y(_09993_));
 AO21x1_ASAP7_75t_R _18303_ (.A1(_09993_),
    .A2(_09546_),
    .B(_08072_),
    .Y(_09994_));
 OAI21x1_ASAP7_75t_R _18304_ (.A1(_09992_),
    .A2(_09994_),
    .B(_00404_),
    .Y(_09995_));
 OAI21x1_ASAP7_75t_R _18305_ (.A1(_09990_),
    .A2(_09995_),
    .B(_09671_),
    .Y(_09996_));
 OAI22x1_ASAP7_75t_R _18306_ (.A1(_09963_),
    .A2(_09976_),
    .B1(_09984_),
    .B2(_09996_),
    .Y(_00022_));
 NAND2x1_ASAP7_75t_R _18307_ (.A(_09567_),
    .B(_09799_),
    .Y(_09997_));
 AO21x1_ASAP7_75t_R _18308_ (.A1(_09997_),
    .A2(_09689_),
    .B(_09526_),
    .Y(_09998_));
 OAI21x1_ASAP7_75t_R _18309_ (.A1(_09950_),
    .A2(_09786_),
    .B(_09564_),
    .Y(_09999_));
 AOI21x1_ASAP7_75t_R _18310_ (.A1(_09998_),
    .A2(_09999_),
    .B(_00402_),
    .Y(_10000_));
 AO21x1_ASAP7_75t_R _18311_ (.A1(_09576_),
    .A2(_09817_),
    .B(_09563_),
    .Y(_10001_));
 AOI211x1_ASAP7_75t_R _18312_ (.A1(_09569_),
    .A2(_09613_),
    .B(_09951_),
    .C(_10001_),
    .Y(_10002_));
 OA21x2_ASAP7_75t_R _18313_ (.A1(_09869_),
    .A2(_09652_),
    .B(_09972_),
    .Y(_10003_));
 AO21x1_ASAP7_75t_R _18314_ (.A1(_10003_),
    .A2(_09526_),
    .B(_09678_),
    .Y(_10004_));
 OAI21x1_ASAP7_75t_R _18315_ (.A1(_10002_),
    .A2(_10004_),
    .B(_09599_),
    .Y(_10005_));
 OAI21x1_ASAP7_75t_R _18316_ (.A1(_10000_),
    .A2(_10005_),
    .B(_00403_),
    .Y(_10006_));
 NOR2x1_ASAP7_75t_R _18317_ (.A(_01137_),
    .B(_00400_),
    .Y(_10007_));
 OAI21x1_ASAP7_75t_R _18318_ (.A1(_10007_),
    .A2(_09960_),
    .B(_00401_),
    .Y(_10008_));
 AO21x1_ASAP7_75t_R _18319_ (.A1(_09700_),
    .A2(_09514_),
    .B(_09536_),
    .Y(_10009_));
 AO21x1_ASAP7_75t_R _18320_ (.A1(_09710_),
    .A2(_09514_),
    .B(_09501_),
    .Y(_10010_));
 AO21x1_ASAP7_75t_R _18321_ (.A1(_10009_),
    .A2(_10010_),
    .B(_09631_),
    .Y(_10011_));
 AOI21x1_ASAP7_75t_R _18322_ (.A1(_10008_),
    .A2(_10011_),
    .B(_00402_),
    .Y(_10012_));
 AO21x1_ASAP7_75t_R _18323_ (.A1(_09522_),
    .A2(net15),
    .B(_09644_),
    .Y(_10013_));
 AO21x1_ASAP7_75t_R _18324_ (.A1(_09538_),
    .A2(_09514_),
    .B(_09547_),
    .Y(_10014_));
 NAND2x1_ASAP7_75t_R _18325_ (.A(_10013_),
    .B(_10014_),
    .Y(_10015_));
 OAI21x1_ASAP7_75t_R _18326_ (.A1(_09546_),
    .A2(_10015_),
    .B(_09595_),
    .Y(_10016_));
 AND3x1_ASAP7_75t_R _18327_ (.A(_09743_),
    .B(_09536_),
    .C(_09889_),
    .Y(_10017_));
 NOR2x1_ASAP7_75t_R _18328_ (.A(_10017_),
    .B(_09876_),
    .Y(_10018_));
 OAI21x1_ASAP7_75t_R _18329_ (.A1(_10016_),
    .A2(_10018_),
    .B(_00404_),
    .Y(_10019_));
 NOR2x1_ASAP7_75t_R _18330_ (.A(_10012_),
    .B(_10019_),
    .Y(_10020_));
 AO21x1_ASAP7_75t_R _18331_ (.A1(_09889_),
    .A2(_09593_),
    .B(_09856_),
    .Y(_10021_));
 OAI22x1_ASAP7_75t_R _18332_ (.A1(_09641_),
    .A2(_09573_),
    .B1(net13),
    .B2(_00400_),
    .Y(_10022_));
 OA21x2_ASAP7_75t_R _18333_ (.A1(_10022_),
    .A2(_09564_),
    .B(_00402_),
    .Y(_10023_));
 AO21x1_ASAP7_75t_R _18334_ (.A1(_09538_),
    .A2(net15),
    .B(_09501_),
    .Y(_10024_));
 AND3x1_ASAP7_75t_R _18335_ (.A(_10024_),
    .B(_09631_),
    .C(_09614_),
    .Y(_10025_));
 AO21x1_ASAP7_75t_R _18336_ (.A1(_09602_),
    .A2(_09654_),
    .B(_09799_),
    .Y(_10026_));
 AO21x1_ASAP7_75t_R _18337_ (.A1(_10026_),
    .A2(_09526_),
    .B(_08072_),
    .Y(_10027_));
 OAI21x1_ASAP7_75t_R _18338_ (.A1(_10025_),
    .A2(_10027_),
    .B(_09599_),
    .Y(_10028_));
 AOI21x1_ASAP7_75t_R _18339_ (.A1(_10021_),
    .A2(_10023_),
    .B(_10028_),
    .Y(_10029_));
 AND3x1_ASAP7_75t_R _18340_ (.A(_09574_),
    .B(_09631_),
    .C(_09621_),
    .Y(_10030_));
 NAND2x1_ASAP7_75t_R _18341_ (.A(net527),
    .B(_08056_),
    .Y(_10031_));
 OA21x2_ASAP7_75t_R _18342_ (.A1(_09501_),
    .A2(_09710_),
    .B(_10031_),
    .Y(_10032_));
 AO21x1_ASAP7_75t_R _18343_ (.A1(_10032_),
    .A2(_09511_),
    .B(_09618_),
    .Y(_10033_));
 AOI21x1_ASAP7_75t_R _18344_ (.A1(_09718_),
    .A2(_10030_),
    .B(_10033_),
    .Y(_10034_));
 AO21x1_ASAP7_75t_R _18345_ (.A1(_09789_),
    .A2(_09629_),
    .B(_09602_),
    .Y(_10035_));
 AO21x1_ASAP7_75t_R _18346_ (.A1(_09867_),
    .A2(_10035_),
    .B(_08072_),
    .Y(_10036_));
 AND3x1_ASAP7_75t_R _18347_ (.A(_09789_),
    .B(_09501_),
    .C(_09499_),
    .Y(_10037_));
 NOR3x1_ASAP7_75t_R _18348_ (.A(_09980_),
    .B(_09788_),
    .C(_10037_),
    .Y(_10038_));
 OAI21x1_ASAP7_75t_R _18349_ (.A1(_10036_),
    .A2(_10038_),
    .B(_00404_),
    .Y(_10039_));
 OAI21x1_ASAP7_75t_R _18350_ (.A1(_10034_),
    .A2(_10039_),
    .B(_09671_),
    .Y(_10040_));
 OAI22x1_ASAP7_75t_R _18351_ (.A1(_10006_),
    .A2(_10020_),
    .B1(_10029_),
    .B2(_10040_),
    .Y(_00023_));
 INVx4_ASAP7_75t_R _18352_ (.A(_15789_),
    .Y(_15783_));
 BUFx12f_ASAP7_75t_R _18353_ (.A(_08208_),
    .Y(_15794_));
 AOI21x1_ASAP7_75t_R _18354_ (.A1(_08183_),
    .A2(net825),
    .B(_15794_),
    .Y(_10041_));
 INVx4_ASAP7_75t_R _18355_ (.A(_10041_),
    .Y(_10042_));
 BUFx4f_ASAP7_75t_R _18356_ (.A(_08207_),
    .Y(_10043_));
 BUFx4f_ASAP7_75t_R _18357_ (.A(_08204_),
    .Y(_10044_));
 AO21x2_ASAP7_75t_R _18358_ (.A1(_10043_),
    .A2(_10044_),
    .B(_01146_),
    .Y(_10045_));
 BUFx6f_ASAP7_75t_R _18359_ (.A(_08216_),
    .Y(_10046_));
 AO21x1_ASAP7_75t_R _18360_ (.A1(_10042_),
    .A2(_10045_),
    .B(_10046_),
    .Y(_10047_));
 INVx3_ASAP7_75t_R _18361_ (.A(_08225_),
    .Y(_10048_));
 BUFx6f_ASAP7_75t_R _18362_ (.A(_10048_),
    .Y(_10049_));
 BUFx10_ASAP7_75t_R _18363_ (.A(_10049_),
    .Y(_10050_));
 INVx2_ASAP7_75t_R _18364_ (.A(_00484_),
    .Y(_10051_));
 AO21x2_ASAP7_75t_R _18365_ (.A1(_10043_),
    .A2(_10044_),
    .B(_10051_),
    .Y(_10052_));
 INVx2_ASAP7_75t_R _18366_ (.A(_10052_),
    .Y(_10053_));
 BUFx16f_ASAP7_75t_R _18367_ (.A(_08208_),
    .Y(_10054_));
 NOR2x2_ASAP7_75t_R _18368_ (.A(_15786_),
    .B(_10054_),
    .Y(_10055_));
 BUFx6f_ASAP7_75t_R _18369_ (.A(_08216_),
    .Y(_10056_));
 OAI21x1_ASAP7_75t_R _18370_ (.A1(_10053_),
    .A2(_10055_),
    .B(_10056_),
    .Y(_10057_));
 NAND3x1_ASAP7_75t_R _18371_ (.A(_10047_),
    .B(_10050_),
    .C(_10057_),
    .Y(_10058_));
 NOR2x2_ASAP7_75t_R _18372_ (.A(_15796_),
    .B(net11),
    .Y(_10059_));
 INVx2_ASAP7_75t_R _18373_ (.A(_10059_),
    .Y(_10060_));
 INVx1_ASAP7_75t_R _18374_ (.A(_00485_),
    .Y(_10061_));
 NOR2x2_ASAP7_75t_R _18375_ (.A(_10061_),
    .B(_10054_),
    .Y(_10062_));
 INVx3_ASAP7_75t_R _18376_ (.A(_10062_),
    .Y(_10063_));
 AO21x1_ASAP7_75t_R _18377_ (.A1(_10060_),
    .A2(_10063_),
    .B(_00395_),
    .Y(_10064_));
 AO21x2_ASAP7_75t_R _18378_ (.A1(_10043_),
    .A2(_10044_),
    .B(_01143_),
    .Y(_10065_));
 INVx2_ASAP7_75t_R _18379_ (.A(_10065_),
    .Y(_10066_));
 NOR2x1_ASAP7_75t_R _18380_ (.A(_10055_),
    .B(_10066_),
    .Y(_10067_));
 INVx1_ASAP7_75t_R _18381_ (.A(_01110_),
    .Y(_10068_));
 XOR2x2_ASAP7_75t_R _18382_ (.A(_08213_),
    .B(_10068_),
    .Y(_10069_));
 NOR2x2_ASAP7_75t_R _18383_ (.A(net114),
    .B(_07956_),
    .Y(_10070_));
 AO21x2_ASAP7_75t_R _18384_ (.A1(_10069_),
    .A2(_07979_),
    .B(_10070_),
    .Y(_10071_));
 BUFx6f_ASAP7_75t_R _18385_ (.A(_10071_),
    .Y(_10072_));
 BUFx6f_ASAP7_75t_R _18386_ (.A(_10072_),
    .Y(_10073_));
 BUFx6f_ASAP7_75t_R _18387_ (.A(_08225_),
    .Y(_10074_));
 OA21x2_ASAP7_75t_R _18388_ (.A1(_10067_),
    .A2(_10073_),
    .B(_10074_),
    .Y(_10075_));
 AOI21x1_ASAP7_75t_R _18389_ (.A1(_10064_),
    .A2(_10075_),
    .B(_00397_),
    .Y(_10076_));
 NOR2x2_ASAP7_75t_R _18390_ (.A(net823),
    .B(_15794_),
    .Y(_10077_));
 BUFx10_ASAP7_75t_R _18391_ (.A(_08216_),
    .Y(_10078_));
 NOR2x1_ASAP7_75t_R _18392_ (.A(_10077_),
    .B(_10078_),
    .Y(_10079_));
 AO21x1_ASAP7_75t_R _18393_ (.A1(_10043_),
    .A2(_10044_),
    .B(_01144_),
    .Y(_10080_));
 INVx1_ASAP7_75t_R _18394_ (.A(_10080_),
    .Y(_10081_));
 BUFx6f_ASAP7_75t_R _18395_ (.A(_10078_),
    .Y(_10082_));
 OA21x2_ASAP7_75t_R _18396_ (.A1(_10062_),
    .A2(_10081_),
    .B(_10082_),
    .Y(_10083_));
 OAI21x1_ASAP7_75t_R _18397_ (.A1(_10079_),
    .A2(_10083_),
    .B(_10050_),
    .Y(_10084_));
 INVx1_ASAP7_75t_R _18398_ (.A(_00483_),
    .Y(_10085_));
 AO21x2_ASAP7_75t_R _18399_ (.A1(_10043_),
    .A2(_10044_),
    .B(_10085_),
    .Y(_10086_));
 INVx4_ASAP7_75t_R _18400_ (.A(_10086_),
    .Y(_10087_));
 NOR2x2_ASAP7_75t_R _18401_ (.A(_07967_),
    .B(_10069_),
    .Y(_10088_));
 INVx1_ASAP7_75t_R _18402_ (.A(_01143_),
    .Y(_10089_));
 NOR2x2_ASAP7_75t_R _18403_ (.A(_10089_),
    .B(_10054_),
    .Y(_10090_));
 INVx1_ASAP7_75t_R _18404_ (.A(_10090_),
    .Y(_10091_));
 OAI21x1_ASAP7_75t_R _18405_ (.A1(_08215_),
    .A2(_10088_),
    .B(_10091_),
    .Y(_10092_));
 NOR2x1_ASAP7_75t_R _18406_ (.A(_10087_),
    .B(_10092_),
    .Y(_10093_));
 NOR2x2_ASAP7_75t_R _18407_ (.A(net822),
    .B(_15796_),
    .Y(_10094_));
 XNOR2x1_ASAP7_75t_R _18408_ (.B(_01110_),
    .Y(_10095_),
    .A(_08211_));
 INVx3_ASAP7_75t_R _18409_ (.A(_01046_),
    .Y(_10096_));
 XOR2x1_ASAP7_75t_R _18410_ (.A(_08210_),
    .Y(_10097_),
    .B(_10096_));
 NAND2x1_ASAP7_75t_R _18411_ (.A(_10095_),
    .B(_10097_),
    .Y(_10098_));
 INVx1_ASAP7_75t_R _18412_ (.A(_10095_),
    .Y(_10099_));
 NAND2x1_ASAP7_75t_R _18413_ (.A(_10099_),
    .B(_08362_),
    .Y(_10100_));
 AO21x1_ASAP7_75t_R _18414_ (.A1(_10098_),
    .A2(_10100_),
    .B(_07967_),
    .Y(_10101_));
 BUFx4f_ASAP7_75t_R _18415_ (.A(_10101_),
    .Y(_10102_));
 CKINVDCx5p33_ASAP7_75t_R _18416_ (.A(_10070_),
    .Y(_10103_));
 NOR2x1_ASAP7_75t_R _18417_ (.A(_00485_),
    .B(_15794_),
    .Y(_10104_));
 AO21x1_ASAP7_75t_R _18418_ (.A1(_10102_),
    .A2(_10103_),
    .B(_10104_),
    .Y(_10105_));
 NOR2x1_ASAP7_75t_R _18419_ (.A(_10094_),
    .B(_10105_),
    .Y(_10106_));
 OAI21x1_ASAP7_75t_R _18420_ (.A1(_10093_),
    .A2(_10106_),
    .B(_00396_),
    .Y(_10107_));
 BUFx6f_ASAP7_75t_R _18421_ (.A(_08234_),
    .Y(_10108_));
 AOI21x1_ASAP7_75t_R _18422_ (.A1(_10084_),
    .A2(_10107_),
    .B(_10108_),
    .Y(_10109_));
 INVx3_ASAP7_75t_R _18423_ (.A(_08243_),
    .Y(_10110_));
 BUFx10_ASAP7_75t_R _18424_ (.A(_10110_),
    .Y(_10111_));
 AOI211x1_ASAP7_75t_R _18425_ (.A1(_10058_),
    .A2(_10076_),
    .B(_10109_),
    .C(_10111_),
    .Y(_10112_));
 AND2x2_ASAP7_75t_R _18426_ (.A(_15794_),
    .B(_00481_),
    .Y(_10113_));
 AO21x2_ASAP7_75t_R _18427_ (.A1(_10043_),
    .A2(_10044_),
    .B(_00483_),
    .Y(_10114_));
 INVx2_ASAP7_75t_R _18428_ (.A(_10114_),
    .Y(_10115_));
 BUFx6f_ASAP7_75t_R _18429_ (.A(_10115_),
    .Y(_10116_));
 NOR2x2_ASAP7_75t_R _18430_ (.A(_10051_),
    .B(_15794_),
    .Y(_10117_));
 BUFx6f_ASAP7_75t_R _18431_ (.A(_10072_),
    .Y(_10118_));
 OA21x2_ASAP7_75t_R _18432_ (.A1(_10116_),
    .A2(_10117_),
    .B(_10118_),
    .Y(_10119_));
 BUFx6f_ASAP7_75t_R _18433_ (.A(_10078_),
    .Y(_10120_));
 INVx1_ASAP7_75t_R _18434_ (.A(_00482_),
    .Y(_10121_));
 NOR2x2_ASAP7_75t_R _18435_ (.A(_10121_),
    .B(_10054_),
    .Y(_10122_));
 AO21x1_ASAP7_75t_R _18436_ (.A1(_10120_),
    .A2(_10122_),
    .B(_08226_),
    .Y(_10123_));
 AOI211x1_ASAP7_75t_R _18437_ (.A1(_00395_),
    .A2(_10113_),
    .B(_10119_),
    .C(_10123_),
    .Y(_10124_));
 BUFx6f_ASAP7_75t_R _18438_ (.A(_10072_),
    .Y(_10125_));
 AOI21x1_ASAP7_75t_R _18439_ (.A1(_08183_),
    .A2(net826),
    .B(net822),
    .Y(_10126_));
 NAND2x2_ASAP7_75t_R _18440_ (.A(net822),
    .B(_08208_),
    .Y(_10127_));
 INVx6_ASAP7_75t_R _18441_ (.A(_10127_),
    .Y(_10128_));
 NOR2x1_ASAP7_75t_R _18442_ (.A(_10126_),
    .B(_10128_),
    .Y(_10129_));
 NAND2x1_ASAP7_75t_R _18443_ (.A(_10125_),
    .B(_10129_),
    .Y(_10130_));
 BUFx6f_ASAP7_75t_R _18444_ (.A(_08225_),
    .Y(_10131_));
 BUFx6f_ASAP7_75t_R _18445_ (.A(_10078_),
    .Y(_10132_));
 OAI21x1_ASAP7_75t_R _18446_ (.A1(_10128_),
    .A2(_10126_),
    .B(_10132_),
    .Y(_10133_));
 BUFx6f_ASAP7_75t_R _18447_ (.A(_08234_),
    .Y(_10134_));
 AO31x2_ASAP7_75t_R _18448_ (.A1(_10130_),
    .A2(_10131_),
    .A3(_10133_),
    .B(_10134_),
    .Y(_10135_));
 OAI21x1_ASAP7_75t_R _18449_ (.A1(_10122_),
    .A2(_10116_),
    .B(_10082_),
    .Y(_10136_));
 AND3x4_ASAP7_75t_R _18450_ (.A(_10043_),
    .B(_00481_),
    .C(_10044_),
    .Y(_10137_));
 AO21x1_ASAP7_75t_R _18451_ (.A1(_10043_),
    .A2(_10044_),
    .B(_10121_),
    .Y(_10138_));
 BUFx6f_ASAP7_75t_R _18452_ (.A(_10138_),
    .Y(_10139_));
 INVx2_ASAP7_75t_R _18453_ (.A(_10139_),
    .Y(_10140_));
 BUFx6f_ASAP7_75t_R _18454_ (.A(_10072_),
    .Y(_10141_));
 OAI21x1_ASAP7_75t_R _18455_ (.A1(_10137_),
    .A2(_10140_),
    .B(_10141_),
    .Y(_10142_));
 AOI21x1_ASAP7_75t_R _18456_ (.A1(_10136_),
    .A2(_10142_),
    .B(_10074_),
    .Y(_10143_));
 NOR2x2_ASAP7_75t_R _18457_ (.A(_10054_),
    .B(_10085_),
    .Y(_10144_));
 NOR2x1_ASAP7_75t_R _18458_ (.A(_07967_),
    .B(_08214_),
    .Y(_10145_));
 OAI21x1_ASAP7_75t_R _18459_ (.A1(_10070_),
    .A2(_10145_),
    .B(_10087_),
    .Y(_10146_));
 OAI21x1_ASAP7_75t_R _18460_ (.A1(_10125_),
    .A2(_10144_),
    .B(_10146_),
    .Y(_10147_));
 BUFx4f_ASAP7_75t_R _18461_ (.A(_10071_),
    .Y(_10148_));
 BUFx6f_ASAP7_75t_R _18462_ (.A(_10048_),
    .Y(_10149_));
 AO21x1_ASAP7_75t_R _18463_ (.A1(_10148_),
    .A2(_10041_),
    .B(_10149_),
    .Y(_10150_));
 NOR2x1_ASAP7_75t_R _18464_ (.A(_10147_),
    .B(_10150_),
    .Y(_10151_));
 OAI21x1_ASAP7_75t_R _18465_ (.A1(_10143_),
    .A2(_10151_),
    .B(_10108_),
    .Y(_10152_));
 OAI21x1_ASAP7_75t_R _18466_ (.A1(_10124_),
    .A2(_10135_),
    .B(_10152_),
    .Y(_10153_));
 INVx2_ASAP7_75t_R _18467_ (.A(_00399_),
    .Y(_10154_));
 BUFx10_ASAP7_75t_R _18468_ (.A(_10154_),
    .Y(_10155_));
 OAI21x1_ASAP7_75t_R _18469_ (.A1(_00398_),
    .A2(_10153_),
    .B(_10155_),
    .Y(_10156_));
 NOR2x2_ASAP7_75t_R _18470_ (.A(_01144_),
    .B(_10054_),
    .Y(_10157_));
 NAND2x1_ASAP7_75t_R _18471_ (.A(_10157_),
    .B(_10148_),
    .Y(_10158_));
 NAND3x1_ASAP7_75t_R _18472_ (.A(_10057_),
    .B(_10049_),
    .C(_10158_),
    .Y(_10159_));
 NOR2x2_ASAP7_75t_R _18473_ (.A(_01145_),
    .B(_15796_),
    .Y(_10160_));
 OAI21x1_ASAP7_75t_R _18474_ (.A1(_10157_),
    .A2(_10160_),
    .B(_10072_),
    .Y(_10161_));
 OAI21x1_ASAP7_75t_R _18475_ (.A1(_08215_),
    .A2(_10088_),
    .B(_10086_),
    .Y(_10162_));
 NAND3x1_ASAP7_75t_R _18476_ (.A(_10161_),
    .B(_10074_),
    .C(_10162_),
    .Y(_10163_));
 BUFx10_ASAP7_75t_R _18477_ (.A(_08235_),
    .Y(_10164_));
 AOI21x1_ASAP7_75t_R _18478_ (.A1(_10159_),
    .A2(_10163_),
    .B(_10164_),
    .Y(_10165_));
 INVx3_ASAP7_75t_R _18479_ (.A(_10137_),
    .Y(_10166_));
 AO21x1_ASAP7_75t_R _18480_ (.A1(_10166_),
    .A2(_10127_),
    .B(_10148_),
    .Y(_10167_));
 NAND2x2_ASAP7_75t_R _18481_ (.A(_10054_),
    .B(net493),
    .Y(_10168_));
 INVx2_ASAP7_75t_R _18482_ (.A(_10144_),
    .Y(_10169_));
 AO21x1_ASAP7_75t_R _18483_ (.A1(_10168_),
    .A2(_10169_),
    .B(_08217_),
    .Y(_10170_));
 AOI21x1_ASAP7_75t_R _18484_ (.A1(_10167_),
    .A2(_10170_),
    .B(_10074_),
    .Y(_10171_));
 BUFx6f_ASAP7_75t_R _18485_ (.A(_10048_),
    .Y(_10172_));
 INVx1_ASAP7_75t_R _18486_ (.A(_10122_),
    .Y(_10173_));
 NAND2x1_ASAP7_75t_R _18487_ (.A(_10045_),
    .B(_10173_),
    .Y(_10174_));
 NAND2x2_ASAP7_75t_R _18488_ (.A(_07980_),
    .B(_08214_),
    .Y(_10175_));
 INVx1_ASAP7_75t_R _18489_ (.A(_08215_),
    .Y(_10176_));
 INVx1_ASAP7_75t_R _18490_ (.A(_01144_),
    .Y(_10177_));
 NOR2x2_ASAP7_75t_R _18491_ (.A(_10177_),
    .B(_15796_),
    .Y(_10178_));
 AOI21x1_ASAP7_75t_R _18492_ (.A1(_10175_),
    .A2(_10176_),
    .B(_10178_),
    .Y(_10179_));
 AOI21x1_ASAP7_75t_R _18493_ (.A1(_10125_),
    .A2(_10174_),
    .B(_10179_),
    .Y(_10180_));
 OAI21x1_ASAP7_75t_R _18494_ (.A1(_10172_),
    .A2(_10180_),
    .B(_08235_),
    .Y(_10181_));
 NOR2x1_ASAP7_75t_R _18495_ (.A(_10171_),
    .B(_10181_),
    .Y(_10182_));
 OAI21x1_ASAP7_75t_R _18496_ (.A1(_10165_),
    .A2(_10182_),
    .B(_00398_),
    .Y(_10183_));
 INVx1_ASAP7_75t_R _18497_ (.A(_10045_),
    .Y(_10184_));
 AOI21x1_ASAP7_75t_R _18498_ (.A1(_10184_),
    .A2(_10056_),
    .B(_10149_),
    .Y(_10185_));
 AO21x2_ASAP7_75t_R _18499_ (.A1(_08207_),
    .A2(_08204_),
    .B(_10061_),
    .Y(_10186_));
 AO21x1_ASAP7_75t_R _18500_ (.A1(_10166_),
    .A2(_10186_),
    .B(_10056_),
    .Y(_10187_));
 NAND2x1_ASAP7_75t_R _18501_ (.A(_10185_),
    .B(_10187_),
    .Y(_10188_));
 AOI21x1_ASAP7_75t_R _18502_ (.A1(_10103_),
    .A2(_10102_),
    .B(_10045_),
    .Y(_10189_));
 INVx1_ASAP7_75t_R _18503_ (.A(_10189_),
    .Y(_10190_));
 NOR2x2_ASAP7_75t_R _18504_ (.A(_01145_),
    .B(_10054_),
    .Y(_10191_));
 INVx2_ASAP7_75t_R _18505_ (.A(_10191_),
    .Y(_10192_));
 NAND2x2_ASAP7_75t_R _18506_ (.A(_10186_),
    .B(_10192_),
    .Y(_10193_));
 BUFx6f_ASAP7_75t_R _18507_ (.A(_08225_),
    .Y(_10194_));
 AOI21x1_ASAP7_75t_R _18508_ (.A1(_10046_),
    .A2(_10193_),
    .B(_10194_),
    .Y(_10195_));
 BUFx6f_ASAP7_75t_R _18509_ (.A(_08234_),
    .Y(_10196_));
 AOI21x1_ASAP7_75t_R _18510_ (.A1(_10190_),
    .A2(_10195_),
    .B(_10196_),
    .Y(_10197_));
 NAND2x1_ASAP7_75t_R _18511_ (.A(_10188_),
    .B(_10197_),
    .Y(_10198_));
 NOR2x2_ASAP7_75t_R _18512_ (.A(net532),
    .B(_10054_),
    .Y(_10199_));
 OAI21x1_ASAP7_75t_R _18513_ (.A1(_08215_),
    .A2(_10088_),
    .B(_01148_),
    .Y(_10200_));
 OAI21x1_ASAP7_75t_R _18514_ (.A1(_10082_),
    .A2(_10199_),
    .B(_10200_),
    .Y(_10201_));
 AOI21x1_ASAP7_75t_R _18515_ (.A1(_10131_),
    .A2(_10201_),
    .B(_10164_),
    .Y(_10202_));
 INVx3_ASAP7_75t_R _18516_ (.A(_10186_),
    .Y(_10203_));
 OAI21x1_ASAP7_75t_R _18517_ (.A1(_10077_),
    .A2(_10203_),
    .B(_10141_),
    .Y(_10204_));
 OAI21x1_ASAP7_75t_R _18518_ (.A1(_10055_),
    .A2(_10140_),
    .B(_10046_),
    .Y(_10205_));
 NAND3x1_ASAP7_75t_R _18519_ (.A(_10204_),
    .B(_10205_),
    .C(_10172_),
    .Y(_10206_));
 AOI21x1_ASAP7_75t_R _18520_ (.A1(_10202_),
    .A2(_10206_),
    .B(_08243_),
    .Y(_10207_));
 AOI21x1_ASAP7_75t_R _18521_ (.A1(_10198_),
    .A2(_10207_),
    .B(_10155_),
    .Y(_10208_));
 NAND2x1_ASAP7_75t_R _18522_ (.A(_10183_),
    .B(_10208_),
    .Y(_10209_));
 OAI21x1_ASAP7_75t_R _18523_ (.A1(_10112_),
    .A2(_10156_),
    .B(_10209_),
    .Y(_00024_));
 NAND2x2_ASAP7_75t_R _18524_ (.A(_10042_),
    .B(_08217_),
    .Y(_10210_));
 NOR2x1_ASAP7_75t_R _18525_ (.A(_10178_),
    .B(_10210_),
    .Y(_10211_));
 BUFx6f_ASAP7_75t_R _18526_ (.A(_10071_),
    .Y(_10212_));
 NOR2x2_ASAP7_75t_R _18527_ (.A(_15794_),
    .B(net11),
    .Y(_10213_));
 INVx1_ASAP7_75t_R _18528_ (.A(_10213_),
    .Y(_10214_));
 AND3x2_ASAP7_75t_R _18529_ (.A(_10212_),
    .B(_10127_),
    .C(_10214_),
    .Y(_10215_));
 BUFx10_ASAP7_75t_R _18530_ (.A(_08234_),
    .Y(_10216_));
 OAI21x1_ASAP7_75t_R _18531_ (.A1(_10211_),
    .A2(_10215_),
    .B(_10216_),
    .Y(_10217_));
 AO21x1_ASAP7_75t_R _18532_ (.A1(_10127_),
    .A2(_10173_),
    .B(_08217_),
    .Y(_10218_));
 AO21x1_ASAP7_75t_R _18533_ (.A1(_10052_),
    .A2(_10063_),
    .B(_10148_),
    .Y(_10219_));
 NAND2x1_ASAP7_75t_R _18534_ (.A(_10218_),
    .B(_10219_),
    .Y(_10220_));
 BUFx6f_ASAP7_75t_R _18535_ (.A(_10149_),
    .Y(_10221_));
 AOI21x1_ASAP7_75t_R _18536_ (.A1(_10164_),
    .A2(_10220_),
    .B(_10221_),
    .Y(_10222_));
 AND3x1_ASAP7_75t_R _18537_ (.A(_10132_),
    .B(_08234_),
    .C(_00486_),
    .Y(_10223_));
 NAND2x2_ASAP7_75t_R _18538_ (.A(_10052_),
    .B(_10166_),
    .Y(_10224_));
 AO21x1_ASAP7_75t_R _18539_ (.A1(_10224_),
    .A2(_10141_),
    .B(_08226_),
    .Y(_10225_));
 OAI21x1_ASAP7_75t_R _18540_ (.A1(_10223_),
    .A2(_10225_),
    .B(_10110_),
    .Y(_10226_));
 AOI21x1_ASAP7_75t_R _18541_ (.A1(_10217_),
    .A2(_10222_),
    .B(_10226_),
    .Y(_10227_));
 OAI21x1_ASAP7_75t_R _18542_ (.A1(_10053_),
    .A2(_10055_),
    .B(_10125_),
    .Y(_10228_));
 AOI21x1_ASAP7_75t_R _18543_ (.A1(_10162_),
    .A2(_10228_),
    .B(_10074_),
    .Y(_10229_));
 NOR2x2_ASAP7_75t_R _18544_ (.A(net500),
    .B(_15794_),
    .Y(_10230_));
 NOR2x2_ASAP7_75t_R _18545_ (.A(_10230_),
    .B(_10115_),
    .Y(_10231_));
 NAND2x2_ASAP7_75t_R _18546_ (.A(_08217_),
    .B(_10231_),
    .Y(_10232_));
 NOR2x2_ASAP7_75t_R _18547_ (.A(_01146_),
    .B(_15794_),
    .Y(_10233_));
 OAI21x1_ASAP7_75t_R _18548_ (.A1(_10066_),
    .A2(_10233_),
    .B(_10125_),
    .Y(_10234_));
 AOI21x1_ASAP7_75t_R _18549_ (.A1(_10232_),
    .A2(_10234_),
    .B(_10172_),
    .Y(_10235_));
 OAI21x1_ASAP7_75t_R _18550_ (.A1(_10229_),
    .A2(_10235_),
    .B(_10216_),
    .Y(_10236_));
 OAI21x1_ASAP7_75t_R _18551_ (.A1(_10122_),
    .A2(_10094_),
    .B(_10212_),
    .Y(_10237_));
 AOI21x1_ASAP7_75t_R _18552_ (.A1(_10042_),
    .A2(_10179_),
    .B(_10194_),
    .Y(_10238_));
 NAND2x1_ASAP7_75t_R _18553_ (.A(_10237_),
    .B(_10238_),
    .Y(_10239_));
 INVx2_ASAP7_75t_R _18554_ (.A(_10199_),
    .Y(_10240_));
 NAND2x1_ASAP7_75t_R _18555_ (.A(_10139_),
    .B(_10240_),
    .Y(_10241_));
 AOI21x1_ASAP7_75t_R _18556_ (.A1(_10132_),
    .A2(_10241_),
    .B(_10189_),
    .Y(_10242_));
 INVx1_ASAP7_75t_R _18557_ (.A(_10055_),
    .Y(_10243_));
 OA21x2_ASAP7_75t_R _18558_ (.A1(_10078_),
    .A2(_10243_),
    .B(_08225_),
    .Y(_10244_));
 AOI21x1_ASAP7_75t_R _18559_ (.A1(_10242_),
    .A2(_10244_),
    .B(_10196_),
    .Y(_10245_));
 NAND2x1_ASAP7_75t_R _18560_ (.A(_10239_),
    .B(_10245_),
    .Y(_10246_));
 AOI21x1_ASAP7_75t_R _18561_ (.A1(_10236_),
    .A2(_10246_),
    .B(_10111_),
    .Y(_10247_));
 OAI21x1_ASAP7_75t_R _18562_ (.A1(_10227_),
    .A2(_10247_),
    .B(_10155_),
    .Y(_10248_));
 AO21x1_ASAP7_75t_R _18563_ (.A1(_10102_),
    .A2(_10103_),
    .B(_10080_),
    .Y(_10249_));
 NAND3x1_ASAP7_75t_R _18564_ (.A(_10232_),
    .B(_10249_),
    .C(_10049_),
    .Y(_10250_));
 BUFx6f_ASAP7_75t_R _18565_ (.A(_08225_),
    .Y(_10251_));
 INVx1_ASAP7_75t_R _18566_ (.A(_10092_),
    .Y(_10252_));
 AOI21x1_ASAP7_75t_R _18567_ (.A1(_10103_),
    .A2(_10102_),
    .B(_10052_),
    .Y(_10253_));
 AOI21x1_ASAP7_75t_R _18568_ (.A1(_10168_),
    .A2(_10252_),
    .B(_10253_),
    .Y(_10254_));
 NAND2x1_ASAP7_75t_R _18569_ (.A(_10251_),
    .B(_10254_),
    .Y(_10255_));
 AOI21x1_ASAP7_75t_R _18570_ (.A1(_10250_),
    .A2(_10255_),
    .B(_10216_),
    .Y(_10256_));
 NOR2x2_ASAP7_75t_R _18571_ (.A(_15786_),
    .B(net11),
    .Y(_10257_));
 OAI21x1_ASAP7_75t_R _18572_ (.A1(_10094_),
    .A2(_10257_),
    .B(_10046_),
    .Y(_10258_));
 AO21x1_ASAP7_75t_R _18573_ (.A1(_10169_),
    .A2(_10127_),
    .B(_08217_),
    .Y(_10259_));
 AOI21x1_ASAP7_75t_R _18574_ (.A1(_10258_),
    .A2(_10259_),
    .B(_10251_),
    .Y(_10260_));
 OAI21x1_ASAP7_75t_R _18575_ (.A1(_10157_),
    .A2(_10162_),
    .B(_10194_),
    .Y(_10261_));
 AND3x1_ASAP7_75t_R _18576_ (.A(_10072_),
    .B(_10243_),
    .C(_10139_),
    .Y(_10262_));
 OAI21x1_ASAP7_75t_R _18577_ (.A1(_10261_),
    .A2(_10262_),
    .B(_08234_),
    .Y(_10263_));
 NOR2x1_ASAP7_75t_R _18578_ (.A(_10260_),
    .B(_10263_),
    .Y(_10264_));
 OAI21x1_ASAP7_75t_R _18579_ (.A1(_10256_),
    .A2(_10264_),
    .B(_08243_),
    .Y(_10265_));
 BUFx6f_ASAP7_75t_R _18580_ (.A(_10071_),
    .Y(_10266_));
 OAI21x1_ASAP7_75t_R _18581_ (.A1(_10077_),
    .A2(_10081_),
    .B(_10266_),
    .Y(_10267_));
 NOR2x2_ASAP7_75t_R _18582_ (.A(_10077_),
    .B(_10087_),
    .Y(_10268_));
 AOI21x1_ASAP7_75t_R _18583_ (.A1(_10046_),
    .A2(_10268_),
    .B(_10149_),
    .Y(_10269_));
 NAND2x1_ASAP7_75t_R _18584_ (.A(_10267_),
    .B(_10269_),
    .Y(_10270_));
 NOR2x1_ASAP7_75t_R _18585_ (.A(_15786_),
    .B(net18),
    .Y(_10271_));
 OAI21x1_ASAP7_75t_R _18586_ (.A1(_10213_),
    .A2(_10271_),
    .B(_10212_),
    .Y(_10272_));
 OA21x2_ASAP7_75t_R _18587_ (.A1(_10072_),
    .A2(_10063_),
    .B(_10048_),
    .Y(_10273_));
 AOI21x1_ASAP7_75t_R _18588_ (.A1(_10272_),
    .A2(_10273_),
    .B(_10196_),
    .Y(_10274_));
 AOI21x1_ASAP7_75t_R _18589_ (.A1(_10270_),
    .A2(_10274_),
    .B(_08243_),
    .Y(_10275_));
 NOR2x1_ASAP7_75t_R _18590_ (.A(_10157_),
    .B(_10203_),
    .Y(_10276_));
 INVx1_ASAP7_75t_R _18591_ (.A(_10276_),
    .Y(_10277_));
 NAND2x2_ASAP7_75t_R _18592_ (.A(_10072_),
    .B(_10277_),
    .Y(_10278_));
 AOI22x1_ASAP7_75t_R _18593_ (.A1(_10240_),
    .A2(_10065_),
    .B1(_10175_),
    .B2(_10176_),
    .Y(_10279_));
 NOR2x1_ASAP7_75t_R _18594_ (.A(_10194_),
    .B(_10279_),
    .Y(_10280_));
 AOI21x1_ASAP7_75t_R _18595_ (.A1(_10278_),
    .A2(_10280_),
    .B(_08235_),
    .Y(_10281_));
 INVx1_ASAP7_75t_R _18596_ (.A(_10157_),
    .Y(_10282_));
 OA21x2_ASAP7_75t_R _18597_ (.A1(_10078_),
    .A2(_10282_),
    .B(_08225_),
    .Y(_10283_));
 NAND2x2_ASAP7_75t_R _18598_ (.A(_00487_),
    .B(_10078_),
    .Y(_10284_));
 OA21x2_ASAP7_75t_R _18599_ (.A1(_08217_),
    .A2(_10168_),
    .B(_10284_),
    .Y(_10285_));
 NAND2x1_ASAP7_75t_R _18600_ (.A(_10283_),
    .B(_10285_),
    .Y(_10286_));
 NAND2x1_ASAP7_75t_R _18601_ (.A(_10281_),
    .B(_10286_),
    .Y(_10287_));
 AOI21x1_ASAP7_75t_R _18602_ (.A1(_10275_),
    .A2(_10287_),
    .B(_10154_),
    .Y(_10288_));
 NAND2x1_ASAP7_75t_R _18603_ (.A(_10265_),
    .B(_10288_),
    .Y(_10289_));
 NAND2x1_ASAP7_75t_R _18604_ (.A(_10248_),
    .B(_10289_),
    .Y(_00025_));
 OAI21x1_ASAP7_75t_R _18605_ (.A1(_10128_),
    .A2(_10191_),
    .B(_10212_),
    .Y(_10290_));
 OAI21x1_ASAP7_75t_R _18606_ (.A1(_10144_),
    .A2(_10116_),
    .B(_10132_),
    .Y(_10291_));
 AOI21x1_ASAP7_75t_R _18607_ (.A1(_10290_),
    .A2(_10291_),
    .B(_10251_),
    .Y(_10292_));
 OAI21x1_ASAP7_75t_R _18608_ (.A1(_10160_),
    .A2(_10041_),
    .B(_10132_),
    .Y(_10293_));
 NOR2x2_ASAP7_75t_R _18609_ (.A(_01143_),
    .B(_10054_),
    .Y(_10294_));
 INVx1_ASAP7_75t_R _18610_ (.A(_10294_),
    .Y(_10295_));
 NAND2x1_ASAP7_75t_R _18611_ (.A(_10127_),
    .B(_10295_),
    .Y(_10296_));
 NAND2x1_ASAP7_75t_R _18612_ (.A(_10212_),
    .B(_10296_),
    .Y(_10297_));
 AOI21x1_ASAP7_75t_R _18613_ (.A1(_10293_),
    .A2(_10297_),
    .B(_10049_),
    .Y(_10298_));
 OAI21x1_ASAP7_75t_R _18614_ (.A1(_10292_),
    .A2(_10298_),
    .B(_10164_),
    .Y(_10299_));
 OAI21x1_ASAP7_75t_R _18615_ (.A1(_10157_),
    .A2(_10128_),
    .B(_10132_),
    .Y(_10300_));
 OAI21x1_ASAP7_75t_R _18616_ (.A1(_10160_),
    .A2(_10294_),
    .B(_10125_),
    .Y(_10301_));
 AOI21x1_ASAP7_75t_R _18617_ (.A1(_10300_),
    .A2(_10301_),
    .B(_10172_),
    .Y(_10302_));
 OAI21x1_ASAP7_75t_R _18618_ (.A1(_10157_),
    .A2(_10059_),
    .B(_10120_),
    .Y(_10303_));
 AOI21x1_ASAP7_75t_R _18619_ (.A1(_10161_),
    .A2(_10303_),
    .B(_10074_),
    .Y(_10304_));
 OAI21x1_ASAP7_75t_R _18620_ (.A1(_10302_),
    .A2(_10304_),
    .B(_10216_),
    .Y(_10305_));
 AOI21x1_ASAP7_75t_R _18621_ (.A1(_10299_),
    .A2(_10305_),
    .B(_10111_),
    .Y(_10306_));
 NOR2x1_ASAP7_75t_R _18622_ (.A(_10116_),
    .B(_10041_),
    .Y(_10307_));
 OAI21x1_ASAP7_75t_R _18623_ (.A1(_10128_),
    .A2(_10233_),
    .B(_10120_),
    .Y(_10308_));
 OAI21x1_ASAP7_75t_R _18624_ (.A1(_00395_),
    .A2(_10307_),
    .B(_10308_),
    .Y(_10309_));
 OAI21x1_ASAP7_75t_R _18625_ (.A1(_10117_),
    .A2(_10066_),
    .B(_10120_),
    .Y(_10310_));
 INVx2_ASAP7_75t_R _18626_ (.A(_10104_),
    .Y(_10311_));
 AOI21x1_ASAP7_75t_R _18627_ (.A1(_10311_),
    .A2(_10148_),
    .B(_10194_),
    .Y(_10312_));
 AOI21x1_ASAP7_75t_R _18628_ (.A1(_10310_),
    .A2(_10312_),
    .B(_10196_),
    .Y(_10313_));
 OAI21x1_ASAP7_75t_R _18629_ (.A1(_10050_),
    .A2(_10309_),
    .B(_10313_),
    .Y(_10314_));
 OAI21x1_ASAP7_75t_R _18630_ (.A1(_10294_),
    .A2(_10081_),
    .B(_10212_),
    .Y(_10315_));
 CKINVDCx5p33_ASAP7_75t_R _18631_ (.A(_10168_),
    .Y(_10316_));
 OAI21x1_ASAP7_75t_R _18632_ (.A1(_10062_),
    .A2(_10316_),
    .B(_10056_),
    .Y(_10317_));
 AOI21x1_ASAP7_75t_R _18633_ (.A1(_10315_),
    .A2(_10317_),
    .B(_10172_),
    .Y(_10318_));
 OA21x2_ASAP7_75t_R _18634_ (.A1(_10316_),
    .A2(_10144_),
    .B(_10072_),
    .Y(_10319_));
 AOI21x1_ASAP7_75t_R _18635_ (.A1(_10078_),
    .A2(_10276_),
    .B(_08225_),
    .Y(_10320_));
 INVx1_ASAP7_75t_R _18636_ (.A(_10320_),
    .Y(_10321_));
 NOR2x1_ASAP7_75t_R _18637_ (.A(_10319_),
    .B(_10321_),
    .Y(_10322_));
 OAI21x1_ASAP7_75t_R _18638_ (.A1(_10318_),
    .A2(_10322_),
    .B(_10216_),
    .Y(_10323_));
 AOI21x1_ASAP7_75t_R _18639_ (.A1(_10314_),
    .A2(_10323_),
    .B(_00398_),
    .Y(_10324_));
 OAI21x1_ASAP7_75t_R _18640_ (.A1(_10306_),
    .A2(_10324_),
    .B(_10155_),
    .Y(_10325_));
 NAND2x1_ASAP7_75t_R _18641_ (.A(_10127_),
    .B(_10056_),
    .Y(_10326_));
 NAND2x1_ASAP7_75t_R _18642_ (.A(_10148_),
    .B(_10224_),
    .Y(_10327_));
 OAI21x1_ASAP7_75t_R _18643_ (.A1(_10326_),
    .A2(_10230_),
    .B(_10327_),
    .Y(_10328_));
 OAI21x1_ASAP7_75t_R _18644_ (.A1(_10157_),
    .A2(_10116_),
    .B(_10120_),
    .Y(_10329_));
 AOI21x1_ASAP7_75t_R _18645_ (.A1(_10140_),
    .A2(_10266_),
    .B(_08226_),
    .Y(_10330_));
 AOI21x1_ASAP7_75t_R _18646_ (.A1(_10329_),
    .A2(_10330_),
    .B(_10196_),
    .Y(_10331_));
 OAI21x1_ASAP7_75t_R _18647_ (.A1(_10221_),
    .A2(_10328_),
    .B(_10331_),
    .Y(_10332_));
 INVx1_ASAP7_75t_R _18648_ (.A(_01149_),
    .Y(_10333_));
 AOI21x1_ASAP7_75t_R _18649_ (.A1(_10333_),
    .A2(_10212_),
    .B(_10149_),
    .Y(_10334_));
 NAND2x1_ASAP7_75t_R _18650_ (.A(_10317_),
    .B(_10334_),
    .Y(_10335_));
 NAND2x1_ASAP7_75t_R _18651_ (.A(_00488_),
    .B(_10056_),
    .Y(_10336_));
 NAND2x1_ASAP7_75t_R _18652_ (.A(_10336_),
    .B(_10312_),
    .Y(_10337_));
 NAND3x1_ASAP7_75t_R _18653_ (.A(_10335_),
    .B(_10337_),
    .C(_10134_),
    .Y(_10338_));
 AOI21x1_ASAP7_75t_R _18654_ (.A1(_10332_),
    .A2(_10338_),
    .B(_08243_),
    .Y(_10339_));
 NOR2x2_ASAP7_75t_R _18655_ (.A(_10094_),
    .B(_10210_),
    .Y(_10340_));
 NAND2x1_ASAP7_75t_R _18656_ (.A(_10251_),
    .B(_10170_),
    .Y(_10341_));
 OAI21x1_ASAP7_75t_R _18657_ (.A1(_10199_),
    .A2(_10203_),
    .B(_10120_),
    .Y(_10342_));
 AOI21x1_ASAP7_75t_R _18658_ (.A1(_10103_),
    .A2(_10102_),
    .B(_01148_),
    .Y(_10343_));
 NOR2x1_ASAP7_75t_R _18659_ (.A(_10194_),
    .B(_10343_),
    .Y(_10344_));
 AOI21x1_ASAP7_75t_R _18660_ (.A1(_10342_),
    .A2(_10344_),
    .B(_10196_),
    .Y(_10345_));
 OAI21x1_ASAP7_75t_R _18661_ (.A1(_10340_),
    .A2(_10341_),
    .B(_10345_),
    .Y(_10346_));
 NAND2x1_ASAP7_75t_R _18662_ (.A(_00486_),
    .B(_10266_),
    .Y(_10347_));
 OAI21x1_ASAP7_75t_R _18663_ (.A1(_10213_),
    .A2(_10271_),
    .B(_10132_),
    .Y(_10348_));
 AOI21x1_ASAP7_75t_R _18664_ (.A1(_10347_),
    .A2(_10348_),
    .B(_10074_),
    .Y(_10349_));
 BUFx6f_ASAP7_75t_R _18665_ (.A(_10078_),
    .Y(_10350_));
 OAI21x1_ASAP7_75t_R _18666_ (.A1(_10199_),
    .A2(_10113_),
    .B(_10350_),
    .Y(_10351_));
 AO21x1_ASAP7_75t_R _18667_ (.A1(_10060_),
    .A2(_10173_),
    .B(_10056_),
    .Y(_10352_));
 AOI21x1_ASAP7_75t_R _18668_ (.A1(_10351_),
    .A2(_10352_),
    .B(_10172_),
    .Y(_10353_));
 OAI21x1_ASAP7_75t_R _18669_ (.A1(_10349_),
    .A2(_10353_),
    .B(_10216_),
    .Y(_10354_));
 AOI21x1_ASAP7_75t_R _18670_ (.A1(_10346_),
    .A2(_10354_),
    .B(_10111_),
    .Y(_10355_));
 OAI21x1_ASAP7_75t_R _18671_ (.A1(_10339_),
    .A2(_10355_),
    .B(_00399_),
    .Y(_10356_));
 NAND2x1_ASAP7_75t_R _18672_ (.A(_10325_),
    .B(_10356_),
    .Y(_00026_));
 BUFx6f_ASAP7_75t_R _18673_ (.A(_10078_),
    .Y(_10357_));
 NOR2x1_ASAP7_75t_R _18674_ (.A(_10126_),
    .B(_10055_),
    .Y(_10358_));
 OAI21x1_ASAP7_75t_R _18675_ (.A1(_10357_),
    .A2(_10358_),
    .B(_10049_),
    .Y(_10359_));
 AOI21x1_ASAP7_75t_R _18676_ (.A1(_00395_),
    .A2(_10311_),
    .B(_10359_),
    .Y(_10360_));
 OA21x2_ASAP7_75t_R _18677_ (.A1(_10087_),
    .A2(_10191_),
    .B(_10073_),
    .Y(_10361_));
 OAI21x1_ASAP7_75t_R _18678_ (.A1(_10316_),
    .A2(_10092_),
    .B(_10131_),
    .Y(_10362_));
 OAI21x1_ASAP7_75t_R _18679_ (.A1(_10361_),
    .A2(_10362_),
    .B(_10108_),
    .Y(_10363_));
 OAI21x1_ASAP7_75t_R _18680_ (.A1(_10360_),
    .A2(_10363_),
    .B(_00398_),
    .Y(_10364_));
 NOR2x1_ASAP7_75t_R _18681_ (.A(_10087_),
    .B(_10137_),
    .Y(_10365_));
 NOR2x1_ASAP7_75t_R _18682_ (.A(_10357_),
    .B(_10365_),
    .Y(_10366_));
 AND2x2_ASAP7_75t_R _18683_ (.A(_10129_),
    .B(_10350_),
    .Y(_10367_));
 OAI21x1_ASAP7_75t_R _18684_ (.A1(_10366_),
    .A2(_10367_),
    .B(_00396_),
    .Y(_10368_));
 OA21x2_ASAP7_75t_R _18685_ (.A1(_10053_),
    .A2(_10199_),
    .B(_10118_),
    .Y(_10369_));
 OA21x2_ASAP7_75t_R _18686_ (.A1(_10113_),
    .A2(_10062_),
    .B(_10357_),
    .Y(_10370_));
 OAI21x1_ASAP7_75t_R _18687_ (.A1(_10369_),
    .A2(_10370_),
    .B(_10050_),
    .Y(_10371_));
 AOI21x1_ASAP7_75t_R _18688_ (.A1(_10368_),
    .A2(_10371_),
    .B(_10108_),
    .Y(_10372_));
 INVx1_ASAP7_75t_R _18689_ (.A(_10162_),
    .Y(_10373_));
 AOI21x1_ASAP7_75t_R _18690_ (.A1(_10373_),
    .A2(_10042_),
    .B(_10359_),
    .Y(_10374_));
 OA21x2_ASAP7_75t_R _18691_ (.A1(_10128_),
    .A2(_10213_),
    .B(_10118_),
    .Y(_10375_));
 AO21x1_ASAP7_75t_R _18692_ (.A1(_10357_),
    .A2(_10169_),
    .B(_10049_),
    .Y(_10376_));
 OAI21x1_ASAP7_75t_R _18693_ (.A1(_10375_),
    .A2(_10376_),
    .B(_10108_),
    .Y(_10377_));
 OAI21x1_ASAP7_75t_R _18694_ (.A1(_10374_),
    .A2(_10377_),
    .B(_10111_),
    .Y(_10378_));
 NAND3x1_ASAP7_75t_R _18695_ (.A(_10357_),
    .B(_10169_),
    .C(_10139_),
    .Y(_10379_));
 AO211x2_ASAP7_75t_R _18696_ (.A1(_10103_),
    .A2(_10102_),
    .B(_10055_),
    .C(_10113_),
    .Y(_10380_));
 AOI21x1_ASAP7_75t_R _18697_ (.A1(_10379_),
    .A2(_10380_),
    .B(_10221_),
    .Y(_10381_));
 NAND2x1_ASAP7_75t_R _18698_ (.A(_10065_),
    .B(_10282_),
    .Y(_10382_));
 AOI21x1_ASAP7_75t_R _18699_ (.A1(_10082_),
    .A2(_10382_),
    .B(_10251_),
    .Y(_10383_));
 NAND2x1_ASAP7_75t_R _18700_ (.A(_10141_),
    .B(_10307_),
    .Y(_10384_));
 AO21x1_ASAP7_75t_R _18701_ (.A1(_10383_),
    .A2(_10384_),
    .B(_10134_),
    .Y(_10385_));
 NOR2x1_ASAP7_75t_R _18702_ (.A(_10381_),
    .B(_10385_),
    .Y(_10386_));
 OAI22x1_ASAP7_75t_R _18703_ (.A1(_10364_),
    .A2(_10372_),
    .B1(_10378_),
    .B2(_10386_),
    .Y(_10387_));
 NAND2x1_ASAP7_75t_R _18704_ (.A(_10144_),
    .B(_10132_),
    .Y(_10388_));
 OAI21x1_ASAP7_75t_R _18705_ (.A1(_10137_),
    .A2(_10316_),
    .B(_10141_),
    .Y(_10389_));
 AOI21x1_ASAP7_75t_R _18706_ (.A1(_10388_),
    .A2(_10389_),
    .B(_08235_),
    .Y(_10390_));
 OAI21x1_ASAP7_75t_R _18707_ (.A1(_10196_),
    .A2(_10146_),
    .B(_10185_),
    .Y(_10391_));
 OAI21x1_ASAP7_75t_R _18708_ (.A1(_10390_),
    .A2(_10391_),
    .B(_10110_),
    .Y(_10392_));
 AOI21x1_ASAP7_75t_R _18709_ (.A1(_10160_),
    .A2(_10120_),
    .B(_08234_),
    .Y(_10393_));
 NAND2x1_ASAP7_75t_R _18710_ (.A(_10290_),
    .B(_10393_),
    .Y(_10394_));
 AOI21x1_ASAP7_75t_R _18711_ (.A1(_10141_),
    .A2(_10268_),
    .B(_08235_),
    .Y(_10395_));
 OAI21x1_ASAP7_75t_R _18712_ (.A1(_10326_),
    .A2(_10090_),
    .B(_10395_),
    .Y(_10396_));
 AOI21x1_ASAP7_75t_R _18713_ (.A1(_10394_),
    .A2(_10396_),
    .B(_00396_),
    .Y(_10397_));
 NOR2x1_ASAP7_75t_R _18714_ (.A(_10392_),
    .B(_10397_),
    .Y(_10398_));
 NAND2x1_ASAP7_75t_R _18715_ (.A(_10205_),
    .B(_10272_),
    .Y(_10399_));
 OAI21x1_ASAP7_75t_R _18716_ (.A1(_10116_),
    .A2(_10294_),
    .B(_10118_),
    .Y(_10400_));
 OAI21x1_ASAP7_75t_R _18717_ (.A1(_10077_),
    .A2(_10160_),
    .B(_10056_),
    .Y(_10401_));
 AOI21x1_ASAP7_75t_R _18718_ (.A1(_10400_),
    .A2(_10401_),
    .B(_10221_),
    .Y(_10402_));
 AOI21x1_ASAP7_75t_R _18719_ (.A1(_10050_),
    .A2(_10399_),
    .B(_10402_),
    .Y(_10403_));
 OAI21x1_ASAP7_75t_R _18720_ (.A1(_10350_),
    .A2(_10296_),
    .B(_08226_),
    .Y(_10404_));
 NAND2x1_ASAP7_75t_R _18721_ (.A(_10196_),
    .B(_10404_),
    .Y(_10405_));
 OAI21x1_ASAP7_75t_R _18722_ (.A1(_10191_),
    .A2(_10094_),
    .B(_10082_),
    .Y(_10406_));
 AOI21x1_ASAP7_75t_R _18723_ (.A1(_10406_),
    .A2(_10327_),
    .B(_10131_),
    .Y(_10407_));
 OAI21x1_ASAP7_75t_R _18724_ (.A1(_10405_),
    .A2(_10407_),
    .B(_08243_),
    .Y(_10408_));
 AOI21x1_ASAP7_75t_R _18725_ (.A1(_00397_),
    .A2(_10403_),
    .B(_10408_),
    .Y(_10409_));
 OAI21x1_ASAP7_75t_R _18726_ (.A1(_10398_),
    .A2(_10409_),
    .B(_10155_),
    .Y(_10410_));
 OAI21x1_ASAP7_75t_R _18727_ (.A1(_10155_),
    .A2(_10387_),
    .B(_10410_),
    .Y(_00027_));
 OA21x2_ASAP7_75t_R _18728_ (.A1(_10059_),
    .A2(_10122_),
    .B(_10357_),
    .Y(_10411_));
 NOR3x1_ASAP7_75t_R _18729_ (.A(_00395_),
    .B(_10316_),
    .C(_10257_),
    .Y(_10412_));
 OAI21x1_ASAP7_75t_R _18730_ (.A1(_10411_),
    .A2(_10412_),
    .B(_00396_),
    .Y(_10413_));
 INVx1_ASAP7_75t_R _18731_ (.A(_10348_),
    .Y(_10414_));
 OAI21x1_ASAP7_75t_R _18732_ (.A1(_10414_),
    .A2(_10215_),
    .B(_10050_),
    .Y(_10415_));
 AOI21x1_ASAP7_75t_R _18733_ (.A1(_10413_),
    .A2(_10415_),
    .B(_00397_),
    .Y(_10416_));
 NAND2x1_ASAP7_75t_R _18734_ (.A(_01145_),
    .B(_15796_),
    .Y(_10417_));
 OAI21x1_ASAP7_75t_R _18735_ (.A1(_08215_),
    .A2(_10088_),
    .B(_10417_),
    .Y(_10418_));
 AND2x2_ASAP7_75t_R _18736_ (.A(_10418_),
    .B(_10045_),
    .Y(_10419_));
 AO21x1_ASAP7_75t_R _18737_ (.A1(_10419_),
    .A2(_10131_),
    .B(_10134_),
    .Y(_10420_));
 OAI21x1_ASAP7_75t_R _18738_ (.A1(_10128_),
    .A2(_10041_),
    .B(_10046_),
    .Y(_10421_));
 AND3x1_ASAP7_75t_R _18739_ (.A(_10218_),
    .B(_10172_),
    .C(_10421_),
    .Y(_10422_));
 OAI21x1_ASAP7_75t_R _18740_ (.A1(_10420_),
    .A2(_10422_),
    .B(_00399_),
    .Y(_10423_));
 OAI21x1_ASAP7_75t_R _18741_ (.A1(_10416_),
    .A2(_10423_),
    .B(_00398_),
    .Y(_10424_));
 NOR2x1_ASAP7_75t_R _18742_ (.A(_10139_),
    .B(_10357_),
    .Y(_10425_));
 OR3x1_ASAP7_75t_R _18743_ (.A(_10211_),
    .B(_10425_),
    .C(_10150_),
    .Y(_10426_));
 AND3x1_ASAP7_75t_R _18744_ (.A(_10073_),
    .B(_10127_),
    .C(_10091_),
    .Y(_10427_));
 AO21x1_ASAP7_75t_R _18745_ (.A1(_00395_),
    .A2(_15796_),
    .B(_10074_),
    .Y(_10428_));
 OA21x2_ASAP7_75t_R _18746_ (.A1(_10427_),
    .A2(_10428_),
    .B(_10108_),
    .Y(_10429_));
 AND3x1_ASAP7_75t_R _18747_ (.A(_10043_),
    .B(_01146_),
    .C(_10044_),
    .Y(_10430_));
 AO21x2_ASAP7_75t_R _18748_ (.A1(_10102_),
    .A2(_10103_),
    .B(_10430_),
    .Y(_10431_));
 OAI21x1_ASAP7_75t_R _18749_ (.A1(_10073_),
    .A2(_10230_),
    .B(_10431_),
    .Y(_10432_));
 OAI21x1_ASAP7_75t_R _18750_ (.A1(_10050_),
    .A2(_10432_),
    .B(_00397_),
    .Y(_10433_));
 AO21x1_ASAP7_75t_R _18751_ (.A1(_10169_),
    .A2(_10080_),
    .B(_10046_),
    .Y(_10434_));
 AND3x1_ASAP7_75t_R _18752_ (.A(_10434_),
    .B(_10172_),
    .C(_10057_),
    .Y(_10435_));
 OAI21x1_ASAP7_75t_R _18753_ (.A1(_10433_),
    .A2(_10435_),
    .B(_10155_),
    .Y(_10436_));
 AOI21x1_ASAP7_75t_R _18754_ (.A1(_10426_),
    .A2(_10429_),
    .B(_10436_),
    .Y(_10437_));
 AO21x1_ASAP7_75t_R _18755_ (.A1(_10240_),
    .A2(_10065_),
    .B(_10056_),
    .Y(_10438_));
 AOI21x1_ASAP7_75t_R _18756_ (.A1(_10195_),
    .A2(_10438_),
    .B(_10196_),
    .Y(_10439_));
 AOI21x1_ASAP7_75t_R _18757_ (.A1(_10160_),
    .A2(_10132_),
    .B(_10149_),
    .Y(_10440_));
 NAND2x2_ASAP7_75t_R _18758_ (.A(_10199_),
    .B(_08217_),
    .Y(_10441_));
 NAND3x1_ASAP7_75t_R _18759_ (.A(_10440_),
    .B(_10161_),
    .C(_10441_),
    .Y(_10442_));
 AOI21x1_ASAP7_75t_R _18760_ (.A1(_10439_),
    .A2(_10442_),
    .B(_10154_),
    .Y(_10443_));
 AO21x1_ASAP7_75t_R _18761_ (.A1(_10214_),
    .A2(_10139_),
    .B(_10148_),
    .Y(_10444_));
 AOI21x1_ASAP7_75t_R _18762_ (.A1(_10278_),
    .A2(_10444_),
    .B(_10074_),
    .Y(_10445_));
 AO21x1_ASAP7_75t_R _18763_ (.A1(_10214_),
    .A2(_10186_),
    .B(_10148_),
    .Y(_10446_));
 AOI21x1_ASAP7_75t_R _18764_ (.A1(_10315_),
    .A2(_10446_),
    .B(_10172_),
    .Y(_10447_));
 OAI21x1_ASAP7_75t_R _18765_ (.A1(_10445_),
    .A2(_10447_),
    .B(_10216_),
    .Y(_10448_));
 NAND2x1_ASAP7_75t_R _18766_ (.A(_10443_),
    .B(_10448_),
    .Y(_10449_));
 AOI21x1_ASAP7_75t_R _18767_ (.A1(_10125_),
    .A2(_10174_),
    .B(_08226_),
    .Y(_10450_));
 AOI21x1_ASAP7_75t_R _18768_ (.A1(_10133_),
    .A2(_10450_),
    .B(_08235_),
    .Y(_10451_));
 OAI21x1_ASAP7_75t_R _18769_ (.A1(_10257_),
    .A2(_10316_),
    .B(_10266_),
    .Y(_10452_));
 OA21x2_ASAP7_75t_R _18770_ (.A1(_10418_),
    .A2(_10128_),
    .B(_10194_),
    .Y(_10453_));
 NAND2x1_ASAP7_75t_R _18771_ (.A(_10452_),
    .B(_10453_),
    .Y(_10454_));
 NAND2x1_ASAP7_75t_R _18772_ (.A(_10451_),
    .B(_10454_),
    .Y(_10455_));
 AO21x1_ASAP7_75t_R _18773_ (.A1(_10060_),
    .A2(_10192_),
    .B(_10148_),
    .Y(_10456_));
 OA21x2_ASAP7_75t_R _18774_ (.A1(_08217_),
    .A2(_10186_),
    .B(_10194_),
    .Y(_10457_));
 NAND2x1_ASAP7_75t_R _18775_ (.A(_10456_),
    .B(_10457_),
    .Y(_10458_));
 AOI21x1_ASAP7_75t_R _18776_ (.A1(_10103_),
    .A2(_10102_),
    .B(_10051_),
    .Y(_10459_));
 AOI21x1_ASAP7_75t_R _18777_ (.A1(_10082_),
    .A2(_10240_),
    .B(_10459_),
    .Y(_10460_));
 AOI21x1_ASAP7_75t_R _18778_ (.A1(_10221_),
    .A2(_10460_),
    .B(_10134_),
    .Y(_10461_));
 AOI21x1_ASAP7_75t_R _18779_ (.A1(_10458_),
    .A2(_10461_),
    .B(_00399_),
    .Y(_10462_));
 AOI21x1_ASAP7_75t_R _18780_ (.A1(_10455_),
    .A2(_10462_),
    .B(_00398_),
    .Y(_10463_));
 NAND2x1_ASAP7_75t_R _18781_ (.A(_10449_),
    .B(_10463_),
    .Y(_10464_));
 OAI21x1_ASAP7_75t_R _18782_ (.A1(_10424_),
    .A2(_10437_),
    .B(_10464_),
    .Y(_00028_));
 OA21x2_ASAP7_75t_R _18783_ (.A1(_10266_),
    .A2(net18),
    .B(_10049_),
    .Y(_10465_));
 NAND2x1_ASAP7_75t_R _18784_ (.A(_10452_),
    .B(_10465_),
    .Y(_10466_));
 INVx1_ASAP7_75t_R _18785_ (.A(_10079_),
    .Y(_10467_));
 OA21x2_ASAP7_75t_R _18786_ (.A1(_10224_),
    .A2(_10141_),
    .B(_10251_),
    .Y(_10468_));
 OAI21x1_ASAP7_75t_R _18787_ (.A1(_10467_),
    .A2(_10257_),
    .B(_10468_),
    .Y(_10469_));
 AOI21x1_ASAP7_75t_R _18788_ (.A1(_10466_),
    .A2(_10469_),
    .B(_10108_),
    .Y(_10470_));
 OA21x2_ASAP7_75t_R _18789_ (.A1(_10350_),
    .A2(_10294_),
    .B(_10162_),
    .Y(_10471_));
 OAI21x1_ASAP7_75t_R _18790_ (.A1(_10123_),
    .A2(_10471_),
    .B(_10216_),
    .Y(_10472_));
 OA211x2_ASAP7_75t_R _18791_ (.A1(_10059_),
    .A2(_10431_),
    .B(_10441_),
    .C(_10251_),
    .Y(_10473_));
 OAI21x1_ASAP7_75t_R _18792_ (.A1(_10472_),
    .A2(_10473_),
    .B(_10111_),
    .Y(_10474_));
 NOR2x1_ASAP7_75t_R _18793_ (.A(_10470_),
    .B(_10474_),
    .Y(_10475_));
 AO21x1_ASAP7_75t_R _18794_ (.A1(_10118_),
    .A2(_10086_),
    .B(_10251_),
    .Y(_10476_));
 INVx1_ASAP7_75t_R _18795_ (.A(_10401_),
    .Y(_10477_));
 OAI21x1_ASAP7_75t_R _18796_ (.A1(_10178_),
    .A2(_00395_),
    .B(_10063_),
    .Y(_10478_));
 OAI22x1_ASAP7_75t_R _18797_ (.A1(_10476_),
    .A2(_10477_),
    .B1(_10478_),
    .B2(_10050_),
    .Y(_10479_));
 OAI21x1_ASAP7_75t_R _18798_ (.A1(_00397_),
    .A2(_10479_),
    .B(_00398_),
    .Y(_10480_));
 OA21x2_ASAP7_75t_R _18799_ (.A1(_10157_),
    .A2(_10094_),
    .B(_10350_),
    .Y(_10481_));
 AOI211x1_ASAP7_75t_R _18800_ (.A1(_10073_),
    .A2(_10193_),
    .B(_10481_),
    .C(_10221_),
    .Y(_10482_));
 OA21x2_ASAP7_75t_R _18801_ (.A1(_10092_),
    .A2(_10178_),
    .B(_10149_),
    .Y(_10483_));
 AO21x1_ASAP7_75t_R _18802_ (.A1(_10483_),
    .A2(_10047_),
    .B(_10134_),
    .Y(_10484_));
 NOR2x1_ASAP7_75t_R _18803_ (.A(_10482_),
    .B(_10484_),
    .Y(_10485_));
 OAI21x1_ASAP7_75t_R _18804_ (.A1(_10480_),
    .A2(_10485_),
    .B(_00399_),
    .Y(_10486_));
 OA21x2_ASAP7_75t_R _18805_ (.A1(_10212_),
    .A2(_15786_),
    .B(_10149_),
    .Y(_10487_));
 AO21x1_ASAP7_75t_R _18806_ (.A1(_10487_),
    .A2(_10130_),
    .B(_10134_),
    .Y(_10488_));
 AO21x1_ASAP7_75t_R _18807_ (.A1(_10114_),
    .A2(_10063_),
    .B(_10212_),
    .Y(_10489_));
 AO21x1_ASAP7_75t_R _18808_ (.A1(_10060_),
    .A2(_10192_),
    .B(_08217_),
    .Y(_10490_));
 AND3x1_ASAP7_75t_R _18809_ (.A(_10489_),
    .B(_10490_),
    .C(_10074_),
    .Y(_10491_));
 NOR2x1_ASAP7_75t_R _18810_ (.A(_10488_),
    .B(_10491_),
    .Y(_10492_));
 AO21x1_ASAP7_75t_R _18811_ (.A1(_10052_),
    .A2(_10295_),
    .B(_10350_),
    .Y(_10493_));
 OA21x2_ASAP7_75t_R _18812_ (.A1(_10125_),
    .A2(_10166_),
    .B(_08226_),
    .Y(_10494_));
 AOI21x1_ASAP7_75t_R _18813_ (.A1(_10493_),
    .A2(_10494_),
    .B(_10164_),
    .Y(_10495_));
 OAI21x1_ASAP7_75t_R _18814_ (.A1(_10157_),
    .A2(_10128_),
    .B(_10073_),
    .Y(_10496_));
 NAND3x1_ASAP7_75t_R _18815_ (.A(_10057_),
    .B(_10496_),
    .C(_10221_),
    .Y(_10497_));
 AO21x1_ASAP7_75t_R _18816_ (.A1(_10495_),
    .A2(_10497_),
    .B(_10111_),
    .Y(_10498_));
 NAND2x1_ASAP7_75t_R _18817_ (.A(_00481_),
    .B(_10350_),
    .Y(_10499_));
 OAI21x1_ASAP7_75t_R _18818_ (.A1(net502),
    .A2(_15796_),
    .B(_10118_),
    .Y(_10500_));
 AOI21x1_ASAP7_75t_R _18819_ (.A1(_10499_),
    .A2(_10500_),
    .B(_10131_),
    .Y(_10501_));
 OAI21x1_ASAP7_75t_R _18820_ (.A1(_10087_),
    .A2(_10294_),
    .B(_10118_),
    .Y(_10502_));
 OAI21x1_ASAP7_75t_R _18821_ (.A1(_10137_),
    .A2(_10116_),
    .B(_10357_),
    .Y(_10503_));
 AOI21x1_ASAP7_75t_R _18822_ (.A1(_10502_),
    .A2(_10503_),
    .B(_10221_),
    .Y(_10504_));
 OAI21x1_ASAP7_75t_R _18823_ (.A1(_10501_),
    .A2(_10504_),
    .B(_10108_),
    .Y(_10505_));
 OAI21x1_ASAP7_75t_R _18824_ (.A1(_10053_),
    .A2(_10062_),
    .B(_10118_),
    .Y(_10506_));
 AOI21x1_ASAP7_75t_R _18825_ (.A1(_10127_),
    .A2(_10082_),
    .B(_08226_),
    .Y(_10507_));
 AOI21x1_ASAP7_75t_R _18826_ (.A1(_10506_),
    .A2(_10507_),
    .B(_10134_),
    .Y(_10508_));
 NAND2x1_ASAP7_75t_R _18827_ (.A(_10092_),
    .B(_10283_),
    .Y(_10509_));
 AOI21x1_ASAP7_75t_R _18828_ (.A1(_10508_),
    .A2(_10509_),
    .B(_08243_),
    .Y(_10510_));
 AOI21x1_ASAP7_75t_R _18829_ (.A1(_10505_),
    .A2(_10510_),
    .B(_00399_),
    .Y(_10511_));
 OAI21x1_ASAP7_75t_R _18830_ (.A1(_10492_),
    .A2(_10498_),
    .B(_10511_),
    .Y(_10512_));
 OAI21x1_ASAP7_75t_R _18831_ (.A1(_10475_),
    .A2(_10486_),
    .B(_10512_),
    .Y(_00029_));
 OA21x2_ASAP7_75t_R _18832_ (.A1(_10072_),
    .A2(_01147_),
    .B(_10048_),
    .Y(_10513_));
 AND2x2_ASAP7_75t_R _18833_ (.A(_10513_),
    .B(_10490_),
    .Y(_10514_));
 AO21x1_ASAP7_75t_R _18834_ (.A1(_10086_),
    .A2(_10295_),
    .B(_10266_),
    .Y(_10515_));
 AO21x1_ASAP7_75t_R _18835_ (.A1(_10244_),
    .A2(_10515_),
    .B(_10134_),
    .Y(_10516_));
 NOR2x1_ASAP7_75t_R _18836_ (.A(_10514_),
    .B(_10516_),
    .Y(_10517_));
 NOR2x1_ASAP7_75t_R _18837_ (.A(_00481_),
    .B(_15794_),
    .Y(_10518_));
 AO21x1_ASAP7_75t_R _18838_ (.A1(_10102_),
    .A2(_10103_),
    .B(_10518_),
    .Y(_10519_));
 OAI21x1_ASAP7_75t_R _18839_ (.A1(_10316_),
    .A2(_10418_),
    .B(_10519_),
    .Y(_10520_));
 AOI21x1_ASAP7_75t_R _18840_ (.A1(_00396_),
    .A2(_10520_),
    .B(_10320_),
    .Y(_10521_));
 OAI21x1_ASAP7_75t_R _18841_ (.A1(_00397_),
    .A2(_10521_),
    .B(_10111_),
    .Y(_10522_));
 OAI21x1_ASAP7_75t_R _18842_ (.A1(_10517_),
    .A2(_10522_),
    .B(_10155_),
    .Y(_10523_));
 AOI21x1_ASAP7_75t_R _18843_ (.A1(_10357_),
    .A2(_10358_),
    .B(_10251_),
    .Y(_10524_));
 OR3x1_ASAP7_75t_R _18844_ (.A(_10046_),
    .B(_10316_),
    .C(_10062_),
    .Y(_10525_));
 NAND2x1_ASAP7_75t_R _18845_ (.A(_10524_),
    .B(_10525_),
    .Y(_10526_));
 NOR2x1_ASAP7_75t_R _18846_ (.A(_10055_),
    .B(_10049_),
    .Y(_10527_));
 AO21x1_ASAP7_75t_R _18847_ (.A1(_10043_),
    .A2(_10044_),
    .B(_10089_),
    .Y(_10528_));
 NAND2x2_ASAP7_75t_R _18848_ (.A(_10528_),
    .B(_10212_),
    .Y(_10529_));
 OAI21x1_ASAP7_75t_R _18849_ (.A1(_10073_),
    .A2(_10126_),
    .B(_10529_),
    .Y(_10530_));
 AOI21x1_ASAP7_75t_R _18850_ (.A1(_10527_),
    .A2(_10530_),
    .B(_10216_),
    .Y(_10531_));
 NAND2x1_ASAP7_75t_R _18851_ (.A(_10526_),
    .B(_10531_),
    .Y(_10532_));
 AO21x1_ASAP7_75t_R _18852_ (.A1(_10102_),
    .A2(_10103_),
    .B(_10114_),
    .Y(_10533_));
 AO21x1_ASAP7_75t_R _18853_ (.A1(_10401_),
    .A2(_10533_),
    .B(_10131_),
    .Y(_10534_));
 OAI21x1_ASAP7_75t_R _18854_ (.A1(_10094_),
    .A2(_10105_),
    .B(_10284_),
    .Y(_10535_));
 AOI21x1_ASAP7_75t_R _18855_ (.A1(_00396_),
    .A2(_10535_),
    .B(_10164_),
    .Y(_10536_));
 NAND2x1_ASAP7_75t_R _18856_ (.A(_10534_),
    .B(_10536_),
    .Y(_10537_));
 AOI21x1_ASAP7_75t_R _18857_ (.A1(_10532_),
    .A2(_10537_),
    .B(_10111_),
    .Y(_10538_));
 OA21x2_ASAP7_75t_R _18858_ (.A1(_10144_),
    .A2(_10094_),
    .B(_10125_),
    .Y(_10539_));
 OAI21x1_ASAP7_75t_R _18859_ (.A1(_10477_),
    .A2(_10539_),
    .B(_00396_),
    .Y(_10540_));
 INVx2_ASAP7_75t_R _18860_ (.A(_10117_),
    .Y(_10541_));
 AO21x1_ASAP7_75t_R _18861_ (.A1(_10045_),
    .A2(_10541_),
    .B(_10266_),
    .Y(_10542_));
 NAND2x1_ASAP7_75t_R _18862_ (.A(_10065_),
    .B(_10192_),
    .Y(_10543_));
 NAND2x1_ASAP7_75t_R _18863_ (.A(_10141_),
    .B(_10543_),
    .Y(_10544_));
 AO21x1_ASAP7_75t_R _18864_ (.A1(_10542_),
    .A2(_10544_),
    .B(_10131_),
    .Y(_10545_));
 AOI21x1_ASAP7_75t_R _18865_ (.A1(_10540_),
    .A2(_10545_),
    .B(_00397_),
    .Y(_10546_));
 OR2x2_ASAP7_75t_R _18866_ (.A(_10233_),
    .B(_10160_),
    .Y(_10547_));
 AOI211x1_ASAP7_75t_R _18867_ (.A1(_10547_),
    .A2(_00395_),
    .B(_10425_),
    .C(_10221_),
    .Y(_10548_));
 OA21x2_ASAP7_75t_R _18868_ (.A1(_10046_),
    .A2(net18),
    .B(_10149_),
    .Y(_10549_));
 OAI21x1_ASAP7_75t_R _18869_ (.A1(_10257_),
    .A2(_10316_),
    .B(_10350_),
    .Y(_10550_));
 AO21x1_ASAP7_75t_R _18870_ (.A1(_10549_),
    .A2(_10550_),
    .B(_10134_),
    .Y(_10551_));
 OAI21x1_ASAP7_75t_R _18871_ (.A1(_10548_),
    .A2(_10551_),
    .B(_00398_),
    .Y(_10552_));
 NOR2x1_ASAP7_75t_R _18872_ (.A(_10546_),
    .B(_10552_),
    .Y(_10553_));
 NOR2x1_ASAP7_75t_R _18873_ (.A(_10166_),
    .B(_00395_),
    .Y(_10554_));
 OA21x2_ASAP7_75t_R _18874_ (.A1(_10041_),
    .A2(_10203_),
    .B(_10082_),
    .Y(_10555_));
 OAI21x1_ASAP7_75t_R _18875_ (.A1(_10554_),
    .A2(_10555_),
    .B(_00396_),
    .Y(_10556_));
 OA21x2_ASAP7_75t_R _18876_ (.A1(_10077_),
    .A2(_10203_),
    .B(_10082_),
    .Y(_10557_));
 OAI21x1_ASAP7_75t_R _18877_ (.A1(_10557_),
    .A2(_10539_),
    .B(_10050_),
    .Y(_10558_));
 AOI21x1_ASAP7_75t_R _18878_ (.A1(_10556_),
    .A2(_10558_),
    .B(_00397_),
    .Y(_10559_));
 NAND2x1_ASAP7_75t_R _18879_ (.A(_10311_),
    .B(_10168_),
    .Y(_10560_));
 OAI21x1_ASAP7_75t_R _18880_ (.A1(_10073_),
    .A2(_10560_),
    .B(_10172_),
    .Y(_10561_));
 NOR2x1_ASAP7_75t_R _18881_ (.A(_10116_),
    .B(_10431_),
    .Y(_10562_));
 NOR2x1_ASAP7_75t_R _18882_ (.A(_10561_),
    .B(_10562_),
    .Y(_10563_));
 OA21x2_ASAP7_75t_R _18883_ (.A1(_10116_),
    .A2(_10062_),
    .B(_10118_),
    .Y(_10564_));
 AO21x1_ASAP7_75t_R _18884_ (.A1(_10357_),
    .A2(_00488_),
    .B(_10049_),
    .Y(_10565_));
 OAI21x1_ASAP7_75t_R _18885_ (.A1(_10564_),
    .A2(_10565_),
    .B(_10164_),
    .Y(_10566_));
 OAI21x1_ASAP7_75t_R _18886_ (.A1(_10563_),
    .A2(_10566_),
    .B(_10111_),
    .Y(_10567_));
 OAI21x1_ASAP7_75t_R _18887_ (.A1(_10559_),
    .A2(_10567_),
    .B(_00399_),
    .Y(_10568_));
 OAI22x1_ASAP7_75t_R _18888_ (.A1(_10523_),
    .A2(_10538_),
    .B1(_10553_),
    .B2(_10568_),
    .Y(_00030_));
 NOR2x2_ASAP7_75t_R _18889_ (.A(net864),
    .B(_15796_),
    .Y(_10569_));
 AO21x1_ASAP7_75t_R _18890_ (.A1(_10139_),
    .A2(_10541_),
    .B(_10125_),
    .Y(_10570_));
 OA21x2_ASAP7_75t_R _18891_ (.A1(_10569_),
    .A2(_10467_),
    .B(_10570_),
    .Y(_10571_));
 AO21x1_ASAP7_75t_R _18892_ (.A1(_10456_),
    .A2(_10529_),
    .B(_10131_),
    .Y(_10572_));
 OAI21x1_ASAP7_75t_R _18893_ (.A1(_10050_),
    .A2(_10571_),
    .B(_10572_),
    .Y(_10573_));
 AOI211x1_ASAP7_75t_R _18894_ (.A1(_10073_),
    .A2(_10268_),
    .B(_10279_),
    .C(_10221_),
    .Y(_10574_));
 AO21x1_ASAP7_75t_R _18895_ (.A1(_10543_),
    .A2(_10118_),
    .B(_10251_),
    .Y(_10575_));
 OAI21x1_ASAP7_75t_R _18896_ (.A1(_10340_),
    .A2(_10575_),
    .B(_10108_),
    .Y(_10576_));
 OAI21x1_ASAP7_75t_R _18897_ (.A1(_10574_),
    .A2(_10576_),
    .B(_00398_),
    .Y(_10577_));
 AOI21x1_ASAP7_75t_R _18898_ (.A1(_00397_),
    .A2(_10573_),
    .B(_10577_),
    .Y(_10578_));
 OA21x2_ASAP7_75t_R _18899_ (.A1(_10266_),
    .A2(_10052_),
    .B(_10049_),
    .Y(_10579_));
 AOI21x1_ASAP7_75t_R _18900_ (.A1(_10146_),
    .A2(_10579_),
    .B(_10164_),
    .Y(_10580_));
 OAI21x1_ASAP7_75t_R _18901_ (.A1(_10569_),
    .A2(_10141_),
    .B(_08226_),
    .Y(_10581_));
 AO21x1_ASAP7_75t_R _18902_ (.A1(_10073_),
    .A2(_10231_),
    .B(_10581_),
    .Y(_10582_));
 AO21x1_ASAP7_75t_R _18903_ (.A1(_10580_),
    .A2(_10582_),
    .B(_08243_),
    .Y(_10583_));
 AO21x1_ASAP7_75t_R _18904_ (.A1(_10060_),
    .A2(_10541_),
    .B(_10120_),
    .Y(_10584_));
 AO21x1_ASAP7_75t_R _18905_ (.A1(_10584_),
    .A2(_10348_),
    .B(_10131_),
    .Y(_10585_));
 OA21x2_ASAP7_75t_R _18906_ (.A1(net824),
    .A2(_10082_),
    .B(_10421_),
    .Y(_10586_));
 NAND2x1_ASAP7_75t_R _18907_ (.A(_00396_),
    .B(_10586_),
    .Y(_10587_));
 AOI21x1_ASAP7_75t_R _18908_ (.A1(_10585_),
    .A2(_10587_),
    .B(_10108_),
    .Y(_10588_));
 OAI21x1_ASAP7_75t_R _18909_ (.A1(_10583_),
    .A2(_10588_),
    .B(_10155_),
    .Y(_10589_));
 INVx1_ASAP7_75t_R _18910_ (.A(_10457_),
    .Y(_10590_));
 NOR2x1_ASAP7_75t_R _18911_ (.A(_10042_),
    .B(_10046_),
    .Y(_10591_));
 AO21x1_ASAP7_75t_R _18912_ (.A1(_10179_),
    .A2(_10042_),
    .B(_10591_),
    .Y(_10592_));
 NAND2x1_ASAP7_75t_R _18913_ (.A(net501),
    .B(_10120_),
    .Y(_10593_));
 AOI21x1_ASAP7_75t_R _18914_ (.A1(_10233_),
    .A2(_10266_),
    .B(_10194_),
    .Y(_10594_));
 AOI21x1_ASAP7_75t_R _18915_ (.A1(_10593_),
    .A2(_10594_),
    .B(_10196_),
    .Y(_10595_));
 OAI21x1_ASAP7_75t_R _18916_ (.A1(_10590_),
    .A2(_10592_),
    .B(_10595_),
    .Y(_10596_));
 NOR2x1_ASAP7_75t_R _18917_ (.A(_10144_),
    .B(_10116_),
    .Y(_10597_));
 AOI21x1_ASAP7_75t_R _18918_ (.A1(_10120_),
    .A2(_10597_),
    .B(_10343_),
    .Y(_10598_));
 NAND2x1_ASAP7_75t_R _18919_ (.A(_10598_),
    .B(_10244_),
    .Y(_10599_));
 AOI21x1_ASAP7_75t_R _18920_ (.A1(_10160_),
    .A2(_10141_),
    .B(_08226_),
    .Y(_10600_));
 OAI21x1_ASAP7_75t_R _18921_ (.A1(_08215_),
    .A2(_10088_),
    .B(_01150_),
    .Y(_10601_));
 OAI21x1_ASAP7_75t_R _18922_ (.A1(_10350_),
    .A2(_10144_),
    .B(_10601_),
    .Y(_10602_));
 AOI21x1_ASAP7_75t_R _18923_ (.A1(_10600_),
    .A2(_10602_),
    .B(_10164_),
    .Y(_10603_));
 AOI21x1_ASAP7_75t_R _18924_ (.A1(_10599_),
    .A2(_10603_),
    .B(_08243_),
    .Y(_10604_));
 AOI21x1_ASAP7_75t_R _18925_ (.A1(_10596_),
    .A2(_10604_),
    .B(_10155_),
    .Y(_10605_));
 AO21x1_ASAP7_75t_R _18926_ (.A1(_10168_),
    .A2(_10541_),
    .B(_10132_),
    .Y(_10606_));
 AND2x2_ASAP7_75t_R _18927_ (.A(_10453_),
    .B(_10606_),
    .Y(_10607_));
 OA21x2_ASAP7_75t_R _18928_ (.A1(_10365_),
    .A2(_10266_),
    .B(_10149_),
    .Y(_10608_));
 AO21x1_ASAP7_75t_R _18929_ (.A1(_10139_),
    .A2(_10541_),
    .B(_10350_),
    .Y(_10609_));
 AO21x1_ASAP7_75t_R _18930_ (.A1(_10608_),
    .A2(_10609_),
    .B(_10216_),
    .Y(_10610_));
 OA21x2_ASAP7_75t_R _18931_ (.A1(_10148_),
    .A2(_10042_),
    .B(_10139_),
    .Y(_10611_));
 NAND2x1_ASAP7_75t_R _18932_ (.A(_10594_),
    .B(_10611_),
    .Y(_10612_));
 OA21x2_ASAP7_75t_R _18933_ (.A1(_10056_),
    .A2(_01144_),
    .B(_10194_),
    .Y(_10613_));
 AOI21x1_ASAP7_75t_R _18934_ (.A1(_10550_),
    .A2(_10613_),
    .B(_10164_),
    .Y(_10614_));
 AOI21x1_ASAP7_75t_R _18935_ (.A1(_10612_),
    .A2(_10614_),
    .B(_10110_),
    .Y(_10615_));
 OAI21x1_ASAP7_75t_R _18936_ (.A1(_10607_),
    .A2(_10610_),
    .B(_10615_),
    .Y(_10616_));
 NAND2x1_ASAP7_75t_R _18937_ (.A(_10605_),
    .B(_10616_),
    .Y(_10617_));
 OAI21x1_ASAP7_75t_R _18938_ (.A1(_10578_),
    .A2(_10589_),
    .B(_10617_),
    .Y(_00031_));
 BUFx6f_ASAP7_75t_R _18939_ (.A(_00731_),
    .Y(_10618_));
 BUFx16f_ASAP7_75t_R _18940_ (.A(_10618_),
    .Y(_10619_));
 BUFx16f_ASAP7_75t_R _18941_ (.A(_10619_),
    .Y(_10620_));
 BUFx16f_ASAP7_75t_R _18942_ (.A(_10620_),
    .Y(_10621_));
 NOR2x2_ASAP7_75t_R _18943_ (.A(_00489_),
    .B(_10621_),
    .Y(_10622_));
 XOR2x2_ASAP7_75t_R _18944_ (.A(_00764_),
    .B(_00771_),
    .Y(_10623_));
 BUFx10_ASAP7_75t_R _18945_ (.A(_00829_),
    .Y(_10624_));
 XOR2x1_ASAP7_75t_R _18946_ (.A(_10623_),
    .Y(_10625_),
    .B(_10624_));
 BUFx6f_ASAP7_75t_R _18947_ (.A(_00739_),
    .Y(_10626_));
 XOR2x2_ASAP7_75t_R _18948_ (.A(_10626_),
    .B(_00732_),
    .Y(_10627_));
 BUFx6f_ASAP7_75t_R _18949_ (.A(_00797_),
    .Y(_10628_));
 XOR2x2_ASAP7_75t_R _18950_ (.A(_00765_),
    .B(_10628_),
    .Y(_10629_));
 XOR2x1_ASAP7_75t_R _18951_ (.A(_10627_),
    .Y(_10630_),
    .B(_10629_));
 NAND2x1_ASAP7_75t_R _18952_ (.A(_10625_),
    .B(_10630_),
    .Y(_10631_));
 INVx3_ASAP7_75t_R _18953_ (.A(_10624_),
    .Y(_10632_));
 XOR2x1_ASAP7_75t_R _18954_ (.A(_10623_),
    .Y(_10633_),
    .B(_10632_));
 BUFx6f_ASAP7_75t_R _18955_ (.A(_00732_),
    .Y(_10634_));
 XNOR2x2_ASAP7_75t_R _18956_ (.A(_10634_),
    .B(_10626_),
    .Y(_10635_));
 XOR2x1_ASAP7_75t_R _18957_ (.A(_10635_),
    .Y(_10636_),
    .B(_10629_));
 NAND2x1_ASAP7_75t_R _18958_ (.A(_10633_),
    .B(_10636_),
    .Y(_10637_));
 INVx6_ASAP7_75t_R _18959_ (.A(_10618_),
    .Y(_10638_));
 BUFx16f_ASAP7_75t_R _18960_ (.A(_10638_),
    .Y(_10639_));
 BUFx12_ASAP7_75t_R _18961_ (.A(_10639_),
    .Y(_10640_));
 AOI21x1_ASAP7_75t_R _18962_ (.A1(_10631_),
    .A2(_10637_),
    .B(_10640_),
    .Y(_10641_));
 OAI21x1_ASAP7_75t_R _18963_ (.A1(_10622_),
    .A2(_10641_),
    .B(_08185_),
    .Y(_10642_));
 BUFx16f_ASAP7_75t_R _18964_ (.A(_10638_),
    .Y(_10643_));
 AND2x2_ASAP7_75t_R _18965_ (.A(_10643_),
    .B(_00489_),
    .Y(_10644_));
 NAND2x1_ASAP7_75t_R _18966_ (.A(_10633_),
    .B(_10630_),
    .Y(_10645_));
 NAND2x1_ASAP7_75t_R _18967_ (.A(_10625_),
    .B(_10636_),
    .Y(_10646_));
 AOI21x1_ASAP7_75t_R _18968_ (.A1(_10645_),
    .A2(_10646_),
    .B(_10640_),
    .Y(_10647_));
 INVx1_ASAP7_75t_R _18969_ (.A(_08185_),
    .Y(_10648_));
 OAI21x1_ASAP7_75t_R _18970_ (.A1(_10644_),
    .A2(_10647_),
    .B(_10648_),
    .Y(_10649_));
 NAND2x2_ASAP7_75t_R _18971_ (.A(_10642_),
    .B(_10649_),
    .Y(_10650_));
 BUFx10_ASAP7_75t_R _18972_ (.A(_10650_),
    .Y(_15804_));
 BUFx6f_ASAP7_75t_R _18973_ (.A(_00828_),
    .Y(_10651_));
 INVx2_ASAP7_75t_R _18974_ (.A(net670),
    .Y(_10652_));
 BUFx6f_ASAP7_75t_R _18975_ (.A(_00771_),
    .Y(_10653_));
 XOR2x2_ASAP7_75t_R _18976_ (.A(_10626_),
    .B(_10653_),
    .Y(_10654_));
 NAND2x1_ASAP7_75t_R _18977_ (.A(_10652_),
    .B(_10654_),
    .Y(_10655_));
 XNOR2x1_ASAP7_75t_R _18978_ (.B(_10653_),
    .Y(_10656_),
    .A(_10626_));
 NAND2x1_ASAP7_75t_R _18979_ (.A(net670),
    .B(_10656_),
    .Y(_10657_));
 BUFx6f_ASAP7_75t_R _18980_ (.A(_00764_),
    .Y(_10658_));
 XNOR2x2_ASAP7_75t_R _18981_ (.A(_10658_),
    .B(_00796_),
    .Y(_10659_));
 AOI21x1_ASAP7_75t_R _18982_ (.A1(_10655_),
    .A2(_10657_),
    .B(_10659_),
    .Y(_10660_));
 NAND2x1_ASAP7_75t_R _18983_ (.A(net670),
    .B(_10654_),
    .Y(_10661_));
 NAND2x1_ASAP7_75t_R _18984_ (.A(_10652_),
    .B(_10656_),
    .Y(_10662_));
 XOR2x2_ASAP7_75t_R _18985_ (.A(_10658_),
    .B(_00796_),
    .Y(_10663_));
 AOI21x1_ASAP7_75t_R _18986_ (.A1(_10661_),
    .A2(_10662_),
    .B(_10663_),
    .Y(_10664_));
 BUFx16f_ASAP7_75t_R _18987_ (.A(_10619_),
    .Y(_10665_));
 BUFx16f_ASAP7_75t_R _18988_ (.A(_10665_),
    .Y(_10666_));
 OAI21x1_ASAP7_75t_R _18989_ (.A1(_10660_),
    .A2(_10664_),
    .B(_10666_),
    .Y(_10667_));
 BUFx16f_ASAP7_75t_R _18990_ (.A(_10619_),
    .Y(_10668_));
 NOR2x2_ASAP7_75t_R _18991_ (.A(_10668_),
    .B(_00490_),
    .Y(_10669_));
 INVx3_ASAP7_75t_R _18992_ (.A(_10669_),
    .Y(_10670_));
 NAND3x2_ASAP7_75t_R _18993_ (.B(_08401_),
    .C(_10670_),
    .Y(_10671_),
    .A(net545));
 AO21x2_ASAP7_75t_R _18994_ (.A1(_10667_),
    .A2(_10670_),
    .B(_08401_),
    .Y(_10672_));
 NAND2x2_ASAP7_75t_R _18995_ (.A(_10671_),
    .B(_10672_),
    .Y(_15806_));
 NOR2x2_ASAP7_75t_R _18996_ (.A(_10619_),
    .B(_00492_),
    .Y(_10673_));
 BUFx6f_ASAP7_75t_R _18997_ (.A(_00766_),
    .Y(_10674_));
 INVx3_ASAP7_75t_R _18998_ (.A(_10674_),
    .Y(_10675_));
 BUFx6f_ASAP7_75t_R _18999_ (.A(_00733_),
    .Y(_10676_));
 XOR2x2_ASAP7_75t_R _19000_ (.A(_00765_),
    .B(_10676_),
    .Y(_10677_));
 NOR2x1_ASAP7_75t_R _19001_ (.A(_10675_),
    .B(_10677_),
    .Y(_10678_));
 XNOR2x2_ASAP7_75t_R _19002_ (.A(_10676_),
    .B(_00765_),
    .Y(_10679_));
 NOR2x1_ASAP7_75t_R _19003_ (.A(_10674_),
    .B(net631),
    .Y(_10680_));
 BUFx10_ASAP7_75t_R _19004_ (.A(_00798_),
    .Y(_10681_));
 BUFx10_ASAP7_75t_R _19005_ (.A(_00830_),
    .Y(_10682_));
 XOR2x2_ASAP7_75t_R _19006_ (.A(_10681_),
    .B(_10682_),
    .Y(_10683_));
 OAI21x1_ASAP7_75t_R _19007_ (.A1(_10678_),
    .A2(_10680_),
    .B(_10683_),
    .Y(_10684_));
 NOR2x1_ASAP7_75t_R _19008_ (.A(_10674_),
    .B(net684),
    .Y(_10685_));
 NOR2x1_ASAP7_75t_R _19009_ (.A(_10675_),
    .B(net631),
    .Y(_10686_));
 XNOR2x2_ASAP7_75t_R _19010_ (.A(_10681_),
    .B(_10682_),
    .Y(_10687_));
 OAI21x1_ASAP7_75t_R _19011_ (.A1(_10685_),
    .A2(_10686_),
    .B(_10687_),
    .Y(_10688_));
 BUFx12f_ASAP7_75t_R _19012_ (.A(_10639_),
    .Y(_10689_));
 AOI21x1_ASAP7_75t_R _19013_ (.A1(_10684_),
    .A2(_10688_),
    .B(_10689_),
    .Y(_10690_));
 OAI21x1_ASAP7_75t_R _19014_ (.A1(_10673_),
    .A2(_10690_),
    .B(_08405_),
    .Y(_10691_));
 NAND2x1_ASAP7_75t_R _19015_ (.A(_10675_),
    .B(net684),
    .Y(_10692_));
 NAND2x1_ASAP7_75t_R _19016_ (.A(_10674_),
    .B(net631),
    .Y(_10693_));
 AOI21x1_ASAP7_75t_R _19017_ (.A1(_10692_),
    .A2(_10693_),
    .B(_10687_),
    .Y(_10694_));
 NAND2x1_ASAP7_75t_R _19018_ (.A(_10674_),
    .B(_10677_),
    .Y(_10695_));
 NAND2x1_ASAP7_75t_R _19019_ (.A(_10675_),
    .B(net631),
    .Y(_10696_));
 AOI21x1_ASAP7_75t_R _19020_ (.A1(_10695_),
    .A2(_10696_),
    .B(_10683_),
    .Y(_10697_));
 OAI21x1_ASAP7_75t_R _19021_ (.A1(_10694_),
    .A2(_10697_),
    .B(net780),
    .Y(_10698_));
 INVx3_ASAP7_75t_R _19022_ (.A(_10673_),
    .Y(_10699_));
 NAND3x2_ASAP7_75t_R _19023_ (.B(_01013_),
    .C(_10699_),
    .Y(_10700_),
    .A(_10698_));
 NAND2x2_ASAP7_75t_R _19024_ (.A(_10691_),
    .B(_10700_),
    .Y(_10701_));
 BUFx10_ASAP7_75t_R _19025_ (.A(_10701_),
    .Y(_15814_));
 NAND3x2_ASAP7_75t_R _19026_ (.B(_01011_),
    .C(_10670_),
    .Y(_10702_),
    .A(net544));
 AO21x1_ASAP7_75t_R _19027_ (.A1(_10667_),
    .A2(_10670_),
    .B(_01011_),
    .Y(_10703_));
 NAND2x2_ASAP7_75t_R _19028_ (.A(_10702_),
    .B(_10703_),
    .Y(_10704_));
 BUFx6f_ASAP7_75t_R _19029_ (.A(_10704_),
    .Y(_15801_));
 NAND3x2_ASAP7_75t_R _19030_ (.B(_08405_),
    .C(_10699_),
    .Y(_10705_),
    .A(_10698_));
 AO21x1_ASAP7_75t_R _19031_ (.A1(_10698_),
    .A2(_10699_),
    .B(_08405_),
    .Y(_10706_));
 BUFx4f_ASAP7_75t_R _19032_ (.A(_10706_),
    .Y(_10707_));
 NAND2x2_ASAP7_75t_R _19033_ (.A(_10705_),
    .B(_10707_),
    .Y(_10708_));
 BUFx10_ASAP7_75t_R _19034_ (.A(_10708_),
    .Y(_10709_));
 BUFx10_ASAP7_75t_R _19035_ (.A(_10709_),
    .Y(_15811_));
 BUFx6f_ASAP7_75t_R _19036_ (.A(_00767_),
    .Y(_10710_));
 BUFx4f_ASAP7_75t_R _19037_ (.A(_00734_),
    .Y(_10711_));
 XOR2x2_ASAP7_75t_R _19038_ (.A(_10711_),
    .B(_10626_),
    .Y(_10712_));
 XNOR2x1_ASAP7_75t_R _19039_ (.B(_10712_),
    .Y(_10713_),
    .A(_10710_));
 BUFx6f_ASAP7_75t_R _19040_ (.A(_00799_),
    .Y(_10714_));
 BUFx6f_ASAP7_75t_R _19041_ (.A(_00831_),
    .Y(_10715_));
 XNOR2x2_ASAP7_75t_R _19042_ (.A(_10714_),
    .B(_10715_),
    .Y(_10716_));
 XOR2x2_ASAP7_75t_R _19043_ (.A(_10674_),
    .B(net726),
    .Y(_10717_));
 XOR2x1_ASAP7_75t_R _19044_ (.A(_10716_),
    .Y(_10718_),
    .B(_10717_));
 NOR2x1_ASAP7_75t_R _19045_ (.A(_10713_),
    .B(_10718_),
    .Y(_10719_));
 XOR2x1_ASAP7_75t_R _19046_ (.A(_10712_),
    .Y(_10720_),
    .B(_10710_));
 XOR2x2_ASAP7_75t_R _19047_ (.A(_10714_),
    .B(_10715_),
    .Y(_10721_));
 XOR2x1_ASAP7_75t_R _19048_ (.A(_10717_),
    .Y(_10722_),
    .B(_10721_));
 BUFx12f_ASAP7_75t_R _19049_ (.A(_10665_),
    .Y(_10723_));
 OAI21x1_ASAP7_75t_R _19050_ (.A1(_10720_),
    .A2(_10722_),
    .B(net651),
    .Y(_10724_));
 NAND2x1_ASAP7_75t_R _19051_ (.A(_00709_),
    .B(_10643_),
    .Y(_10725_));
 OAI21x1_ASAP7_75t_R _19052_ (.A1(_10719_),
    .A2(_10724_),
    .B(_10725_),
    .Y(_10726_));
 XNOR2x2_ASAP7_75t_R _19053_ (.A(_01014_),
    .B(_10726_),
    .Y(_10727_));
 BUFx6f_ASAP7_75t_R _19054_ (.A(_10727_),
    .Y(_10728_));
 AOI21x1_ASAP7_75t_R _19055_ (.A1(_15801_),
    .A2(_15814_),
    .B(_10728_),
    .Y(_10729_));
 INVx1_ASAP7_75t_R _19056_ (.A(_01154_),
    .Y(_10730_));
 AO21x1_ASAP7_75t_R _19057_ (.A1(_10707_),
    .A2(_10705_),
    .B(_10730_),
    .Y(_10731_));
 BUFx4f_ASAP7_75t_R _19058_ (.A(_10731_),
    .Y(_10732_));
 BUFx16f_ASAP7_75t_R _19059_ (.A(_10668_),
    .Y(_10733_));
 BUFx12_ASAP7_75t_R _19060_ (.A(_10733_),
    .Y(_10734_));
 XNOR2x2_ASAP7_75t_R _19061_ (.A(_10710_),
    .B(net726),
    .Y(_10735_));
 XOR2x2_ASAP7_75t_R _19062_ (.A(_00800_),
    .B(_00832_),
    .Y(_10736_));
 XOR2x1_ASAP7_75t_R _19063_ (.A(_10735_),
    .Y(_10737_),
    .B(_10736_));
 XOR2x2_ASAP7_75t_R _19064_ (.A(_00735_),
    .B(net50),
    .Y(_10738_));
 XOR2x1_ASAP7_75t_R _19065_ (.A(_10738_),
    .Y(_10739_),
    .B(_00768_));
 XOR2x1_ASAP7_75t_R _19066_ (.A(_10737_),
    .Y(_10740_),
    .B(_10739_));
 BUFx16f_ASAP7_75t_R _19067_ (.A(_10618_),
    .Y(_10741_));
 BUFx16f_ASAP7_75t_R _19068_ (.A(_10741_),
    .Y(_10742_));
 BUFx16f_ASAP7_75t_R _19069_ (.A(_10742_),
    .Y(_10743_));
 NOR2x1_ASAP7_75t_R _19070_ (.A(_10743_),
    .B(_00708_),
    .Y(_10744_));
 AOI21x1_ASAP7_75t_R _19071_ (.A1(_10734_),
    .A2(_10740_),
    .B(_10744_),
    .Y(_10745_));
 XNOR2x2_ASAP7_75t_R _19072_ (.A(_01015_),
    .B(_10745_),
    .Y(_10746_));
 BUFx6f_ASAP7_75t_R _19073_ (.A(_10746_),
    .Y(_10747_));
 AO21x1_ASAP7_75t_R _19074_ (.A1(_10729_),
    .A2(_10732_),
    .B(_10747_),
    .Y(_10748_));
 NAND2x2_ASAP7_75t_R _19075_ (.A(_10709_),
    .B(net3),
    .Y(_10749_));
 AO21x1_ASAP7_75t_R _19076_ (.A1(_15804_),
    .A2(net65),
    .B(_15811_),
    .Y(_10750_));
 XOR2x2_ASAP7_75t_R _19077_ (.A(_10726_),
    .B(_01014_),
    .Y(_10751_));
 BUFx6f_ASAP7_75t_R _19078_ (.A(_10751_),
    .Y(_10752_));
 BUFx6f_ASAP7_75t_R _19079_ (.A(_10752_),
    .Y(_10753_));
 AOI21x1_ASAP7_75t_R _19080_ (.A1(_10749_),
    .A2(_10750_),
    .B(_10753_),
    .Y(_10754_));
 XOR2x2_ASAP7_75t_R _19081_ (.A(_00769_),
    .B(_00801_),
    .Y(_10755_));
 BUFx4f_ASAP7_75t_R _19082_ (.A(_00736_),
    .Y(_10756_));
 XOR2x2_ASAP7_75t_R _19083_ (.A(_10756_),
    .B(_00768_),
    .Y(_10757_));
 BUFx6f_ASAP7_75t_R _19084_ (.A(_00833_),
    .Y(_10758_));
 XOR2x1_ASAP7_75t_R _19085_ (.A(_10757_),
    .Y(_10759_),
    .B(_10758_));
 XNOR2x1_ASAP7_75t_R _19086_ (.B(_10759_),
    .Y(_10760_),
    .A(_10755_));
 BUFx12f_ASAP7_75t_R _19087_ (.A(_10666_),
    .Y(_10761_));
 BUFx16f_ASAP7_75t_R _19088_ (.A(_10741_),
    .Y(_10762_));
 BUFx12f_ASAP7_75t_R _19089_ (.A(_10762_),
    .Y(_10763_));
 NOR2x1_ASAP7_75t_R _19090_ (.A(_10763_),
    .B(_00707_),
    .Y(_10764_));
 AO21x1_ASAP7_75t_R _19091_ (.A1(_10760_),
    .A2(_10761_),
    .B(_10764_),
    .Y(_10765_));
 XOR2x2_ASAP7_75t_R _19092_ (.A(_10765_),
    .B(_01016_),
    .Y(_10766_));
 BUFx10_ASAP7_75t_R _19093_ (.A(_10766_),
    .Y(_10767_));
 OAI21x1_ASAP7_75t_R _19094_ (.A1(_10748_),
    .A2(_10754_),
    .B(_10767_),
    .Y(_10768_));
 BUFx12_ASAP7_75t_R _19095_ (.A(_10701_),
    .Y(_10769_));
 NOR2x2_ASAP7_75t_R _19096_ (.A(_01151_),
    .B(_10769_),
    .Y(_10770_));
 NOR2x2_ASAP7_75t_R _19097_ (.A(_10708_),
    .B(_10650_),
    .Y(_10771_));
 NOR2x1_ASAP7_75t_R _19098_ (.A(_10770_),
    .B(_10771_),
    .Y(_10772_));
 NOR2x1_ASAP7_75t_R _19099_ (.A(_10753_),
    .B(_10772_),
    .Y(_10773_));
 NOR2x2_ASAP7_75t_R _19100_ (.A(_10701_),
    .B(net784),
    .Y(_10774_));
 NAND2x2_ASAP7_75t_R _19101_ (.A(_15804_),
    .B(_10774_),
    .Y(_10775_));
 XOR2x2_ASAP7_75t_R _19102_ (.A(_10745_),
    .B(_01015_),
    .Y(_10776_));
 BUFx6f_ASAP7_75t_R _19103_ (.A(_10776_),
    .Y(_10777_));
 BUFx6f_ASAP7_75t_R _19104_ (.A(_10777_),
    .Y(_10778_));
 AO21x1_ASAP7_75t_R _19105_ (.A1(_10775_),
    .A2(_10729_),
    .B(_10778_),
    .Y(_10779_));
 NOR2x1_ASAP7_75t_R _19106_ (.A(_10773_),
    .B(_10779_),
    .Y(_10780_));
 XOR2x2_ASAP7_75t_R _19107_ (.A(_00770_),
    .B(_00802_),
    .Y(_10781_));
 XOR2x1_ASAP7_75t_R _19108_ (.A(_10781_),
    .Y(_10782_),
    .B(_00834_));
 BUFx6f_ASAP7_75t_R _19109_ (.A(_00737_),
    .Y(_10783_));
 XNOR2x2_ASAP7_75t_R _19110_ (.A(_10783_),
    .B(_00769_),
    .Y(_10784_));
 XOR2x1_ASAP7_75t_R _19111_ (.A(_10782_),
    .Y(_10785_),
    .B(_10784_));
 BUFx12f_ASAP7_75t_R _19112_ (.A(_10761_),
    .Y(_10786_));
 BUFx12f_ASAP7_75t_R _19113_ (.A(_10763_),
    .Y(_10787_));
 NOR2x1_ASAP7_75t_R _19114_ (.A(_10787_),
    .B(_00706_),
    .Y(_10788_));
 AO21x1_ASAP7_75t_R _19115_ (.A1(_10785_),
    .A2(_10786_),
    .B(_10788_),
    .Y(_10789_));
 XOR2x2_ASAP7_75t_R _19116_ (.A(_10789_),
    .B(_01018_),
    .Y(_10790_));
 CKINVDCx6p67_ASAP7_75t_R _19117_ (.A(_10790_),
    .Y(_10791_));
 BUFx10_ASAP7_75t_R _19118_ (.A(_10791_),
    .Y(_10792_));
 OAI21x1_ASAP7_75t_R _19119_ (.A1(_10768_),
    .A2(_10780_),
    .B(_10792_),
    .Y(_10793_));
 INVx2_ASAP7_75t_R _19120_ (.A(_01152_),
    .Y(_10794_));
 AOI21x1_ASAP7_75t_R _19121_ (.A1(_10705_),
    .A2(_10707_),
    .B(_10794_),
    .Y(_10795_));
 NOR2x2_ASAP7_75t_R _19122_ (.A(_10727_),
    .B(_10795_),
    .Y(_10796_));
 NOR2x2_ASAP7_75t_R _19123_ (.A(_15806_),
    .B(_10708_),
    .Y(_10797_));
 NAND2x2_ASAP7_75t_R _19124_ (.A(net3),
    .B(_10797_),
    .Y(_10798_));
 NAND2x1_ASAP7_75t_R _19125_ (.A(_10796_),
    .B(_10798_),
    .Y(_10799_));
 AOI21x1_ASAP7_75t_R _19126_ (.A1(net784),
    .A2(_10769_),
    .B(_10751_),
    .Y(_10800_));
 INVx2_ASAP7_75t_R _19127_ (.A(_10800_),
    .Y(_10801_));
 BUFx6f_ASAP7_75t_R _19128_ (.A(_10776_),
    .Y(_10802_));
 BUFx6f_ASAP7_75t_R _19129_ (.A(_10802_),
    .Y(_10803_));
 AO21x1_ASAP7_75t_R _19130_ (.A1(_10799_),
    .A2(_10801_),
    .B(_10803_),
    .Y(_10804_));
 BUFx6f_ASAP7_75t_R _19131_ (.A(_10751_),
    .Y(_10805_));
 NOR2x2_ASAP7_75t_R _19132_ (.A(_10701_),
    .B(_15806_),
    .Y(_10806_));
 NOR2x1_ASAP7_75t_R _19133_ (.A(_10805_),
    .B(_10806_),
    .Y(_10807_));
 NAND2x1_ASAP7_75t_R _19134_ (.A(_10807_),
    .B(_10798_),
    .Y(_10808_));
 BUFx6f_ASAP7_75t_R _19135_ (.A(_10700_),
    .Y(_10809_));
 BUFx4f_ASAP7_75t_R _19136_ (.A(_10691_),
    .Y(_10810_));
 AO21x1_ASAP7_75t_R _19137_ (.A1(_10809_),
    .A2(_10810_),
    .B(_10730_),
    .Y(_10811_));
 BUFx4f_ASAP7_75t_R _19138_ (.A(_10811_),
    .Y(_10812_));
 INVx3_ASAP7_75t_R _19139_ (.A(net466),
    .Y(_10813_));
 AOI21x1_ASAP7_75t_R _19140_ (.A1(_10705_),
    .A2(_10707_),
    .B(_10813_),
    .Y(_10814_));
 NOR2x2_ASAP7_75t_R _19141_ (.A(net486),
    .B(_10727_),
    .Y(_10815_));
 NAND2x1_ASAP7_75t_R _19142_ (.A(_10812_),
    .B(net1),
    .Y(_10816_));
 BUFx6f_ASAP7_75t_R _19143_ (.A(_10746_),
    .Y(_10817_));
 BUFx6f_ASAP7_75t_R _19144_ (.A(_10817_),
    .Y(_10818_));
 AO21x1_ASAP7_75t_R _19145_ (.A1(_10808_),
    .A2(_10816_),
    .B(_10818_),
    .Y(_10819_));
 AOI21x1_ASAP7_75t_R _19146_ (.A1(_10804_),
    .A2(_10819_),
    .B(_10767_),
    .Y(_10820_));
 XNOR2x2_ASAP7_75t_R _19147_ (.A(_00738_),
    .B(_00770_),
    .Y(_10821_));
 BUFx6f_ASAP7_75t_R _19148_ (.A(_00835_),
    .Y(_10822_));
 INVx4_ASAP7_75t_R _19149_ (.A(net682),
    .Y(_10823_));
 XOR2x1_ASAP7_75t_R _19150_ (.A(_10821_),
    .Y(_10824_),
    .B(_10823_));
 BUFx10_ASAP7_75t_R _19151_ (.A(_10653_),
    .Y(_10825_));
 BUFx6f_ASAP7_75t_R _19152_ (.A(_00803_),
    .Y(_10826_));
 XNOR2x2_ASAP7_75t_R _19153_ (.A(_10825_),
    .B(net58),
    .Y(_10827_));
 XOR2x1_ASAP7_75t_R _19154_ (.A(_10824_),
    .Y(_10828_),
    .B(_10827_));
 BUFx12f_ASAP7_75t_R _19155_ (.A(_10743_),
    .Y(_10829_));
 BUFx10_ASAP7_75t_R _19156_ (.A(_10829_),
    .Y(_10830_));
 BUFx12_ASAP7_75t_R _19157_ (.A(_10787_),
    .Y(_10831_));
 NOR2x1_ASAP7_75t_R _19158_ (.A(_10831_),
    .B(_00705_),
    .Y(_10832_));
 AO21x1_ASAP7_75t_R _19159_ (.A1(_10828_),
    .A2(_10830_),
    .B(_10832_),
    .Y(_10833_));
 XOR2x2_ASAP7_75t_R _19160_ (.A(_10833_),
    .B(_01019_),
    .Y(_10834_));
 BUFx10_ASAP7_75t_R _19161_ (.A(_10834_),
    .Y(_10835_));
 OAI21x1_ASAP7_75t_R _19162_ (.A1(_10793_),
    .A2(_10820_),
    .B(_10835_),
    .Y(_10836_));
 AOI21x1_ASAP7_75t_R _19163_ (.A1(_15806_),
    .A2(_10709_),
    .B(_10805_),
    .Y(_10837_));
 INVx4_ASAP7_75t_R _19164_ (.A(_10650_),
    .Y(_10838_));
 BUFx6f_ASAP7_75t_R _19165_ (.A(_10838_),
    .Y(_15802_));
 NAND2x2_ASAP7_75t_R _19166_ (.A(net65),
    .B(_15802_),
    .Y(_10839_));
 NAND2x1_ASAP7_75t_R _19167_ (.A(_10837_),
    .B(_10839_),
    .Y(_10840_));
 AOI22x1_ASAP7_75t_R _19168_ (.A1(_10672_),
    .A2(_10671_),
    .B1(_10809_),
    .B2(_10691_),
    .Y(_10841_));
 INVx5_ASAP7_75t_R _19169_ (.A(_10841_),
    .Y(_10842_));
 BUFx10_ASAP7_75t_R _19170_ (.A(_10727_),
    .Y(_10843_));
 AOI21x1_ASAP7_75t_R _19171_ (.A1(_15801_),
    .A2(_15804_),
    .B(_10843_),
    .Y(_10844_));
 NAND2x1_ASAP7_75t_R _19172_ (.A(_10842_),
    .B(_10844_),
    .Y(_10845_));
 AO21x1_ASAP7_75t_R _19173_ (.A1(_10840_),
    .A2(_10845_),
    .B(_10818_),
    .Y(_10846_));
 NAND2x2_ASAP7_75t_R _19174_ (.A(_15806_),
    .B(net550),
    .Y(_10847_));
 INVx2_ASAP7_75t_R _19175_ (.A(_10847_),
    .Y(_10848_));
 NOR2x2_ASAP7_75t_R _19176_ (.A(net486),
    .B(_10751_),
    .Y(_10849_));
 INVx1_ASAP7_75t_R _19177_ (.A(_10849_),
    .Y(_10850_));
 AO21x1_ASAP7_75t_R _19178_ (.A1(_15814_),
    .A2(_10848_),
    .B(_10850_),
    .Y(_10851_));
 INVx2_ASAP7_75t_R _19179_ (.A(_00491_),
    .Y(_10852_));
 NOR2x2_ASAP7_75t_R _19180_ (.A(_10852_),
    .B(_10769_),
    .Y(_10853_));
 INVx3_ASAP7_75t_R _19181_ (.A(_00493_),
    .Y(_10854_));
 NOR2x1_ASAP7_75t_R _19182_ (.A(_10854_),
    .B(_15811_),
    .Y(_10855_));
 OAI21x1_ASAP7_75t_R _19183_ (.A1(_10853_),
    .A2(_10855_),
    .B(_10753_),
    .Y(_10856_));
 BUFx6f_ASAP7_75t_R _19184_ (.A(_10777_),
    .Y(_10857_));
 AO21x1_ASAP7_75t_R _19185_ (.A1(_10851_),
    .A2(_10856_),
    .B(_10857_),
    .Y(_10858_));
 AOI21x1_ASAP7_75t_R _19186_ (.A1(_10846_),
    .A2(_10858_),
    .B(_10767_),
    .Y(_10859_));
 INVx6_ASAP7_75t_R _19187_ (.A(_10766_),
    .Y(_10860_));
 BUFx10_ASAP7_75t_R _19188_ (.A(_10860_),
    .Y(_10861_));
 AOI21x1_ASAP7_75t_R _19189_ (.A1(_10691_),
    .A2(_10700_),
    .B(_10813_),
    .Y(_10862_));
 NOR2x2_ASAP7_75t_R _19190_ (.A(_10727_),
    .B(_10862_),
    .Y(_10863_));
 NOR2x2_ASAP7_75t_R _19191_ (.A(_10817_),
    .B(_10863_),
    .Y(_10864_));
 OA21x2_ASAP7_75t_R _19192_ (.A1(_10641_),
    .A2(_10622_),
    .B(_10648_),
    .Y(_10865_));
 OA21x2_ASAP7_75t_R _19193_ (.A1(_10647_),
    .A2(_10644_),
    .B(_08185_),
    .Y(_10866_));
 OAI21x1_ASAP7_75t_R _19194_ (.A1(_10865_),
    .A2(_10866_),
    .B(_10701_),
    .Y(_10867_));
 INVx2_ASAP7_75t_R _19195_ (.A(net486),
    .Y(_10868_));
 BUFx4f_ASAP7_75t_R _19196_ (.A(_10751_),
    .Y(_10869_));
 BUFx6f_ASAP7_75t_R _19197_ (.A(_10869_),
    .Y(_10870_));
 AO21x1_ASAP7_75t_R _19198_ (.A1(_10867_),
    .A2(_10868_),
    .B(_10870_),
    .Y(_10871_));
 AO21x1_ASAP7_75t_R _19199_ (.A1(_10707_),
    .A2(_10705_),
    .B(_10854_),
    .Y(_10872_));
 BUFx4f_ASAP7_75t_R _19200_ (.A(_10872_),
    .Y(_10873_));
 AO21x2_ASAP7_75t_R _19201_ (.A1(_10809_),
    .A2(_10810_),
    .B(_10852_),
    .Y(_10874_));
 BUFx6f_ASAP7_75t_R _19202_ (.A(_10751_),
    .Y(_10875_));
 AO21x1_ASAP7_75t_R _19203_ (.A1(_10873_),
    .A2(_10874_),
    .B(_10875_),
    .Y(_10876_));
 AO21x2_ASAP7_75t_R _19204_ (.A1(_10707_),
    .A2(_10705_),
    .B(net466),
    .Y(_10877_));
 AO21x2_ASAP7_75t_R _19205_ (.A1(_10809_),
    .A2(_10810_),
    .B(_10854_),
    .Y(_10878_));
 BUFx6f_ASAP7_75t_R _19206_ (.A(_10843_),
    .Y(_10879_));
 AO21x1_ASAP7_75t_R _19207_ (.A1(_10877_),
    .A2(_10878_),
    .B(_10879_),
    .Y(_10880_));
 AOI21x1_ASAP7_75t_R _19208_ (.A1(_10876_),
    .A2(_10880_),
    .B(_10857_),
    .Y(_10881_));
 AOI21x1_ASAP7_75t_R _19209_ (.A1(_10864_),
    .A2(_10871_),
    .B(_10881_),
    .Y(_10882_));
 BUFx10_ASAP7_75t_R _19210_ (.A(_10790_),
    .Y(_10883_));
 BUFx10_ASAP7_75t_R _19211_ (.A(_10883_),
    .Y(_10884_));
 OAI21x1_ASAP7_75t_R _19212_ (.A1(_10861_),
    .A2(_10882_),
    .B(_10884_),
    .Y(_10885_));
 NOR2x1_ASAP7_75t_R _19213_ (.A(_10885_),
    .B(_10859_),
    .Y(_10886_));
 NAND2x2_ASAP7_75t_R _19214_ (.A(net783),
    .B(net559),
    .Y(_10887_));
 NOR2x2_ASAP7_75t_R _19215_ (.A(_15814_),
    .B(_10887_),
    .Y(_10888_));
 AO21x2_ASAP7_75t_R _19216_ (.A1(_10809_),
    .A2(_10810_),
    .B(_00491_),
    .Y(_10889_));
 NAND2x2_ASAP7_75t_R _19217_ (.A(_10728_),
    .B(_10889_),
    .Y(_10890_));
 NAND2x1_ASAP7_75t_R _19218_ (.A(_10870_),
    .B(_10770_),
    .Y(_10891_));
 OA21x2_ASAP7_75t_R _19219_ (.A1(_10888_),
    .A2(_10890_),
    .B(_10891_),
    .Y(_10892_));
 BUFx6f_ASAP7_75t_R _19220_ (.A(_10887_),
    .Y(_10893_));
 AOI21x1_ASAP7_75t_R _19221_ (.A1(_01153_),
    .A2(_10769_),
    .B(_10727_),
    .Y(_10894_));
 OAI21x1_ASAP7_75t_R _19222_ (.A1(_15814_),
    .A2(_10893_),
    .B(_10894_),
    .Y(_10895_));
 INVx2_ASAP7_75t_R _19223_ (.A(_01151_),
    .Y(_10896_));
 NAND3x2_ASAP7_75t_R _19224_ (.B(_10896_),
    .C(_10810_),
    .Y(_10897_),
    .A(_10809_));
 OA21x2_ASAP7_75t_R _19225_ (.A1(_10897_),
    .A2(_10875_),
    .B(_10747_),
    .Y(_10898_));
 BUFx6f_ASAP7_75t_R _19226_ (.A(_10766_),
    .Y(_10899_));
 AO21x1_ASAP7_75t_R _19227_ (.A1(_10895_),
    .A2(_10898_),
    .B(_10899_),
    .Y(_10900_));
 AOI21x1_ASAP7_75t_R _19228_ (.A1(_10803_),
    .A2(_10892_),
    .B(_10900_),
    .Y(_10901_));
 AOI21x1_ASAP7_75t_R _19229_ (.A1(_10691_),
    .A2(_10700_),
    .B(_01152_),
    .Y(_10902_));
 AOI21x1_ASAP7_75t_R _19230_ (.A1(net784),
    .A2(net3),
    .B(_10769_),
    .Y(_10903_));
 OAI21x1_ASAP7_75t_R _19231_ (.A1(_10902_),
    .A2(_10903_),
    .B(_10879_),
    .Y(_10904_));
 NAND2x1_ASAP7_75t_R _19232_ (.A(_10873_),
    .B(_10842_),
    .Y(_10905_));
 AO21x1_ASAP7_75t_R _19233_ (.A1(_10809_),
    .A2(_10810_),
    .B(_01151_),
    .Y(_10906_));
 BUFx6f_ASAP7_75t_R _19234_ (.A(_10746_),
    .Y(_10907_));
 OAI21x1_ASAP7_75t_R _19235_ (.A1(_10752_),
    .A2(_10906_),
    .B(_10907_),
    .Y(_10908_));
 AOI21x1_ASAP7_75t_R _19236_ (.A1(_10753_),
    .A2(_10905_),
    .B(_10908_),
    .Y(_10909_));
 NAND2x1_ASAP7_75t_R _19237_ (.A(_10904_),
    .B(_10909_),
    .Y(_10910_));
 AOI21x1_ASAP7_75t_R _19238_ (.A1(_10691_),
    .A2(_10700_),
    .B(net466),
    .Y(_10911_));
 AO21x1_ASAP7_75t_R _19239_ (.A1(_10728_),
    .A2(net537),
    .B(_10907_),
    .Y(_10912_));
 BUFx6f_ASAP7_75t_R _19240_ (.A(_10843_),
    .Y(_10913_));
 NOR2x1_ASAP7_75t_R _19241_ (.A(_01156_),
    .B(_10913_),
    .Y(_10914_));
 OA21x2_ASAP7_75t_R _19242_ (.A1(_10912_),
    .A2(_10914_),
    .B(_10899_),
    .Y(_10915_));
 AO21x1_ASAP7_75t_R _19243_ (.A1(_10910_),
    .A2(_10915_),
    .B(_10792_),
    .Y(_10916_));
 NOR2x2_ASAP7_75t_R _19244_ (.A(_01153_),
    .B(_10769_),
    .Y(_10917_));
 OAI21x1_ASAP7_75t_R _19245_ (.A1(_10902_),
    .A2(_10917_),
    .B(_10913_),
    .Y(_10918_));
 NOR2x1_ASAP7_75t_R _19246_ (.A(_10747_),
    .B(_10815_),
    .Y(_10919_));
 BUFx6f_ASAP7_75t_R _19247_ (.A(_10860_),
    .Y(_10920_));
 AOI21x1_ASAP7_75t_R _19248_ (.A1(_10918_),
    .A2(_10919_),
    .B(_10920_),
    .Y(_10921_));
 INVx1_ASAP7_75t_R _19249_ (.A(_10902_),
    .Y(_10922_));
 OAI21x1_ASAP7_75t_R _19250_ (.A1(_10875_),
    .A2(_10922_),
    .B(_10907_),
    .Y(_10923_));
 AO21x1_ASAP7_75t_R _19251_ (.A1(_10775_),
    .A2(_10729_),
    .B(_10923_),
    .Y(_10924_));
 AOI21x1_ASAP7_75t_R _19252_ (.A1(_10921_),
    .A2(_10924_),
    .B(_10884_),
    .Y(_10925_));
 NOR2x2_ASAP7_75t_R _19253_ (.A(net784),
    .B(_10843_),
    .Y(_10926_));
 NOR2x2_ASAP7_75t_R _19254_ (.A(_10708_),
    .B(_10727_),
    .Y(_10927_));
 OAI21x1_ASAP7_75t_R _19255_ (.A1(_10926_),
    .A2(_10927_),
    .B(_10889_),
    .Y(_10928_));
 INVx2_ASAP7_75t_R _19256_ (.A(net538),
    .Y(_10929_));
 AOI21x1_ASAP7_75t_R _19257_ (.A1(_10709_),
    .A2(net3),
    .B(_10751_),
    .Y(_10930_));
 NAND2x2_ASAP7_75t_R _19258_ (.A(_10929_),
    .B(_10930_),
    .Y(_10931_));
 AOI21x1_ASAP7_75t_R _19259_ (.A1(_10928_),
    .A2(_10931_),
    .B(_10857_),
    .Y(_10932_));
 AOI21x1_ASAP7_75t_R _19260_ (.A1(_10897_),
    .A2(_10878_),
    .B(_10869_),
    .Y(_10933_));
 BUFx6f_ASAP7_75t_R _19261_ (.A(_10777_),
    .Y(_10934_));
 OA21x2_ASAP7_75t_R _19262_ (.A1(_10933_),
    .A2(_10796_),
    .B(_10934_),
    .Y(_10935_));
 OAI21x1_ASAP7_75t_R _19263_ (.A1(_10932_),
    .A2(_10935_),
    .B(_10861_),
    .Y(_10936_));
 AOI21x1_ASAP7_75t_R _19264_ (.A1(_10925_),
    .A2(_10936_),
    .B(_10835_),
    .Y(_10937_));
 OAI21x1_ASAP7_75t_R _19265_ (.A1(_10901_),
    .A2(_10916_),
    .B(_10937_),
    .Y(_10938_));
 OAI21x1_ASAP7_75t_R _19266_ (.A1(_10836_),
    .A2(_10886_),
    .B(_10938_),
    .Y(_00032_));
 INVx2_ASAP7_75t_R _19267_ (.A(_10877_),
    .Y(_10939_));
 OAI21x1_ASAP7_75t_R _19268_ (.A1(_15811_),
    .A2(_10847_),
    .B(_10875_),
    .Y(_10940_));
 AOI21x1_ASAP7_75t_R _19269_ (.A1(_10705_),
    .A2(_10707_),
    .B(_01152_),
    .Y(_10941_));
 AOI21x1_ASAP7_75t_R _19270_ (.A1(_10913_),
    .A2(_10941_),
    .B(_10778_),
    .Y(_10942_));
 OAI21x1_ASAP7_75t_R _19271_ (.A1(_10939_),
    .A2(_10940_),
    .B(_10942_),
    .Y(_10943_));
 OAI21x1_ASAP7_75t_R _19272_ (.A1(net65),
    .A2(net24),
    .B(_15811_),
    .Y(_10944_));
 AOI21x1_ASAP7_75t_R _19273_ (.A1(_01154_),
    .A2(_10701_),
    .B(_10727_),
    .Y(_10945_));
 NAND2x2_ASAP7_75t_R _19274_ (.A(_10709_),
    .B(net604),
    .Y(_10946_));
 AOI21x1_ASAP7_75t_R _19275_ (.A1(_10945_),
    .A2(_10946_),
    .B(_10817_),
    .Y(_10947_));
 OAI21x1_ASAP7_75t_R _19276_ (.A1(_10753_),
    .A2(_10944_),
    .B(_10947_),
    .Y(_10948_));
 NAND2x1_ASAP7_75t_R _19277_ (.A(_10943_),
    .B(_10948_),
    .Y(_10949_));
 OAI21x1_ASAP7_75t_R _19278_ (.A1(_10902_),
    .A2(net486),
    .B(_10870_),
    .Y(_10950_));
 NOR2x2_ASAP7_75t_R _19279_ (.A(_10854_),
    .B(_10701_),
    .Y(_10951_));
 OAI21x1_ASAP7_75t_R _19280_ (.A1(_10951_),
    .A2(_10841_),
    .B(_10913_),
    .Y(_10952_));
 BUFx6f_ASAP7_75t_R _19281_ (.A(_10907_),
    .Y(_10953_));
 AOI21x1_ASAP7_75t_R _19282_ (.A1(_10950_),
    .A2(_10952_),
    .B(_10953_),
    .Y(_10954_));
 NOR2x2_ASAP7_75t_R _19283_ (.A(_10805_),
    .B(net537),
    .Y(_10955_));
 INVx2_ASAP7_75t_R _19284_ (.A(_10806_),
    .Y(_10956_));
 NAND2x1_ASAP7_75t_R _19285_ (.A(_10955_),
    .B(_10956_),
    .Y(_10957_));
 NAND2x1_ASAP7_75t_R _19286_ (.A(_15806_),
    .B(net24),
    .Y(_10958_));
 NAND2x1_ASAP7_75t_R _19287_ (.A(_10729_),
    .B(_10958_),
    .Y(_10959_));
 AOI21x1_ASAP7_75t_R _19288_ (.A1(_10957_),
    .A2(_10959_),
    .B(_10857_),
    .Y(_10960_));
 OAI21x1_ASAP7_75t_R _19289_ (.A1(_10954_),
    .A2(_10960_),
    .B(_10767_),
    .Y(_10961_));
 OAI21x1_ASAP7_75t_R _19290_ (.A1(_10767_),
    .A2(_10949_),
    .B(_10961_),
    .Y(_10962_));
 NAND2x2_ASAP7_75t_R _19291_ (.A(_10769_),
    .B(net784),
    .Y(_10963_));
 NAND2x1_ASAP7_75t_R _19292_ (.A(_10963_),
    .B(net1),
    .Y(_10964_));
 NOR2x1_ASAP7_75t_R _19293_ (.A(_10869_),
    .B(_10795_),
    .Y(_10965_));
 AOI21x1_ASAP7_75t_R _19294_ (.A1(_10842_),
    .A2(_10965_),
    .B(_10817_),
    .Y(_10966_));
 NAND2x1_ASAP7_75t_R _19295_ (.A(_10964_),
    .B(_10966_),
    .Y(_10967_));
 AOI21x1_ASAP7_75t_R _19296_ (.A1(_10927_),
    .A2(_10893_),
    .B(_10778_),
    .Y(_10968_));
 NAND2x1_ASAP7_75t_R _19297_ (.A(_10930_),
    .B(_10839_),
    .Y(_10969_));
 BUFx6f_ASAP7_75t_R _19298_ (.A(_10766_),
    .Y(_10970_));
 AOI21x1_ASAP7_75t_R _19299_ (.A1(_10968_),
    .A2(_10969_),
    .B(_10970_),
    .Y(_10971_));
 NAND2x1_ASAP7_75t_R _19300_ (.A(_10967_),
    .B(_10971_),
    .Y(_10972_));
 AOI21x1_ASAP7_75t_R _19301_ (.A1(_10732_),
    .A2(_10863_),
    .B(_10802_),
    .Y(_10973_));
 NAND2x1_ASAP7_75t_R _19302_ (.A(_10973_),
    .B(_10904_),
    .Y(_10974_));
 OA21x2_ASAP7_75t_R _19303_ (.A1(_10922_),
    .A2(_10869_),
    .B(_10777_),
    .Y(_10975_));
 NOR2x1_ASAP7_75t_R _19304_ (.A(_15814_),
    .B(_15804_),
    .Y(_10976_));
 AOI21x1_ASAP7_75t_R _19305_ (.A1(_10769_),
    .A2(net3),
    .B(_10727_),
    .Y(_10977_));
 NOR2x1_ASAP7_75t_R _19306_ (.A(_10976_),
    .B(_10977_),
    .Y(_10978_));
 AOI21x1_ASAP7_75t_R _19307_ (.A1(_10975_),
    .A2(_10978_),
    .B(_10920_),
    .Y(_10979_));
 NAND2x1_ASAP7_75t_R _19308_ (.A(_10974_),
    .B(_10979_),
    .Y(_10980_));
 AOI21x1_ASAP7_75t_R _19309_ (.A1(_10972_),
    .A2(_10980_),
    .B(_10792_),
    .Y(_10981_));
 AOI21x1_ASAP7_75t_R _19310_ (.A1(_10792_),
    .A2(_10962_),
    .B(_10981_),
    .Y(_10982_));
 OAI21x1_ASAP7_75t_R _19311_ (.A1(net538),
    .A2(_10951_),
    .B(_10870_),
    .Y(_10983_));
 OAI21x1_ASAP7_75t_R _19312_ (.A1(_10770_),
    .A2(_10841_),
    .B(_10913_),
    .Y(_10984_));
 AOI21x1_ASAP7_75t_R _19313_ (.A1(_10983_),
    .A2(_10984_),
    .B(_10953_),
    .Y(_10985_));
 NAND2x2_ASAP7_75t_R _19314_ (.A(_10867_),
    .B(_10796_),
    .Y(_10986_));
 BUFx6f_ASAP7_75t_R _19315_ (.A(_10843_),
    .Y(_10987_));
 OAI21x1_ASAP7_75t_R _19316_ (.A1(_10855_),
    .A2(_10806_),
    .B(_10987_),
    .Y(_10988_));
 AOI21x1_ASAP7_75t_R _19317_ (.A1(_10986_),
    .A2(_10988_),
    .B(_10857_),
    .Y(_10989_));
 OAI21x1_ASAP7_75t_R _19318_ (.A1(_10985_),
    .A2(_10989_),
    .B(_10861_),
    .Y(_10990_));
 NOR2x1_ASAP7_75t_R _19319_ (.A(_10939_),
    .B(_10940_),
    .Y(_10991_));
 AOI21x1_ASAP7_75t_R _19320_ (.A1(_01154_),
    .A2(_10709_),
    .B(_10805_),
    .Y(_10992_));
 AO21x2_ASAP7_75t_R _19321_ (.A1(_10809_),
    .A2(_10810_),
    .B(_10896_),
    .Y(_10993_));
 AO21x1_ASAP7_75t_R _19322_ (.A1(_10992_),
    .A2(_10993_),
    .B(_10953_),
    .Y(_10994_));
 NOR2x1_ASAP7_75t_R _19323_ (.A(_10778_),
    .B(_10815_),
    .Y(_10995_));
 OAI21x1_ASAP7_75t_R _19324_ (.A1(_15814_),
    .A2(_10847_),
    .B(_10800_),
    .Y(_10996_));
 AOI21x1_ASAP7_75t_R _19325_ (.A1(_10995_),
    .A2(_10996_),
    .B(_10920_),
    .Y(_10997_));
 OAI21x1_ASAP7_75t_R _19326_ (.A1(_10991_),
    .A2(_10994_),
    .B(_10997_),
    .Y(_10998_));
 AOI21x1_ASAP7_75t_R _19327_ (.A1(_10990_),
    .A2(_10998_),
    .B(_10884_),
    .Y(_10999_));
 AOI21x1_ASAP7_75t_R _19328_ (.A1(_10944_),
    .A2(_10750_),
    .B(_10987_),
    .Y(_11000_));
 AO21x1_ASAP7_75t_R _19329_ (.A1(_10854_),
    .A2(_15814_),
    .B(_10875_),
    .Y(_11001_));
 OAI21x1_ASAP7_75t_R _19330_ (.A1(_10806_),
    .A2(_11001_),
    .B(_10920_),
    .Y(_11002_));
 INVx1_ASAP7_75t_R _19331_ (.A(_10986_),
    .Y(_11003_));
 NOR2x2_ASAP7_75t_R _19332_ (.A(_10709_),
    .B(net604),
    .Y(_11004_));
 INVx1_ASAP7_75t_R _19333_ (.A(_10837_),
    .Y(_11005_));
 OAI21x1_ASAP7_75t_R _19334_ (.A1(_11004_),
    .A2(_11005_),
    .B(_10766_),
    .Y(_11006_));
 OAI22x1_ASAP7_75t_R _19335_ (.A1(_11000_),
    .A2(_11002_),
    .B1(_11003_),
    .B2(_11006_),
    .Y(_11007_));
 INVx1_ASAP7_75t_R _19336_ (.A(_00495_),
    .Y(_11008_));
 NOR2x1_ASAP7_75t_R _19337_ (.A(_11008_),
    .B(_10879_),
    .Y(_11009_));
 AO21x1_ASAP7_75t_R _19338_ (.A1(_10766_),
    .A2(_11009_),
    .B(_10934_),
    .Y(_11010_));
 NAND2x2_ASAP7_75t_R _19339_ (.A(_15806_),
    .B(_10708_),
    .Y(_11011_));
 NOR2x2_ASAP7_75t_R _19340_ (.A(net24),
    .B(_11011_),
    .Y(_11012_));
 NOR2x1_ASAP7_75t_R _19341_ (.A(_10890_),
    .B(_11012_),
    .Y(_11013_));
 OAI21x1_ASAP7_75t_R _19342_ (.A1(_11010_),
    .A2(_11013_),
    .B(_10884_),
    .Y(_11014_));
 AOI21x1_ASAP7_75t_R _19343_ (.A1(_10803_),
    .A2(_11007_),
    .B(_11014_),
    .Y(_11015_));
 OAI21x1_ASAP7_75t_R _19344_ (.A1(_10999_),
    .A2(_11015_),
    .B(_10835_),
    .Y(_11016_));
 OAI21x1_ASAP7_75t_R _19345_ (.A1(_10835_),
    .A2(_10982_),
    .B(_11016_),
    .Y(_00033_));
 AO21x2_ASAP7_75t_R _19346_ (.A1(_10700_),
    .A2(_10810_),
    .B(_10794_),
    .Y(_11017_));
 OA21x2_ASAP7_75t_R _19347_ (.A1(_15804_),
    .A2(_10769_),
    .B(_10805_),
    .Y(_11018_));
 NAND2x1_ASAP7_75t_R _19348_ (.A(_10953_),
    .B(_10918_),
    .Y(_11019_));
 AO21x1_ASAP7_75t_R _19349_ (.A1(_11017_),
    .A2(_11018_),
    .B(_11019_),
    .Y(_11020_));
 NAND2x2_ASAP7_75t_R _19350_ (.A(_10805_),
    .B(_11017_),
    .Y(_11021_));
 OAI21x1_ASAP7_75t_R _19351_ (.A1(_10806_),
    .A2(_11021_),
    .B(_10857_),
    .Y(_11022_));
 AOI21x1_ASAP7_75t_R _19352_ (.A1(_10810_),
    .A2(_10809_),
    .B(_01154_),
    .Y(_11023_));
 OA21x2_ASAP7_75t_R _19353_ (.A1(_10917_),
    .A2(_11023_),
    .B(_10913_),
    .Y(_11024_));
 OA21x2_ASAP7_75t_R _19354_ (.A1(_11022_),
    .A2(_11024_),
    .B(_10899_),
    .Y(_11025_));
 AO21x2_ASAP7_75t_R _19355_ (.A1(_10707_),
    .A2(_10705_),
    .B(_01153_),
    .Y(_11026_));
 NAND2x1_ASAP7_75t_R _19356_ (.A(_10752_),
    .B(_11026_),
    .Y(_11027_));
 NOR2x2_ASAP7_75t_R _19357_ (.A(_10752_),
    .B(_11023_),
    .Y(_11028_));
 AOI21x1_ASAP7_75t_R _19358_ (.A1(_11011_),
    .A2(_11028_),
    .B(_10747_),
    .Y(_11029_));
 OAI21x1_ASAP7_75t_R _19359_ (.A1(_10771_),
    .A2(_11027_),
    .B(_11029_),
    .Y(_11030_));
 AND2x2_ASAP7_75t_R _19360_ (.A(_10815_),
    .B(_10929_),
    .Y(_11031_));
 AOI21x1_ASAP7_75t_R _19361_ (.A1(_01153_),
    .A2(_10769_),
    .B(_10805_),
    .Y(_11032_));
 INVx1_ASAP7_75t_R _19362_ (.A(_11032_),
    .Y(_11033_));
 NOR2x2_ASAP7_75t_R _19363_ (.A(_10806_),
    .B(_11033_),
    .Y(_11034_));
 OAI21x1_ASAP7_75t_R _19364_ (.A1(_11031_),
    .A2(_11034_),
    .B(_10818_),
    .Y(_11035_));
 AOI21x1_ASAP7_75t_R _19365_ (.A1(_11035_),
    .A2(_11030_),
    .B(_10767_),
    .Y(_11036_));
 AOI211x1_ASAP7_75t_R _19366_ (.A1(_11020_),
    .A2(_11025_),
    .B(_10884_),
    .C(_11036_),
    .Y(_11037_));
 INVx1_ASAP7_75t_R _19367_ (.A(_10940_),
    .Y(_11038_));
 OAI21x1_ASAP7_75t_R _19368_ (.A1(net24),
    .A2(_10963_),
    .B(_10879_),
    .Y(_11039_));
 NAND2x1_ASAP7_75t_R _19369_ (.A(_10747_),
    .B(_11039_),
    .Y(_11040_));
 AOI21x1_ASAP7_75t_R _19370_ (.A1(_10732_),
    .A2(_11038_),
    .B(_11040_),
    .Y(_11041_));
 OA21x2_ASAP7_75t_R _19371_ (.A1(_10709_),
    .A2(_01151_),
    .B(_10869_),
    .Y(_11042_));
 OA21x2_ASAP7_75t_R _19372_ (.A1(_10701_),
    .A2(_00494_),
    .B(_10727_),
    .Y(_11043_));
 AOI22x1_ASAP7_75t_R _19373_ (.A1(_11042_),
    .A2(_11011_),
    .B1(_11043_),
    .B2(_10867_),
    .Y(_11044_));
 OAI21x1_ASAP7_75t_R _19374_ (.A1(_10818_),
    .A2(_11044_),
    .B(_10861_),
    .Y(_11045_));
 NOR2x1_ASAP7_75t_R _19375_ (.A(_11041_),
    .B(_11045_),
    .Y(_11046_));
 INVx1_ASAP7_75t_R _19376_ (.A(_10749_),
    .Y(_11047_));
 INVx1_ASAP7_75t_R _19377_ (.A(_10844_),
    .Y(_11048_));
 OAI21x1_ASAP7_75t_R _19378_ (.A1(_11023_),
    .A2(_10941_),
    .B(_10879_),
    .Y(_11049_));
 OAI21x1_ASAP7_75t_R _19379_ (.A1(_11047_),
    .A2(_11048_),
    .B(_11049_),
    .Y(_11050_));
 NOR2x1_ASAP7_75t_R _19380_ (.A(_10728_),
    .B(_10902_),
    .Y(_11051_));
 INVx1_ASAP7_75t_R _19381_ (.A(_10903_),
    .Y(_11052_));
 AOI21x1_ASAP7_75t_R _19382_ (.A1(_11051_),
    .A2(_11052_),
    .B(_10778_),
    .Y(_11053_));
 AOI22x1_ASAP7_75t_R _19383_ (.A1(_11050_),
    .A2(_10803_),
    .B1(_11053_),
    .B2(_10931_),
    .Y(_11054_));
 OAI21x1_ASAP7_75t_R _19384_ (.A1(_10861_),
    .A2(_11054_),
    .B(_10884_),
    .Y(_11055_));
 OAI21x1_ASAP7_75t_R _19385_ (.A1(_11046_),
    .A2(_11055_),
    .B(_10835_),
    .Y(_11056_));
 OAI21x1_ASAP7_75t_R _19386_ (.A1(_10926_),
    .A2(_10927_),
    .B(_10867_),
    .Y(_11057_));
 AOI21x1_ASAP7_75t_R _19387_ (.A1(_10929_),
    .A2(_10930_),
    .B(_10817_),
    .Y(_11058_));
 NAND2x1_ASAP7_75t_R _19388_ (.A(_11057_),
    .B(_11058_),
    .Y(_11059_));
 OA21x2_ASAP7_75t_R _19389_ (.A1(_01156_),
    .A2(_10875_),
    .B(_10907_),
    .Y(_11060_));
 OAI21x1_ASAP7_75t_R _19390_ (.A1(_15814_),
    .A2(_10893_),
    .B(_10863_),
    .Y(_11061_));
 AOI21x1_ASAP7_75t_R _19391_ (.A1(_11060_),
    .A2(_11061_),
    .B(_10899_),
    .Y(_11062_));
 AOI21x1_ASAP7_75t_R _19392_ (.A1(_11059_),
    .A2(_11062_),
    .B(_10883_),
    .Y(_11063_));
 NOR3x1_ASAP7_75t_R _19393_ (.A(_10853_),
    .B(_10879_),
    .C(net537),
    .Y(_11064_));
 AND2x2_ASAP7_75t_R _19394_ (.A(_10930_),
    .B(_10878_),
    .Y(_11065_));
 OAI21x1_ASAP7_75t_R _19395_ (.A1(_11064_),
    .A2(_11065_),
    .B(_10857_),
    .Y(_11066_));
 AOI21x1_ASAP7_75t_R _19396_ (.A1(_15801_),
    .A2(net604),
    .B(_10843_),
    .Y(_11067_));
 NOR2x1_ASAP7_75t_R _19397_ (.A(_11008_),
    .B(_10752_),
    .Y(_11068_));
 AOI21x1_ASAP7_75t_R _19398_ (.A1(_10749_),
    .A2(_11067_),
    .B(_11068_),
    .Y(_11069_));
 AOI21x1_ASAP7_75t_R _19399_ (.A1(_10953_),
    .A2(_11069_),
    .B(_10860_),
    .Y(_11070_));
 NAND2x1_ASAP7_75t_R _19400_ (.A(_11066_),
    .B(_11070_),
    .Y(_11071_));
 AOI21x1_ASAP7_75t_R _19401_ (.A1(_11063_),
    .A2(_11071_),
    .B(_10834_),
    .Y(_11072_));
 OA21x2_ASAP7_75t_R _19402_ (.A1(_10875_),
    .A2(_10873_),
    .B(_10860_),
    .Y(_11073_));
 NAND2x1_ASAP7_75t_R _19403_ (.A(_11017_),
    .B(net1),
    .Y(_11074_));
 AO21x1_ASAP7_75t_R _19404_ (.A1(_11073_),
    .A2(_11074_),
    .B(_10803_),
    .Y(_11075_));
 INVx1_ASAP7_75t_R _19405_ (.A(_00496_),
    .Y(_11076_));
 OA211x2_ASAP7_75t_R _19406_ (.A1(_11076_),
    .A2(_10987_),
    .B(_11039_),
    .C(_10970_),
    .Y(_11077_));
 NAND2x1_ASAP7_75t_R _19407_ (.A(_10749_),
    .B(_10844_),
    .Y(_11078_));
 OA21x2_ASAP7_75t_R _19408_ (.A1(_01158_),
    .A2(_10875_),
    .B(_10766_),
    .Y(_11079_));
 AOI21x1_ASAP7_75t_R _19409_ (.A1(_11078_),
    .A2(_11079_),
    .B(_10953_),
    .Y(_11080_));
 AND2x2_ASAP7_75t_R _19410_ (.A(_01152_),
    .B(_01151_),
    .Y(_11081_));
 INVx1_ASAP7_75t_R _19411_ (.A(_11081_),
    .Y(_11082_));
 NOR2x2_ASAP7_75t_R _19412_ (.A(_11082_),
    .B(_10701_),
    .Y(_11083_));
 NOR2x2_ASAP7_75t_R _19413_ (.A(_10728_),
    .B(_11083_),
    .Y(_11084_));
 OAI21x1_ASAP7_75t_R _19414_ (.A1(_15811_),
    .A2(_10847_),
    .B(_11084_),
    .Y(_11085_));
 OA21x2_ASAP7_75t_R _19415_ (.A1(_10709_),
    .A2(_00491_),
    .B(_10728_),
    .Y(_11086_));
 AOI21x1_ASAP7_75t_R _19416_ (.A1(_11086_),
    .A2(_10775_),
    .B(_10766_),
    .Y(_11087_));
 NAND2x1_ASAP7_75t_R _19417_ (.A(_11085_),
    .B(_11087_),
    .Y(_11088_));
 AOI21x1_ASAP7_75t_R _19418_ (.A1(_11080_),
    .A2(_11088_),
    .B(_10791_),
    .Y(_11089_));
 OAI21x1_ASAP7_75t_R _19419_ (.A1(_11075_),
    .A2(_11077_),
    .B(_11089_),
    .Y(_11090_));
 NAND2x1_ASAP7_75t_R _19420_ (.A(_11072_),
    .B(_11090_),
    .Y(_11091_));
 OAI21x1_ASAP7_75t_R _19421_ (.A1(_11056_),
    .A2(_11037_),
    .B(_11091_),
    .Y(_00034_));
 AO21x1_ASAP7_75t_R _19422_ (.A1(_10963_),
    .A2(_11026_),
    .B(_10728_),
    .Y(_11092_));
 NAND2x1_ASAP7_75t_R _19423_ (.A(_10812_),
    .B(_10849_),
    .Y(_11093_));
 AO21x1_ASAP7_75t_R _19424_ (.A1(_11092_),
    .A2(_11093_),
    .B(_10953_),
    .Y(_11094_));
 AO21x1_ASAP7_75t_R _19425_ (.A1(_10842_),
    .A2(_10873_),
    .B(_10913_),
    .Y(_11095_));
 AO21x1_ASAP7_75t_R _19426_ (.A1(_11095_),
    .A2(_10969_),
    .B(_10857_),
    .Y(_11096_));
 AOI21x1_ASAP7_75t_R _19427_ (.A1(_11094_),
    .A2(_11096_),
    .B(_10767_),
    .Y(_11097_));
 INVx1_ASAP7_75t_R _19428_ (.A(_10894_),
    .Y(_11098_));
 OAI22x1_ASAP7_75t_R _19429_ (.A1(_11012_),
    .A2(_10890_),
    .B1(_11098_),
    .B2(_11083_),
    .Y(_11099_));
 AOI21x1_ASAP7_75t_R _19430_ (.A1(_10818_),
    .A2(_11099_),
    .B(_11029_),
    .Y(_11100_));
 OAI21x1_ASAP7_75t_R _19431_ (.A1(_10861_),
    .A2(_11100_),
    .B(_10792_),
    .Y(_11101_));
 NOR2x1_ASAP7_75t_R _19432_ (.A(_11097_),
    .B(_11101_),
    .Y(_11102_));
 AO21x1_ASAP7_75t_R _19433_ (.A1(_10870_),
    .A2(_10917_),
    .B(_10766_),
    .Y(_11103_));
 OAI21x1_ASAP7_75t_R _19434_ (.A1(_11034_),
    .A2(_11103_),
    .B(_10818_),
    .Y(_11104_));
 NOR2x1_ASAP7_75t_R _19435_ (.A(net488),
    .B(_10801_),
    .Y(_11105_));
 AOI211x1_ASAP7_75t_R _19436_ (.A1(_10812_),
    .A2(_11084_),
    .B(_11105_),
    .C(_10861_),
    .Y(_11106_));
 NOR2x1_ASAP7_75t_R _19437_ (.A(_11104_),
    .B(_11106_),
    .Y(_11107_));
 AO21x1_ASAP7_75t_R _19438_ (.A1(_10749_),
    .A2(_10889_),
    .B(_10753_),
    .Y(_11108_));
 NOR2x1_ASAP7_75t_R _19439_ (.A(_10863_),
    .B(_10920_),
    .Y(_11109_));
 NAND2x1_ASAP7_75t_R _19440_ (.A(_10843_),
    .B(net486),
    .Y(_11110_));
 OAI21x1_ASAP7_75t_R _19441_ (.A1(_10899_),
    .A2(_11110_),
    .B(_10891_),
    .Y(_11111_));
 AOI21x1_ASAP7_75t_R _19442_ (.A1(_11108_),
    .A2(_11109_),
    .B(_11111_),
    .Y(_11112_));
 OAI21x1_ASAP7_75t_R _19443_ (.A1(_10818_),
    .A2(_11112_),
    .B(_10884_),
    .Y(_11113_));
 OAI21x1_ASAP7_75t_R _19444_ (.A1(_11107_),
    .A2(_11113_),
    .B(_10835_),
    .Y(_11114_));
 NOR2x1_ASAP7_75t_R _19445_ (.A(_10853_),
    .B(_10841_),
    .Y(_11115_));
 NOR2x2_ASAP7_75t_R _19446_ (.A(_10843_),
    .B(_10771_),
    .Y(_11116_));
 NAND2x1_ASAP7_75t_R _19447_ (.A(_11115_),
    .B(_11116_),
    .Y(_11117_));
 AOI21x1_ASAP7_75t_R _19448_ (.A1(_10955_),
    .A2(_10944_),
    .B(_10934_),
    .Y(_11118_));
 AOI21x1_ASAP7_75t_R _19449_ (.A1(_10874_),
    .A2(_10849_),
    .B(_10953_),
    .Y(_11119_));
 AOI22x1_ASAP7_75t_R _19450_ (.A1(_11117_),
    .A2(_11118_),
    .B1(_10845_),
    .B2(_11119_),
    .Y(_11120_));
 AND3x1_ASAP7_75t_R _19451_ (.A(_10707_),
    .B(_10705_),
    .C(_01153_),
    .Y(_11121_));
 INVx2_ASAP7_75t_R _19452_ (.A(_11043_),
    .Y(_11122_));
 OAI21x1_ASAP7_75t_R _19453_ (.A1(_11121_),
    .A2(_11122_),
    .B(_10947_),
    .Y(_11123_));
 NAND2x1_ASAP7_75t_R _19454_ (.A(_10709_),
    .B(_10869_),
    .Y(_11124_));
 AOI211x1_ASAP7_75t_R _19455_ (.A1(net24),
    .A2(net65),
    .B(_10841_),
    .C(_10777_),
    .Y(_11125_));
 AOI21x1_ASAP7_75t_R _19456_ (.A1(_11124_),
    .A2(_11125_),
    .B(_10920_),
    .Y(_11126_));
 AOI21x1_ASAP7_75t_R _19457_ (.A1(_11123_),
    .A2(_11126_),
    .B(_10884_),
    .Y(_11127_));
 OAI21x1_ASAP7_75t_R _19458_ (.A1(_10767_),
    .A2(_11120_),
    .B(_11127_),
    .Y(_11128_));
 AND2x2_ASAP7_75t_R _19459_ (.A(_10873_),
    .B(_10863_),
    .Y(_11129_));
 NOR3x1_ASAP7_75t_R _19460_ (.A(_10841_),
    .B(_10853_),
    .C(_10875_),
    .Y(_11130_));
 OAI21x1_ASAP7_75t_R _19461_ (.A1(_11129_),
    .A2(_11130_),
    .B(_10857_),
    .Y(_11131_));
 INVx1_ASAP7_75t_R _19462_ (.A(_11021_),
    .Y(_11132_));
 NAND2x1_ASAP7_75t_R _19463_ (.A(_10732_),
    .B(_11132_),
    .Y(_11133_));
 AOI21x1_ASAP7_75t_R _19464_ (.A1(_10867_),
    .A2(_11043_),
    .B(_10778_),
    .Y(_11134_));
 AOI21x1_ASAP7_75t_R _19465_ (.A1(_11133_),
    .A2(_11134_),
    .B(_10970_),
    .Y(_11135_));
 NAND2x1_ASAP7_75t_R _19466_ (.A(_11131_),
    .B(_11135_),
    .Y(_11136_));
 NAND2x1_ASAP7_75t_R _19467_ (.A(_10893_),
    .B(_10837_),
    .Y(_11137_));
 AOI21x1_ASAP7_75t_R _19468_ (.A1(_10867_),
    .A2(net1),
    .B(_10778_),
    .Y(_11138_));
 NAND2x1_ASAP7_75t_R _19469_ (.A(_11138_),
    .B(_11137_),
    .Y(_11139_));
 OAI21x1_ASAP7_75t_R _19470_ (.A1(_10774_),
    .A2(_11004_),
    .B(_10987_),
    .Y(_11140_));
 AOI21x1_ASAP7_75t_R _19471_ (.A1(_10864_),
    .A2(_11140_),
    .B(_10920_),
    .Y(_11141_));
 AOI21x1_ASAP7_75t_R _19472_ (.A1(_11141_),
    .A2(_11139_),
    .B(_10792_),
    .Y(_11142_));
 AOI21x1_ASAP7_75t_R _19473_ (.A1(_11142_),
    .A2(_11136_),
    .B(_10835_),
    .Y(_11143_));
 NAND2x1_ASAP7_75t_R _19474_ (.A(_11143_),
    .B(_11128_),
    .Y(_11144_));
 OAI21x1_ASAP7_75t_R _19475_ (.A1(_11102_),
    .A2(_11114_),
    .B(_11144_),
    .Y(_00035_));
 INVx1_ASAP7_75t_R _19476_ (.A(_10862_),
    .Y(_11145_));
 AOI21x1_ASAP7_75t_R _19477_ (.A1(_11145_),
    .A2(_10992_),
    .B(_10802_),
    .Y(_11146_));
 NAND2x1_ASAP7_75t_R _19478_ (.A(_10895_),
    .B(_11146_),
    .Y(_11147_));
 NAND2x2_ASAP7_75t_R _19479_ (.A(_10751_),
    .B(net538),
    .Y(_11148_));
 AND2x2_ASAP7_75t_R _19480_ (.A(_11026_),
    .B(_11148_),
    .Y(_11149_));
 AOI21x1_ASAP7_75t_R _19481_ (.A1(_10975_),
    .A2(_11149_),
    .B(_10970_),
    .Y(_11150_));
 AOI21x1_ASAP7_75t_R _19482_ (.A1(_11147_),
    .A2(_11150_),
    .B(_10791_),
    .Y(_11151_));
 OAI21x1_ASAP7_75t_R _19483_ (.A1(_10951_),
    .A2(_11004_),
    .B(_10870_),
    .Y(_11152_));
 AOI21x1_ASAP7_75t_R _19484_ (.A1(_10904_),
    .A2(_11152_),
    .B(_10934_),
    .Y(_11153_));
 OAI21x1_ASAP7_75t_R _19485_ (.A1(_10903_),
    .A2(_11004_),
    .B(_10870_),
    .Y(_11154_));
 AOI21x1_ASAP7_75t_R _19486_ (.A1(_11049_),
    .A2(_11154_),
    .B(_10953_),
    .Y(_11155_));
 OAI21x1_ASAP7_75t_R _19487_ (.A1(_11153_),
    .A2(_11155_),
    .B(_10899_),
    .Y(_11156_));
 AOI21x1_ASAP7_75t_R _19488_ (.A1(_11151_),
    .A2(_11156_),
    .B(_10834_),
    .Y(_11157_));
 AO21x1_ASAP7_75t_R _19489_ (.A1(net24),
    .A2(_15811_),
    .B(_10869_),
    .Y(_11158_));
 NOR2x1_ASAP7_75t_R _19490_ (.A(_10907_),
    .B(_10860_),
    .Y(_11159_));
 OAI21x1_ASAP7_75t_R _19491_ (.A1(_10848_),
    .A2(_11158_),
    .B(_11159_),
    .Y(_11160_));
 AO21x1_ASAP7_75t_R _19492_ (.A1(_10809_),
    .A2(_10810_),
    .B(_00493_),
    .Y(_11161_));
 AND2x2_ASAP7_75t_R _19493_ (.A(_11018_),
    .B(_11161_),
    .Y(_11162_));
 AO21x1_ASAP7_75t_R _19494_ (.A1(_11067_),
    .A2(_10749_),
    .B(_10802_),
    .Y(_11163_));
 OAI22x1_ASAP7_75t_R _19495_ (.A1(_11160_),
    .A2(_11162_),
    .B1(_11163_),
    .B2(_11006_),
    .Y(_11164_));
 OR3x1_ASAP7_75t_R _19496_ (.A(_10894_),
    .B(_10770_),
    .C(_10817_),
    .Y(_11165_));
 NAND2x1_ASAP7_75t_R _19497_ (.A(_10956_),
    .B(_10977_),
    .Y(_11166_));
 AOI21x1_ASAP7_75t_R _19498_ (.A1(_11161_),
    .A2(_10807_),
    .B(_10802_),
    .Y(_11167_));
 NAND2x1_ASAP7_75t_R _19499_ (.A(_11166_),
    .B(_11167_),
    .Y(_11168_));
 AOI21x1_ASAP7_75t_R _19500_ (.A1(_11165_),
    .A2(_11168_),
    .B(_10899_),
    .Y(_11169_));
 OAI21x1_ASAP7_75t_R _19501_ (.A1(_11164_),
    .A2(_11169_),
    .B(_10792_),
    .Y(_11170_));
 NAND2x1_ASAP7_75t_R _19502_ (.A(_11157_),
    .B(_11170_),
    .Y(_11171_));
 AO21x1_ASAP7_75t_R _19503_ (.A1(_10951_),
    .A2(_10843_),
    .B(_10746_),
    .Y(_11172_));
 OAI21x1_ASAP7_75t_R _19504_ (.A1(_10753_),
    .A2(_10867_),
    .B(_10986_),
    .Y(_11173_));
 NOR2x1_ASAP7_75t_R _19505_ (.A(_10802_),
    .B(_10927_),
    .Y(_11174_));
 NAND2x1_ASAP7_75t_R _19506_ (.A(_10812_),
    .B(_10837_),
    .Y(_11175_));
 AOI21x1_ASAP7_75t_R _19507_ (.A1(_11174_),
    .A2(_11175_),
    .B(_10860_),
    .Y(_11176_));
 OAI21x1_ASAP7_75t_R _19508_ (.A1(_11172_),
    .A2(_11173_),
    .B(_11176_),
    .Y(_11177_));
 INVx1_ASAP7_75t_R _19509_ (.A(_10965_),
    .Y(_11178_));
 NOR2x1_ASAP7_75t_R _19510_ (.A(net538),
    .B(_11178_),
    .Y(_11179_));
 AOI21x1_ASAP7_75t_R _19511_ (.A1(_10913_),
    .A2(_10993_),
    .B(_10817_),
    .Y(_11180_));
 AOI21x1_ASAP7_75t_R _19512_ (.A1(_11180_),
    .A2(_10940_),
    .B(_10970_),
    .Y(_11181_));
 OAI21x1_ASAP7_75t_R _19513_ (.A1(_11179_),
    .A2(_10779_),
    .B(_11181_),
    .Y(_11182_));
 AOI21x1_ASAP7_75t_R _19514_ (.A1(_11177_),
    .A2(_11182_),
    .B(_10884_),
    .Y(_11183_));
 NAND2x1_ASAP7_75t_R _19515_ (.A(_10879_),
    .B(_10903_),
    .Y(_11184_));
 NAND2x2_ASAP7_75t_R _19516_ (.A(_10894_),
    .B(_10946_),
    .Y(_11185_));
 AOI21x1_ASAP7_75t_R _19517_ (.A1(_11184_),
    .A2(_11185_),
    .B(_10953_),
    .Y(_11186_));
 OA21x2_ASAP7_75t_R _19518_ (.A1(_00497_),
    .A2(_10869_),
    .B(_10746_),
    .Y(_11187_));
 AO21x1_ASAP7_75t_R _19519_ (.A1(_11187_),
    .A2(_11148_),
    .B(_10766_),
    .Y(_11188_));
 OAI21x1_ASAP7_75t_R _19520_ (.A1(_11186_),
    .A2(_11188_),
    .B(_10883_),
    .Y(_11189_));
 NAND2x1_ASAP7_75t_R _19521_ (.A(_11011_),
    .B(_10894_),
    .Y(_11190_));
 AO21x1_ASAP7_75t_R _19522_ (.A1(_10946_),
    .A2(_10847_),
    .B(_10752_),
    .Y(_11191_));
 AOI21x1_ASAP7_75t_R _19523_ (.A1(_11190_),
    .A2(_11191_),
    .B(_10747_),
    .Y(_11192_));
 AOI21x1_ASAP7_75t_R _19524_ (.A1(_10842_),
    .A2(_10844_),
    .B(_10933_),
    .Y(_11193_));
 OAI21x1_ASAP7_75t_R _19525_ (.A1(_10934_),
    .A2(_11193_),
    .B(_10970_),
    .Y(_11194_));
 NOR2x1_ASAP7_75t_R _19526_ (.A(_11192_),
    .B(_11194_),
    .Y(_11195_));
 NOR2x1_ASAP7_75t_R _19527_ (.A(_11189_),
    .B(_11195_),
    .Y(_11196_));
 OAI21x1_ASAP7_75t_R _19528_ (.A1(_11183_),
    .A2(_11196_),
    .B(_10835_),
    .Y(_11197_));
 NAND2x1_ASAP7_75t_R _19529_ (.A(_11197_),
    .B(_11171_),
    .Y(_00036_));
 NAND2x1_ASAP7_75t_R _19530_ (.A(_10913_),
    .B(_10993_),
    .Y(_11198_));
 OAI21x1_ASAP7_75t_R _19531_ (.A1(_11047_),
    .A2(_11198_),
    .B(_11148_),
    .Y(_11199_));
 AOI211x1_ASAP7_75t_R _19532_ (.A1(net1),
    .A2(_10878_),
    .B(_11028_),
    .C(_10934_),
    .Y(_11200_));
 AOI21x1_ASAP7_75t_R _19533_ (.A1(_10803_),
    .A2(_11199_),
    .B(_11200_),
    .Y(_11201_));
 AOI21x1_ASAP7_75t_R _19534_ (.A1(_10927_),
    .A2(_10893_),
    .B(_10817_),
    .Y(_11202_));
 NAND2x1_ASAP7_75t_R _19535_ (.A(_11178_),
    .B(_11202_),
    .Y(_11203_));
 NOR2x1_ASAP7_75t_R _19536_ (.A(_10802_),
    .B(_10849_),
    .Y(_11204_));
 AOI21x1_ASAP7_75t_R _19537_ (.A1(_11204_),
    .A2(_11092_),
    .B(_10883_),
    .Y(_11205_));
 NAND2x1_ASAP7_75t_R _19538_ (.A(_11203_),
    .B(_11205_),
    .Y(_11206_));
 OAI21x1_ASAP7_75t_R _19539_ (.A1(_10792_),
    .A2(_11201_),
    .B(_11206_),
    .Y(_11207_));
 AOI21x1_ASAP7_75t_R _19540_ (.A1(_10767_),
    .A2(_11207_),
    .B(_10835_),
    .Y(_11208_));
 NAND2x1_ASAP7_75t_R _19541_ (.A(_10812_),
    .B(_10796_),
    .Y(_11209_));
 OAI21x1_ASAP7_75t_R _19542_ (.A1(_10753_),
    .A2(_10772_),
    .B(_11209_),
    .Y(_11210_));
 OAI21x1_ASAP7_75t_R _19543_ (.A1(_10803_),
    .A2(_11210_),
    .B(_10791_),
    .Y(_11211_));
 OA21x2_ASAP7_75t_R _19544_ (.A1(_11021_),
    .A2(_11081_),
    .B(_10778_),
    .Y(_11212_));
 OA21x2_ASAP7_75t_R _19545_ (.A1(_10888_),
    .A2(_11033_),
    .B(_11212_),
    .Y(_11213_));
 NOR2x1_ASAP7_75t_R _19546_ (.A(_11211_),
    .B(_11213_),
    .Y(_11214_));
 AO21x1_ASAP7_75t_R _19547_ (.A1(_10775_),
    .A2(_10889_),
    .B(_10987_),
    .Y(_11215_));
 OAI21x1_ASAP7_75t_R _19548_ (.A1(_10848_),
    .A2(_10801_),
    .B(_11215_),
    .Y(_11216_));
 AO21x1_ASAP7_75t_R _19549_ (.A1(_10893_),
    .A2(_10867_),
    .B(_10870_),
    .Y(_11217_));
 OA21x2_ASAP7_75t_R _19550_ (.A1(net24),
    .A2(_10879_),
    .B(_10817_),
    .Y(_11218_));
 AO21x1_ASAP7_75t_R _19551_ (.A1(_11217_),
    .A2(_11218_),
    .B(_10791_),
    .Y(_11219_));
 AOI21x1_ASAP7_75t_R _19552_ (.A1(_10803_),
    .A2(_11216_),
    .B(_11219_),
    .Y(_11220_));
 OAI21x1_ASAP7_75t_R _19553_ (.A1(_11214_),
    .A2(_11220_),
    .B(_10861_),
    .Y(_11221_));
 AND2x2_ASAP7_75t_R _19554_ (.A(_10815_),
    .B(_10889_),
    .Y(_11222_));
 AO21x1_ASAP7_75t_R _19555_ (.A1(_11043_),
    .A2(_10812_),
    .B(_10747_),
    .Y(_11223_));
 OA21x2_ASAP7_75t_R _19556_ (.A1(_10852_),
    .A2(_10728_),
    .B(_10907_),
    .Y(_11224_));
 NOR2x2_ASAP7_75t_R _19557_ (.A(_15806_),
    .B(_10805_),
    .Y(_11225_));
 NOR2x1_ASAP7_75t_R _19558_ (.A(_11225_),
    .B(_10930_),
    .Y(_11226_));
 AOI21x1_ASAP7_75t_R _19559_ (.A1(_11224_),
    .A2(_11226_),
    .B(_10860_),
    .Y(_11227_));
 OAI21x1_ASAP7_75t_R _19560_ (.A1(_11222_),
    .A2(_11223_),
    .B(_11227_),
    .Y(_11228_));
 INVx1_ASAP7_75t_R _19561_ (.A(_10945_),
    .Y(_11229_));
 AOI21x1_ASAP7_75t_R _19562_ (.A1(_11229_),
    .A2(_10975_),
    .B(_10970_),
    .Y(_11230_));
 INVx1_ASAP7_75t_R _19563_ (.A(_11083_),
    .Y(_11231_));
 AOI21x1_ASAP7_75t_R _19564_ (.A1(_10870_),
    .A2(_11231_),
    .B(_10778_),
    .Y(_11232_));
 OAI21x1_ASAP7_75t_R _19565_ (.A1(_11012_),
    .A2(_11039_),
    .B(_11232_),
    .Y(_11233_));
 AOI21x1_ASAP7_75t_R _19566_ (.A1(_11230_),
    .A2(_11233_),
    .B(_10791_),
    .Y(_11234_));
 NAND2x1_ASAP7_75t_R _19567_ (.A(_11228_),
    .B(_11234_),
    .Y(_11235_));
 OAI21x1_ASAP7_75t_R _19568_ (.A1(_15811_),
    .A2(_10893_),
    .B(_10815_),
    .Y(_11236_));
 AOI21x1_ASAP7_75t_R _19569_ (.A1(_11032_),
    .A2(_10946_),
    .B(_10817_),
    .Y(_11237_));
 NAND2x1_ASAP7_75t_R _19570_ (.A(_11237_),
    .B(_11236_),
    .Y(_11238_));
 NOR2x1_ASAP7_75t_R _19571_ (.A(_10802_),
    .B(_10926_),
    .Y(_11239_));
 AOI21x1_ASAP7_75t_R _19572_ (.A1(_11239_),
    .A2(_10840_),
    .B(_10970_),
    .Y(_11240_));
 AOI21x1_ASAP7_75t_R _19573_ (.A1(_11238_),
    .A2(_11240_),
    .B(_10883_),
    .Y(_11241_));
 NOR2x1_ASAP7_75t_R _19574_ (.A(_10752_),
    .B(_11011_),
    .Y(_11242_));
 OA21x2_ASAP7_75t_R _19575_ (.A1(_10874_),
    .A2(_10728_),
    .B(_10777_),
    .Y(_11243_));
 OAI21x1_ASAP7_75t_R _19576_ (.A1(_11225_),
    .A2(_10930_),
    .B(_10812_),
    .Y(_11244_));
 AOI21x1_ASAP7_75t_R _19577_ (.A1(_11243_),
    .A2(_11244_),
    .B(_10860_),
    .Y(_11245_));
 OAI21x1_ASAP7_75t_R _19578_ (.A1(_10924_),
    .A2(_11242_),
    .B(_11245_),
    .Y(_11246_));
 NAND2x1_ASAP7_75t_R _19579_ (.A(_11246_),
    .B(_11241_),
    .Y(_11247_));
 INVx2_ASAP7_75t_R _19580_ (.A(_10834_),
    .Y(_11248_));
 AOI21x1_ASAP7_75t_R _19581_ (.A1(_11235_),
    .A2(_11247_),
    .B(_11248_),
    .Y(_11249_));
 AOI21x1_ASAP7_75t_R _19582_ (.A1(_11208_),
    .A2(_11221_),
    .B(_11249_),
    .Y(_00037_));
 AOI21x1_ASAP7_75t_R _19583_ (.A1(_10890_),
    .A2(_11185_),
    .B(_10747_),
    .Y(_11250_));
 OAI21x1_ASAP7_75t_R _19584_ (.A1(_11053_),
    .A2(_11250_),
    .B(_10883_),
    .Y(_11251_));
 NOR2x1_ASAP7_75t_R _19585_ (.A(_10907_),
    .B(_10977_),
    .Y(_11252_));
 AOI21x1_ASAP7_75t_R _19586_ (.A1(_11252_),
    .A2(_10808_),
    .B(_10883_),
    .Y(_11253_));
 AO21x1_ASAP7_75t_R _19587_ (.A1(_10927_),
    .A2(net65),
    .B(_10777_),
    .Y(_11254_));
 AO21x1_ASAP7_75t_R _19588_ (.A1(_11027_),
    .A2(_11122_),
    .B(_11254_),
    .Y(_11255_));
 AOI21x1_ASAP7_75t_R _19589_ (.A1(_11253_),
    .A2(_11255_),
    .B(_10920_),
    .Y(_11256_));
 NAND2x1_ASAP7_75t_R _19590_ (.A(_11251_),
    .B(_11256_),
    .Y(_11257_));
 OAI21x1_ASAP7_75t_R _19591_ (.A1(_10992_),
    .A2(_11067_),
    .B(_10842_),
    .Y(_11258_));
 NAND2x1_ASAP7_75t_R _19592_ (.A(_10934_),
    .B(_11258_),
    .Y(_11259_));
 NAND2x1_ASAP7_75t_R _19593_ (.A(_10879_),
    .B(net24),
    .Y(_11260_));
 AOI21x1_ASAP7_75t_R _19594_ (.A1(_11260_),
    .A2(_11125_),
    .B(_10883_),
    .Y(_11261_));
 AOI21x1_ASAP7_75t_R _19595_ (.A1(_11259_),
    .A2(_11261_),
    .B(_10899_),
    .Y(_11262_));
 AO21x1_ASAP7_75t_R _19596_ (.A1(_00498_),
    .A2(_10869_),
    .B(_10777_),
    .Y(_11263_));
 AO21x1_ASAP7_75t_R _19597_ (.A1(_10946_),
    .A2(_11032_),
    .B(_11263_),
    .Y(_11264_));
 NOR2x1_ASAP7_75t_R _19598_ (.A(_10939_),
    .B(_11229_),
    .Y(_11265_));
 AO21x1_ASAP7_75t_R _19599_ (.A1(_10841_),
    .A2(_10843_),
    .B(_10746_),
    .Y(_11266_));
 OA21x2_ASAP7_75t_R _19600_ (.A1(_11265_),
    .A2(_11266_),
    .B(_10790_),
    .Y(_11267_));
 NAND2x1_ASAP7_75t_R _19601_ (.A(_11264_),
    .B(_11267_),
    .Y(_11268_));
 AOI21x1_ASAP7_75t_R _19602_ (.A1(_11262_),
    .A2(_11268_),
    .B(_11248_),
    .Y(_11269_));
 NAND2x1_ASAP7_75t_R _19603_ (.A(_11257_),
    .B(_11269_),
    .Y(_11270_));
 NOR2x1_ASAP7_75t_R _19604_ (.A(_10902_),
    .B(_10917_),
    .Y(_11271_));
 AOI211x1_ASAP7_75t_R _19605_ (.A1(_11271_),
    .A2(_11042_),
    .B(_11242_),
    .C(_10912_),
    .Y(_11272_));
 NAND2x2_ASAP7_75t_R _19606_ (.A(_10732_),
    .B(_11032_),
    .Y(_11273_));
 AOI22x1_ASAP7_75t_R _19607_ (.A1(_10847_),
    .A2(_10927_),
    .B1(_10875_),
    .B2(_10770_),
    .Y(_11274_));
 AOI21x1_ASAP7_75t_R _19608_ (.A1(_11273_),
    .A2(_11274_),
    .B(_10934_),
    .Y(_11275_));
 OAI21x1_ASAP7_75t_R _19609_ (.A1(_11272_),
    .A2(_11275_),
    .B(_10899_),
    .Y(_11276_));
 NAND2x1_ASAP7_75t_R _19610_ (.A(_10906_),
    .B(_11026_),
    .Y(_11277_));
 AO21x1_ASAP7_75t_R _19611_ (.A1(_10870_),
    .A2(_11277_),
    .B(_11172_),
    .Y(_11278_));
 AO21x1_ASAP7_75t_R _19612_ (.A1(_01157_),
    .A2(_01155_),
    .B(_10805_),
    .Y(_11279_));
 AND2x2_ASAP7_75t_R _19613_ (.A(_11279_),
    .B(_10907_),
    .Y(_11280_));
 NAND2x1_ASAP7_75t_R _19614_ (.A(_10893_),
    .B(_11116_),
    .Y(_11281_));
 AOI21x1_ASAP7_75t_R _19615_ (.A1(_11280_),
    .A2(_11281_),
    .B(_10970_),
    .Y(_11282_));
 AOI21x1_ASAP7_75t_R _19616_ (.A1(_11278_),
    .A2(_11282_),
    .B(_10883_),
    .Y(_11283_));
 NAND2x1_ASAP7_75t_R _19617_ (.A(_11276_),
    .B(_11283_),
    .Y(_11284_));
 NAND2x1_ASAP7_75t_R _19618_ (.A(_10893_),
    .B(_10977_),
    .Y(_11285_));
 OA21x2_ASAP7_75t_R _19619_ (.A1(_10874_),
    .A2(_10752_),
    .B(_10777_),
    .Y(_11286_));
 AOI21x1_ASAP7_75t_R _19620_ (.A1(_11285_),
    .A2(_11286_),
    .B(_10860_),
    .Y(_11287_));
 AOI21x1_ASAP7_75t_R _19621_ (.A1(_10842_),
    .A2(_10844_),
    .B(_10802_),
    .Y(_11288_));
 AOI22x1_ASAP7_75t_R _19622_ (.A1(_11231_),
    .A2(_10955_),
    .B1(net65),
    .B2(_10927_),
    .Y(_11289_));
 NAND2x1_ASAP7_75t_R _19623_ (.A(_11288_),
    .B(_11289_),
    .Y(_11290_));
 AOI21x1_ASAP7_75t_R _19624_ (.A1(_11287_),
    .A2(_11290_),
    .B(_10791_),
    .Y(_11291_));
 AOI21x1_ASAP7_75t_R _19625_ (.A1(_15804_),
    .A2(_10797_),
    .B(net487),
    .Y(_11292_));
 AND2x2_ASAP7_75t_R _19626_ (.A(_10805_),
    .B(_00496_),
    .Y(_11293_));
 AOI21x1_ASAP7_75t_R _19627_ (.A1(_10879_),
    .A2(_11292_),
    .B(_11293_),
    .Y(_11294_));
 NAND2x1_ASAP7_75t_R _19628_ (.A(_10934_),
    .B(_11294_),
    .Y(_11295_));
 AO21x1_ASAP7_75t_R _19629_ (.A1(_10906_),
    .A2(_10868_),
    .B(_10752_),
    .Y(_11296_));
 AOI21x1_ASAP7_75t_R _19630_ (.A1(_10798_),
    .A2(_11018_),
    .B(_10802_),
    .Y(_11297_));
 AOI21x1_ASAP7_75t_R _19631_ (.A1(_11296_),
    .A2(_11297_),
    .B(_10970_),
    .Y(_11298_));
 NAND2x1_ASAP7_75t_R _19632_ (.A(_11295_),
    .B(_11298_),
    .Y(_11299_));
 AOI21x1_ASAP7_75t_R _19633_ (.A1(_11291_),
    .A2(_11299_),
    .B(_10834_),
    .Y(_11300_));
 NAND2x1_ASAP7_75t_R _19634_ (.A(_11300_),
    .B(_11284_),
    .Y(_11301_));
 NAND2x1_ASAP7_75t_R _19635_ (.A(_11270_),
    .B(_11301_),
    .Y(_00038_));
 AND2x2_ASAP7_75t_R _19636_ (.A(_10863_),
    .B(_10732_),
    .Y(_11302_));
 OAI21x1_ASAP7_75t_R _19637_ (.A1(_11302_),
    .A2(_11105_),
    .B(_10803_),
    .Y(_11303_));
 AO21x1_ASAP7_75t_R _19638_ (.A1(_11057_),
    .A2(_11273_),
    .B(_10803_),
    .Y(_11304_));
 AOI21x1_ASAP7_75t_R _19639_ (.A1(_11303_),
    .A2(_11304_),
    .B(_10861_),
    .Y(_11305_));
 NOR2x1_ASAP7_75t_R _19640_ (.A(_10778_),
    .B(_10992_),
    .Y(_11306_));
 AO21x1_ASAP7_75t_R _19641_ (.A1(_11185_),
    .A2(_11306_),
    .B(_10899_),
    .Y(_11307_));
 AO21x1_ASAP7_75t_R _19642_ (.A1(_15804_),
    .A2(_15806_),
    .B(_15811_),
    .Y(_11308_));
 AOI21x1_ASAP7_75t_R _19643_ (.A1(_10873_),
    .A2(_11308_),
    .B(_10987_),
    .Y(_11309_));
 OAI21x1_ASAP7_75t_R _19644_ (.A1(_10801_),
    .A2(_10888_),
    .B(_10857_),
    .Y(_11310_));
 NOR2x1_ASAP7_75t_R _19645_ (.A(_11309_),
    .B(_11310_),
    .Y(_11311_));
 OAI21x1_ASAP7_75t_R _19646_ (.A1(_11307_),
    .A2(_11311_),
    .B(_10792_),
    .Y(_11312_));
 OAI21x1_ASAP7_75t_R _19647_ (.A1(_11305_),
    .A2(_11312_),
    .B(_10835_),
    .Y(_11313_));
 AOI21x1_ASAP7_75t_R _19648_ (.A1(_10956_),
    .A2(_10977_),
    .B(_11225_),
    .Y(_11314_));
 OAI21x1_ASAP7_75t_R _19649_ (.A1(_10818_),
    .A2(_11314_),
    .B(_10920_),
    .Y(_11315_));
 NOR2x1_ASAP7_75t_R _19650_ (.A(_15811_),
    .B(_10847_),
    .Y(_11316_));
 NOR2x1_ASAP7_75t_R _19651_ (.A(_11316_),
    .B(_11158_),
    .Y(_11317_));
 NOR2x1_ASAP7_75t_R _19652_ (.A(_11317_),
    .B(_11163_),
    .Y(_11318_));
 NOR2x1_ASAP7_75t_R _19653_ (.A(_11315_),
    .B(_11318_),
    .Y(_11319_));
 NOR2x1_ASAP7_75t_R _19654_ (.A(_11122_),
    .B(_11316_),
    .Y(_11320_));
 OAI21x1_ASAP7_75t_R _19655_ (.A1(_10987_),
    .A2(_10888_),
    .B(_10934_),
    .Y(_11321_));
 NOR2x1_ASAP7_75t_R _19656_ (.A(_11320_),
    .B(_11321_),
    .Y(_11322_));
 AO21x1_ASAP7_75t_R _19657_ (.A1(_15804_),
    .A2(_15806_),
    .B(_11124_),
    .Y(_11323_));
 AND2x2_ASAP7_75t_R _19658_ (.A(_11110_),
    .B(_10907_),
    .Y(_11324_));
 AO21x1_ASAP7_75t_R _19659_ (.A1(_11323_),
    .A2(_11324_),
    .B(_10920_),
    .Y(_11325_));
 OAI21x1_ASAP7_75t_R _19660_ (.A1(_11322_),
    .A2(_11325_),
    .B(_10884_),
    .Y(_11326_));
 NOR2x1_ASAP7_75t_R _19661_ (.A(_11319_),
    .B(_11326_),
    .Y(_11327_));
 OA21x2_ASAP7_75t_R _19662_ (.A1(_15804_),
    .A2(_10752_),
    .B(_10777_),
    .Y(_11328_));
 OAI21x1_ASAP7_75t_R _19663_ (.A1(_10753_),
    .A2(_11011_),
    .B(_11328_),
    .Y(_11329_));
 AND2x2_ASAP7_75t_R _19664_ (.A(_10869_),
    .B(_00497_),
    .Y(_11330_));
 OA21x2_ASAP7_75t_R _19665_ (.A1(_10908_),
    .A2(_11330_),
    .B(_10883_),
    .Y(_11331_));
 OA21x2_ASAP7_75t_R _19666_ (.A1(_11003_),
    .A2(_11329_),
    .B(_11331_),
    .Y(_11332_));
 AOI21x1_ASAP7_75t_R _19667_ (.A1(_10873_),
    .A2(_11308_),
    .B(_10753_),
    .Y(_11333_));
 AO21x1_ASAP7_75t_R _19668_ (.A1(_10874_),
    .A2(_10868_),
    .B(_10728_),
    .Y(_11334_));
 NAND2x1_ASAP7_75t_R _19669_ (.A(_10747_),
    .B(_11334_),
    .Y(_11335_));
 NOR2x1_ASAP7_75t_R _19670_ (.A(_11333_),
    .B(_11335_),
    .Y(_11336_));
 NOR2x1_ASAP7_75t_R _19671_ (.A(_11083_),
    .B(_11098_),
    .Y(_11337_));
 NAND2x1_ASAP7_75t_R _19672_ (.A(_15814_),
    .B(_11225_),
    .Y(_11338_));
 NAND2x1_ASAP7_75t_R _19673_ (.A(_11338_),
    .B(_11328_),
    .Y(_11339_));
 OAI21x1_ASAP7_75t_R _19674_ (.A1(_11337_),
    .A2(_11339_),
    .B(_10791_),
    .Y(_11340_));
 OAI21x1_ASAP7_75t_R _19675_ (.A1(_11336_),
    .A2(_11340_),
    .B(_10861_),
    .Y(_11341_));
 NOR2x1_ASAP7_75t_R _19676_ (.A(_11332_),
    .B(_11341_),
    .Y(_11342_));
 AO21x1_ASAP7_75t_R _19677_ (.A1(_10794_),
    .A2(_10913_),
    .B(_10747_),
    .Y(_11343_));
 AOI21x1_ASAP7_75t_R _19678_ (.A1(_10893_),
    .A2(_11116_),
    .B(_11343_),
    .Y(_11344_));
 OAI21x1_ASAP7_75t_R _19679_ (.A1(_10987_),
    .A2(_10867_),
    .B(_10873_),
    .Y(_11345_));
 OAI21x1_ASAP7_75t_R _19680_ (.A1(_10908_),
    .A2(_11345_),
    .B(_10791_),
    .Y(_11346_));
 OAI21x1_ASAP7_75t_R _19681_ (.A1(_11344_),
    .A2(_11346_),
    .B(_10767_),
    .Y(_11347_));
 NOR2x1_ASAP7_75t_R _19682_ (.A(_01157_),
    .B(_10987_),
    .Y(_11348_));
 OA21x2_ASAP7_75t_R _19683_ (.A1(_10917_),
    .A2(_10862_),
    .B(_10987_),
    .Y(_11349_));
 OAI21x1_ASAP7_75t_R _19684_ (.A1(_11348_),
    .A2(_11349_),
    .B(_10818_),
    .Y(_11350_));
 NAND2x1_ASAP7_75t_R _19685_ (.A(_10800_),
    .B(_10946_),
    .Y(_11351_));
 NAND2x1_ASAP7_75t_R _19686_ (.A(_10877_),
    .B(_10863_),
    .Y(_11352_));
 AO21x1_ASAP7_75t_R _19687_ (.A1(_11351_),
    .A2(_11352_),
    .B(_10818_),
    .Y(_11353_));
 AOI21x1_ASAP7_75t_R _19688_ (.A1(_11350_),
    .A2(_11353_),
    .B(_10792_),
    .Y(_11354_));
 OAI21x1_ASAP7_75t_R _19689_ (.A1(_11347_),
    .A2(_11354_),
    .B(_11248_),
    .Y(_11355_));
 OAI22x1_ASAP7_75t_R _19690_ (.A1(_11313_),
    .A2(_11327_),
    .B1(_11342_),
    .B2(_11355_),
    .Y(_00039_));
 BUFx16f_ASAP7_75t_R _19691_ (.A(_10762_),
    .Y(_11356_));
 NOR2x2_ASAP7_75t_R _19692_ (.A(net641),
    .B(_00499_),
    .Y(_11357_));
 BUFx2_ASAP7_75t_R rebuffer252 (.A(_00772_),
    .Y(net705));
 XOR2x2_ASAP7_75t_R _19694_ (.A(_00779_),
    .B(_00772_),
    .Y(_11359_));
 BUFx6f_ASAP7_75t_R _19695_ (.A(_00837_),
    .Y(_11360_));
 XOR2x2_ASAP7_75t_R _19696_ (.A(_11360_),
    .B(_11359_),
    .Y(_11361_));
 BUFx6f_ASAP7_75t_R _19697_ (.A(_00740_),
    .Y(_11362_));
 BUFx6f_ASAP7_75t_R _19698_ (.A(_00747_),
    .Y(_11363_));
 XOR2x2_ASAP7_75t_R _19699_ (.A(_11362_),
    .B(_11363_),
    .Y(_11364_));
 BUFx4f_ASAP7_75t_R _19700_ (.A(_00805_),
    .Y(_11365_));
 XOR2x2_ASAP7_75t_R _19701_ (.A(_00773_),
    .B(_11365_),
    .Y(_11366_));
 XOR2x2_ASAP7_75t_R _19702_ (.A(_11364_),
    .B(_11366_),
    .Y(_11367_));
 NAND2x1_ASAP7_75t_R _19703_ (.A(_11361_),
    .B(net853),
    .Y(_11368_));
 OR2x2_ASAP7_75t_R _19704_ (.A(_11361_),
    .B(net853),
    .Y(_11369_));
 BUFx12f_ASAP7_75t_R _19705_ (.A(_10643_),
    .Y(_11370_));
 AOI21x1_ASAP7_75t_R _19706_ (.A1(_11368_),
    .A2(_11369_),
    .B(_11370_),
    .Y(_11371_));
 OAI21x1_ASAP7_75t_R _19707_ (.A1(_11357_),
    .A2(_11371_),
    .B(_08186_),
    .Y(_11372_));
 BUFx12f_ASAP7_75t_R _19708_ (.A(_10638_),
    .Y(_11373_));
 BUFx12f_ASAP7_75t_R _19709_ (.A(_11373_),
    .Y(_11374_));
 AND2x2_ASAP7_75t_R _19710_ (.A(_11374_),
    .B(_00499_),
    .Y(_11375_));
 XNOR2x2_ASAP7_75t_R _19711_ (.A(_11367_),
    .B(_11361_),
    .Y(_11376_));
 NOR2x2_ASAP7_75t_R _19712_ (.A(_11370_),
    .B(_11376_),
    .Y(_11377_));
 INVx2_ASAP7_75t_R _19713_ (.A(_08186_),
    .Y(_11378_));
 OAI21x1_ASAP7_75t_R _19714_ (.A1(_11377_),
    .A2(_11375_),
    .B(_11378_),
    .Y(_11379_));
 NAND2x2_ASAP7_75t_R _19715_ (.A(_11372_),
    .B(_11379_),
    .Y(_11380_));
 BUFx6f_ASAP7_75t_R _19716_ (.A(_11380_),
    .Y(_15821_));
 BUFx6f_ASAP7_75t_R _19717_ (.A(_00836_),
    .Y(_11381_));
 INVx2_ASAP7_75t_R _19718_ (.A(net776),
    .Y(_11382_));
 BUFx10_ASAP7_75t_R _19719_ (.A(_00779_),
    .Y(_11383_));
 XOR2x2_ASAP7_75t_R _19720_ (.A(_11363_),
    .B(_11383_),
    .Y(_11384_));
 NAND2x1_ASAP7_75t_R _19721_ (.A(_11382_),
    .B(_11384_),
    .Y(_11385_));
 XNOR2x1_ASAP7_75t_R _19722_ (.B(_11383_),
    .Y(_11386_),
    .A(_11363_));
 NAND2x1_ASAP7_75t_R _19723_ (.A(net777),
    .B(_11386_),
    .Y(_11387_));
 BUFx6f_ASAP7_75t_R _19724_ (.A(_00804_),
    .Y(_11388_));
 XNOR2x2_ASAP7_75t_R _19725_ (.A(_00772_),
    .B(_11388_),
    .Y(_11389_));
 AOI21x1_ASAP7_75t_R _19726_ (.A1(_11385_),
    .A2(_11387_),
    .B(_11389_),
    .Y(_11390_));
 NAND2x1_ASAP7_75t_R _19727_ (.A(net777),
    .B(_11384_),
    .Y(_11391_));
 NAND2x1_ASAP7_75t_R _19728_ (.A(_11382_),
    .B(_11386_),
    .Y(_11392_));
 XOR2x2_ASAP7_75t_R _19729_ (.A(_11388_),
    .B(_00772_),
    .Y(_11393_));
 AOI21x1_ASAP7_75t_R _19730_ (.A1(_11391_),
    .A2(_11392_),
    .B(_11393_),
    .Y(_11394_));
 OAI21x1_ASAP7_75t_R _19731_ (.A1(_11390_),
    .A2(_11394_),
    .B(net651),
    .Y(_11395_));
 INVx2_ASAP7_75t_R _19732_ (.A(_01043_),
    .Y(_11396_));
 NOR2x1_ASAP7_75t_R _19733_ (.A(_10620_),
    .B(_00500_),
    .Y(_11397_));
 INVx3_ASAP7_75t_R _19734_ (.A(_11397_),
    .Y(_11398_));
 NAND3x2_ASAP7_75t_R _19735_ (.B(_11396_),
    .C(_11398_),
    .Y(_11399_),
    .A(net687));
 AO21x1_ASAP7_75t_R _19736_ (.A1(net687),
    .A2(_11398_),
    .B(_11396_),
    .Y(_11400_));
 NAND2x2_ASAP7_75t_R _19737_ (.A(_11399_),
    .B(_11400_),
    .Y(_11401_));
 BUFx12_ASAP7_75t_R _19738_ (.A(_11401_),
    .Y(_15823_));
 BUFx4f_ASAP7_75t_R _19739_ (.A(_00774_),
    .Y(_11402_));
 INVx1_ASAP7_75t_R _19740_ (.A(_11402_),
    .Y(_11403_));
 BUFx6f_ASAP7_75t_R _19741_ (.A(_00741_),
    .Y(_11404_));
 XOR2x2_ASAP7_75t_R _19742_ (.A(_00773_),
    .B(_11404_),
    .Y(_11405_));
 NAND2x1_ASAP7_75t_R _19743_ (.A(_11403_),
    .B(_11405_),
    .Y(_11406_));
 XNOR2x2_ASAP7_75t_R _19744_ (.A(_11404_),
    .B(_00773_),
    .Y(_11407_));
 NAND2x1_ASAP7_75t_R _19745_ (.A(_11402_),
    .B(net629),
    .Y(_11408_));
 BUFx6f_ASAP7_75t_R _19746_ (.A(_00806_),
    .Y(_11409_));
 BUFx6f_ASAP7_75t_R _19747_ (.A(_00838_),
    .Y(_11410_));
 XNOR2x2_ASAP7_75t_R _19748_ (.A(_11409_),
    .B(_11410_),
    .Y(_11411_));
 AOI21x1_ASAP7_75t_R _19749_ (.A1(_11406_),
    .A2(_11408_),
    .B(_11411_),
    .Y(_11412_));
 NAND2x1_ASAP7_75t_R _19750_ (.A(_11402_),
    .B(_11405_),
    .Y(_11413_));
 NAND2x1_ASAP7_75t_R _19751_ (.A(_11403_),
    .B(net629),
    .Y(_11414_));
 XOR2x2_ASAP7_75t_R _19752_ (.A(_11409_),
    .B(_11410_),
    .Y(_11415_));
 AOI21x1_ASAP7_75t_R _19753_ (.A1(_11413_),
    .A2(_11414_),
    .B(_11415_),
    .Y(_11416_));
 OAI21x1_ASAP7_75t_R _19754_ (.A1(_11412_),
    .A2(_11416_),
    .B(net680),
    .Y(_11417_));
 OR2x4_ASAP7_75t_R _19755_ (.A(_10619_),
    .B(_00502_),
    .Y(_11418_));
 NAND3x2_ASAP7_75t_R _19756_ (.B(_01045_),
    .C(_11418_),
    .Y(_11419_),
    .A(_11417_));
 AO21x1_ASAP7_75t_R _19757_ (.A1(_11417_),
    .A2(_11418_),
    .B(_01045_),
    .Y(_11420_));
 BUFx6f_ASAP7_75t_R _19758_ (.A(_11420_),
    .Y(_11421_));
 NAND2x2_ASAP7_75t_R _19759_ (.A(_11419_),
    .B(_11421_),
    .Y(_11422_));
 BUFx10_ASAP7_75t_R _19760_ (.A(_11422_),
    .Y(_15831_));
 NAND3x2_ASAP7_75t_R _19761_ (.B(_01043_),
    .C(_11398_),
    .Y(_11423_),
    .A(net690));
 AO21x1_ASAP7_75t_R _19762_ (.A1(_11395_),
    .A2(_11398_),
    .B(_01043_),
    .Y(_11424_));
 NAND2x2_ASAP7_75t_R _19763_ (.A(_11423_),
    .B(_11424_),
    .Y(_11425_));
 BUFx10_ASAP7_75t_R _19764_ (.A(_11425_),
    .Y(_15818_));
 INVx2_ASAP7_75t_R _19765_ (.A(_01045_),
    .Y(_11426_));
 NAND3x2_ASAP7_75t_R _19766_ (.B(_11426_),
    .C(_11418_),
    .Y(_11427_),
    .A(_11417_));
 AO21x1_ASAP7_75t_R _19767_ (.A1(_11417_),
    .A2(_11418_),
    .B(_11426_),
    .Y(_11428_));
 BUFx6f_ASAP7_75t_R _19768_ (.A(_11428_),
    .Y(_11429_));
 NAND2x2_ASAP7_75t_R _19769_ (.A(_11427_),
    .B(_11429_),
    .Y(_11430_));
 BUFx10_ASAP7_75t_R _19770_ (.A(_11430_),
    .Y(_11431_));
 BUFx10_ASAP7_75t_R _19771_ (.A(_11431_),
    .Y(_15828_));
 BUFx6f_ASAP7_75t_R _19772_ (.A(_11430_),
    .Y(_11432_));
 BUFx6f_ASAP7_75t_R _19773_ (.A(_00742_),
    .Y(_11433_));
 XOR2x2_ASAP7_75t_R _19774_ (.A(_11433_),
    .B(_11363_),
    .Y(_11434_));
 XOR2x1_ASAP7_75t_R _19775_ (.A(_11434_),
    .Y(_11435_),
    .B(_00775_));
 XOR2x2_ASAP7_75t_R _19776_ (.A(_11402_),
    .B(_11383_),
    .Y(_11436_));
 XOR2x2_ASAP7_75t_R _19777_ (.A(_00807_),
    .B(_00839_),
    .Y(_11437_));
 XOR2x1_ASAP7_75t_R _19778_ (.A(_11436_),
    .Y(_11438_),
    .B(_11437_));
 OAI21x1_ASAP7_75t_R _19779_ (.A1(_11435_),
    .A2(_11438_),
    .B(net867),
    .Y(_11439_));
 AND2x2_ASAP7_75t_R _19780_ (.A(_11438_),
    .B(_11435_),
    .Y(_11440_));
 BUFx12f_ASAP7_75t_R _19781_ (.A(_10639_),
    .Y(_11441_));
 NAND2x1_ASAP7_75t_R _19782_ (.A(_00650_),
    .B(_11441_),
    .Y(_11442_));
 OAI21x1_ASAP7_75t_R _19783_ (.A1(_11439_),
    .A2(_11440_),
    .B(_11442_),
    .Y(_11443_));
 XOR2x2_ASAP7_75t_R _19784_ (.A(_11443_),
    .B(_01046_),
    .Y(_11444_));
 BUFx6f_ASAP7_75t_R _19785_ (.A(_11444_),
    .Y(_11445_));
 AO21x1_ASAP7_75t_R _19786_ (.A1(_15818_),
    .A2(_11432_),
    .B(_11445_),
    .Y(_11446_));
 INVx1_ASAP7_75t_R _19787_ (.A(_11357_),
    .Y(_11447_));
 NAND2x1_ASAP7_75t_R _19788_ (.A(_10786_),
    .B(_11376_),
    .Y(_11448_));
 AOI21x1_ASAP7_75t_R _19789_ (.A1(_11447_),
    .A2(_11448_),
    .B(_11378_),
    .Y(_11449_));
 BUFx12f_ASAP7_75t_R _19790_ (.A(_10666_),
    .Y(_11450_));
 BUFx10_ASAP7_75t_R _19791_ (.A(_11450_),
    .Y(_11451_));
 AOI211x1_ASAP7_75t_R _19792_ (.A1(_11376_),
    .A2(_11451_),
    .B(_11357_),
    .C(_08186_),
    .Y(_11452_));
 OAI21x1_ASAP7_75t_R _19793_ (.A1(_11449_),
    .A2(_11452_),
    .B(_15818_),
    .Y(_11453_));
 NOR2x2_ASAP7_75t_R _19794_ (.A(_11431_),
    .B(_11453_),
    .Y(_11454_));
 NOR2x1_ASAP7_75t_R _19795_ (.A(_11446_),
    .B(_11454_),
    .Y(_11455_));
 BUFx6f_ASAP7_75t_R _19796_ (.A(_11422_),
    .Y(_11456_));
 XOR2x2_ASAP7_75t_R _19797_ (.A(_11443_),
    .B(_10096_),
    .Y(_11457_));
 BUFx6f_ASAP7_75t_R _19798_ (.A(_11457_),
    .Y(_11458_));
 AOI21x1_ASAP7_75t_R _19799_ (.A1(_01162_),
    .A2(_11456_),
    .B(_11458_),
    .Y(_11459_));
 INVx2_ASAP7_75t_R _19800_ (.A(net582),
    .Y(_11460_));
 AOI21x1_ASAP7_75t_R _19801_ (.A1(_11427_),
    .A2(_11429_),
    .B(_11460_),
    .Y(_11461_));
 INVx3_ASAP7_75t_R _19802_ (.A(net508),
    .Y(_11462_));
 XOR2x2_ASAP7_75t_R _19803_ (.A(_00743_),
    .B(_11363_),
    .Y(_11463_));
 XNOR2x1_ASAP7_75t_R _19804_ (.B(_11463_),
    .Y(_11464_),
    .A(_00776_));
 XOR2x2_ASAP7_75t_R _19805_ (.A(_00775_),
    .B(_11383_),
    .Y(_11465_));
 XOR2x2_ASAP7_75t_R _19806_ (.A(_00808_),
    .B(_00840_),
    .Y(_11466_));
 XOR2x1_ASAP7_75t_R _19807_ (.A(_11465_),
    .Y(_11467_),
    .B(_11466_));
 XOR2x1_ASAP7_75t_R _19808_ (.A(_11464_),
    .Y(_11468_),
    .B(_11467_));
 NOR2x1_ASAP7_75t_R _19809_ (.A(_10743_),
    .B(_00649_),
    .Y(_11469_));
 AOI21x1_ASAP7_75t_R _19810_ (.A1(_10734_),
    .A2(_11468_),
    .B(_11469_),
    .Y(_11470_));
 XNOR2x2_ASAP7_75t_R _19811_ (.A(_08220_),
    .B(_11470_),
    .Y(_11471_));
 BUFx6f_ASAP7_75t_R _19812_ (.A(_11471_),
    .Y(_11472_));
 AO21x1_ASAP7_75t_R _19813_ (.A1(_11459_),
    .A2(_11462_),
    .B(_11472_),
    .Y(_11473_));
 NOR2x1_ASAP7_75t_R _19814_ (.A(_11455_),
    .B(_11473_),
    .Y(_11474_));
 BUFx6f_ASAP7_75t_R _19815_ (.A(_11471_),
    .Y(_11475_));
 AO21x1_ASAP7_75t_R _19816_ (.A1(_15818_),
    .A2(_11422_),
    .B(_11444_),
    .Y(_11476_));
 BUFx4f_ASAP7_75t_R _19817_ (.A(_11476_),
    .Y(_11477_));
 NAND2x1_ASAP7_75t_R _19818_ (.A(_11475_),
    .B(_11477_),
    .Y(_11478_));
 INVx1_ASAP7_75t_R _19819_ (.A(_01160_),
    .Y(_11479_));
 BUFx6f_ASAP7_75t_R _19820_ (.A(_11444_),
    .Y(_11480_));
 OA21x2_ASAP7_75t_R _19821_ (.A1(_11456_),
    .A2(_11479_),
    .B(_11480_),
    .Y(_11481_));
 INVx1_ASAP7_75t_R _19822_ (.A(_11481_),
    .Y(_11482_));
 NOR2x1_ASAP7_75t_R _19823_ (.A(_11454_),
    .B(_11482_),
    .Y(_11483_));
 XOR2x2_ASAP7_75t_R _19824_ (.A(_00744_),
    .B(_00776_),
    .Y(_11484_));
 INVx3_ASAP7_75t_R _19825_ (.A(_00841_),
    .Y(_11485_));
 XOR2x1_ASAP7_75t_R _19826_ (.A(_11484_),
    .Y(_11486_),
    .B(_11485_));
 XOR2x2_ASAP7_75t_R _19827_ (.A(_00777_),
    .B(_00809_),
    .Y(_11487_));
 XOR2x1_ASAP7_75t_R _19828_ (.A(_11486_),
    .Y(_11488_),
    .B(_11487_));
 NOR2x1_ASAP7_75t_R _19829_ (.A(net585),
    .B(_00648_),
    .Y(_11489_));
 AO21x1_ASAP7_75t_R _19830_ (.A1(_11488_),
    .A2(_10761_),
    .B(_11489_),
    .Y(_11490_));
 XOR2x2_ASAP7_75t_R _19831_ (.A(_11490_),
    .B(_01048_),
    .Y(_11491_));
 INVx1_ASAP7_75t_R _19832_ (.A(_11491_),
    .Y(_11492_));
 BUFx6f_ASAP7_75t_R _19833_ (.A(_11492_),
    .Y(_11493_));
 BUFx6f_ASAP7_75t_R _19834_ (.A(_11493_),
    .Y(_11494_));
 OAI21x1_ASAP7_75t_R _19835_ (.A1(_11478_),
    .A2(_11483_),
    .B(_11494_),
    .Y(_11495_));
 XOR2x2_ASAP7_75t_R _19836_ (.A(_00745_),
    .B(_00777_),
    .Y(_11496_));
 XOR2x2_ASAP7_75t_R _19837_ (.A(_00778_),
    .B(_00810_),
    .Y(_11497_));
 XOR2x1_ASAP7_75t_R _19838_ (.A(_11497_),
    .Y(_11498_),
    .B(_00842_));
 XNOR2x1_ASAP7_75t_R _19839_ (.B(_11498_),
    .Y(_11499_),
    .A(_11496_));
 NOR2x1_ASAP7_75t_R _19840_ (.A(_10829_),
    .B(_00647_),
    .Y(_11500_));
 AO21x1_ASAP7_75t_R _19841_ (.A1(_11499_),
    .A2(_11451_),
    .B(_11500_),
    .Y(_11501_));
 XOR2x2_ASAP7_75t_R _19842_ (.A(_11501_),
    .B(_01050_),
    .Y(_11502_));
 CKINVDCx9p33_ASAP7_75t_R _19843_ (.A(_11502_),
    .Y(_11503_));
 BUFx10_ASAP7_75t_R _19844_ (.A(_11503_),
    .Y(_11504_));
 OAI21x1_ASAP7_75t_R _19845_ (.A1(_11474_),
    .A2(_11495_),
    .B(_11504_),
    .Y(_11505_));
 XOR2x2_ASAP7_75t_R _19846_ (.A(_11470_),
    .B(_08220_),
    .Y(_11506_));
 BUFx6f_ASAP7_75t_R _19847_ (.A(_11506_),
    .Y(_11507_));
 BUFx6f_ASAP7_75t_R _19848_ (.A(_11507_),
    .Y(_11508_));
 INVx1_ASAP7_75t_R _19849_ (.A(_11454_),
    .Y(_11509_));
 BUFx6f_ASAP7_75t_R _19850_ (.A(_11480_),
    .Y(_11510_));
 OAI21x1_ASAP7_75t_R _19851_ (.A1(_11371_),
    .A2(_11357_),
    .B(_11378_),
    .Y(_11511_));
 OAI21x1_ASAP7_75t_R _19852_ (.A1(_11375_),
    .A2(_11377_),
    .B(_08186_),
    .Y(_11512_));
 AOI21x1_ASAP7_75t_R _19853_ (.A1(_11511_),
    .A2(_11512_),
    .B(_11422_),
    .Y(_11513_));
 NOR2x2_ASAP7_75t_R _19854_ (.A(_11510_),
    .B(_11513_),
    .Y(_11514_));
 OA21x2_ASAP7_75t_R _19855_ (.A1(_15823_),
    .A2(_11431_),
    .B(_11480_),
    .Y(_11515_));
 INVx1_ASAP7_75t_R _19856_ (.A(_01162_),
    .Y(_11516_));
 AO21x2_ASAP7_75t_R _19857_ (.A1(_11429_),
    .A2(_11427_),
    .B(_11516_),
    .Y(_11517_));
 AOI22x1_ASAP7_75t_R _19858_ (.A1(_11509_),
    .A2(_11514_),
    .B1(_11515_),
    .B2(_11517_),
    .Y(_11518_));
 BUFx4f_ASAP7_75t_R _19859_ (.A(_11444_),
    .Y(_11519_));
 BUFx6f_ASAP7_75t_R _19860_ (.A(_11519_),
    .Y(_11520_));
 INVx1_ASAP7_75t_R _19861_ (.A(_11511_),
    .Y(_11521_));
 INVx1_ASAP7_75t_R _19862_ (.A(net686),
    .Y(_11522_));
 OAI21x1_ASAP7_75t_R _19863_ (.A1(_11521_),
    .A2(_11522_),
    .B(_11422_),
    .Y(_11523_));
 BUFx6f_ASAP7_75t_R _19864_ (.A(_11457_),
    .Y(_11524_));
 AOI21x1_ASAP7_75t_R _19865_ (.A1(_11427_),
    .A2(_11429_),
    .B(_01159_),
    .Y(_11525_));
 AOI21x1_ASAP7_75t_R _19866_ (.A1(_11524_),
    .A2(_11525_),
    .B(_11506_),
    .Y(_11526_));
 OAI21x1_ASAP7_75t_R _19867_ (.A1(_11520_),
    .A2(_11523_),
    .B(_11526_),
    .Y(_11527_));
 NOR2x2_ASAP7_75t_R _19868_ (.A(_11425_),
    .B(_11422_),
    .Y(_11528_));
 NAND2x2_ASAP7_75t_R _19869_ (.A(net564),
    .B(_11528_),
    .Y(_11529_));
 AND2x2_ASAP7_75t_R _19870_ (.A(_11529_),
    .B(_11515_),
    .Y(_11530_));
 BUFx6f_ASAP7_75t_R _19871_ (.A(_11491_),
    .Y(_11531_));
 BUFx10_ASAP7_75t_R _19872_ (.A(_11531_),
    .Y(_11532_));
 OAI21x1_ASAP7_75t_R _19873_ (.A1(_11527_),
    .A2(_11530_),
    .B(_11532_),
    .Y(_11533_));
 AOI21x1_ASAP7_75t_R _19874_ (.A1(_11508_),
    .A2(_11518_),
    .B(_11533_),
    .Y(_11534_));
 XNOR2x2_ASAP7_75t_R _19875_ (.A(_00746_),
    .B(_00778_),
    .Y(_11535_));
 BUFx6f_ASAP7_75t_R _19876_ (.A(_00843_),
    .Y(_11536_));
 INVx4_ASAP7_75t_R _19877_ (.A(net616),
    .Y(_11537_));
 XOR2x1_ASAP7_75t_R _19878_ (.A(_11535_),
    .Y(_11538_),
    .B(_11537_));
 BUFx6f_ASAP7_75t_R _19879_ (.A(_00811_),
    .Y(_11539_));
 XNOR2x2_ASAP7_75t_R _19880_ (.A(_11383_),
    .B(net28),
    .Y(_11540_));
 XOR2x1_ASAP7_75t_R _19881_ (.A(_11538_),
    .Y(_11541_),
    .B(_11540_));
 NOR2x1_ASAP7_75t_R _19882_ (.A(_10830_),
    .B(_00646_),
    .Y(_11542_));
 AO21x1_ASAP7_75t_R _19883_ (.A1(_11541_),
    .A2(_10830_),
    .B(_11542_),
    .Y(_11543_));
 XOR2x2_ASAP7_75t_R _19884_ (.A(_11543_),
    .B(_01051_),
    .Y(_11544_));
 BUFx10_ASAP7_75t_R _19885_ (.A(_11544_),
    .Y(_11545_));
 OAI21x1_ASAP7_75t_R _19886_ (.A1(_11505_),
    .A2(_11534_),
    .B(_11545_),
    .Y(_11546_));
 NOR2x2_ASAP7_75t_R _19887_ (.A(_15823_),
    .B(net566),
    .Y(_11547_));
 AO21x2_ASAP7_75t_R _19888_ (.A1(_15823_),
    .A2(_11431_),
    .B(_11480_),
    .Y(_11548_));
 BUFx4f_ASAP7_75t_R _19889_ (.A(_11480_),
    .Y(_11549_));
 OAI21x1_ASAP7_75t_R _19890_ (.A1(_11528_),
    .A2(_11547_),
    .B(_11549_),
    .Y(_11550_));
 OA21x2_ASAP7_75t_R _19891_ (.A1(_11547_),
    .A2(_11548_),
    .B(_11550_),
    .Y(_11551_));
 OAI21x1_ASAP7_75t_R _19892_ (.A1(_11449_),
    .A2(_11452_),
    .B(_15823_),
    .Y(_11552_));
 NOR2x2_ASAP7_75t_R _19893_ (.A(_11432_),
    .B(_11552_),
    .Y(_11553_));
 NOR2x2_ASAP7_75t_R _19894_ (.A(_11445_),
    .B(net508),
    .Y(_11554_));
 INVx1_ASAP7_75t_R _19895_ (.A(_11554_),
    .Y(_11555_));
 INVx1_ASAP7_75t_R _19896_ (.A(_00501_),
    .Y(_11556_));
 AO21x1_ASAP7_75t_R _19897_ (.A1(_11429_),
    .A2(_11427_),
    .B(_11556_),
    .Y(_11557_));
 INVx2_ASAP7_75t_R _19898_ (.A(_00503_),
    .Y(_11558_));
 AOI21x1_ASAP7_75t_R _19899_ (.A1(_11419_),
    .A2(_11421_),
    .B(_11558_),
    .Y(_11559_));
 INVx1_ASAP7_75t_R _19900_ (.A(_11559_),
    .Y(_11560_));
 BUFx6f_ASAP7_75t_R _19901_ (.A(_11457_),
    .Y(_11561_));
 AO21x1_ASAP7_75t_R _19902_ (.A1(_11557_),
    .A2(_11560_),
    .B(_11561_),
    .Y(_11562_));
 OAI21x1_ASAP7_75t_R _19903_ (.A1(_11553_),
    .A2(_11555_),
    .B(_11562_),
    .Y(_11563_));
 BUFx6f_ASAP7_75t_R _19904_ (.A(_11492_),
    .Y(_11564_));
 OAI21x1_ASAP7_75t_R _19905_ (.A1(_11508_),
    .A2(_11563_),
    .B(_11564_),
    .Y(_11565_));
 AOI21x1_ASAP7_75t_R _19906_ (.A1(_11508_),
    .A2(_11551_),
    .B(_11565_),
    .Y(_11566_));
 AO21x1_ASAP7_75t_R _19907_ (.A1(_11429_),
    .A2(_11427_),
    .B(net461),
    .Y(_11567_));
 BUFx4f_ASAP7_75t_R _19908_ (.A(_11567_),
    .Y(_11568_));
 AO21x1_ASAP7_75t_R _19909_ (.A1(_11568_),
    .A2(_11560_),
    .B(_11561_),
    .Y(_11569_));
 AO21x2_ASAP7_75t_R _19910_ (.A1(_11421_),
    .A2(_11419_),
    .B(_11556_),
    .Y(_11570_));
 AOI21x1_ASAP7_75t_R _19911_ (.A1(_11427_),
    .A2(_11429_),
    .B(_11558_),
    .Y(_11571_));
 INVx2_ASAP7_75t_R _19912_ (.A(_11571_),
    .Y(_11572_));
 BUFx6f_ASAP7_75t_R _19913_ (.A(_11480_),
    .Y(_11573_));
 AO21x1_ASAP7_75t_R _19914_ (.A1(_11570_),
    .A2(_11572_),
    .B(_11573_),
    .Y(_11574_));
 AND3x1_ASAP7_75t_R _19915_ (.A(_11569_),
    .B(_11574_),
    .C(_11475_),
    .Y(_11575_));
 BUFx6f_ASAP7_75t_R _19916_ (.A(_11491_),
    .Y(_11576_));
 BUFx6f_ASAP7_75t_R _19917_ (.A(_11480_),
    .Y(_11577_));
 NOR2x1_ASAP7_75t_R _19918_ (.A(_11577_),
    .B(_11523_),
    .Y(_11578_));
 AOI21x1_ASAP7_75t_R _19919_ (.A1(_11419_),
    .A2(_11421_),
    .B(_11460_),
    .Y(_11579_));
 NOR2x2_ASAP7_75t_R _19920_ (.A(_11457_),
    .B(_11579_),
    .Y(_11580_));
 AO21x1_ASAP7_75t_R _19921_ (.A1(_11561_),
    .A2(net508),
    .B(_11580_),
    .Y(_11581_));
 BUFx6f_ASAP7_75t_R _19922_ (.A(_11506_),
    .Y(_11582_));
 OAI21x1_ASAP7_75t_R _19923_ (.A1(_11578_),
    .A2(_11581_),
    .B(_11582_),
    .Y(_11583_));
 NAND2x1_ASAP7_75t_R _19924_ (.A(_11576_),
    .B(_11583_),
    .Y(_11584_));
 BUFx6f_ASAP7_75t_R _19925_ (.A(_11502_),
    .Y(_11585_));
 BUFx10_ASAP7_75t_R _19926_ (.A(_11585_),
    .Y(_11586_));
 OAI21x1_ASAP7_75t_R _19927_ (.A1(_11575_),
    .A2(_11584_),
    .B(_11586_),
    .Y(_11587_));
 NOR2x1_ASAP7_75t_R _19928_ (.A(_11566_),
    .B(_11587_),
    .Y(_11588_));
 BUFx6f_ASAP7_75t_R _19929_ (.A(_11458_),
    .Y(_11589_));
 OAI21x1_ASAP7_75t_R _19930_ (.A1(_11559_),
    .A2(_11525_),
    .B(_11589_),
    .Y(_11590_));
 AOI21x1_ASAP7_75t_R _19931_ (.A1(_11590_),
    .A2(_11482_),
    .B(_11475_),
    .Y(_11591_));
 NAND2x2_ASAP7_75t_R _19932_ (.A(_11401_),
    .B(_11430_),
    .Y(_11592_));
 AO21x1_ASAP7_75t_R _19933_ (.A1(_11592_),
    .A2(_11570_),
    .B(_11524_),
    .Y(_11593_));
 AOI21x1_ASAP7_75t_R _19934_ (.A1(_11419_),
    .A2(_11421_),
    .B(net460),
    .Y(_11594_));
 INVx3_ASAP7_75t_R _19935_ (.A(_11594_),
    .Y(_11595_));
 AOI21x1_ASAP7_75t_R _19936_ (.A1(_11432_),
    .A2(net565),
    .B(_11445_),
    .Y(_11596_));
 NAND2x1_ASAP7_75t_R _19937_ (.A(_11595_),
    .B(_11596_),
    .Y(_11597_));
 BUFx10_ASAP7_75t_R _19938_ (.A(_11506_),
    .Y(_11598_));
 AOI21x1_ASAP7_75t_R _19939_ (.A1(_11593_),
    .A2(_11597_),
    .B(_11598_),
    .Y(_11599_));
 OAI21x1_ASAP7_75t_R _19940_ (.A1(_11591_),
    .A2(_11599_),
    .B(_11503_),
    .Y(_11600_));
 INVx2_ASAP7_75t_R _19941_ (.A(_01161_),
    .Y(_11601_));
 OAI21x1_ASAP7_75t_R _19942_ (.A1(_11431_),
    .A2(_11601_),
    .B(_11445_),
    .Y(_11602_));
 NOR2x2_ASAP7_75t_R _19943_ (.A(_11456_),
    .B(_11453_),
    .Y(_11603_));
 OAI21x1_ASAP7_75t_R _19944_ (.A1(_11602_),
    .A2(_11603_),
    .B(_11526_),
    .Y(_11604_));
 BUFx6f_ASAP7_75t_R _19945_ (.A(_11471_),
    .Y(_11605_));
 AOI21x1_ASAP7_75t_R _19946_ (.A1(_11577_),
    .A2(_11525_),
    .B(_11605_),
    .Y(_11606_));
 BUFx6f_ASAP7_75t_R _19947_ (.A(_11453_),
    .Y(_11607_));
 OA21x2_ASAP7_75t_R _19948_ (.A1(_11430_),
    .A2(_00501_),
    .B(_11457_),
    .Y(_11608_));
 BUFx4f_ASAP7_75t_R _19949_ (.A(_11608_),
    .Y(_11609_));
 OAI21x1_ASAP7_75t_R _19950_ (.A1(_15831_),
    .A2(_11607_),
    .B(_11609_),
    .Y(_11610_));
 AOI21x1_ASAP7_75t_R _19951_ (.A1(_11606_),
    .A2(_11610_),
    .B(_11503_),
    .Y(_11611_));
 AOI21x1_ASAP7_75t_R _19952_ (.A1(_11604_),
    .A2(_11611_),
    .B(_11532_),
    .Y(_11612_));
 NAND2x1_ASAP7_75t_R _19953_ (.A(_11600_),
    .B(_11612_),
    .Y(_11613_));
 OAI21x1_ASAP7_75t_R _19954_ (.A1(_11521_),
    .A2(_11522_),
    .B(_11431_),
    .Y(_11614_));
 AOI21x1_ASAP7_75t_R _19955_ (.A1(_11419_),
    .A2(_11421_),
    .B(_01160_),
    .Y(_11615_));
 NOR2x1_ASAP7_75t_R _19956_ (.A(net894),
    .B(_11528_),
    .Y(_11616_));
 AOI21x1_ASAP7_75t_R _19957_ (.A1(_11614_),
    .A2(_11616_),
    .B(_11520_),
    .Y(_11617_));
 AO21x2_ASAP7_75t_R _19958_ (.A1(_11421_),
    .A2(_11419_),
    .B(_01159_),
    .Y(_11618_));
 OAI21x1_ASAP7_75t_R _19959_ (.A1(_11519_),
    .A2(_11618_),
    .B(_11471_),
    .Y(_11619_));
 INVx1_ASAP7_75t_R _19960_ (.A(_11619_),
    .Y(_11620_));
 NAND2x2_ASAP7_75t_R _19961_ (.A(_11401_),
    .B(_11422_),
    .Y(_11621_));
 AO21x1_ASAP7_75t_R _19962_ (.A1(_11621_),
    .A2(_11572_),
    .B(_11561_),
    .Y(_11622_));
 NAND2x1_ASAP7_75t_R _19963_ (.A(_11620_),
    .B(_11622_),
    .Y(_11623_));
 BUFx6f_ASAP7_75t_R _19964_ (.A(_11457_),
    .Y(_11624_));
 AO21x1_ASAP7_75t_R _19965_ (.A1(_11624_),
    .A2(_11594_),
    .B(_11471_),
    .Y(_11625_));
 NOR2x1_ASAP7_75t_R _19966_ (.A(_01164_),
    .B(_11561_),
    .Y(_11626_));
 OA21x2_ASAP7_75t_R _19967_ (.A1(_11625_),
    .A2(_11626_),
    .B(_11585_),
    .Y(_11627_));
 OAI21x1_ASAP7_75t_R _19968_ (.A1(_11617_),
    .A2(_11623_),
    .B(_11627_),
    .Y(_11628_));
 AO21x1_ASAP7_75t_R _19969_ (.A1(_11624_),
    .A2(net894),
    .B(_11506_),
    .Y(_11629_));
 AO21x1_ASAP7_75t_R _19970_ (.A1(_11515_),
    .A2(_11529_),
    .B(_11629_),
    .Y(_11630_));
 AOI21x1_ASAP7_75t_R _19971_ (.A1(_11615_),
    .A2(_11524_),
    .B(_11605_),
    .Y(_11631_));
 NOR2x2_ASAP7_75t_R _19972_ (.A(_11461_),
    .B(_11457_),
    .Y(_11632_));
 AO21x2_ASAP7_75t_R _19973_ (.A1(_11429_),
    .A2(_11427_),
    .B(_01161_),
    .Y(_11633_));
 NOR2x2_ASAP7_75t_R _19974_ (.A(_11480_),
    .B(_11633_),
    .Y(_11634_));
 NOR2x1_ASAP7_75t_R _19975_ (.A(_11632_),
    .B(_11634_),
    .Y(_11635_));
 AOI21x1_ASAP7_75t_R _19976_ (.A1(net898),
    .A2(_11635_),
    .B(_11585_),
    .Y(_11636_));
 AOI21x1_ASAP7_75t_R _19977_ (.A1(_11630_),
    .A2(_11636_),
    .B(_11494_),
    .Y(_11637_));
 AOI21x1_ASAP7_75t_R _19978_ (.A1(_11628_),
    .A2(_11637_),
    .B(_11545_),
    .Y(_11638_));
 NAND2x1_ASAP7_75t_R _19979_ (.A(_11613_),
    .B(_11638_),
    .Y(_11639_));
 OAI21x1_ASAP7_75t_R _19980_ (.A1(_11546_),
    .A2(_11588_),
    .B(_11639_),
    .Y(_00040_));
 BUFx6f_ASAP7_75t_R _19981_ (.A(_11458_),
    .Y(_11640_));
 AOI21x1_ASAP7_75t_R _19982_ (.A1(_15831_),
    .A2(_11552_),
    .B(net509),
    .Y(_11641_));
 AO21x1_ASAP7_75t_R _19983_ (.A1(_11429_),
    .A2(_11427_),
    .B(_01160_),
    .Y(_11642_));
 OA21x2_ASAP7_75t_R _19984_ (.A1(_11642_),
    .A2(_11519_),
    .B(_11471_),
    .Y(_11643_));
 OAI21x1_ASAP7_75t_R _19985_ (.A1(_11641_),
    .A2(_11640_),
    .B(_11643_),
    .Y(_11644_));
 NAND2x2_ASAP7_75t_R _19986_ (.A(_15818_),
    .B(_11430_),
    .Y(_11645_));
 INVx1_ASAP7_75t_R _19987_ (.A(_11645_),
    .Y(_11646_));
 OAI21x1_ASAP7_75t_R _19988_ (.A1(_11513_),
    .A2(_11646_),
    .B(_11589_),
    .Y(_11647_));
 AOI21x1_ASAP7_75t_R _19989_ (.A1(_11614_),
    .A2(_11459_),
    .B(_11605_),
    .Y(_11648_));
 AOI21x1_ASAP7_75t_R _19990_ (.A1(_11647_),
    .A2(_11648_),
    .B(_11531_),
    .Y(_11649_));
 AOI21x1_ASAP7_75t_R _19991_ (.A1(_11649_),
    .A2(_11644_),
    .B(_11585_),
    .Y(_11650_));
 INVx2_ASAP7_75t_R _19992_ (.A(net893),
    .Y(_11651_));
 AO21x1_ASAP7_75t_R _19993_ (.A1(_11651_),
    .A2(_11462_),
    .B(_11624_),
    .Y(_11652_));
 AO21x1_ASAP7_75t_R _19994_ (.A1(_11621_),
    .A2(_11572_),
    .B(_11519_),
    .Y(_11653_));
 BUFx6f_ASAP7_75t_R _19995_ (.A(_11471_),
    .Y(_11654_));
 AOI21x1_ASAP7_75t_R _19996_ (.A1(_11653_),
    .A2(_11652_),
    .B(_11654_),
    .Y(_11655_));
 NOR2x2_ASAP7_75t_R _19997_ (.A(_11480_),
    .B(_11594_),
    .Y(_11656_));
 NAND2x1_ASAP7_75t_R _19998_ (.A(_11645_),
    .B(_11656_),
    .Y(_11657_));
 NAND2x2_ASAP7_75t_R _19999_ (.A(_11511_),
    .B(_11512_),
    .Y(_15819_));
 NAND2x2_ASAP7_75t_R _20000_ (.A(_15823_),
    .B(net4),
    .Y(_11658_));
 NAND2x1_ASAP7_75t_R _20001_ (.A(_11658_),
    .B(_11515_),
    .Y(_11659_));
 AOI21x1_ASAP7_75t_R _20002_ (.A1(_11657_),
    .A2(_11659_),
    .B(_11598_),
    .Y(_11660_));
 OAI21x1_ASAP7_75t_R _20003_ (.A1(_11655_),
    .A2(_11660_),
    .B(_11576_),
    .Y(_11661_));
 NAND2x1_ASAP7_75t_R _20004_ (.A(_11661_),
    .B(_11650_),
    .Y(_11662_));
 INVx3_ASAP7_75t_R _20005_ (.A(_11621_),
    .Y(_11663_));
 AO21x2_ASAP7_75t_R _20006_ (.A1(_11432_),
    .A2(_01160_),
    .B(_11445_),
    .Y(_11664_));
 NAND2x2_ASAP7_75t_R _20007_ (.A(_15818_),
    .B(_11422_),
    .Y(_11665_));
 AOI21x1_ASAP7_75t_R _20008_ (.A1(_11665_),
    .A2(_11632_),
    .B(_11472_),
    .Y(_11666_));
 OA21x2_ASAP7_75t_R _20009_ (.A1(_11663_),
    .A2(_11664_),
    .B(_11666_),
    .Y(_11667_));
 NAND2x1_ASAP7_75t_R _20010_ (.A(_15818_),
    .B(net4),
    .Y(_11668_));
 AOI21x1_ASAP7_75t_R _20011_ (.A1(_11668_),
    .A2(_11596_),
    .B(_11507_),
    .Y(_11669_));
 NOR2x2_ASAP7_75t_R _20012_ (.A(_11431_),
    .B(_11458_),
    .Y(_11670_));
 NAND2x1_ASAP7_75t_R _20013_ (.A(_11670_),
    .B(_11607_),
    .Y(_11671_));
 AO21x1_ASAP7_75t_R _20014_ (.A1(_11669_),
    .A2(_11671_),
    .B(_11576_),
    .Y(_11672_));
 AOI21x1_ASAP7_75t_R _20015_ (.A1(_15828_),
    .A2(_11607_),
    .B(net895),
    .Y(_11673_));
 AOI21x1_ASAP7_75t_R _20016_ (.A1(_11517_),
    .A2(_11580_),
    .B(_11507_),
    .Y(_11674_));
 OAI21x1_ASAP7_75t_R _20017_ (.A1(_11520_),
    .A2(_11673_),
    .B(_11674_),
    .Y(_11675_));
 OAI21x1_ASAP7_75t_R _20018_ (.A1(_11449_),
    .A2(_11452_),
    .B(_11456_),
    .Y(_11676_));
 AOI21x1_ASAP7_75t_R _20019_ (.A1(_11676_),
    .A2(_11510_),
    .B(_11513_),
    .Y(_11677_));
 AOI21x1_ASAP7_75t_R _20020_ (.A1(net898),
    .A2(_11677_),
    .B(_11493_),
    .Y(_11678_));
 AOI21x1_ASAP7_75t_R _20021_ (.A1(_11675_),
    .A2(_11678_),
    .B(_11503_),
    .Y(_11679_));
 OAI21x1_ASAP7_75t_R _20022_ (.A1(_11667_),
    .A2(_11672_),
    .B(_11679_),
    .Y(_11680_));
 AOI21x1_ASAP7_75t_R _20023_ (.A1(_11680_),
    .A2(_11662_),
    .B(_11545_),
    .Y(_11681_));
 INVx1_ASAP7_75t_R _20024_ (.A(_11676_),
    .Y(_11682_));
 OAI21x1_ASAP7_75t_R _20025_ (.A1(_11682_),
    .A2(_11548_),
    .B(_11531_),
    .Y(_11683_));
 AOI21x1_ASAP7_75t_R _20026_ (.A1(_11523_),
    .A2(_11481_),
    .B(_11605_),
    .Y(_11684_));
 INVx1_ASAP7_75t_R _20027_ (.A(_11684_),
    .Y(_11685_));
 OAI21x1_ASAP7_75t_R _20028_ (.A1(_11683_),
    .A2(_11685_),
    .B(_11585_),
    .Y(_11686_));
 AO21x1_ASAP7_75t_R _20029_ (.A1(_11529_),
    .A2(_11609_),
    .B(_11507_),
    .Y(_11687_));
 AOI21x1_ASAP7_75t_R _20030_ (.A1(_11670_),
    .A2(_11607_),
    .B(_11605_),
    .Y(_11688_));
 OAI21x1_ASAP7_75t_R _20031_ (.A1(_11559_),
    .A2(_11528_),
    .B(_11561_),
    .Y(_11689_));
 NOR2x1_ASAP7_75t_R _20032_ (.A(_11422_),
    .B(_11458_),
    .Y(_11690_));
 NAND2x1_ASAP7_75t_R _20033_ (.A(_11690_),
    .B(_11552_),
    .Y(_11691_));
 NAND3x1_ASAP7_75t_R _20034_ (.A(_11688_),
    .B(_11689_),
    .C(_11691_),
    .Y(_11692_));
 AO21x1_ASAP7_75t_R _20035_ (.A1(_00505_),
    .A2(_11445_),
    .B(_11506_),
    .Y(_11693_));
 AND2x2_ASAP7_75t_R _20036_ (.A(_11693_),
    .B(_11531_),
    .Y(_11694_));
 AOI21x1_ASAP7_75t_R _20037_ (.A1(_11687_),
    .A2(_11692_),
    .B(_11694_),
    .Y(_11695_));
 OAI21x1_ASAP7_75t_R _20038_ (.A1(_11686_),
    .A2(_11695_),
    .B(_11544_),
    .Y(_11696_));
 AO21x1_ASAP7_75t_R _20039_ (.A1(_11572_),
    .A2(_11595_),
    .B(_11624_),
    .Y(_11697_));
 OAI21x1_ASAP7_75t_R _20040_ (.A1(_11525_),
    .A2(_11663_),
    .B(_11589_),
    .Y(_11698_));
 AOI21x1_ASAP7_75t_R _20041_ (.A1(_11697_),
    .A2(_11698_),
    .B(_11654_),
    .Y(_11699_));
 NAND2x1_ASAP7_75t_R _20042_ (.A(_11523_),
    .B(_11481_),
    .Y(_11700_));
 AO21x1_ASAP7_75t_R _20043_ (.A1(_11645_),
    .A2(_11560_),
    .B(_11577_),
    .Y(_11701_));
 AOI21x1_ASAP7_75t_R _20044_ (.A1(_11700_),
    .A2(_11701_),
    .B(_11598_),
    .Y(_11702_));
 OAI21x1_ASAP7_75t_R _20045_ (.A1(_11699_),
    .A2(_11702_),
    .B(_11564_),
    .Y(_11703_));
 NOR2x2_ASAP7_75t_R _20046_ (.A(_11401_),
    .B(_11430_),
    .Y(_11704_));
 NOR2x1_ASAP7_75t_R _20047_ (.A(_11445_),
    .B(_11704_),
    .Y(_11705_));
 AOI21x1_ASAP7_75t_R _20048_ (.A1(_11529_),
    .A2(_11705_),
    .B(_11632_),
    .Y(_11706_));
 NAND2x1_ASAP7_75t_R _20049_ (.A(_11654_),
    .B(_11706_),
    .Y(_11707_));
 AOI21x1_ASAP7_75t_R _20050_ (.A1(_11427_),
    .A2(_11429_),
    .B(_01162_),
    .Y(_11708_));
 INVx1_ASAP7_75t_R _20051_ (.A(_11708_),
    .Y(_11709_));
 NAND2x1_ASAP7_75t_R _20052_ (.A(_11709_),
    .B(_11618_),
    .Y(_11710_));
 AOI21x1_ASAP7_75t_R _20053_ (.A1(_11589_),
    .A2(_11710_),
    .B(_11472_),
    .Y(_11711_));
 AOI21x1_ASAP7_75t_R _20054_ (.A1(_15823_),
    .A2(net564),
    .B(_11432_),
    .Y(_11712_));
 OAI21x1_ASAP7_75t_R _20055_ (.A1(net509),
    .A2(_11712_),
    .B(_11510_),
    .Y(_11713_));
 AOI21x1_ASAP7_75t_R _20056_ (.A1(_11711_),
    .A2(_11713_),
    .B(_11493_),
    .Y(_11714_));
 NAND2x1_ASAP7_75t_R _20057_ (.A(_11714_),
    .B(_11707_),
    .Y(_11715_));
 AOI21x1_ASAP7_75t_R _20058_ (.A1(_11703_),
    .A2(_11715_),
    .B(_11586_),
    .Y(_11716_));
 NOR2x1_ASAP7_75t_R _20059_ (.A(_11696_),
    .B(_11716_),
    .Y(_11717_));
 NOR2x1_ASAP7_75t_R _20060_ (.A(_11717_),
    .B(_11681_),
    .Y(_00041_));
 AO21x1_ASAP7_75t_R _20061_ (.A1(_11568_),
    .A2(_11651_),
    .B(_11624_),
    .Y(_11718_));
 NAND2x1_ASAP7_75t_R _20062_ (.A(_11457_),
    .B(_11571_),
    .Y(_11719_));
 INVx1_ASAP7_75t_R _20063_ (.A(_11719_),
    .Y(_11720_));
 NOR2x1_ASAP7_75t_R _20064_ (.A(_11491_),
    .B(_11720_),
    .Y(_11721_));
 BUFx4f_ASAP7_75t_R _20065_ (.A(_11506_),
    .Y(_11722_));
 AOI21x1_ASAP7_75t_R _20066_ (.A1(_11718_),
    .A2(_11721_),
    .B(_11722_),
    .Y(_11723_));
 OAI21x1_ASAP7_75t_R _20067_ (.A1(net4),
    .A2(_11665_),
    .B(_11524_),
    .Y(_11724_));
 NAND2x1_ASAP7_75t_R _20068_ (.A(_00506_),
    .B(_11519_),
    .Y(_11725_));
 NAND3x1_ASAP7_75t_R _20069_ (.A(_11724_),
    .B(_11531_),
    .C(_11725_),
    .Y(_11726_));
 AOI21x1_ASAP7_75t_R _20070_ (.A1(_11723_),
    .A2(_11726_),
    .B(_11503_),
    .Y(_11727_));
 AO21x1_ASAP7_75t_R _20071_ (.A1(_11529_),
    .A2(_11609_),
    .B(_11531_),
    .Y(_11728_));
 AND2x4_ASAP7_75t_R _20072_ (.A(net505),
    .B(_01159_),
    .Y(_11729_));
 NAND2x2_ASAP7_75t_R _20073_ (.A(_11431_),
    .B(_11729_),
    .Y(_11730_));
 OA211x2_ASAP7_75t_R _20074_ (.A1(_11552_),
    .A2(_15828_),
    .B(_11577_),
    .C(_11730_),
    .Y(_11731_));
 OA21x2_ASAP7_75t_R _20075_ (.A1(_01166_),
    .A2(_11519_),
    .B(_11491_),
    .Y(_11732_));
 OAI21x1_ASAP7_75t_R _20076_ (.A1(_15818_),
    .A2(_11432_),
    .B(_11380_),
    .Y(_11733_));
 NAND2x1_ASAP7_75t_R _20077_ (.A(_11573_),
    .B(_11733_),
    .Y(_11734_));
 AOI21x1_ASAP7_75t_R _20078_ (.A1(_11732_),
    .A2(_11734_),
    .B(_11654_),
    .Y(_11735_));
 OAI21x1_ASAP7_75t_R _20079_ (.A1(_11728_),
    .A2(_11731_),
    .B(_11735_),
    .Y(_11736_));
 NAND2x1_ASAP7_75t_R _20080_ (.A(_11727_),
    .B(_11736_),
    .Y(_11737_));
 OA21x2_ASAP7_75t_R _20081_ (.A1(_01164_),
    .A2(_11519_),
    .B(_11471_),
    .Y(_11738_));
 OAI21x1_ASAP7_75t_R _20082_ (.A1(_15831_),
    .A2(_11607_),
    .B(_11580_),
    .Y(_11739_));
 AOI21x1_ASAP7_75t_R _20083_ (.A1(_11738_),
    .A2(_11739_),
    .B(_11531_),
    .Y(_11740_));
 AOI21x1_ASAP7_75t_R _20084_ (.A1(_11456_),
    .A2(net4),
    .B(_11458_),
    .Y(_11741_));
 NAND2x1_ASAP7_75t_R _20085_ (.A(_11645_),
    .B(_11741_),
    .Y(_11742_));
 AOI21x1_ASAP7_75t_R _20086_ (.A1(_11595_),
    .A2(_11596_),
    .B(_11605_),
    .Y(_11743_));
 NAND2x1_ASAP7_75t_R _20087_ (.A(_11742_),
    .B(_11743_),
    .Y(_11744_));
 AOI21x1_ASAP7_75t_R _20088_ (.A1(_11740_),
    .A2(_11744_),
    .B(_11585_),
    .Y(_11745_));
 AND3x1_ASAP7_75t_R _20089_ (.A(_11557_),
    .B(_11595_),
    .C(_11519_),
    .Y(_11746_));
 AOI21x1_ASAP7_75t_R _20090_ (.A1(_11372_),
    .A2(_11379_),
    .B(_11456_),
    .Y(_11747_));
 NOR3x1_ASAP7_75t_R _20091_ (.A(_11747_),
    .B(_11577_),
    .C(_11559_),
    .Y(_11748_));
 OAI21x1_ASAP7_75t_R _20092_ (.A1(_11746_),
    .A2(_11748_),
    .B(_11598_),
    .Y(_11749_));
 AOI21x1_ASAP7_75t_R _20093_ (.A1(_11432_),
    .A2(_11380_),
    .B(_11624_),
    .Y(_11750_));
 AND2x2_ASAP7_75t_R _20094_ (.A(_11458_),
    .B(_00505_),
    .Y(_11751_));
 AOI21x1_ASAP7_75t_R _20095_ (.A1(_11668_),
    .A2(_11750_),
    .B(_11751_),
    .Y(_11752_));
 AOI21x1_ASAP7_75t_R _20096_ (.A1(_11475_),
    .A2(_11752_),
    .B(_11493_),
    .Y(_11753_));
 NAND2x1_ASAP7_75t_R _20097_ (.A(_11749_),
    .B(_11753_),
    .Y(_11754_));
 NAND2x1_ASAP7_75t_R _20098_ (.A(_11745_),
    .B(_11754_),
    .Y(_11755_));
 AOI21x1_ASAP7_75t_R _20099_ (.A1(_11737_),
    .A2(_11755_),
    .B(_11545_),
    .Y(_11756_));
 NAND2x1_ASAP7_75t_R _20100_ (.A(_11632_),
    .B(_11595_),
    .Y(_11757_));
 OA21x2_ASAP7_75t_R _20101_ (.A1(_11431_),
    .A2(_11601_),
    .B(_11458_),
    .Y(_11758_));
 NAND2x1_ASAP7_75t_R _20102_ (.A(_11645_),
    .B(_11758_),
    .Y(_11759_));
 AOI21x1_ASAP7_75t_R _20103_ (.A1(_11759_),
    .A2(_11757_),
    .B(_11722_),
    .Y(_11760_));
 NOR2x2_ASAP7_75t_R _20104_ (.A(_01161_),
    .B(_11456_),
    .Y(_11761_));
 AOI211x1_ASAP7_75t_R _20105_ (.A1(net4),
    .A2(_15831_),
    .B(_11761_),
    .C(_11561_),
    .Y(_11762_));
 AO21x2_ASAP7_75t_R _20106_ (.A1(_11421_),
    .A2(_11419_),
    .B(_01162_),
    .Y(_11763_));
 NAND2x1_ASAP7_75t_R _20107_ (.A(_11624_),
    .B(_11763_),
    .Y(_11764_));
 OAI21x1_ASAP7_75t_R _20108_ (.A1(_11528_),
    .A2(_11764_),
    .B(_11506_),
    .Y(_11765_));
 OAI21x1_ASAP7_75t_R _20109_ (.A1(_11762_),
    .A2(_11765_),
    .B(_11493_),
    .Y(_11766_));
 NOR2x1_ASAP7_75t_R _20110_ (.A(_11766_),
    .B(_11760_),
    .Y(_11767_));
 AOI21x1_ASAP7_75t_R _20111_ (.A1(_11573_),
    .A2(_11747_),
    .B(net893),
    .Y(_11768_));
 NOR2x1_ASAP7_75t_R _20112_ (.A(_11493_),
    .B(_11634_),
    .Y(_11769_));
 OAI21x1_ASAP7_75t_R _20113_ (.A1(_11598_),
    .A2(_11768_),
    .B(_11769_),
    .Y(_11770_));
 OR3x1_ASAP7_75t_R _20114_ (.A(_11519_),
    .B(_11432_),
    .C(_01162_),
    .Y(_11771_));
 OA21x2_ASAP7_75t_R _20115_ (.A1(_11431_),
    .A2(_11479_),
    .B(_11480_),
    .Y(_11772_));
 NAND2x1_ASAP7_75t_R _20116_ (.A(_11645_),
    .B(_11772_),
    .Y(_11773_));
 AOI21x1_ASAP7_75t_R _20117_ (.A1(_11771_),
    .A2(_11773_),
    .B(_11654_),
    .Y(_11774_));
 OAI21x1_ASAP7_75t_R _20118_ (.A1(_11770_),
    .A2(_11774_),
    .B(_11503_),
    .Y(_11775_));
 OAI21x1_ASAP7_75t_R _20119_ (.A1(_11775_),
    .A2(_11767_),
    .B(_11544_),
    .Y(_11776_));
 OAI21x1_ASAP7_75t_R _20120_ (.A1(_11594_),
    .A2(_11747_),
    .B(_11561_),
    .Y(_11777_));
 NAND2x1_ASAP7_75t_R _20121_ (.A(_11592_),
    .B(_11651_),
    .Y(_11778_));
 OAI21x1_ASAP7_75t_R _20122_ (.A1(_11513_),
    .A2(_11778_),
    .B(_11573_),
    .Y(_11779_));
 AOI21x1_ASAP7_75t_R _20123_ (.A1(_11779_),
    .A2(_11777_),
    .B(_11722_),
    .Y(_11780_));
 AOI21x1_ASAP7_75t_R _20124_ (.A1(_11763_),
    .A2(_11642_),
    .B(_11445_),
    .Y(_11781_));
 AOI21x1_ASAP7_75t_R _20125_ (.A1(_11573_),
    .A2(_11733_),
    .B(_11781_),
    .Y(_11782_));
 OAI21x1_ASAP7_75t_R _20126_ (.A1(_11654_),
    .A2(_11782_),
    .B(_11531_),
    .Y(_11783_));
 NOR2x1_ASAP7_75t_R _20127_ (.A(_11783_),
    .B(_11780_),
    .Y(_11784_));
 INVx2_ASAP7_75t_R _20128_ (.A(_11523_),
    .Y(_11785_));
 NAND2x2_ASAP7_75t_R _20129_ (.A(_11458_),
    .B(_11568_),
    .Y(_11786_));
 NOR2x1_ASAP7_75t_R _20130_ (.A(_11785_),
    .B(_11786_),
    .Y(_11787_));
 NAND2x1_ASAP7_75t_R _20131_ (.A(_11519_),
    .B(_11618_),
    .Y(_11788_));
 OAI21x1_ASAP7_75t_R _20132_ (.A1(_11528_),
    .A2(_11788_),
    .B(_11507_),
    .Y(_11789_));
 OAI21x1_ASAP7_75t_R _20133_ (.A1(_11787_),
    .A2(_11789_),
    .B(_11493_),
    .Y(_11790_));
 OAI21x1_ASAP7_75t_R _20134_ (.A1(_11708_),
    .A2(_11712_),
    .B(_11510_),
    .Y(_11791_));
 AOI21x1_ASAP7_75t_R _20135_ (.A1(_11724_),
    .A2(_11791_),
    .B(_11598_),
    .Y(_11792_));
 OAI21x1_ASAP7_75t_R _20136_ (.A1(_11790_),
    .A2(_11792_),
    .B(_11585_),
    .Y(_11793_));
 NOR2x1_ASAP7_75t_R _20137_ (.A(_11793_),
    .B(_11784_),
    .Y(_11794_));
 NOR2x1_ASAP7_75t_R _20138_ (.A(_11776_),
    .B(_11794_),
    .Y(_11795_));
 NOR2x1_ASAP7_75t_R _20139_ (.A(_11756_),
    .B(_11795_),
    .Y(_00042_));
 NOR2x1_ASAP7_75t_R _20140_ (.A(_11528_),
    .B(_11764_),
    .Y(_11796_));
 AO21x1_ASAP7_75t_R _20141_ (.A1(_11796_),
    .A2(_11582_),
    .B(_11564_),
    .Y(_11797_));
 AOI21x1_ASAP7_75t_R _20142_ (.A1(_15828_),
    .A2(_11729_),
    .B(_11602_),
    .Y(_11798_));
 AOI211x1_ASAP7_75t_R _20143_ (.A1(_11529_),
    .A2(_11609_),
    .B(_11798_),
    .C(_11582_),
    .Y(_11799_));
 OAI21x1_ASAP7_75t_R _20144_ (.A1(_11797_),
    .A2(_11799_),
    .B(_11503_),
    .Y(_11800_));
 NOR2x1_ASAP7_75t_R _20145_ (.A(_11516_),
    .B(_11432_),
    .Y(_11801_));
 INVx1_ASAP7_75t_R _20146_ (.A(_11801_),
    .Y(_11802_));
 OA21x2_ASAP7_75t_R _20147_ (.A1(_11704_),
    .A2(_11761_),
    .B(_11573_),
    .Y(_11803_));
 BUFx6f_ASAP7_75t_R _20148_ (.A(_11605_),
    .Y(_11804_));
 AOI211x1_ASAP7_75t_R _20149_ (.A1(_11554_),
    .A2(_11802_),
    .B(_11803_),
    .C(_11804_),
    .Y(_11805_));
 AO21x1_ASAP7_75t_R _20150_ (.A1(_11669_),
    .A2(_11622_),
    .B(_11531_),
    .Y(_11806_));
 NOR2x1_ASAP7_75t_R _20151_ (.A(_11805_),
    .B(_11806_),
    .Y(_11807_));
 NOR2x1_ASAP7_75t_R _20152_ (.A(_11800_),
    .B(_11807_),
    .Y(_11808_));
 NAND2x1_ASAP7_75t_R _20153_ (.A(_11458_),
    .B(_11461_),
    .Y(_11809_));
 AO21x1_ASAP7_75t_R _20154_ (.A1(_11606_),
    .A2(_11809_),
    .B(_11576_),
    .Y(_11810_));
 OA21x2_ASAP7_75t_R _20155_ (.A1(_11633_),
    .A2(_11524_),
    .B(_11605_),
    .Y(_11811_));
 AND2x2_ASAP7_75t_R _20156_ (.A(_11759_),
    .B(_11811_),
    .Y(_11812_));
 OAI21x1_ASAP7_75t_R _20157_ (.A1(_11810_),
    .A2(_11812_),
    .B(_11586_),
    .Y(_11813_));
 NOR2x2_ASAP7_75t_R _20158_ (.A(net510),
    .B(_11477_),
    .Y(_11814_));
 AO21x1_ASAP7_75t_R _20159_ (.A1(_11459_),
    .A2(_11730_),
    .B(_11722_),
    .Y(_11815_));
 OAI21x1_ASAP7_75t_R _20160_ (.A1(_11814_),
    .A2(_11815_),
    .B(_11576_),
    .Y(_11816_));
 INVx1_ASAP7_75t_R _20161_ (.A(_11747_),
    .Y(_11817_));
 INVx1_ASAP7_75t_R _20162_ (.A(_11670_),
    .Y(_11818_));
 OAI21x1_ASAP7_75t_R _20163_ (.A1(_11460_),
    .A2(_11818_),
    .B(_11606_),
    .Y(_11819_));
 AOI21x1_ASAP7_75t_R _20164_ (.A1(_11817_),
    .A2(_11609_),
    .B(_11819_),
    .Y(_11820_));
 NOR2x1_ASAP7_75t_R _20165_ (.A(_11816_),
    .B(_11820_),
    .Y(_11821_));
 OAI21x1_ASAP7_75t_R _20166_ (.A1(_11813_),
    .A2(_11821_),
    .B(_11545_),
    .Y(_11822_));
 OAI21x1_ASAP7_75t_R _20167_ (.A1(_15828_),
    .A2(_15821_),
    .B(_11573_),
    .Y(_11823_));
 NAND2x1_ASAP7_75t_R _20168_ (.A(_11557_),
    .B(_11621_),
    .Y(_11824_));
 NOR2x1_ASAP7_75t_R _20169_ (.A(_11823_),
    .B(_11824_),
    .Y(_11825_));
 NAND2x1_ASAP7_75t_R _20170_ (.A(_15828_),
    .B(_11552_),
    .Y(_11826_));
 AO21x1_ASAP7_75t_R _20171_ (.A1(_11826_),
    .A2(_11656_),
    .B(_11582_),
    .Y(_11827_));
 AOI21x1_ASAP7_75t_R _20172_ (.A1(_11570_),
    .A2(_11554_),
    .B(_11475_),
    .Y(_11828_));
 AOI21x1_ASAP7_75t_R _20173_ (.A1(_11828_),
    .A2(_11550_),
    .B(_11585_),
    .Y(_11829_));
 OAI21x1_ASAP7_75t_R _20174_ (.A1(_11825_),
    .A2(_11827_),
    .B(_11829_),
    .Y(_11830_));
 OAI21x1_ASAP7_75t_R _20175_ (.A1(_11785_),
    .A2(_11786_),
    .B(_11475_),
    .Y(_11831_));
 AND2x2_ASAP7_75t_R _20176_ (.A(_11772_),
    .B(_11517_),
    .Y(_11832_));
 NOR2x1_ASAP7_75t_R _20177_ (.A(_11831_),
    .B(_11832_),
    .Y(_11833_));
 BUFx6f_ASAP7_75t_R _20178_ (.A(_11624_),
    .Y(_11834_));
 OA21x2_ASAP7_75t_R _20179_ (.A1(net757),
    .A2(_11571_),
    .B(_11549_),
    .Y(_11835_));
 AOI211x1_ASAP7_75t_R _20180_ (.A1(_11824_),
    .A2(_11834_),
    .B(_11835_),
    .C(_11804_),
    .Y(_11836_));
 OAI21x1_ASAP7_75t_R _20181_ (.A1(_11833_),
    .A2(_11836_),
    .B(_11586_),
    .Y(_11837_));
 AOI21x1_ASAP7_75t_R _20182_ (.A1(_11830_),
    .A2(_11837_),
    .B(_11532_),
    .Y(_11838_));
 AO21x1_ASAP7_75t_R _20183_ (.A1(_11421_),
    .A2(_11419_),
    .B(_01161_),
    .Y(_11839_));
 AO21x1_ASAP7_75t_R _20184_ (.A1(_11839_),
    .A2(_11462_),
    .B(_11577_),
    .Y(_11840_));
 AND2x2_ASAP7_75t_R _20185_ (.A(_11648_),
    .B(_11840_),
    .Y(_11841_));
 AOI21x1_ASAP7_75t_R _20186_ (.A1(_11592_),
    .A2(_11607_),
    .B(_11690_),
    .Y(_11842_));
 AO21x1_ASAP7_75t_R _20187_ (.A1(_11842_),
    .A2(_11475_),
    .B(_11585_),
    .Y(_11843_));
 NOR2x1_ASAP7_75t_R _20188_ (.A(_11843_),
    .B(_11841_),
    .Y(_11844_));
 OAI21x1_ASAP7_75t_R _20189_ (.A1(_11834_),
    .A2(net757),
    .B(_11582_),
    .Y(_11845_));
 NOR2x1_ASAP7_75t_R _20190_ (.A(_11785_),
    .B(_11446_),
    .Y(_11846_));
 OAI21x1_ASAP7_75t_R _20191_ (.A1(_11845_),
    .A2(_11846_),
    .B(_11586_),
    .Y(_11847_));
 INVx1_ASAP7_75t_R _20192_ (.A(_11453_),
    .Y(_11848_));
 NOR2x1_ASAP7_75t_R _20193_ (.A(_11848_),
    .B(_11548_),
    .Y(_11849_));
 AO21x1_ASAP7_75t_R _20194_ (.A1(_11523_),
    .A2(_11632_),
    .B(_11722_),
    .Y(_11850_));
 NOR2x1_ASAP7_75t_R _20195_ (.A(_11849_),
    .B(_11850_),
    .Y(_11851_));
 OAI21x1_ASAP7_75t_R _20196_ (.A1(_11847_),
    .A2(_11851_),
    .B(_11532_),
    .Y(_11852_));
 INVx3_ASAP7_75t_R _20197_ (.A(_11544_),
    .Y(_11853_));
 OAI21x1_ASAP7_75t_R _20198_ (.A1(_11844_),
    .A2(_11852_),
    .B(_11853_),
    .Y(_11854_));
 OAI22x1_ASAP7_75t_R _20199_ (.A1(_11808_),
    .A2(_11822_),
    .B1(_11854_),
    .B2(_11838_),
    .Y(_00043_));
 OAI21x1_ASAP7_75t_R _20200_ (.A1(_11708_),
    .A2(_11594_),
    .B(_11640_),
    .Y(_11855_));
 NAND2x1_ASAP7_75t_R _20201_ (.A(_11475_),
    .B(_11855_),
    .Y(_11856_));
 AOI21x1_ASAP7_75t_R _20202_ (.A1(_15818_),
    .A2(_11747_),
    .B(_11602_),
    .Y(_11857_));
 AOI22x1_ASAP7_75t_R _20203_ (.A1(_11594_),
    .A2(_11510_),
    .B1(_11601_),
    .B2(_15828_),
    .Y(_11858_));
 NAND2x1_ASAP7_75t_R _20204_ (.A(_11631_),
    .B(_11858_),
    .Y(_11859_));
 OAI21x1_ASAP7_75t_R _20205_ (.A1(_11856_),
    .A2(_11857_),
    .B(_11859_),
    .Y(_11860_));
 AOI21x1_ASAP7_75t_R _20206_ (.A1(_11494_),
    .A2(_11860_),
    .B(_11504_),
    .Y(_11861_));
 OAI21x1_ASAP7_75t_R _20207_ (.A1(_11801_),
    .A2(_11664_),
    .B(_11598_),
    .Y(_11862_));
 NOR2x1_ASAP7_75t_R _20208_ (.A(_11823_),
    .B(_11603_),
    .Y(_11863_));
 NOR2x1_ASAP7_75t_R _20209_ (.A(_11862_),
    .B(_11863_),
    .Y(_11864_));
 AOI21x1_ASAP7_75t_R _20210_ (.A1(_15831_),
    .A2(net41),
    .B(_11571_),
    .Y(_11865_));
 OAI21x1_ASAP7_75t_R _20211_ (.A1(_11834_),
    .A2(_11865_),
    .B(_11475_),
    .Y(_11866_));
 NOR2x1_ASAP7_75t_R _20212_ (.A(_11866_),
    .B(_11617_),
    .Y(_11867_));
 OAI21x1_ASAP7_75t_R _20213_ (.A1(_11864_),
    .A2(_11867_),
    .B(_11532_),
    .Y(_11868_));
 AOI21x1_ASAP7_75t_R _20214_ (.A1(_11861_),
    .A2(_11868_),
    .B(_11545_),
    .Y(_11869_));
 AO21x1_ASAP7_75t_R _20215_ (.A1(_11523_),
    .A2(_11592_),
    .B(_11834_),
    .Y(_11870_));
 AND2x2_ASAP7_75t_R _20216_ (.A(_11689_),
    .B(_11475_),
    .Y(_11871_));
 NOR2x1_ASAP7_75t_R _20217_ (.A(_11525_),
    .B(_11472_),
    .Y(_11872_));
 AO21x1_ASAP7_75t_R _20218_ (.A1(_11872_),
    .A2(_11602_),
    .B(_11576_),
    .Y(_11873_));
 AOI21x1_ASAP7_75t_R _20219_ (.A1(_11870_),
    .A2(_11871_),
    .B(_11873_),
    .Y(_11874_));
 AOI21x1_ASAP7_75t_R _20220_ (.A1(_11607_),
    .A2(_11523_),
    .B(_11520_),
    .Y(_11875_));
 AO21x1_ASAP7_75t_R _20221_ (.A1(_15831_),
    .A2(_11558_),
    .B(_11524_),
    .Y(_11876_));
 NOR2x1_ASAP7_75t_R _20222_ (.A(_11513_),
    .B(_11876_),
    .Y(_11877_));
 OAI21x1_ASAP7_75t_R _20223_ (.A1(_11875_),
    .A2(_11877_),
    .B(_11508_),
    .Y(_11878_));
 NOR2x1_ASAP7_75t_R _20224_ (.A(_11682_),
    .B(_11548_),
    .Y(_11879_));
 AOI21x1_ASAP7_75t_R _20225_ (.A1(_11676_),
    .A2(_11658_),
    .B(_11640_),
    .Y(_11880_));
 OAI21x1_ASAP7_75t_R _20226_ (.A1(_11879_),
    .A2(_11880_),
    .B(_11804_),
    .Y(_11881_));
 AOI21x1_ASAP7_75t_R _20227_ (.A1(_11878_),
    .A2(_11881_),
    .B(_11494_),
    .Y(_11882_));
 OAI21x1_ASAP7_75t_R _20228_ (.A1(_11874_),
    .A2(_11882_),
    .B(_11504_),
    .Y(_11883_));
 OAI21x1_ASAP7_75t_R _20229_ (.A1(_00507_),
    .A2(_11549_),
    .B(_11654_),
    .Y(_11884_));
 NOR2x1_ASAP7_75t_R _20230_ (.A(_11589_),
    .B(_11595_),
    .Y(_11885_));
 OA21x2_ASAP7_75t_R _20231_ (.A1(_11884_),
    .A2(_11885_),
    .B(_11564_),
    .Y(_11886_));
 NOR2x2_ASAP7_75t_R _20232_ (.A(_11602_),
    .B(_11513_),
    .Y(_11887_));
 AOI21x1_ASAP7_75t_R _20233_ (.A1(_11592_),
    .A2(_11614_),
    .B(_11520_),
    .Y(_11888_));
 OAI21x1_ASAP7_75t_R _20234_ (.A1(_11887_),
    .A2(_11888_),
    .B(_11508_),
    .Y(_11889_));
 AOI21x1_ASAP7_75t_R _20235_ (.A1(_11886_),
    .A2(_11889_),
    .B(_11504_),
    .Y(_11890_));
 NOR2x1_ASAP7_75t_R _20236_ (.A(_11528_),
    .B(_11602_),
    .Y(_11891_));
 OAI21x1_ASAP7_75t_R _20237_ (.A1(_15828_),
    .A2(net41),
    .B(_11640_),
    .Y(_11892_));
 OAI21x1_ASAP7_75t_R _20238_ (.A1(_11848_),
    .A2(_11892_),
    .B(_11598_),
    .Y(_11893_));
 NOR2x1_ASAP7_75t_R _20239_ (.A(_11891_),
    .B(_11893_),
    .Y(_11894_));
 OAI21x1_ASAP7_75t_R _20240_ (.A1(_15823_),
    .A2(net4),
    .B(_11577_),
    .Y(_11895_));
 OAI21x1_ASAP7_75t_R _20241_ (.A1(_11663_),
    .A2(_11895_),
    .B(_11590_),
    .Y(_11896_));
 NOR2x1_ASAP7_75t_R _20242_ (.A(_11508_),
    .B(_11896_),
    .Y(_11897_));
 OAI21x1_ASAP7_75t_R _20243_ (.A1(_11894_),
    .A2(_11897_),
    .B(_11532_),
    .Y(_11898_));
 AOI21x1_ASAP7_75t_R _20244_ (.A1(_11890_),
    .A2(_11898_),
    .B(_11853_),
    .Y(_11899_));
 INVx1_ASAP7_75t_R _20245_ (.A(_01159_),
    .Y(_11900_));
 AO21x1_ASAP7_75t_R _20246_ (.A1(_11421_),
    .A2(_11419_),
    .B(_11900_),
    .Y(_11901_));
 AO21x1_ASAP7_75t_R _20247_ (.A1(_11901_),
    .A2(_11640_),
    .B(_11472_),
    .Y(_11902_));
 OA21x2_ASAP7_75t_R _20248_ (.A1(_11676_),
    .A2(_15818_),
    .B(_11510_),
    .Y(_11903_));
 OAI21x1_ASAP7_75t_R _20249_ (.A1(_11902_),
    .A2(_11903_),
    .B(_11564_),
    .Y(_11904_));
 OAI21x1_ASAP7_75t_R _20250_ (.A1(net897),
    .A2(_11664_),
    .B(_11654_),
    .Y(_11905_));
 NOR2x1_ASAP7_75t_R _20251_ (.A(_11905_),
    .B(_11530_),
    .Y(_11906_));
 NOR2x1_ASAP7_75t_R _20252_ (.A(_11904_),
    .B(_11906_),
    .Y(_11907_));
 NAND2x1_ASAP7_75t_R _20253_ (.A(_11507_),
    .B(_11719_),
    .Y(_11908_));
 AOI211x1_ASAP7_75t_R _20254_ (.A1(_11481_),
    .A2(_11523_),
    .B(_11908_),
    .C(_11578_),
    .Y(_11909_));
 AO21x1_ASAP7_75t_R _20255_ (.A1(_11645_),
    .A2(_11763_),
    .B(_11573_),
    .Y(_11910_));
 NOR2x1_ASAP7_75t_R _20256_ (.A(_11507_),
    .B(_11670_),
    .Y(_11911_));
 AO21x1_ASAP7_75t_R _20257_ (.A1(_11910_),
    .A2(_11911_),
    .B(_11564_),
    .Y(_11912_));
 NOR2x1_ASAP7_75t_R _20258_ (.A(_11909_),
    .B(_11912_),
    .Y(_11913_));
 OAI21x1_ASAP7_75t_R _20259_ (.A1(_11907_),
    .A2(_11913_),
    .B(_11504_),
    .Y(_11914_));
 AOI22x1_ASAP7_75t_R _20260_ (.A1(_11869_),
    .A2(_11883_),
    .B1(_11899_),
    .B2(_11914_),
    .Y(_00044_));
 AO21x1_ASAP7_75t_R _20261_ (.A1(_15823_),
    .A2(_11549_),
    .B(_11722_),
    .Y(_11915_));
 NOR2x1_ASAP7_75t_R _20262_ (.A(_11547_),
    .B(_11548_),
    .Y(_11916_));
 OAI21x1_ASAP7_75t_R _20263_ (.A1(_11915_),
    .A2(_11916_),
    .B(_11494_),
    .Y(_11917_));
 AO21x2_ASAP7_75t_R _20264_ (.A1(_11456_),
    .A2(_01161_),
    .B(_11445_),
    .Y(_11918_));
 OAI21x1_ASAP7_75t_R _20265_ (.A1(_11513_),
    .A2(_11918_),
    .B(_11598_),
    .Y(_11919_));
 INVx2_ASAP7_75t_R _20266_ (.A(_11632_),
    .Y(_11920_));
 NOR2x1_ASAP7_75t_R _20267_ (.A(_11920_),
    .B(_11454_),
    .Y(_11921_));
 NOR2x1_ASAP7_75t_R _20268_ (.A(_11919_),
    .B(_11921_),
    .Y(_11922_));
 OAI21x1_ASAP7_75t_R _20269_ (.A1(_11917_),
    .A2(_11922_),
    .B(_11504_),
    .Y(_11923_));
 NOR2x1_ASAP7_75t_R _20270_ (.A(_11577_),
    .B(_11592_),
    .Y(_11924_));
 AOI211x1_ASAP7_75t_R _20271_ (.A1(_11529_),
    .A2(_11515_),
    .B(_11924_),
    .C(_11629_),
    .Y(_11925_));
 INVx1_ASAP7_75t_R _20272_ (.A(_11570_),
    .Y(_11926_));
 AO21x1_ASAP7_75t_R _20273_ (.A1(_11926_),
    .A2(_11549_),
    .B(_11472_),
    .Y(_11927_));
 AOI21x1_ASAP7_75t_R _20274_ (.A1(_11763_),
    .A2(_11826_),
    .B(_11520_),
    .Y(_11928_));
 OAI21x1_ASAP7_75t_R _20275_ (.A1(_11927_),
    .A2(_11928_),
    .B(_11532_),
    .Y(_11929_));
 NOR2x1_ASAP7_75t_R _20276_ (.A(_11925_),
    .B(_11929_),
    .Y(_11930_));
 OAI21x1_ASAP7_75t_R _20277_ (.A1(_11923_),
    .A2(_11930_),
    .B(_11545_),
    .Y(_11931_));
 INVx1_ASAP7_75t_R _20278_ (.A(_11459_),
    .Y(_11932_));
 AO21x1_ASAP7_75t_R _20279_ (.A1(_11631_),
    .A2(_11932_),
    .B(_11531_),
    .Y(_11933_));
 INVx1_ASAP7_75t_R _20280_ (.A(_11724_),
    .Y(_11934_));
 AO21x1_ASAP7_75t_R _20281_ (.A1(_11730_),
    .A2(_11510_),
    .B(_11507_),
    .Y(_11935_));
 AOI21x1_ASAP7_75t_R _20282_ (.A1(_11529_),
    .A2(_11934_),
    .B(_11935_),
    .Y(_11936_));
 OAI21x1_ASAP7_75t_R _20283_ (.A1(_11933_),
    .A2(_11936_),
    .B(_11586_),
    .Y(_11937_));
 AO21x1_ASAP7_75t_R _20284_ (.A1(_11528_),
    .A2(net41),
    .B(_11573_),
    .Y(_11938_));
 OA21x2_ASAP7_75t_R _20285_ (.A1(_11556_),
    .A2(_11524_),
    .B(_11605_),
    .Y(_11939_));
 AO21x1_ASAP7_75t_R _20286_ (.A1(_11938_),
    .A2(_11939_),
    .B(_11493_),
    .Y(_11940_));
 AND2x2_ASAP7_75t_R _20287_ (.A(_11809_),
    .B(_11506_),
    .Y(_11941_));
 AO21x1_ASAP7_75t_R _20288_ (.A1(_11568_),
    .A2(_11570_),
    .B(_11524_),
    .Y(_11942_));
 AND3x1_ASAP7_75t_R _20289_ (.A(_11941_),
    .B(_11942_),
    .C(_11771_),
    .Y(_11943_));
 NOR2x1_ASAP7_75t_R _20290_ (.A(_11940_),
    .B(_11943_),
    .Y(_11944_));
 NOR2x1_ASAP7_75t_R _20291_ (.A(_11937_),
    .B(_11944_),
    .Y(_11945_));
 AO21x1_ASAP7_75t_R _20292_ (.A1(_11552_),
    .A2(_15828_),
    .B(_11926_),
    .Y(_11946_));
 NOR2x1_ASAP7_75t_R _20293_ (.A(_11834_),
    .B(_11946_),
    .Y(_11947_));
 AO21x1_ASAP7_75t_R _20294_ (.A1(_11705_),
    .A2(_11552_),
    .B(_11804_),
    .Y(_11948_));
 OA21x2_ASAP7_75t_R _20295_ (.A1(net41),
    .A2(_11640_),
    .B(_11654_),
    .Y(_11949_));
 AO21x1_ASAP7_75t_R _20296_ (.A1(_11614_),
    .A2(_11552_),
    .B(_11549_),
    .Y(_11950_));
 AOI21x1_ASAP7_75t_R _20297_ (.A1(_11949_),
    .A2(_11950_),
    .B(_11532_),
    .Y(_11951_));
 OAI21x1_ASAP7_75t_R _20298_ (.A1(_11947_),
    .A2(_11948_),
    .B(_11951_),
    .Y(_11952_));
 AND2x2_ASAP7_75t_R _20299_ (.A(_11901_),
    .B(_11524_),
    .Y(_11953_));
 AO21x1_ASAP7_75t_R _20300_ (.A1(_11953_),
    .A2(_11817_),
    .B(_11885_),
    .Y(_11954_));
 AO21x1_ASAP7_75t_R _20301_ (.A1(_11763_),
    .A2(_11589_),
    .B(_11507_),
    .Y(_11955_));
 NOR2x1_ASAP7_75t_R _20302_ (.A(_11559_),
    .B(_11920_),
    .Y(_11956_));
 OAI21x1_ASAP7_75t_R _20303_ (.A1(_11955_),
    .A2(_11956_),
    .B(_11576_),
    .Y(_11957_));
 AO21x1_ASAP7_75t_R _20304_ (.A1(_11954_),
    .A2(_11508_),
    .B(_11957_),
    .Y(_11958_));
 AOI21x1_ASAP7_75t_R _20305_ (.A1(_11952_),
    .A2(_11958_),
    .B(_11504_),
    .Y(_11959_));
 AO21x1_ASAP7_75t_R _20306_ (.A1(_11456_),
    .A2(net507),
    .B(_11624_),
    .Y(_11960_));
 OAI21x1_ASAP7_75t_R _20307_ (.A1(_11729_),
    .A2(_11960_),
    .B(_11598_),
    .Y(_11961_));
 NOR2x1_ASAP7_75t_R _20308_ (.A(_11918_),
    .B(_11603_),
    .Y(_11962_));
 NOR2x1_ASAP7_75t_R _20309_ (.A(_11961_),
    .B(_11962_),
    .Y(_11963_));
 OA21x2_ASAP7_75t_R _20310_ (.A1(_11479_),
    .A2(_15831_),
    .B(_11459_),
    .Y(_11964_));
 OAI21x1_ASAP7_75t_R _20311_ (.A1(_11964_),
    .A2(_11527_),
    .B(_11564_),
    .Y(_11965_));
 NOR2x1_ASAP7_75t_R _20312_ (.A(_11963_),
    .B(_11965_),
    .Y(_11966_));
 AO21x1_ASAP7_75t_R _20313_ (.A1(_11462_),
    .A2(_11640_),
    .B(_11722_),
    .Y(_11967_));
 NOR2x1_ASAP7_75t_R _20314_ (.A(_11967_),
    .B(_11803_),
    .Y(_11968_));
 AO21x1_ASAP7_75t_R _20315_ (.A1(_11688_),
    .A2(_11664_),
    .B(_11564_),
    .Y(_11969_));
 OAI21x1_ASAP7_75t_R _20316_ (.A1(_11968_),
    .A2(_11969_),
    .B(_11504_),
    .Y(_11970_));
 OAI21x1_ASAP7_75t_R _20317_ (.A1(_11966_),
    .A2(_11970_),
    .B(_11853_),
    .Y(_11971_));
 OAI22x1_ASAP7_75t_R _20318_ (.A1(_11931_),
    .A2(_11945_),
    .B1(_11959_),
    .B2(_11971_),
    .Y(_00045_));
 AOI21x1_ASAP7_75t_R _20319_ (.A1(_11618_),
    .A2(_11633_),
    .B(_11834_),
    .Y(_11972_));
 OAI21x1_ASAP7_75t_R _20320_ (.A1(_11972_),
    .A2(_11908_),
    .B(_11494_),
    .Y(_11973_));
 AOI21x1_ASAP7_75t_R _20321_ (.A1(_01165_),
    .A2(_01163_),
    .B(_11520_),
    .Y(_11974_));
 AOI211x1_ASAP7_75t_R _20322_ (.A1(_11741_),
    .A2(_11607_),
    .B(_11974_),
    .C(_11508_),
    .Y(_11975_));
 OAI21x1_ASAP7_75t_R _20323_ (.A1(_11973_),
    .A2(_11975_),
    .B(_11504_),
    .Y(_11976_));
 AOI21x1_ASAP7_75t_R _20324_ (.A1(_11709_),
    .A2(_11839_),
    .B(_11549_),
    .Y(_11977_));
 INVx1_ASAP7_75t_R _20325_ (.A(_11552_),
    .Y(_11978_));
 NAND2x1_ASAP7_75t_R _20326_ (.A(_11510_),
    .B(_11525_),
    .Y(_11979_));
 OAI21x1_ASAP7_75t_R _20327_ (.A1(_11818_),
    .A2(_11978_),
    .B(_11979_),
    .Y(_11980_));
 OAI21x1_ASAP7_75t_R _20328_ (.A1(_11977_),
    .A2(_11980_),
    .B(_11804_),
    .Y(_11981_));
 NOR2x2_ASAP7_75t_R _20329_ (.A(_11561_),
    .B(_11761_),
    .Y(_11982_));
 OAI21x1_ASAP7_75t_R _20330_ (.A1(_15828_),
    .A2(_11729_),
    .B(_11982_),
    .Y(_11983_));
 NOR2x1_ASAP7_75t_R _20331_ (.A(_11924_),
    .B(_11625_),
    .Y(_11984_));
 NAND2x1_ASAP7_75t_R _20332_ (.A(_11983_),
    .B(_11984_),
    .Y(_11985_));
 AOI21x1_ASAP7_75t_R _20333_ (.A1(_11981_),
    .A2(_11985_),
    .B(_11494_),
    .Y(_11986_));
 OAI21x1_ASAP7_75t_R _20334_ (.A1(_11976_),
    .A2(_11986_),
    .B(_11853_),
    .Y(_11987_));
 AO21x1_ASAP7_75t_R _20335_ (.A1(_11926_),
    .A2(_11640_),
    .B(_11472_),
    .Y(_11988_));
 OA21x2_ASAP7_75t_R _20336_ (.A1(_11528_),
    .A2(net4),
    .B(_11549_),
    .Y(_11989_));
 OAI21x1_ASAP7_75t_R _20337_ (.A1(_11988_),
    .A2(_11989_),
    .B(_11576_),
    .Y(_11990_));
 OAI21x1_ASAP7_75t_R _20338_ (.A1(_11663_),
    .A2(_11895_),
    .B(_11654_),
    .Y(_11991_));
 NAND2x1_ASAP7_75t_R _20339_ (.A(_11730_),
    .B(_11656_),
    .Y(_11992_));
 OAI21x1_ASAP7_75t_R _20340_ (.A1(_11640_),
    .A2(_11665_),
    .B(_11992_),
    .Y(_11993_));
 NOR2x1_ASAP7_75t_R _20341_ (.A(_11991_),
    .B(_11993_),
    .Y(_11994_));
 OAI21x1_ASAP7_75t_R _20342_ (.A1(_11990_),
    .A2(_11994_),
    .B(_11586_),
    .Y(_11995_));
 INVx1_ASAP7_75t_R _20343_ (.A(_11725_),
    .Y(_11996_));
 OAI21x1_ASAP7_75t_R _20344_ (.A1(_11996_),
    .A2(_11934_),
    .B(_11941_),
    .Y(_11997_));
 AND3x1_ASAP7_75t_R _20345_ (.A(_11568_),
    .B(_11901_),
    .C(_11589_),
    .Y(_11998_));
 OAI21x1_ASAP7_75t_R _20346_ (.A1(_15831_),
    .A2(net41),
    .B(_11573_),
    .Y(_11999_));
 NOR2x1_ASAP7_75t_R _20347_ (.A(_11999_),
    .B(_11454_),
    .Y(_12000_));
 OAI21x1_ASAP7_75t_R _20348_ (.A1(_11998_),
    .A2(_12000_),
    .B(_11804_),
    .Y(_12001_));
 AOI21x1_ASAP7_75t_R _20349_ (.A1(_11997_),
    .A2(_12001_),
    .B(_11532_),
    .Y(_12002_));
 NOR2x1_ASAP7_75t_R _20350_ (.A(_12002_),
    .B(_11995_),
    .Y(_12003_));
 OAI21x1_ASAP7_75t_R _20351_ (.A1(_11609_),
    .A2(_11887_),
    .B(_11508_),
    .Y(_12004_));
 AO21x1_ASAP7_75t_R _20352_ (.A1(_11673_),
    .A2(_11520_),
    .B(_11582_),
    .Y(_12005_));
 AOI21x1_ASAP7_75t_R _20353_ (.A1(_12004_),
    .A2(_12005_),
    .B(_11504_),
    .Y(_12006_));
 AO21x1_ASAP7_75t_R _20354_ (.A1(_11676_),
    .A2(_11549_),
    .B(_11472_),
    .Y(_12007_));
 NOR2x1_ASAP7_75t_R _20355_ (.A(_12007_),
    .B(_11455_),
    .Y(_12008_));
 AO21x1_ASAP7_75t_R _20356_ (.A1(_11704_),
    .A2(_11549_),
    .B(_11722_),
    .Y(_12009_));
 OA21x2_ASAP7_75t_R _20357_ (.A1(_11456_),
    .A2(net462),
    .B(_11524_),
    .Y(_12010_));
 NOR2x1_ASAP7_75t_R _20358_ (.A(_12010_),
    .B(_11982_),
    .Y(_12011_));
 OAI21x1_ASAP7_75t_R _20359_ (.A1(_12009_),
    .A2(_12011_),
    .B(_11503_),
    .Y(_12012_));
 OAI21x1_ASAP7_75t_R _20360_ (.A1(_12008_),
    .A2(_12012_),
    .B(_11532_),
    .Y(_12013_));
 OAI21x1_ASAP7_75t_R _20361_ (.A1(_12006_),
    .A2(_12013_),
    .B(_11545_),
    .Y(_12014_));
 AOI22x1_ASAP7_75t_R _20362_ (.A1(_11459_),
    .A2(_11568_),
    .B1(_11834_),
    .B2(_11663_),
    .Y(_12015_));
 AO21x1_ASAP7_75t_R _20363_ (.A1(_00508_),
    .A2(_11510_),
    .B(_11507_),
    .Y(_12016_));
 NOR2x1_ASAP7_75t_R _20364_ (.A(_11513_),
    .B(_11918_),
    .Y(_12017_));
 OAI21x1_ASAP7_75t_R _20365_ (.A1(_12016_),
    .A2(_12017_),
    .B(_11585_),
    .Y(_12018_));
 AOI21x1_ASAP7_75t_R _20366_ (.A1(_11508_),
    .A2(_12015_),
    .B(_12018_),
    .Y(_12019_));
 NOR2x1_ASAP7_75t_R _20367_ (.A(_11520_),
    .B(net41),
    .Y(_12020_));
 AO21x1_ASAP7_75t_R _20368_ (.A1(_11607_),
    .A2(_11592_),
    .B(_11722_),
    .Y(_12021_));
 OAI21x1_ASAP7_75t_R _20369_ (.A1(_12020_),
    .A2(_12021_),
    .B(_11503_),
    .Y(_12022_));
 NAND2x1_ASAP7_75t_R _20370_ (.A(_11589_),
    .B(_11517_),
    .Y(_12023_));
 OAI21x1_ASAP7_75t_R _20371_ (.A1(_11834_),
    .A2(_11547_),
    .B(_12023_),
    .Y(_12024_));
 AOI21x1_ASAP7_75t_R _20372_ (.A1(_11621_),
    .A2(_12024_),
    .B(_11804_),
    .Y(_12025_));
 OAI21x1_ASAP7_75t_R _20373_ (.A1(_12022_),
    .A2(_12025_),
    .B(_11494_),
    .Y(_12026_));
 NOR2x1_ASAP7_75t_R _20374_ (.A(_12019_),
    .B(_12026_),
    .Y(_12027_));
 OAI22x1_ASAP7_75t_R _20375_ (.A1(_12003_),
    .A2(_11987_),
    .B1(_12014_),
    .B2(_12027_),
    .Y(_00046_));
 AO21x1_ASAP7_75t_R _20376_ (.A1(_11552_),
    .A2(_15831_),
    .B(_11571_),
    .Y(_12028_));
 OAI21x1_ASAP7_75t_R _20377_ (.A1(_11477_),
    .A2(_11603_),
    .B(_11582_),
    .Y(_12029_));
 AO21x1_ASAP7_75t_R _20378_ (.A1(_11520_),
    .A2(_12028_),
    .B(_12029_),
    .Y(_12030_));
 AO21x1_ASAP7_75t_R _20379_ (.A1(_11517_),
    .A2(_11640_),
    .B(_11722_),
    .Y(_12031_));
 OA21x2_ASAP7_75t_R _20380_ (.A1(_12031_),
    .A2(_11887_),
    .B(_11494_),
    .Y(_12032_));
 AOI211x1_ASAP7_75t_R _20381_ (.A1(_11741_),
    .A2(_11645_),
    .B(_11977_),
    .C(_11582_),
    .Y(_12033_));
 AO21x1_ASAP7_75t_R _20382_ (.A1(_11580_),
    .A2(_11517_),
    .B(_11472_),
    .Y(_12034_));
 OAI21x1_ASAP7_75t_R _20383_ (.A1(_11814_),
    .A2(_12034_),
    .B(_11576_),
    .Y(_12035_));
 NOR2x1_ASAP7_75t_R _20384_ (.A(_12033_),
    .B(_12035_),
    .Y(_12036_));
 AOI211x1_ASAP7_75t_R _20385_ (.A1(_12030_),
    .A2(_12032_),
    .B(_12036_),
    .C(_11586_),
    .Y(_12037_));
 AND2x2_ASAP7_75t_R _20386_ (.A(_11809_),
    .B(_11605_),
    .Y(_12038_));
 AO21x1_ASAP7_75t_R _20387_ (.A1(_12038_),
    .A2(_11691_),
    .B(_11564_),
    .Y(_12039_));
 INVx1_ASAP7_75t_R _20388_ (.A(_11553_),
    .Y(_12040_));
 OAI21x1_ASAP7_75t_R _20389_ (.A1(_11834_),
    .A2(_11603_),
    .B(_11582_),
    .Y(_12041_));
 AOI21x1_ASAP7_75t_R _20390_ (.A1(_12040_),
    .A2(_12010_),
    .B(_12041_),
    .Y(_12042_));
 OAI21x1_ASAP7_75t_R _20391_ (.A1(_12039_),
    .A2(_12042_),
    .B(_11586_),
    .Y(_12043_));
 AOI211x1_ASAP7_75t_R _20392_ (.A1(_12040_),
    .A2(_11514_),
    .B(_11880_),
    .C(_11582_),
    .Y(_12044_));
 NAND2x1_ASAP7_75t_R _20393_ (.A(_15823_),
    .B(_11589_),
    .Y(_12045_));
 AO21x1_ASAP7_75t_R _20394_ (.A1(_11676_),
    .A2(_11645_),
    .B(_11561_),
    .Y(_12046_));
 NAND2x1_ASAP7_75t_R _20395_ (.A(_12045_),
    .B(_12046_),
    .Y(_12047_));
 OAI21x1_ASAP7_75t_R _20396_ (.A1(_11804_),
    .A2(_12047_),
    .B(_11494_),
    .Y(_12048_));
 NOR2x1_ASAP7_75t_R _20397_ (.A(_12044_),
    .B(_12048_),
    .Y(_12049_));
 OAI21x1_ASAP7_75t_R _20398_ (.A1(_12043_),
    .A2(_12049_),
    .B(_11545_),
    .Y(_12050_));
 AOI21x1_ASAP7_75t_R _20399_ (.A1(_11568_),
    .A2(_11580_),
    .B(_11472_),
    .Y(_12051_));
 OAI21x1_ASAP7_75t_R _20400_ (.A1(_11513_),
    .A2(_11477_),
    .B(_12051_),
    .Y(_12052_));
 NAND2x1_ASAP7_75t_R _20401_ (.A(_11589_),
    .B(_11579_),
    .Y(_12053_));
 OAI21x1_ASAP7_75t_R _20402_ (.A1(_01165_),
    .A2(_11624_),
    .B(_11471_),
    .Y(_12054_));
 NOR2x1_ASAP7_75t_R _20403_ (.A(_11634_),
    .B(_12054_),
    .Y(_12055_));
 AOI21x1_ASAP7_75t_R _20404_ (.A1(_12053_),
    .A2(_12055_),
    .B(_11493_),
    .Y(_12056_));
 NAND2x1_ASAP7_75t_R _20405_ (.A(_12052_),
    .B(_12056_),
    .Y(_12057_));
 AND2x2_ASAP7_75t_R _20406_ (.A(_11445_),
    .B(_00507_),
    .Y(_12058_));
 OA21x2_ASAP7_75t_R _20407_ (.A1(_11619_),
    .A2(_12058_),
    .B(_11493_),
    .Y(_12059_));
 AO21x1_ASAP7_75t_R _20408_ (.A1(_11592_),
    .A2(_15821_),
    .B(_11577_),
    .Y(_12060_));
 NAND2x1_ASAP7_75t_R _20409_ (.A(_12060_),
    .B(_11684_),
    .Y(_12061_));
 AOI21x1_ASAP7_75t_R _20410_ (.A1(_12059_),
    .A2(_12061_),
    .B(_11503_),
    .Y(_12062_));
 AOI21x1_ASAP7_75t_R _20411_ (.A1(_12057_),
    .A2(_12062_),
    .B(_11545_),
    .Y(_12063_));
 NAND2x1_ASAP7_75t_R _20412_ (.A(net41),
    .B(_11665_),
    .Y(_12064_));
 AOI211x1_ASAP7_75t_R _20413_ (.A1(_11834_),
    .A2(_12064_),
    .B(_11798_),
    .C(_11804_),
    .Y(_12065_));
 OAI21x1_ASAP7_75t_R _20414_ (.A1(_11432_),
    .A2(_11380_),
    .B(_11572_),
    .Y(_12066_));
 NAND2x1_ASAP7_75t_R _20415_ (.A(_11632_),
    .B(_11570_),
    .Y(_12067_));
 OAI21x1_ASAP7_75t_R _20416_ (.A1(_11477_),
    .A2(_12066_),
    .B(_12067_),
    .Y(_12068_));
 AO21x1_ASAP7_75t_R _20417_ (.A1(_12068_),
    .A2(_11804_),
    .B(_11576_),
    .Y(_12069_));
 NAND2x1_ASAP7_75t_R _20418_ (.A(_11510_),
    .B(_12066_),
    .Y(_12070_));
 NOR2x1_ASAP7_75t_R _20419_ (.A(_11720_),
    .B(_11619_),
    .Y(_12071_));
 NAND2x1_ASAP7_75t_R _20420_ (.A(_12070_),
    .B(_12071_),
    .Y(_12072_));
 OA21x2_ASAP7_75t_R _20421_ (.A1(net506),
    .A2(_11577_),
    .B(_11506_),
    .Y(_12073_));
 NAND2x1_ASAP7_75t_R _20422_ (.A(_11607_),
    .B(_11741_),
    .Y(_12074_));
 AOI21x1_ASAP7_75t_R _20423_ (.A1(_12073_),
    .A2(_12074_),
    .B(_11564_),
    .Y(_12075_));
 AOI21x1_ASAP7_75t_R _20424_ (.A1(_12072_),
    .A2(_12075_),
    .B(_11586_),
    .Y(_12076_));
 OAI21x1_ASAP7_75t_R _20425_ (.A1(_12065_),
    .A2(_12069_),
    .B(_12076_),
    .Y(_12077_));
 NAND2x1_ASAP7_75t_R _20426_ (.A(_12063_),
    .B(_12077_),
    .Y(_12078_));
 OAI21x1_ASAP7_75t_R _20427_ (.A1(_12037_),
    .A2(_12050_),
    .B(_12078_),
    .Y(_00047_));
 NOR2x2_ASAP7_75t_R _20428_ (.A(_10743_),
    .B(_00509_),
    .Y(_12079_));
 BUFx6f_ASAP7_75t_R _20429_ (.A(_00787_),
    .Y(_12080_));
 XOR2x2_ASAP7_75t_R _20430_ (.A(_12080_),
    .B(_00780_),
    .Y(_12081_));
 BUFx12f_ASAP7_75t_R _20431_ (.A(_00845_),
    .Y(_12082_));
 XOR2x1_ASAP7_75t_R _20432_ (.A(_12081_),
    .Y(_12083_),
    .B(net905));
 BUFx6f_ASAP7_75t_R _20433_ (.A(_00748_),
    .Y(_12084_));
 BUFx6f_ASAP7_75t_R _20434_ (.A(_00755_),
    .Y(_12085_));
 XOR2x2_ASAP7_75t_R _20435_ (.A(_12084_),
    .B(_12085_),
    .Y(_12086_));
 BUFx6f_ASAP7_75t_R _20436_ (.A(_00813_),
    .Y(_12087_));
 XOR2x2_ASAP7_75t_R _20437_ (.A(_12087_),
    .B(_00781_),
    .Y(_12088_));
 XOR2x2_ASAP7_75t_R _20438_ (.A(_12086_),
    .B(_12088_),
    .Y(_12089_));
 NAND2x1_ASAP7_75t_R _20439_ (.A(_12083_),
    .B(_12089_),
    .Y(_12090_));
 OR2x2_ASAP7_75t_R _20440_ (.A(_12083_),
    .B(_12089_),
    .Y(_12091_));
 BUFx12f_ASAP7_75t_R _20441_ (.A(_10689_),
    .Y(_12092_));
 AOI21x1_ASAP7_75t_R _20442_ (.A1(_12090_),
    .A2(_12091_),
    .B(_12092_),
    .Y(_12093_));
 OAI21x1_ASAP7_75t_R _20443_ (.A1(_12079_),
    .A2(_12093_),
    .B(_08190_),
    .Y(_12094_));
 BUFx12_ASAP7_75t_R _20444_ (.A(_11373_),
    .Y(_12095_));
 AND2x2_ASAP7_75t_R _20445_ (.A(_12095_),
    .B(_00509_),
    .Y(_12096_));
 INVx3_ASAP7_75t_R _20446_ (.A(net905),
    .Y(_12097_));
 XOR2x1_ASAP7_75t_R _20447_ (.A(_12081_),
    .Y(_12098_),
    .B(_12097_));
 XOR2x2_ASAP7_75t_R _20448_ (.A(_12089_),
    .B(_12098_),
    .Y(_12099_));
 NOR2x2_ASAP7_75t_R _20449_ (.A(_12092_),
    .B(_12099_),
    .Y(_12100_));
 INVx2_ASAP7_75t_R _20450_ (.A(_08190_),
    .Y(_12101_));
 OAI21x1_ASAP7_75t_R _20451_ (.A1(_12096_),
    .A2(_12100_),
    .B(_12101_),
    .Y(_12102_));
 NAND2x2_ASAP7_75t_R _20452_ (.A(_12102_),
    .B(_12094_),
    .Y(_12103_));
 BUFx10_ASAP7_75t_R _20453_ (.A(_12103_),
    .Y(_15838_));
 BUFx6f_ASAP7_75t_R _20454_ (.A(_00844_),
    .Y(_12104_));
 INVx2_ASAP7_75t_R _20455_ (.A(_12104_),
    .Y(_12105_));
 XOR2x2_ASAP7_75t_R _20456_ (.A(_12085_),
    .B(_12080_),
    .Y(_12106_));
 NAND2x1_ASAP7_75t_R _20457_ (.A(_12105_),
    .B(_12106_),
    .Y(_12107_));
 BUFx10_ASAP7_75t_R _20458_ (.A(_12080_),
    .Y(_12108_));
 XNOR2x1_ASAP7_75t_R _20459_ (.B(_12108_),
    .Y(_12109_),
    .A(_12085_));
 NAND2x1_ASAP7_75t_R _20460_ (.A(_12104_),
    .B(_12109_),
    .Y(_12110_));
 XNOR2x2_ASAP7_75t_R _20461_ (.A(net618),
    .B(_00812_),
    .Y(_12111_));
 AOI21x1_ASAP7_75t_R _20462_ (.A1(_12107_),
    .A2(_12110_),
    .B(_12111_),
    .Y(_12112_));
 NAND2x1_ASAP7_75t_R _20463_ (.A(_12104_),
    .B(_12106_),
    .Y(_12113_));
 NAND2x1_ASAP7_75t_R _20464_ (.A(_12105_),
    .B(_12109_),
    .Y(_12114_));
 BUFx6f_ASAP7_75t_R _20465_ (.A(_00780_),
    .Y(_12115_));
 XOR2x2_ASAP7_75t_R _20466_ (.A(_12115_),
    .B(_00812_),
    .Y(_12116_));
 AOI21x1_ASAP7_75t_R _20467_ (.A1(_12113_),
    .A2(_12114_),
    .B(net635),
    .Y(_12117_));
 OAI21x1_ASAP7_75t_R _20468_ (.A1(_12112_),
    .A2(_12117_),
    .B(_10621_),
    .Y(_12118_));
 INVx2_ASAP7_75t_R _20469_ (.A(_08177_),
    .Y(_12119_));
 NOR2x1_ASAP7_75t_R _20470_ (.A(_10762_),
    .B(_00510_),
    .Y(_12120_));
 INVx3_ASAP7_75t_R _20471_ (.A(_12120_),
    .Y(_12121_));
 NAND3x2_ASAP7_75t_R _20472_ (.B(_12119_),
    .C(_12121_),
    .Y(_12122_),
    .A(net611));
 AO21x1_ASAP7_75t_R _20473_ (.A1(net611),
    .A2(_12121_),
    .B(_12119_),
    .Y(_12123_));
 NAND2x2_ASAP7_75t_R _20474_ (.A(_12122_),
    .B(_12123_),
    .Y(_12124_));
 BUFx12_ASAP7_75t_R _20475_ (.A(_12124_),
    .Y(_15840_));
 BUFx6f_ASAP7_75t_R _20476_ (.A(_00782_),
    .Y(_12125_));
 INVx2_ASAP7_75t_R _20477_ (.A(_12125_),
    .Y(_12126_));
 BUFx6f_ASAP7_75t_R _20478_ (.A(_00749_),
    .Y(_12127_));
 XOR2x2_ASAP7_75t_R _20479_ (.A(_12127_),
    .B(_00781_),
    .Y(_12128_));
 NAND2x1_ASAP7_75t_R _20480_ (.A(_12126_),
    .B(_12128_),
    .Y(_12129_));
 XNOR2x2_ASAP7_75t_R _20481_ (.A(_12127_),
    .B(_00781_),
    .Y(_12130_));
 NAND2x1_ASAP7_75t_R _20482_ (.A(_12125_),
    .B(net834),
    .Y(_12131_));
 BUFx10_ASAP7_75t_R _20483_ (.A(_00814_),
    .Y(_12132_));
 BUFx10_ASAP7_75t_R _20484_ (.A(_00846_),
    .Y(_12133_));
 XNOR2x2_ASAP7_75t_R _20485_ (.A(_12132_),
    .B(_12133_),
    .Y(_12134_));
 AOI21x1_ASAP7_75t_R _20486_ (.A1(_12129_),
    .A2(_12131_),
    .B(_12134_),
    .Y(_12135_));
 NAND2x1_ASAP7_75t_R _20487_ (.A(_12125_),
    .B(_12128_),
    .Y(_12136_));
 NAND2x1_ASAP7_75t_R _20488_ (.A(_12126_),
    .B(net834),
    .Y(_12137_));
 XOR2x2_ASAP7_75t_R _20489_ (.A(_12132_),
    .B(_12133_),
    .Y(_12138_));
 AOI21x1_ASAP7_75t_R _20490_ (.A1(_12136_),
    .A2(_12137_),
    .B(_12138_),
    .Y(_12139_));
 OAI21x1_ASAP7_75t_R _20491_ (.A1(_12135_),
    .A2(_12139_),
    .B(_10665_),
    .Y(_12140_));
 NOR2x2_ASAP7_75t_R _20492_ (.A(net786),
    .B(_00512_),
    .Y(_12141_));
 INVx3_ASAP7_75t_R _20493_ (.A(_12141_),
    .Y(_12142_));
 NAND3x2_ASAP7_75t_R _20494_ (.B(_08197_),
    .C(_12142_),
    .Y(_12143_),
    .A(_12140_));
 AO21x2_ASAP7_75t_R _20495_ (.A1(_12140_),
    .A2(_12142_),
    .B(_08197_),
    .Y(_12144_));
 NAND2x2_ASAP7_75t_R _20496_ (.A(_12143_),
    .B(_12144_),
    .Y(_12145_));
 BUFx10_ASAP7_75t_R _20497_ (.A(_12145_),
    .Y(_15848_));
 NAND3x2_ASAP7_75t_R _20498_ (.B(_08177_),
    .C(_12121_),
    .Y(_12146_),
    .A(_12118_));
 AO21x1_ASAP7_75t_R _20499_ (.A1(_12121_),
    .A2(_12118_),
    .B(_08177_),
    .Y(_12147_));
 NAND2x2_ASAP7_75t_R _20500_ (.A(_12146_),
    .B(_12147_),
    .Y(_12148_));
 BUFx6f_ASAP7_75t_R _20501_ (.A(_12148_),
    .Y(_15835_));
 NAND3x2_ASAP7_75t_R _20502_ (.B(_08314_),
    .C(_12142_),
    .Y(_12149_),
    .A(_12140_));
 AO21x1_ASAP7_75t_R _20503_ (.A1(_12140_),
    .A2(_12142_),
    .B(_08314_),
    .Y(_12150_));
 BUFx4f_ASAP7_75t_R _20504_ (.A(_12150_),
    .Y(_12151_));
 NAND2x2_ASAP7_75t_R _20505_ (.A(_12149_),
    .B(_12151_),
    .Y(_12152_));
 BUFx12_ASAP7_75t_R _20506_ (.A(_12152_),
    .Y(_12153_));
 BUFx10_ASAP7_75t_R _20507_ (.A(_12153_),
    .Y(_15845_));
 NOR2x1_ASAP7_75t_R _20508_ (.A(_12126_),
    .B(_12128_),
    .Y(_12154_));
 NOR2x1_ASAP7_75t_R _20509_ (.A(_12125_),
    .B(_12130_),
    .Y(_12155_));
 OAI21x1_ASAP7_75t_R _20510_ (.A1(_12154_),
    .A2(_12155_),
    .B(_12138_),
    .Y(_12156_));
 NOR2x1_ASAP7_75t_R _20511_ (.A(_12125_),
    .B(_12128_),
    .Y(_12157_));
 NOR2x1_ASAP7_75t_R _20512_ (.A(_12126_),
    .B(_12130_),
    .Y(_12158_));
 OAI21x1_ASAP7_75t_R _20513_ (.A1(_12157_),
    .A2(_12158_),
    .B(_12134_),
    .Y(_12159_));
 BUFx12f_ASAP7_75t_R _20514_ (.A(_10639_),
    .Y(_12160_));
 BUFx16f_ASAP7_75t_R _20515_ (.A(_12160_),
    .Y(_12161_));
 AOI21x1_ASAP7_75t_R _20516_ (.A1(_12156_),
    .A2(_12159_),
    .B(_12161_),
    .Y(_12162_));
 NOR3x2_ASAP7_75t_R _20517_ (.B(_08314_),
    .C(_12141_),
    .Y(_12163_),
    .A(_12162_));
 OA21x2_ASAP7_75t_R _20518_ (.A1(_12162_),
    .A2(_12141_),
    .B(_08314_),
    .Y(_12164_));
 BUFx4f_ASAP7_75t_R _20519_ (.A(_01168_),
    .Y(_12165_));
 INVx2_ASAP7_75t_R _20520_ (.A(_12165_),
    .Y(_12166_));
 OAI21x1_ASAP7_75t_R _20521_ (.A1(_12163_),
    .A2(_12164_),
    .B(_12166_),
    .Y(_12167_));
 INVx2_ASAP7_75t_R _20522_ (.A(_12167_),
    .Y(_12168_));
 BUFx4f_ASAP7_75t_R _20523_ (.A(_00750_),
    .Y(_12169_));
 XOR2x2_ASAP7_75t_R _20524_ (.A(_12169_),
    .B(_12085_),
    .Y(_12170_));
 XNOR2x1_ASAP7_75t_R _20525_ (.B(_12170_),
    .Y(_12171_),
    .A(_00783_));
 XNOR2x2_ASAP7_75t_R _20526_ (.A(_00815_),
    .B(_00847_),
    .Y(_12172_));
 XOR2x2_ASAP7_75t_R _20527_ (.A(_12125_),
    .B(_12080_),
    .Y(_12173_));
 XOR2x1_ASAP7_75t_R _20528_ (.A(_12172_),
    .Y(_12174_),
    .B(_12173_));
 NOR2x1_ASAP7_75t_R _20529_ (.A(_12171_),
    .B(_12174_),
    .Y(_12175_));
 AO21x1_ASAP7_75t_R _20530_ (.A1(_12174_),
    .A2(_12171_),
    .B(_10643_),
    .Y(_12176_));
 AND2x2_ASAP7_75t_R _20531_ (.A(net866),
    .B(_00673_),
    .Y(_12177_));
 INVx1_ASAP7_75t_R _20532_ (.A(_12177_),
    .Y(_12178_));
 OAI21x1_ASAP7_75t_R _20533_ (.A1(_12175_),
    .A2(_12176_),
    .B(_12178_),
    .Y(_12179_));
 INVx1_ASAP7_75t_R _20534_ (.A(_08211_),
    .Y(_12180_));
 XOR2x2_ASAP7_75t_R _20535_ (.A(_12179_),
    .B(_12180_),
    .Y(_12181_));
 BUFx12_ASAP7_75t_R _20536_ (.A(_12181_),
    .Y(_12182_));
 BUFx6f_ASAP7_75t_R _20537_ (.A(_12182_),
    .Y(_12183_));
 XOR2x2_ASAP7_75t_R _20538_ (.A(_00751_),
    .B(_12085_),
    .Y(_12184_));
 INVx1_ASAP7_75t_R _20539_ (.A(_00784_),
    .Y(_12185_));
 XOR2x1_ASAP7_75t_R _20540_ (.A(_12184_),
    .Y(_12186_),
    .B(_12185_));
 XNOR2x2_ASAP7_75t_R _20541_ (.A(_00783_),
    .B(_12080_),
    .Y(_12187_));
 XOR2x2_ASAP7_75t_R _20542_ (.A(_00816_),
    .B(_00848_),
    .Y(_12188_));
 XOR2x1_ASAP7_75t_R _20543_ (.A(_12187_),
    .Y(_12189_),
    .B(_12188_));
 NOR2x1_ASAP7_75t_R _20544_ (.A(_12186_),
    .B(_12189_),
    .Y(_12190_));
 AO21x1_ASAP7_75t_R _20545_ (.A1(_12189_),
    .A2(_12186_),
    .B(_11374_),
    .Y(_12191_));
 NAND2x1_ASAP7_75t_R _20546_ (.A(_00671_),
    .B(_12095_),
    .Y(_12192_));
 OAI21x1_ASAP7_75t_R _20547_ (.A1(_12190_),
    .A2(_12191_),
    .B(_12192_),
    .Y(_12193_));
 XOR2x2_ASAP7_75t_R _20548_ (.A(_12193_),
    .B(_01079_),
    .Y(_12194_));
 BUFx6f_ASAP7_75t_R _20549_ (.A(_12194_),
    .Y(_12195_));
 AO21x1_ASAP7_75t_R _20550_ (.A1(_12168_),
    .A2(_12183_),
    .B(_12195_),
    .Y(_12196_));
 INVx1_ASAP7_75t_R _20551_ (.A(_12079_),
    .Y(_12197_));
 NAND2x1_ASAP7_75t_R _20552_ (.A(_10829_),
    .B(net848),
    .Y(_12198_));
 AOI21x1_ASAP7_75t_R _20553_ (.A1(_12197_),
    .A2(_12198_),
    .B(_12101_),
    .Y(_12199_));
 AOI211x1_ASAP7_75t_R _20554_ (.A1(net848),
    .A2(_10786_),
    .B(_12079_),
    .C(_08190_),
    .Y(_12200_));
 OAI21x1_ASAP7_75t_R _20555_ (.A1(_12199_),
    .A2(_12200_),
    .B(_12124_),
    .Y(_12201_));
 INVx3_ASAP7_75t_R _20556_ (.A(_12201_),
    .Y(_12202_));
 XOR2x2_ASAP7_75t_R _20557_ (.A(_12179_),
    .B(_08211_),
    .Y(_12203_));
 OAI21x1_ASAP7_75t_R _20558_ (.A1(_15840_),
    .A2(_12153_),
    .B(_12203_),
    .Y(_12204_));
 AOI21x1_ASAP7_75t_R _20559_ (.A1(_15845_),
    .A2(_12202_),
    .B(_12204_),
    .Y(_12205_));
 NOR2x1_ASAP7_75t_R _20560_ (.A(_12196_),
    .B(_12205_),
    .Y(_12206_));
 BUFx6f_ASAP7_75t_R _20561_ (.A(_12203_),
    .Y(_12207_));
 OA21x2_ASAP7_75t_R _20562_ (.A1(_12207_),
    .A2(_12167_),
    .B(_12194_),
    .Y(_12208_));
 INVx1_ASAP7_75t_R _20563_ (.A(_12208_),
    .Y(_12209_));
 BUFx6f_ASAP7_75t_R _20564_ (.A(_12203_),
    .Y(_12210_));
 INVx3_ASAP7_75t_R _20565_ (.A(net497),
    .Y(_12211_));
 AO21x2_ASAP7_75t_R _20566_ (.A1(_12151_),
    .A2(_12149_),
    .B(_12211_),
    .Y(_12212_));
 NOR3x1_ASAP7_75t_R _20567_ (.A(_12162_),
    .B(_08197_),
    .C(_12141_),
    .Y(_12213_));
 OA21x2_ASAP7_75t_R _20568_ (.A1(_12162_),
    .A2(_12141_),
    .B(_08197_),
    .Y(_12214_));
 INVx2_ASAP7_75t_R _20569_ (.A(_01169_),
    .Y(_12215_));
 OAI21x1_ASAP7_75t_R _20570_ (.A1(_12213_),
    .A2(_12214_),
    .B(_12215_),
    .Y(_12216_));
 NOR2x1_ASAP7_75t_R _20571_ (.A(_12216_),
    .B(_12207_),
    .Y(_12217_));
 AO21x1_ASAP7_75t_R _20572_ (.A1(_12210_),
    .A2(_12212_),
    .B(_12217_),
    .Y(_12218_));
 XOR2x2_ASAP7_75t_R _20573_ (.A(_00753_),
    .B(_00785_),
    .Y(_12219_));
 XOR2x2_ASAP7_75t_R _20574_ (.A(_00786_),
    .B(_00818_),
    .Y(_12220_));
 XOR2x1_ASAP7_75t_R _20575_ (.A(_12220_),
    .Y(_12221_),
    .B(_00850_));
 XNOR2x1_ASAP7_75t_R _20576_ (.B(_12221_),
    .Y(_12222_),
    .A(_12219_));
 NOR2x1_ASAP7_75t_R _20577_ (.A(_10787_),
    .B(_00669_),
    .Y(_12223_));
 AO21x1_ASAP7_75t_R _20578_ (.A1(_12222_),
    .A2(_10786_),
    .B(_12223_),
    .Y(_12224_));
 XNOR2x2_ASAP7_75t_R _20579_ (.A(_01082_),
    .B(_12224_),
    .Y(_12225_));
 BUFx10_ASAP7_75t_R _20580_ (.A(_12225_),
    .Y(_12226_));
 OAI21x1_ASAP7_75t_R _20581_ (.A1(_12209_),
    .A2(_12218_),
    .B(_12226_),
    .Y(_12227_));
 NOR2x1_ASAP7_75t_R _20582_ (.A(_12206_),
    .B(_12227_),
    .Y(_12228_));
 BUFx10_ASAP7_75t_R _20583_ (.A(_12181_),
    .Y(_12229_));
 BUFx6f_ASAP7_75t_R _20584_ (.A(_12229_),
    .Y(_12230_));
 NOR2x1_ASAP7_75t_R _20585_ (.A(_01172_),
    .B(_12230_),
    .Y(_12231_));
 BUFx4f_ASAP7_75t_R _20586_ (.A(_12143_),
    .Y(_12232_));
 BUFx4f_ASAP7_75t_R _20587_ (.A(_12144_),
    .Y(_12233_));
 AOI21x1_ASAP7_75t_R _20588_ (.A1(_12232_),
    .A2(_12233_),
    .B(net498),
    .Y(_12234_));
 XOR2x2_ASAP7_75t_R _20589_ (.A(_12193_),
    .B(_08323_),
    .Y(_12235_));
 AO21x1_ASAP7_75t_R _20590_ (.A1(_12229_),
    .A2(_12234_),
    .B(_12235_),
    .Y(_12236_));
 INVx8_ASAP7_75t_R _20591_ (.A(_12225_),
    .Y(_12237_));
 OAI21x1_ASAP7_75t_R _20592_ (.A1(_12231_),
    .A2(_12236_),
    .B(_12237_),
    .Y(_12238_));
 OAI21x1_ASAP7_75t_R _20593_ (.A1(_12093_),
    .A2(_12079_),
    .B(_12101_),
    .Y(_12239_));
 INVx1_ASAP7_75t_R _20594_ (.A(_12239_),
    .Y(_12240_));
 OAI21x1_ASAP7_75t_R _20595_ (.A1(_12096_),
    .A2(_12100_),
    .B(_08190_),
    .Y(_12241_));
 INVx1_ASAP7_75t_R _20596_ (.A(_12241_),
    .Y(_12242_));
 OAI21x1_ASAP7_75t_R _20597_ (.A1(_12240_),
    .A2(_12242_),
    .B(_12153_),
    .Y(_12243_));
 OAI21x1_ASAP7_75t_R _20598_ (.A1(_15835_),
    .A2(_15848_),
    .B(_12167_),
    .Y(_12244_));
 INVx1_ASAP7_75t_R _20599_ (.A(_12244_),
    .Y(_12245_));
 BUFx6f_ASAP7_75t_R _20600_ (.A(_12207_),
    .Y(_12246_));
 AOI21x1_ASAP7_75t_R _20601_ (.A1(_12243_),
    .A2(_12245_),
    .B(_12246_),
    .Y(_12247_));
 INVx2_ASAP7_75t_R _20602_ (.A(_00513_),
    .Y(_12248_));
 AOI21x1_ASAP7_75t_R _20603_ (.A1(_12149_),
    .A2(_12151_),
    .B(_12248_),
    .Y(_12249_));
 NOR2x2_ASAP7_75t_R _20604_ (.A(net529),
    .B(_12152_),
    .Y(_12250_));
 NOR2x1_ASAP7_75t_R _20605_ (.A(_12249_),
    .B(_12250_),
    .Y(_12251_));
 AOI21x1_ASAP7_75t_R _20606_ (.A1(_12232_),
    .A2(_12233_),
    .B(_01167_),
    .Y(_12252_));
 AOI21x1_ASAP7_75t_R _20607_ (.A1(_12252_),
    .A2(_12182_),
    .B(_12194_),
    .Y(_12253_));
 OAI21x1_ASAP7_75t_R _20608_ (.A1(_12230_),
    .A2(_12251_),
    .B(_12253_),
    .Y(_12254_));
 NOR2x1_ASAP7_75t_R _20609_ (.A(_12247_),
    .B(_12254_),
    .Y(_12255_));
 XOR2x2_ASAP7_75t_R _20610_ (.A(_00752_),
    .B(_00784_),
    .Y(_12256_));
 INVx1_ASAP7_75t_R _20611_ (.A(_12256_),
    .Y(_12257_));
 XOR2x2_ASAP7_75t_R _20612_ (.A(_00785_),
    .B(_00817_),
    .Y(_12258_));
 BUFx6f_ASAP7_75t_R _20613_ (.A(_00849_),
    .Y(_12259_));
 INVx3_ASAP7_75t_R _20614_ (.A(_12259_),
    .Y(_12260_));
 XOR2x1_ASAP7_75t_R _20615_ (.A(_12258_),
    .Y(_12261_),
    .B(_12260_));
 NAND2x1_ASAP7_75t_R _20616_ (.A(_12257_),
    .B(_12261_),
    .Y(_12262_));
 XOR2x1_ASAP7_75t_R _20617_ (.A(_12258_),
    .Y(_12263_),
    .B(_12259_));
 NAND2x1_ASAP7_75t_R _20618_ (.A(_12256_),
    .B(_12263_),
    .Y(_12264_));
 AOI21x1_ASAP7_75t_R _20619_ (.A1(_12262_),
    .A2(_12264_),
    .B(_12161_),
    .Y(_12265_));
 NOR2x1_ASAP7_75t_R _20620_ (.A(_10787_),
    .B(_00670_),
    .Y(_12266_));
 OA21x2_ASAP7_75t_R _20621_ (.A1(_12265_),
    .A2(_12266_),
    .B(_01080_),
    .Y(_12267_));
 INVx1_ASAP7_75t_R _20622_ (.A(_00670_),
    .Y(_12268_));
 AOI211x1_ASAP7_75t_R _20623_ (.A1(_12161_),
    .A2(_12268_),
    .B(_12265_),
    .C(_01080_),
    .Y(_12269_));
 NOR2x2_ASAP7_75t_R _20624_ (.A(_12267_),
    .B(_12269_),
    .Y(_12270_));
 BUFx6f_ASAP7_75t_R _20625_ (.A(_12270_),
    .Y(_12271_));
 BUFx10_ASAP7_75t_R _20626_ (.A(_12271_),
    .Y(_12272_));
 OAI21x1_ASAP7_75t_R _20627_ (.A1(_12238_),
    .A2(_12255_),
    .B(_12272_),
    .Y(_12273_));
 XNOR2x2_ASAP7_75t_R _20628_ (.A(_00754_),
    .B(_00786_),
    .Y(_12274_));
 BUFx12f_ASAP7_75t_R _20629_ (.A(_00851_),
    .Y(_12275_));
 INVx5_ASAP7_75t_R _20630_ (.A(_12275_),
    .Y(_12276_));
 XOR2x1_ASAP7_75t_R _20631_ (.A(_12274_),
    .Y(_12277_),
    .B(_12276_));
 BUFx2_ASAP7_75t_R rebuffer381 (.A(_12130_),
    .Y(net834));
 XNOR2x2_ASAP7_75t_R _20633_ (.A(_12108_),
    .B(net40),
    .Y(_12279_));
 XOR2x1_ASAP7_75t_R _20634_ (.A(_12277_),
    .Y(_12280_),
    .B(_12279_));
 NOR2x1_ASAP7_75t_R _20635_ (.A(_10831_),
    .B(_00668_),
    .Y(_12281_));
 AO21x1_ASAP7_75t_R _20636_ (.A1(_12280_),
    .A2(_10830_),
    .B(_12281_),
    .Y(_12282_));
 XOR2x2_ASAP7_75t_R _20637_ (.A(_12282_),
    .B(_01083_),
    .Y(_12283_));
 INVx4_ASAP7_75t_R _20638_ (.A(_12283_),
    .Y(_12284_));
 OAI21x1_ASAP7_75t_R _20639_ (.A1(_12228_),
    .A2(_12273_),
    .B(_12284_),
    .Y(_12285_));
 BUFx12_ASAP7_75t_R _20640_ (.A(_12145_),
    .Y(_12286_));
 OAI21x1_ASAP7_75t_R _20641_ (.A1(_12199_),
    .A2(_12200_),
    .B(_12148_),
    .Y(_12287_));
 NOR2x2_ASAP7_75t_R _20642_ (.A(_12286_),
    .B(_12287_),
    .Y(_12288_));
 AOI21x1_ASAP7_75t_R _20643_ (.A1(_12232_),
    .A2(_12233_),
    .B(_12215_),
    .Y(_12289_));
 NOR2x2_ASAP7_75t_R _20644_ (.A(_12182_),
    .B(_12289_),
    .Y(_12290_));
 INVx1_ASAP7_75t_R _20645_ (.A(_12290_),
    .Y(_12291_));
 AOI21x1_ASAP7_75t_R _20646_ (.A1(_12149_),
    .A2(_12151_),
    .B(_01167_),
    .Y(_12292_));
 BUFx6f_ASAP7_75t_R _20647_ (.A(_12194_),
    .Y(_12293_));
 AOI21x1_ASAP7_75t_R _20648_ (.A1(_12292_),
    .A2(_12183_),
    .B(_12293_),
    .Y(_12294_));
 OA21x2_ASAP7_75t_R _20649_ (.A1(_12288_),
    .A2(_12291_),
    .B(_12294_),
    .Y(_12295_));
 BUFx6f_ASAP7_75t_R _20650_ (.A(_12203_),
    .Y(_12296_));
 AO21x1_ASAP7_75t_R _20651_ (.A1(_12296_),
    .A2(_12292_),
    .B(_12235_),
    .Y(_12297_));
 INVx2_ASAP7_75t_R _20652_ (.A(_00511_),
    .Y(_12298_));
 AOI21x1_ASAP7_75t_R _20653_ (.A1(_12298_),
    .A2(_12286_),
    .B(_12203_),
    .Y(_12299_));
 INVx1_ASAP7_75t_R _20654_ (.A(_12299_),
    .Y(_12300_));
 NOR2x1_ASAP7_75t_R _20655_ (.A(_12300_),
    .B(_12288_),
    .Y(_12301_));
 OAI21x1_ASAP7_75t_R _20656_ (.A1(_12297_),
    .A2(_12301_),
    .B(_12237_),
    .Y(_12302_));
 INVx6_ASAP7_75t_R _20657_ (.A(_12270_),
    .Y(_12303_));
 BUFx10_ASAP7_75t_R _20658_ (.A(_12303_),
    .Y(_12304_));
 OAI21x1_ASAP7_75t_R _20659_ (.A1(_12295_),
    .A2(_12302_),
    .B(_12304_),
    .Y(_12305_));
 AOI21x1_ASAP7_75t_R _20660_ (.A1(_12165_),
    .A2(_12153_),
    .B(_12229_),
    .Y(_12306_));
 BUFx10_ASAP7_75t_R _20661_ (.A(_12152_),
    .Y(_12307_));
 NOR2x2_ASAP7_75t_R _20662_ (.A(_12248_),
    .B(_12307_),
    .Y(_12308_));
 BUFx6f_ASAP7_75t_R _20663_ (.A(_12182_),
    .Y(_12309_));
 OA21x2_ASAP7_75t_R _20664_ (.A1(_12308_),
    .A2(_12292_),
    .B(_12309_),
    .Y(_12310_));
 BUFx6f_ASAP7_75t_R _20665_ (.A(_12194_),
    .Y(_12311_));
 OAI21x1_ASAP7_75t_R _20666_ (.A1(_12306_),
    .A2(_12310_),
    .B(_12311_),
    .Y(_12312_));
 AO21x2_ASAP7_75t_R _20667_ (.A1(_12233_),
    .A2(_12232_),
    .B(_12298_),
    .Y(_12313_));
 INVx1_ASAP7_75t_R _20668_ (.A(_12313_),
    .Y(_12314_));
 NOR2x2_ASAP7_75t_R _20669_ (.A(_12148_),
    .B(_12145_),
    .Y(_12315_));
 OA21x2_ASAP7_75t_R _20670_ (.A1(_12314_),
    .A2(_12315_),
    .B(_12210_),
    .Y(_12316_));
 AOI21x1_ASAP7_75t_R _20671_ (.A1(_12153_),
    .A2(net865),
    .B(_12296_),
    .Y(_12317_));
 INVx2_ASAP7_75t_R _20672_ (.A(_12234_),
    .Y(_12318_));
 AND2x2_ASAP7_75t_R _20673_ (.A(_12317_),
    .B(_12318_),
    .Y(_12319_));
 BUFx6f_ASAP7_75t_R _20674_ (.A(_12235_),
    .Y(_12320_));
 BUFx10_ASAP7_75t_R _20675_ (.A(_12320_),
    .Y(_12321_));
 OAI21x1_ASAP7_75t_R _20676_ (.A1(_12316_),
    .A2(_12319_),
    .B(_12321_),
    .Y(_12322_));
 BUFx10_ASAP7_75t_R _20677_ (.A(_12237_),
    .Y(_12323_));
 AOI21x1_ASAP7_75t_R _20678_ (.A1(_12312_),
    .A2(_12322_),
    .B(_12323_),
    .Y(_12324_));
 NOR2x1_ASAP7_75t_R _20679_ (.A(_12305_),
    .B(_12324_),
    .Y(_12325_));
 AO21x2_ASAP7_75t_R _20680_ (.A1(_12233_),
    .A2(_12232_),
    .B(_12248_),
    .Y(_12326_));
 AOI21x1_ASAP7_75t_R _20681_ (.A1(_12149_),
    .A2(_12151_),
    .B(net498),
    .Y(_12327_));
 INVx2_ASAP7_75t_R _20682_ (.A(_12327_),
    .Y(_12328_));
 AO21x1_ASAP7_75t_R _20683_ (.A1(_12326_),
    .A2(_12328_),
    .B(_12309_),
    .Y(_12329_));
 INVx2_ASAP7_75t_R _20684_ (.A(_12249_),
    .Y(_12330_));
 BUFx6f_ASAP7_75t_R _20685_ (.A(_12203_),
    .Y(_12331_));
 AO21x1_ASAP7_75t_R _20686_ (.A1(_12313_),
    .A2(_12330_),
    .B(_12331_),
    .Y(_12332_));
 AO21x1_ASAP7_75t_R _20687_ (.A1(_12332_),
    .A2(_12329_),
    .B(_12311_),
    .Y(_12333_));
 BUFx6f_ASAP7_75t_R _20688_ (.A(_12235_),
    .Y(_12334_));
 AOI21x1_ASAP7_75t_R _20689_ (.A1(_12232_),
    .A2(_12233_),
    .B(_12211_),
    .Y(_12335_));
 NOR2x2_ASAP7_75t_R _20690_ (.A(_12181_),
    .B(_12335_),
    .Y(_12336_));
 NOR2x2_ASAP7_75t_R _20691_ (.A(_12336_),
    .B(_12334_),
    .Y(_12337_));
 NAND2x2_ASAP7_75t_R _20692_ (.A(_12239_),
    .B(_12241_),
    .Y(_12338_));
 NAND2x2_ASAP7_75t_R _20693_ (.A(_12286_),
    .B(net847),
    .Y(_12339_));
 AO21x1_ASAP7_75t_R _20694_ (.A1(_12339_),
    .A2(_12212_),
    .B(_12246_),
    .Y(_12340_));
 AOI21x1_ASAP7_75t_R _20695_ (.A1(_12340_),
    .A2(_12337_),
    .B(_12304_),
    .Y(_12341_));
 NAND2x1_ASAP7_75t_R _20696_ (.A(_12333_),
    .B(_12341_),
    .Y(_12342_));
 NAND2x2_ASAP7_75t_R _20697_ (.A(_12229_),
    .B(_12212_),
    .Y(_12343_));
 NOR2x2_ASAP7_75t_R _20698_ (.A(_12307_),
    .B(_12201_),
    .Y(_12344_));
 NOR2x1_ASAP7_75t_R _20699_ (.A(_12343_),
    .B(_12344_),
    .Y(_12345_));
 BUFx10_ASAP7_75t_R _20700_ (.A(_12235_),
    .Y(_12346_));
 NOR2x2_ASAP7_75t_R _20701_ (.A(_12298_),
    .B(_12286_),
    .Y(_12347_));
 BUFx6f_ASAP7_75t_R _20702_ (.A(_12296_),
    .Y(_12348_));
 OAI21x1_ASAP7_75t_R _20703_ (.A1(_12308_),
    .A2(_12347_),
    .B(_12348_),
    .Y(_12349_));
 NAND2x1_ASAP7_75t_R _20704_ (.A(_12346_),
    .B(_12349_),
    .Y(_12350_));
 NOR2x1_ASAP7_75t_R _20705_ (.A(_12345_),
    .B(_12350_),
    .Y(_12351_));
 NAND2x2_ASAP7_75t_R _20706_ (.A(_12124_),
    .B(_12145_),
    .Y(_12352_));
 AOI21x1_ASAP7_75t_R _20707_ (.A1(_12148_),
    .A2(_12103_),
    .B(_12182_),
    .Y(_12353_));
 BUFx6f_ASAP7_75t_R _20708_ (.A(_12287_),
    .Y(_12354_));
 AOI21x1_ASAP7_75t_R _20709_ (.A1(_12352_),
    .A2(_12354_),
    .B(_12246_),
    .Y(_12355_));
 AOI211x1_ASAP7_75t_R _20710_ (.A1(_12352_),
    .A2(_12353_),
    .B(_12355_),
    .C(_12321_),
    .Y(_12356_));
 OAI21x1_ASAP7_75t_R _20711_ (.A1(_12351_),
    .A2(_12356_),
    .B(_12304_),
    .Y(_12357_));
 AOI21x1_ASAP7_75t_R _20712_ (.A1(_12357_),
    .A2(_12342_),
    .B(_12226_),
    .Y(_12358_));
 NOR2x1_ASAP7_75t_R _20713_ (.A(_15845_),
    .B(_12354_),
    .Y(_12359_));
 INVx1_ASAP7_75t_R _20714_ (.A(_12359_),
    .Y(_12360_));
 AOI21x1_ASAP7_75t_R _20715_ (.A1(_12239_),
    .A2(_12241_),
    .B(_12145_),
    .Y(_12361_));
 NOR2x2_ASAP7_75t_R _20716_ (.A(_12210_),
    .B(_12361_),
    .Y(_12362_));
 INVx3_ASAP7_75t_R _20717_ (.A(_01170_),
    .Y(_12363_));
 NOR2x2_ASAP7_75t_R _20718_ (.A(_12363_),
    .B(_12145_),
    .Y(_12364_));
 BUFx10_ASAP7_75t_R _20719_ (.A(_12194_),
    .Y(_12365_));
 OAI21x1_ASAP7_75t_R _20720_ (.A1(_12364_),
    .A2(_12204_),
    .B(_12365_),
    .Y(_12366_));
 AOI21x1_ASAP7_75t_R _20721_ (.A1(_12360_),
    .A2(_12362_),
    .B(_12366_),
    .Y(_12367_));
 OAI21x1_ASAP7_75t_R _20722_ (.A1(_12246_),
    .A2(_12339_),
    .B(_12294_),
    .Y(_12368_));
 BUFx6f_ASAP7_75t_R _20723_ (.A(_12271_),
    .Y(_12369_));
 OAI21x1_ASAP7_75t_R _20724_ (.A1(_12368_),
    .A2(_12205_),
    .B(_12369_),
    .Y(_12370_));
 NOR2x1_ASAP7_75t_R _20725_ (.A(_12367_),
    .B(_12370_),
    .Y(_12371_));
 NOR2x2_ASAP7_75t_R _20726_ (.A(_12211_),
    .B(_12145_),
    .Y(_12372_));
 AOI21x1_ASAP7_75t_R _20727_ (.A1(_12232_),
    .A2(_12233_),
    .B(_12363_),
    .Y(_12373_));
 NOR2x2_ASAP7_75t_R _20728_ (.A(_12373_),
    .B(_12182_),
    .Y(_12374_));
 INVx2_ASAP7_75t_R _20729_ (.A(_12374_),
    .Y(_12375_));
 OAI21x1_ASAP7_75t_R _20730_ (.A1(_12372_),
    .A2(_12375_),
    .B(_12365_),
    .Y(_12376_));
 BUFx6f_ASAP7_75t_R _20731_ (.A(_12181_),
    .Y(_12377_));
 NAND2x2_ASAP7_75t_R _20732_ (.A(net529),
    .B(_12152_),
    .Y(_12378_));
 NAND2x1_ASAP7_75t_R _20733_ (.A(_12377_),
    .B(_12378_),
    .Y(_12379_));
 NOR2x1_ASAP7_75t_R _20734_ (.A(_12379_),
    .B(_12359_),
    .Y(_12380_));
 NOR2x1_ASAP7_75t_R _20735_ (.A(_12376_),
    .B(_12380_),
    .Y(_12381_));
 NAND2x2_ASAP7_75t_R _20736_ (.A(net592),
    .B(_12145_),
    .Y(_12382_));
 BUFx6f_ASAP7_75t_R _20737_ (.A(_12229_),
    .Y(_12383_));
 BUFx6f_ASAP7_75t_R _20738_ (.A(_12194_),
    .Y(_12384_));
 AO21x1_ASAP7_75t_R _20739_ (.A1(_12382_),
    .A2(_12383_),
    .B(_12384_),
    .Y(_12385_));
 INVx1_ASAP7_75t_R _20740_ (.A(_12354_),
    .Y(_12386_));
 OAI21x1_ASAP7_75t_R _20741_ (.A1(_12166_),
    .A2(_12286_),
    .B(_12296_),
    .Y(_12387_));
 AOI21x1_ASAP7_75t_R _20742_ (.A1(_15848_),
    .A2(_12386_),
    .B(_12387_),
    .Y(_12388_));
 OAI21x1_ASAP7_75t_R _20743_ (.A1(_12385_),
    .A2(_12388_),
    .B(_12304_),
    .Y(_12389_));
 OAI21x1_ASAP7_75t_R _20744_ (.A1(_12381_),
    .A2(_12389_),
    .B(_12226_),
    .Y(_12390_));
 BUFx10_ASAP7_75t_R _20745_ (.A(_12283_),
    .Y(_12391_));
 OAI21x1_ASAP7_75t_R _20746_ (.A1(_12371_),
    .A2(_12390_),
    .B(_12391_),
    .Y(_12392_));
 OAI22x1_ASAP7_75t_R _20747_ (.A1(_12285_),
    .A2(_12325_),
    .B1(_12358_),
    .B2(_12392_),
    .Y(_00048_));
 OAI21x1_ASAP7_75t_R _20748_ (.A1(_12307_),
    .A2(_12201_),
    .B(_12331_),
    .Y(_12393_));
 AO21x1_ASAP7_75t_R _20749_ (.A1(_12151_),
    .A2(_12149_),
    .B(_12165_),
    .Y(_12394_));
 OA21x2_ASAP7_75t_R _20750_ (.A1(_12394_),
    .A2(_12207_),
    .B(_12235_),
    .Y(_12395_));
 OAI21x1_ASAP7_75t_R _20751_ (.A1(_12327_),
    .A2(_12393_),
    .B(_12395_),
    .Y(_12396_));
 NOR2x2_ASAP7_75t_R _20752_ (.A(_15840_),
    .B(_12286_),
    .Y(_12397_));
 OAI21x1_ASAP7_75t_R _20753_ (.A1(_12397_),
    .A2(_12361_),
    .B(_12309_),
    .Y(_12398_));
 AOI21x1_ASAP7_75t_R _20754_ (.A1(_12243_),
    .A2(_12374_),
    .B(_12334_),
    .Y(_12399_));
 AOI21x1_ASAP7_75t_R _20755_ (.A1(_12398_),
    .A2(_12399_),
    .B(_12271_),
    .Y(_12400_));
 AOI21x1_ASAP7_75t_R _20756_ (.A1(_12396_),
    .A2(_12400_),
    .B(_12237_),
    .Y(_12401_));
 OAI21x1_ASAP7_75t_R _20757_ (.A1(_12249_),
    .A2(_12250_),
    .B(_12309_),
    .Y(_12402_));
 AO21x1_ASAP7_75t_R _20758_ (.A1(_12212_),
    .A2(_12167_),
    .B(_12377_),
    .Y(_12403_));
 AOI21x1_ASAP7_75t_R _20759_ (.A1(_12402_),
    .A2(_12403_),
    .B(_12346_),
    .Y(_12404_));
 NOR2x1_ASAP7_75t_R _20760_ (.A(_12234_),
    .B(_12296_),
    .Y(_12405_));
 NAND2x1_ASAP7_75t_R _20761_ (.A(_12378_),
    .B(_12405_),
    .Y(_12406_));
 OAI21x1_ASAP7_75t_R _20762_ (.A1(_12397_),
    .A2(_12202_),
    .B(_12348_),
    .Y(_12407_));
 AOI21x1_ASAP7_75t_R _20763_ (.A1(_12406_),
    .A2(_12407_),
    .B(_12384_),
    .Y(_12408_));
 OAI21x1_ASAP7_75t_R _20764_ (.A1(_12404_),
    .A2(_12408_),
    .B(_12369_),
    .Y(_12409_));
 NAND2x1_ASAP7_75t_R _20765_ (.A(_12401_),
    .B(_12409_),
    .Y(_12410_));
 AOI21x1_ASAP7_75t_R _20766_ (.A1(_15845_),
    .A2(_12354_),
    .B(_12168_),
    .Y(_12411_));
 AO21x2_ASAP7_75t_R _20767_ (.A1(_12151_),
    .A2(_12149_),
    .B(_12363_),
    .Y(_12412_));
 AOI21x1_ASAP7_75t_R _20768_ (.A1(_12336_),
    .A2(_12412_),
    .B(_12293_),
    .Y(_12413_));
 OAI21x1_ASAP7_75t_R _20769_ (.A1(_12246_),
    .A2(_12411_),
    .B(_12413_),
    .Y(_12414_));
 NAND2x2_ASAP7_75t_R _20770_ (.A(_12286_),
    .B(net865),
    .Y(_12415_));
 AOI21x1_ASAP7_75t_R _20771_ (.A1(_12331_),
    .A2(_12415_),
    .B(_12361_),
    .Y(_12416_));
 AOI21x1_ASAP7_75t_R _20772_ (.A1(_12208_),
    .A2(_12416_),
    .B(_12303_),
    .Y(_12417_));
 AOI21x1_ASAP7_75t_R _20773_ (.A1(_12417_),
    .A2(_12414_),
    .B(_12225_),
    .Y(_12418_));
 AO21x1_ASAP7_75t_R _20774_ (.A1(_12382_),
    .A2(_12394_),
    .B(_12207_),
    .Y(_12419_));
 OA21x2_ASAP7_75t_R _20775_ (.A1(_12204_),
    .A2(_12372_),
    .B(_12194_),
    .Y(_12420_));
 NAND2x1_ASAP7_75t_R _20776_ (.A(_12419_),
    .B(_12420_),
    .Y(_12421_));
 NOR2x2_ASAP7_75t_R _20777_ (.A(_12153_),
    .B(_12182_),
    .Y(_12422_));
 NAND2x1_ASAP7_75t_R _20778_ (.A(_12354_),
    .B(_12422_),
    .Y(_12423_));
 BUFx6f_ASAP7_75t_R _20779_ (.A(_12338_),
    .Y(_15836_));
 NAND2x1_ASAP7_75t_R _20780_ (.A(net529),
    .B(_15836_),
    .Y(_12424_));
 AOI21x1_ASAP7_75t_R _20781_ (.A1(_12424_),
    .A2(_12317_),
    .B(_12293_),
    .Y(_12425_));
 BUFx10_ASAP7_75t_R _20782_ (.A(_12270_),
    .Y(_12426_));
 AOI21x1_ASAP7_75t_R _20783_ (.A1(_12423_),
    .A2(_12425_),
    .B(_12426_),
    .Y(_12427_));
 NAND2x1_ASAP7_75t_R _20784_ (.A(_12421_),
    .B(_12427_),
    .Y(_12428_));
 NAND2x1_ASAP7_75t_R _20785_ (.A(_12428_),
    .B(_12418_),
    .Y(_12429_));
 AOI21x1_ASAP7_75t_R _20786_ (.A1(_12410_),
    .A2(_12429_),
    .B(_12391_),
    .Y(_12430_));
 INVx1_ASAP7_75t_R _20787_ (.A(_12252_),
    .Y(_12431_));
 AO21x1_ASAP7_75t_R _20788_ (.A1(_12151_),
    .A2(_12149_),
    .B(_01170_),
    .Y(_12432_));
 NAND2x1_ASAP7_75t_R _20789_ (.A(_12431_),
    .B(_12432_),
    .Y(_12433_));
 AOI21x1_ASAP7_75t_R _20790_ (.A1(_12183_),
    .A2(_12433_),
    .B(_12334_),
    .Y(_12434_));
 OAI21x1_ASAP7_75t_R _20791_ (.A1(_12327_),
    .A2(_12393_),
    .B(_12434_),
    .Y(_12435_));
 NOR2x2_ASAP7_75t_R _20792_ (.A(_12372_),
    .B(_12181_),
    .Y(_12436_));
 NOR2x1_ASAP7_75t_R _20793_ (.A(_12293_),
    .B(_12436_),
    .Y(_12437_));
 NAND2x2_ASAP7_75t_R _20794_ (.A(_12103_),
    .B(_12315_),
    .Y(_12438_));
 OA21x2_ASAP7_75t_R _20795_ (.A1(_15840_),
    .A2(_12152_),
    .B(_12182_),
    .Y(_12439_));
 NAND2x2_ASAP7_75t_R _20796_ (.A(_12438_),
    .B(_12439_),
    .Y(_12440_));
 AOI21x1_ASAP7_75t_R _20797_ (.A1(_12437_),
    .A2(_12440_),
    .B(_12303_),
    .Y(_12441_));
 NAND2x1_ASAP7_75t_R _20798_ (.A(_12435_),
    .B(_12441_),
    .Y(_12442_));
 AO21x1_ASAP7_75t_R _20799_ (.A1(_12318_),
    .A2(_12330_),
    .B(_12377_),
    .Y(_12443_));
 INVx1_ASAP7_75t_R _20800_ (.A(_12292_),
    .Y(_12444_));
 AO21x1_ASAP7_75t_R _20801_ (.A1(_12352_),
    .A2(_12444_),
    .B(_12331_),
    .Y(_12445_));
 AOI21x1_ASAP7_75t_R _20802_ (.A1(_12443_),
    .A2(_12445_),
    .B(_12346_),
    .Y(_12446_));
 NAND2x1_ASAP7_75t_R _20803_ (.A(_12339_),
    .B(_12306_),
    .Y(_12447_));
 AO21x1_ASAP7_75t_R _20804_ (.A1(_12378_),
    .A2(_12326_),
    .B(_12331_),
    .Y(_12448_));
 AOI21x1_ASAP7_75t_R _20805_ (.A1(_12447_),
    .A2(_12448_),
    .B(_12365_),
    .Y(_12449_));
 BUFx10_ASAP7_75t_R _20806_ (.A(_12303_),
    .Y(_12450_));
 OAI21x1_ASAP7_75t_R _20807_ (.A1(_12446_),
    .A2(_12449_),
    .B(_12450_),
    .Y(_12451_));
 AOI21x1_ASAP7_75t_R _20808_ (.A1(_12442_),
    .A2(_12451_),
    .B(_12237_),
    .Y(_12452_));
 NOR2x2_ASAP7_75t_R _20809_ (.A(_12153_),
    .B(net865),
    .Y(_12453_));
 OA21x2_ASAP7_75t_R _20810_ (.A1(_12387_),
    .A2(_12453_),
    .B(_12293_),
    .Y(_12454_));
 NOR2x1_ASAP7_75t_R _20811_ (.A(_12296_),
    .B(_12315_),
    .Y(_12455_));
 AOI21x1_ASAP7_75t_R _20812_ (.A1(_12415_),
    .A2(_12455_),
    .B(_12303_),
    .Y(_12456_));
 AO21x1_ASAP7_75t_R _20813_ (.A1(_12454_),
    .A2(_12456_),
    .B(_12225_),
    .Y(_12457_));
 NAND2x2_ASAP7_75t_R _20814_ (.A(_12299_),
    .B(_12438_),
    .Y(_12458_));
 AO21x1_ASAP7_75t_R _20815_ (.A1(_12296_),
    .A2(_00515_),
    .B(_12194_),
    .Y(_12459_));
 NAND2x1_ASAP7_75t_R _20816_ (.A(_12271_),
    .B(_12459_),
    .Y(_12460_));
 OAI21x1_ASAP7_75t_R _20817_ (.A1(_12384_),
    .A2(_12458_),
    .B(_12460_),
    .Y(_12461_));
 NAND2x2_ASAP7_75t_R _20818_ (.A(_12124_),
    .B(_12152_),
    .Y(_12462_));
 BUFx6f_ASAP7_75t_R _20819_ (.A(_12203_),
    .Y(_12463_));
 AO21x1_ASAP7_75t_R _20820_ (.A1(_12462_),
    .A2(_12326_),
    .B(_12463_),
    .Y(_12464_));
 AOI21x1_ASAP7_75t_R _20821_ (.A1(_15840_),
    .A2(_15838_),
    .B(_15848_),
    .Y(_12465_));
 AOI21x1_ASAP7_75t_R _20822_ (.A1(net53),
    .A2(_15838_),
    .B(_12307_),
    .Y(_12466_));
 OAI21x1_ASAP7_75t_R _20823_ (.A1(_12465_),
    .A2(_12466_),
    .B(_12348_),
    .Y(_12467_));
 AOI21x1_ASAP7_75t_R _20824_ (.A1(_12464_),
    .A2(_12467_),
    .B(_12346_),
    .Y(_12468_));
 NOR2x1_ASAP7_75t_R _20825_ (.A(_12461_),
    .B(_12468_),
    .Y(_12469_));
 OAI21x1_ASAP7_75t_R _20826_ (.A1(_12457_),
    .A2(_12469_),
    .B(_12391_),
    .Y(_12470_));
 NOR2x1_ASAP7_75t_R _20827_ (.A(_12452_),
    .B(_12470_),
    .Y(_12471_));
 NOR2x1_ASAP7_75t_R _20828_ (.A(_12471_),
    .B(_12430_),
    .Y(_00049_));
 AND2x2_ASAP7_75t_R _20829_ (.A(_12165_),
    .B(_01167_),
    .Y(_12472_));
 NAND2x2_ASAP7_75t_R _20830_ (.A(_12472_),
    .B(_12153_),
    .Y(_12473_));
 NAND2x1_ASAP7_75t_R _20831_ (.A(_12331_),
    .B(_12473_),
    .Y(_12474_));
 NOR2x1_ASAP7_75t_R _20832_ (.A(_12474_),
    .B(_12344_),
    .Y(_12475_));
 AO21x1_ASAP7_75t_R _20833_ (.A1(_12438_),
    .A2(_12299_),
    .B(_12271_),
    .Y(_12476_));
 OA21x2_ASAP7_75t_R _20834_ (.A1(_01174_),
    .A2(_12463_),
    .B(_12271_),
    .Y(_12477_));
 NAND2x2_ASAP7_75t_R _20835_ (.A(_12153_),
    .B(_12103_),
    .Y(_12478_));
 NAND2x1_ASAP7_75t_R _20836_ (.A(_12478_),
    .B(_12353_),
    .Y(_12479_));
 AOI21x1_ASAP7_75t_R _20837_ (.A1(_12477_),
    .A2(_12479_),
    .B(_12346_),
    .Y(_12480_));
 OAI21x1_ASAP7_75t_R _20838_ (.A1(_12475_),
    .A2(_12476_),
    .B(_12480_),
    .Y(_12481_));
 OAI21x1_ASAP7_75t_R _20839_ (.A1(net10),
    .A2(_12382_),
    .B(_12377_),
    .Y(_12482_));
 NAND2x2_ASAP7_75t_R _20840_ (.A(_00516_),
    .B(_12207_),
    .Y(_12483_));
 NAND3x1_ASAP7_75t_R _20841_ (.A(_12482_),
    .B(_12271_),
    .C(_12483_),
    .Y(_12484_));
 AO21x1_ASAP7_75t_R _20842_ (.A1(_12328_),
    .A2(_12167_),
    .B(_12377_),
    .Y(_12485_));
 NAND2x1_ASAP7_75t_R _20843_ (.A(_12249_),
    .B(_12181_),
    .Y(_12486_));
 INVx2_ASAP7_75t_R _20844_ (.A(_12486_),
    .Y(_12487_));
 NOR2x1_ASAP7_75t_R _20845_ (.A(_12271_),
    .B(_12487_),
    .Y(_12488_));
 AOI21x1_ASAP7_75t_R _20846_ (.A1(_12485_),
    .A2(_12488_),
    .B(_12365_),
    .Y(_12489_));
 AOI21x1_ASAP7_75t_R _20847_ (.A1(_12484_),
    .A2(_12489_),
    .B(_12225_),
    .Y(_12490_));
 AOI21x1_ASAP7_75t_R _20848_ (.A1(_12490_),
    .A2(_12481_),
    .B(_12283_),
    .Y(_12491_));
 NAND2x1_ASAP7_75t_R _20849_ (.A(_12326_),
    .B(_12317_),
    .Y(_12492_));
 OR3x1_ASAP7_75t_R _20850_ (.A(_12347_),
    .B(_12234_),
    .C(_12183_),
    .Y(_12493_));
 BUFx6f_ASAP7_75t_R _20851_ (.A(_12334_),
    .Y(_12494_));
 AOI21x1_ASAP7_75t_R _20852_ (.A1(_12492_),
    .A2(_12493_),
    .B(_12494_),
    .Y(_12495_));
 AOI21x1_ASAP7_75t_R _20853_ (.A1(net53),
    .A2(net10),
    .B(_12229_),
    .Y(_12496_));
 AOI21x1_ASAP7_75t_R _20854_ (.A1(_12478_),
    .A2(_12496_),
    .B(_12195_),
    .Y(_12497_));
 NAND2x1_ASAP7_75t_R _20855_ (.A(_00515_),
    .B(_12383_),
    .Y(_12498_));
 AO21x1_ASAP7_75t_R _20856_ (.A1(_12497_),
    .A2(_12498_),
    .B(_12450_),
    .Y(_12499_));
 OA21x2_ASAP7_75t_R _20857_ (.A1(_12463_),
    .A2(_01172_),
    .B(_12334_),
    .Y(_12500_));
 OAI21x1_ASAP7_75t_R _20858_ (.A1(_15848_),
    .A2(_12354_),
    .B(_12336_),
    .Y(_12501_));
 AOI21x1_ASAP7_75t_R _20859_ (.A1(_12500_),
    .A2(_12501_),
    .B(_12426_),
    .Y(_12502_));
 AOI21x1_ASAP7_75t_R _20860_ (.A1(_12318_),
    .A2(_12317_),
    .B(_12334_),
    .Y(_12503_));
 AOI21x1_ASAP7_75t_R _20861_ (.A1(_12462_),
    .A2(_12415_),
    .B(_12229_),
    .Y(_12504_));
 INVx1_ASAP7_75t_R _20862_ (.A(_12504_),
    .Y(_12505_));
 NAND2x1_ASAP7_75t_R _20863_ (.A(_12503_),
    .B(_12505_),
    .Y(_12506_));
 AOI21x1_ASAP7_75t_R _20864_ (.A1(_12506_),
    .A2(_12502_),
    .B(_12237_),
    .Y(_12507_));
 OAI21x1_ASAP7_75t_R _20865_ (.A1(_12495_),
    .A2(_12499_),
    .B(_12507_),
    .Y(_12508_));
 NAND2x1_ASAP7_75t_R _20866_ (.A(_12508_),
    .B(_12491_),
    .Y(_12509_));
 NOR2x2_ASAP7_75t_R _20867_ (.A(_12203_),
    .B(_12327_),
    .Y(_12510_));
 OAI21x1_ASAP7_75t_R _20868_ (.A1(_15835_),
    .A2(_12286_),
    .B(_12296_),
    .Y(_12511_));
 NOR2x1_ASAP7_75t_R _20869_ (.A(_12252_),
    .B(_12511_),
    .Y(_12512_));
 AOI21x1_ASAP7_75t_R _20870_ (.A1(_12339_),
    .A2(_12510_),
    .B(_12512_),
    .Y(_12513_));
 OAI21x1_ASAP7_75t_R _20871_ (.A1(_12494_),
    .A2(_12513_),
    .B(_12450_),
    .Y(_12514_));
 OA211x2_ASAP7_75t_R _20872_ (.A1(_12364_),
    .A2(_12393_),
    .B(_12482_),
    .C(_12320_),
    .Y(_12515_));
 NOR2x1_ASAP7_75t_R _20873_ (.A(_12514_),
    .B(_12515_),
    .Y(_12516_));
 OAI21x1_ASAP7_75t_R _20874_ (.A1(_12163_),
    .A2(_12164_),
    .B(_12363_),
    .Y(_12517_));
 INVx1_ASAP7_75t_R _20875_ (.A(_12517_),
    .Y(_12518_));
 NOR2x1_ASAP7_75t_R _20876_ (.A(_12165_),
    .B(_12286_),
    .Y(_12519_));
 OAI21x1_ASAP7_75t_R _20877_ (.A1(_12518_),
    .A2(_12519_),
    .B(_12183_),
    .Y(_12520_));
 AOI21x1_ASAP7_75t_R _20878_ (.A1(_12520_),
    .A2(_12479_),
    .B(_12346_),
    .Y(_12521_));
 OAI21x1_ASAP7_75t_R _20879_ (.A1(_12361_),
    .A2(_12244_),
    .B(_12210_),
    .Y(_12522_));
 NOR2x1_ASAP7_75t_R _20880_ (.A(_12286_),
    .B(net10),
    .Y(_12523_));
 OAI21x1_ASAP7_75t_R _20881_ (.A1(_12234_),
    .A2(_12523_),
    .B(_12383_),
    .Y(_12524_));
 AOI21x1_ASAP7_75t_R _20882_ (.A1(_12522_),
    .A2(_12524_),
    .B(_12365_),
    .Y(_12525_));
 OAI21x1_ASAP7_75t_R _20883_ (.A1(_12521_),
    .A2(_12525_),
    .B(_12272_),
    .Y(_12526_));
 NAND2x1_ASAP7_75t_R _20884_ (.A(_12323_),
    .B(_12526_),
    .Y(_12527_));
 NAND2x1_ASAP7_75t_R _20885_ (.A(_12216_),
    .B(_12207_),
    .Y(_12528_));
 NOR2x1_ASAP7_75t_R _20886_ (.A(_12528_),
    .B(_12453_),
    .Y(_12529_));
 NAND2x1_ASAP7_75t_R _20887_ (.A(_12517_),
    .B(_12182_),
    .Y(_12530_));
 OAI21x1_ASAP7_75t_R _20888_ (.A1(_12315_),
    .A2(_12530_),
    .B(_12293_),
    .Y(_12531_));
 OAI21x1_ASAP7_75t_R _20889_ (.A1(_12529_),
    .A2(_12531_),
    .B(_12450_),
    .Y(_12532_));
 INVx2_ASAP7_75t_R _20890_ (.A(_12335_),
    .Y(_12533_));
 AO21x1_ASAP7_75t_R _20891_ (.A1(_12533_),
    .A2(_12328_),
    .B(_12183_),
    .Y(_12534_));
 AO21x1_ASAP7_75t_R _20892_ (.A1(_12233_),
    .A2(_12232_),
    .B(_01169_),
    .Y(_12535_));
 AO21x1_ASAP7_75t_R _20893_ (.A1(_12462_),
    .A2(_12535_),
    .B(_12463_),
    .Y(_12536_));
 AOI21x1_ASAP7_75t_R _20894_ (.A1(_12534_),
    .A2(_12536_),
    .B(_12311_),
    .Y(_12537_));
 AOI21x1_ASAP7_75t_R _20895_ (.A1(_12517_),
    .A2(_12377_),
    .B(_12235_),
    .Y(_12538_));
 OAI21x1_ASAP7_75t_R _20896_ (.A1(_12168_),
    .A2(_12511_),
    .B(_12538_),
    .Y(_12539_));
 OAI21x1_ASAP7_75t_R _20897_ (.A1(_12377_),
    .A2(net10),
    .B(_12307_),
    .Y(_12540_));
 AOI21x1_ASAP7_75t_R _20898_ (.A1(_12165_),
    .A2(_15848_),
    .B(_12194_),
    .Y(_12541_));
 OAI21x1_ASAP7_75t_R _20899_ (.A1(_12463_),
    .A2(_12216_),
    .B(_12271_),
    .Y(_12542_));
 AOI21x1_ASAP7_75t_R _20900_ (.A1(_12540_),
    .A2(_12541_),
    .B(_12542_),
    .Y(_12543_));
 NAND2x1_ASAP7_75t_R _20901_ (.A(_12539_),
    .B(_12543_),
    .Y(_12544_));
 OAI21x1_ASAP7_75t_R _20902_ (.A1(_12532_),
    .A2(_12537_),
    .B(_12544_),
    .Y(_12545_));
 AOI21x1_ASAP7_75t_R _20903_ (.A1(_12226_),
    .A2(_12545_),
    .B(_12284_),
    .Y(_12546_));
 OAI21x1_ASAP7_75t_R _20904_ (.A1(_12516_),
    .A2(_12527_),
    .B(_12546_),
    .Y(_12547_));
 NAND2x1_ASAP7_75t_R _20905_ (.A(_12547_),
    .B(_12509_),
    .Y(_00050_));
 NAND2x2_ASAP7_75t_R _20906_ (.A(_12473_),
    .B(_12290_),
    .Y(_12548_));
 OAI21x1_ASAP7_75t_R _20907_ (.A1(_12384_),
    .A2(_12548_),
    .B(_12531_),
    .Y(_12549_));
 NOR2x1_ASAP7_75t_R _20908_ (.A(_12384_),
    .B(_12458_),
    .Y(_12550_));
 NOR2x1_ASAP7_75t_R _20909_ (.A(_12549_),
    .B(_12550_),
    .Y(_12551_));
 OAI21x1_ASAP7_75t_R _20910_ (.A1(_12304_),
    .A2(_12551_),
    .B(_12226_),
    .Y(_12552_));
 INVx1_ASAP7_75t_R _20911_ (.A(_12343_),
    .Y(_12553_));
 INVx1_ASAP7_75t_R _20912_ (.A(_12373_),
    .Y(_12554_));
 BUFx6f_ASAP7_75t_R _20913_ (.A(_12182_),
    .Y(_12555_));
 AOI21x1_ASAP7_75t_R _20914_ (.A1(_12216_),
    .A2(_12382_),
    .B(_12555_),
    .Y(_12556_));
 AO21x1_ASAP7_75t_R _20915_ (.A1(_12553_),
    .A2(_12554_),
    .B(_12556_),
    .Y(_12557_));
 AO21x1_ASAP7_75t_R _20916_ (.A1(_12352_),
    .A2(_12330_),
    .B(_12309_),
    .Y(_12558_));
 AOI21x1_ASAP7_75t_R _20917_ (.A1(_12558_),
    .A2(_12425_),
    .B(_12369_),
    .Y(_12559_));
 OA21x2_ASAP7_75t_R _20918_ (.A1(_12321_),
    .A2(_12557_),
    .B(_12559_),
    .Y(_12560_));
 OA21x2_ASAP7_75t_R _20919_ (.A1(_12229_),
    .A2(_12216_),
    .B(_12235_),
    .Y(_12561_));
 NAND2x1_ASAP7_75t_R _20920_ (.A(_12561_),
    .B(_12536_),
    .Y(_12562_));
 NOR2x2_ASAP7_75t_R _20921_ (.A(_12296_),
    .B(_12212_),
    .Y(_12563_));
 INVx1_ASAP7_75t_R _20922_ (.A(_12563_),
    .Y(_12564_));
 INVx1_ASAP7_75t_R _20923_ (.A(_12297_),
    .Y(_12565_));
 AOI21x1_ASAP7_75t_R _20924_ (.A1(_12564_),
    .A2(_12565_),
    .B(_12426_),
    .Y(_12566_));
 AOI21x1_ASAP7_75t_R _20925_ (.A1(_12562_),
    .A2(_12566_),
    .B(_12225_),
    .Y(_12567_));
 OAI21x1_ASAP7_75t_R _20926_ (.A1(net560),
    .A2(_12250_),
    .B(_12309_),
    .Y(_12568_));
 NAND2x1_ASAP7_75t_R _20927_ (.A(_12473_),
    .B(_12374_),
    .Y(_12569_));
 AOI21x1_ASAP7_75t_R _20928_ (.A1(_12568_),
    .A2(_12569_),
    .B(_12365_),
    .Y(_12570_));
 AO21x1_ASAP7_75t_R _20929_ (.A1(_12444_),
    .A2(_12533_),
    .B(_12555_),
    .Y(_12571_));
 NAND2x1_ASAP7_75t_R _20930_ (.A(_12478_),
    .B(_12299_),
    .Y(_12572_));
 AOI21x1_ASAP7_75t_R _20931_ (.A1(_12571_),
    .A2(_12572_),
    .B(_12494_),
    .Y(_12573_));
 OAI21x1_ASAP7_75t_R _20932_ (.A1(_12570_),
    .A2(_12573_),
    .B(_12272_),
    .Y(_12574_));
 AOI21x1_ASAP7_75t_R _20933_ (.A1(_12567_),
    .A2(_12574_),
    .B(_12284_),
    .Y(_12575_));
 OAI21x1_ASAP7_75t_R _20934_ (.A1(_12552_),
    .A2(_12560_),
    .B(_12575_),
    .Y(_12576_));
 NOR2x2_ASAP7_75t_R _20935_ (.A(_12347_),
    .B(_12250_),
    .Y(_12577_));
 NOR2x1_ASAP7_75t_R _20936_ (.A(_12555_),
    .B(_12453_),
    .Y(_12578_));
 NAND2x1_ASAP7_75t_R _20937_ (.A(_12577_),
    .B(_12578_),
    .Y(_12579_));
 NAND2x2_ASAP7_75t_R _20938_ (.A(_15845_),
    .B(_12201_),
    .Y(_12580_));
 AOI21x1_ASAP7_75t_R _20939_ (.A1(_12405_),
    .A2(_12580_),
    .B(_12384_),
    .Y(_12581_));
 OA21x2_ASAP7_75t_R _20940_ (.A1(_12343_),
    .A2(_12314_),
    .B(_12195_),
    .Y(_12582_));
 AOI21x1_ASAP7_75t_R _20941_ (.A1(_12462_),
    .A2(_12424_),
    .B(_12183_),
    .Y(_12583_));
 INVx1_ASAP7_75t_R _20942_ (.A(_12583_),
    .Y(_12584_));
 AOI22x1_ASAP7_75t_R _20943_ (.A1(_12579_),
    .A2(_12581_),
    .B1(_12582_),
    .B2(_12584_),
    .Y(_12585_));
 INVx2_ASAP7_75t_R _20944_ (.A(_12510_),
    .Y(_12586_));
 OAI21x1_ASAP7_75t_R _20945_ (.A1(net922),
    .A2(_12586_),
    .B(_12399_),
    .Y(_12587_));
 NAND2x1_ASAP7_75t_R _20946_ (.A(_15845_),
    .B(_12331_),
    .Y(_12588_));
 OAI21x1_ASAP7_75t_R _20947_ (.A1(_15835_),
    .A2(_12307_),
    .B(_12235_),
    .Y(_12589_));
 NOR2x1_ASAP7_75t_R _20948_ (.A(_15840_),
    .B(_12103_),
    .Y(_12590_));
 NOR2x2_ASAP7_75t_R _20949_ (.A(_12589_),
    .B(_12590_),
    .Y(_12591_));
 AOI21x1_ASAP7_75t_R _20950_ (.A1(_12588_),
    .A2(_12591_),
    .B(_12303_),
    .Y(_12592_));
 AOI21x1_ASAP7_75t_R _20951_ (.A1(_12587_),
    .A2(_12592_),
    .B(_12237_),
    .Y(_12593_));
 OAI21x1_ASAP7_75t_R _20952_ (.A1(_12272_),
    .A2(_12585_),
    .B(_12593_),
    .Y(_12594_));
 AOI22x1_ASAP7_75t_R _20953_ (.A1(_12577_),
    .A2(_12230_),
    .B1(_12330_),
    .B2(_12336_),
    .Y(_12595_));
 AO21x1_ASAP7_75t_R _20954_ (.A1(_12432_),
    .A2(_12167_),
    .B(_12555_),
    .Y(_12596_));
 AOI21x1_ASAP7_75t_R _20955_ (.A1(_12510_),
    .A2(_12339_),
    .B(_12195_),
    .Y(_12597_));
 AOI21x1_ASAP7_75t_R _20956_ (.A1(_12596_),
    .A2(_12597_),
    .B(_12426_),
    .Y(_12598_));
 OAI21x1_ASAP7_75t_R _20957_ (.A1(_12321_),
    .A2(_12595_),
    .B(_12598_),
    .Y(_12599_));
 NAND2x1_ASAP7_75t_R _20958_ (.A(_12354_),
    .B(_12455_),
    .Y(_12600_));
 AOI21x1_ASAP7_75t_R _20959_ (.A1(_12339_),
    .A2(_12436_),
    .B(_12195_),
    .Y(_12601_));
 NAND2x1_ASAP7_75t_R _20960_ (.A(_12600_),
    .B(_12601_),
    .Y(_12602_));
 NOR2x1_ASAP7_75t_R _20961_ (.A(_12207_),
    .B(_12397_),
    .Y(_12603_));
 NAND2x1_ASAP7_75t_R _20962_ (.A(_12339_),
    .B(_12603_),
    .Y(_12604_));
 AOI21x1_ASAP7_75t_R _20963_ (.A1(_12337_),
    .A2(_12604_),
    .B(_12450_),
    .Y(_12605_));
 AOI21x1_ASAP7_75t_R _20964_ (.A1(_12602_),
    .A2(_12605_),
    .B(_12225_),
    .Y(_12606_));
 AOI21x1_ASAP7_75t_R _20965_ (.A1(_12599_),
    .A2(_12606_),
    .B(_12391_),
    .Y(_12607_));
 NAND2x1_ASAP7_75t_R _20966_ (.A(_12594_),
    .B(_12607_),
    .Y(_12608_));
 NAND2x1_ASAP7_75t_R _20967_ (.A(_12576_),
    .B(_12608_),
    .Y(_00051_));
 NAND2x1_ASAP7_75t_R _20968_ (.A(_12555_),
    .B(_12412_),
    .Y(_12609_));
 OAI21x1_ASAP7_75t_R _20969_ (.A1(_12335_),
    .A2(_12609_),
    .B(_12346_),
    .Y(_12610_));
 NOR2x1_ASAP7_75t_R _20970_ (.A(_12291_),
    .B(_12288_),
    .Y(_12611_));
 NOR2x1_ASAP7_75t_R _20971_ (.A(_12610_),
    .B(_12611_),
    .Y(_12612_));
 OA21x2_ASAP7_75t_R _20972_ (.A1(_12318_),
    .A2(_12183_),
    .B(_12216_),
    .Y(_12613_));
 AO21x1_ASAP7_75t_R _20973_ (.A1(_12613_),
    .A2(_12208_),
    .B(_12369_),
    .Y(_12614_));
 OAI21x1_ASAP7_75t_R _20974_ (.A1(_12612_),
    .A2(_12614_),
    .B(_12323_),
    .Y(_12615_));
 AOI21x1_ASAP7_75t_R _20975_ (.A1(_15848_),
    .A2(_15838_),
    .B(_12249_),
    .Y(_12616_));
 OAI21x1_ASAP7_75t_R _20976_ (.A1(_12230_),
    .A2(_12616_),
    .B(_12494_),
    .Y(_12617_));
 OAI21x1_ASAP7_75t_R _20977_ (.A1(_12617_),
    .A2(_12247_),
    .B(_12369_),
    .Y(_12618_));
 NOR2x1_ASAP7_75t_R _20978_ (.A(_12230_),
    .B(_12288_),
    .Y(_12619_));
 NAND2x1_ASAP7_75t_R _20979_ (.A(_12365_),
    .B(_12520_),
    .Y(_12620_));
 AOI21x1_ASAP7_75t_R _20980_ (.A1(_12339_),
    .A2(_12619_),
    .B(_12620_),
    .Y(_12621_));
 NOR2x1_ASAP7_75t_R _20981_ (.A(_12618_),
    .B(_12621_),
    .Y(_12622_));
 OAI21x1_ASAP7_75t_R _20982_ (.A1(_12615_),
    .A2(_12622_),
    .B(_12284_),
    .Y(_12623_));
 NAND2x1_ASAP7_75t_R _20983_ (.A(_12384_),
    .B(_12426_),
    .Y(_12624_));
 AOI21x1_ASAP7_75t_R _20984_ (.A1(_12201_),
    .A2(_12362_),
    .B(_12624_),
    .Y(_12625_));
 AO21x1_ASAP7_75t_R _20985_ (.A1(_12478_),
    .A2(_12326_),
    .B(_12230_),
    .Y(_12626_));
 AOI22x1_ASAP7_75t_R _20986_ (.A1(_12625_),
    .A2(_12626_),
    .B1(_12456_),
    .B2(_12497_),
    .Y(_12627_));
 AND3x1_ASAP7_75t_R _20987_ (.A(_12291_),
    .B(_12365_),
    .C(_12444_),
    .Y(_12628_));
 AOI21x1_ASAP7_75t_R _20988_ (.A1(_12462_),
    .A2(_12339_),
    .B(_12183_),
    .Y(_12629_));
 NOR2x1_ASAP7_75t_R _20989_ (.A(_00513_),
    .B(_15845_),
    .Y(_12630_));
 OAI21x1_ASAP7_75t_R _20990_ (.A1(_12630_),
    .A2(_12379_),
    .B(_12494_),
    .Y(_12631_));
 NOR2x1_ASAP7_75t_R _20991_ (.A(_12629_),
    .B(_12631_),
    .Y(_12632_));
 OAI21x1_ASAP7_75t_R _20992_ (.A1(_12628_),
    .A2(_12632_),
    .B(_12304_),
    .Y(_12633_));
 AOI21x1_ASAP7_75t_R _20993_ (.A1(_12627_),
    .A2(_12633_),
    .B(_12323_),
    .Y(_12634_));
 AOI21x1_ASAP7_75t_R _20994_ (.A1(_12201_),
    .A2(_12243_),
    .B(_12246_),
    .Y(_12635_));
 NOR2x1_ASAP7_75t_R _20995_ (.A(net922),
    .B(_12511_),
    .Y(_12636_));
 OAI21x1_ASAP7_75t_R _20996_ (.A1(_12635_),
    .A2(_12636_),
    .B(_12311_),
    .Y(_12637_));
 OAI21x1_ASAP7_75t_R _20997_ (.A1(_12310_),
    .A2(_12583_),
    .B(_12321_),
    .Y(_12638_));
 AOI21x1_ASAP7_75t_R _20998_ (.A1(_12637_),
    .A2(_12638_),
    .B(_12304_),
    .Y(_12639_));
 NAND2x1_ASAP7_75t_R _20999_ (.A(_00517_),
    .B(_12309_),
    .Y(_12640_));
 OAI21x1_ASAP7_75t_R _21000_ (.A1(_12234_),
    .A2(_12230_),
    .B(_12640_),
    .Y(_12641_));
 OAI21x1_ASAP7_75t_R _21001_ (.A1(_12311_),
    .A2(_12641_),
    .B(_12304_),
    .Y(_12642_));
 AO21x1_ASAP7_75t_R _21002_ (.A1(_12290_),
    .A2(_12243_),
    .B(_12320_),
    .Y(_12643_));
 AND3x1_ASAP7_75t_R _21003_ (.A(_12354_),
    .B(_15845_),
    .C(_12309_),
    .Y(_12644_));
 NOR2x1_ASAP7_75t_R _21004_ (.A(_12643_),
    .B(_12644_),
    .Y(_12645_));
 OAI21x1_ASAP7_75t_R _21005_ (.A1(_12642_),
    .A2(_12645_),
    .B(_12323_),
    .Y(_12646_));
 OAI21x1_ASAP7_75t_R _21006_ (.A1(_12639_),
    .A2(_12646_),
    .B(_12391_),
    .Y(_12647_));
 OAI21x1_ASAP7_75t_R _21007_ (.A1(_12166_),
    .A2(_15848_),
    .B(_12183_),
    .Y(_12648_));
 OAI21x1_ASAP7_75t_R _21008_ (.A1(net577),
    .A2(_12648_),
    .B(_12346_),
    .Y(_12649_));
 NOR2x1_ASAP7_75t_R _21009_ (.A(_12649_),
    .B(_12205_),
    .Y(_12650_));
 NAND2x1_ASAP7_75t_R _21010_ (.A(_01167_),
    .B(_15848_),
    .Y(_12651_));
 AOI21x1_ASAP7_75t_R _21011_ (.A1(_12383_),
    .A2(_12651_),
    .B(_12320_),
    .Y(_12652_));
 AO21x1_ASAP7_75t_R _21012_ (.A1(_12393_),
    .A2(_12652_),
    .B(_12369_),
    .Y(_12653_));
 OAI21x1_ASAP7_75t_R _21013_ (.A1(_12650_),
    .A2(_12653_),
    .B(_12226_),
    .Y(_12654_));
 AO21x1_ASAP7_75t_R _21014_ (.A1(_12306_),
    .A2(_12339_),
    .B(_12487_),
    .Y(_12655_));
 AO21x1_ASAP7_75t_R _21015_ (.A1(_12453_),
    .A2(_12383_),
    .B(_12320_),
    .Y(_12656_));
 NOR2x1_ASAP7_75t_R _21016_ (.A(_12195_),
    .B(_12422_),
    .Y(_12657_));
 AO21x1_ASAP7_75t_R _21017_ (.A1(_12378_),
    .A2(_12517_),
    .B(_12348_),
    .Y(_12658_));
 AOI21x1_ASAP7_75t_R _21018_ (.A1(_12657_),
    .A2(_12658_),
    .B(_12450_),
    .Y(_12659_));
 OA21x2_ASAP7_75t_R _21019_ (.A1(_12655_),
    .A2(_12656_),
    .B(_12659_),
    .Y(_12660_));
 NOR2x1_ASAP7_75t_R _21020_ (.A(_12654_),
    .B(_12660_),
    .Y(_12661_));
 OAI22x1_ASAP7_75t_R _21021_ (.A1(_12623_),
    .A2(_12634_),
    .B1(_12647_),
    .B2(_12661_),
    .Y(_00052_));
 AO21x1_ASAP7_75t_R _21022_ (.A1(_12210_),
    .A2(_15840_),
    .B(_12384_),
    .Y(_12662_));
 OAI21x1_ASAP7_75t_R _21023_ (.A1(_12662_),
    .A2(_12355_),
    .B(_12304_),
    .Y(_12663_));
 OAI21x1_ASAP7_75t_R _21024_ (.A1(_12215_),
    .A2(_12152_),
    .B(_12181_),
    .Y(_12664_));
 OAI21x1_ASAP7_75t_R _21025_ (.A1(_12361_),
    .A2(_12664_),
    .B(_12311_),
    .Y(_12665_));
 AOI21x1_ASAP7_75t_R _21026_ (.A1(_12436_),
    .A2(_12360_),
    .B(_12665_),
    .Y(_12666_));
 OAI21x1_ASAP7_75t_R _21027_ (.A1(_12663_),
    .A2(_12666_),
    .B(_12226_),
    .Y(_12667_));
 AOI21x1_ASAP7_75t_R _21028_ (.A1(net53),
    .A2(_15848_),
    .B(_12383_),
    .Y(_12668_));
 NOR2x2_ASAP7_75t_R _21029_ (.A(_12463_),
    .B(_12462_),
    .Y(_12669_));
 AOI211x1_ASAP7_75t_R _21030_ (.A1(_12438_),
    .A2(_12668_),
    .B(_12669_),
    .C(_12196_),
    .Y(_12670_));
 AO21x1_ASAP7_75t_R _21031_ (.A1(_12314_),
    .A2(_12210_),
    .B(_12320_),
    .Y(_12671_));
 AOI21x1_ASAP7_75t_R _21032_ (.A1(_12517_),
    .A2(_12580_),
    .B(_12246_),
    .Y(_12672_));
 OAI21x1_ASAP7_75t_R _21033_ (.A1(_12671_),
    .A2(_12672_),
    .B(_12272_),
    .Y(_12673_));
 NOR2x1_ASAP7_75t_R _21034_ (.A(_12670_),
    .B(_12673_),
    .Y(_12674_));
 OAI21x1_ASAP7_75t_R _21035_ (.A1(_12667_),
    .A2(_12674_),
    .B(_12391_),
    .Y(_12675_));
 NAND2x1_ASAP7_75t_R _21036_ (.A(_12555_),
    .B(net10),
    .Y(_12676_));
 AND3x1_ASAP7_75t_R _21037_ (.A(_12474_),
    .B(_12346_),
    .C(_12676_),
    .Y(_12677_));
 AO21x1_ASAP7_75t_R _21038_ (.A1(_12208_),
    .A2(_12375_),
    .B(_12426_),
    .Y(_12678_));
 AOI21x1_ASAP7_75t_R _21039_ (.A1(_12440_),
    .A2(_12677_),
    .B(_12678_),
    .Y(_12679_));
 AO21x1_ASAP7_75t_R _21040_ (.A1(_12210_),
    .A2(_00511_),
    .B(_12195_),
    .Y(_12680_));
 OA21x2_ASAP7_75t_R _21041_ (.A1(_12462_),
    .A2(net10),
    .B(_12383_),
    .Y(_12681_));
 OAI21x1_ASAP7_75t_R _21042_ (.A1(_12680_),
    .A2(_12681_),
    .B(_12369_),
    .Y(_12682_));
 AO21x1_ASAP7_75t_R _21043_ (.A1(_12233_),
    .A2(_12232_),
    .B(_00511_),
    .Y(_12683_));
 AO21x1_ASAP7_75t_R _21044_ (.A1(_12554_),
    .A2(_12510_),
    .B(_12320_),
    .Y(_12684_));
 AOI21x1_ASAP7_75t_R _21045_ (.A1(_12683_),
    .A2(_12436_),
    .B(_12684_),
    .Y(_12685_));
 OAI21x1_ASAP7_75t_R _21046_ (.A1(_12682_),
    .A2(_12685_),
    .B(_12323_),
    .Y(_12686_));
 NOR2x1_ASAP7_75t_R _21047_ (.A(_12679_),
    .B(_12686_),
    .Y(_12687_));
 NAND2x1_ASAP7_75t_R _21048_ (.A(_12326_),
    .B(_12436_),
    .Y(_12688_));
 AOI21x1_ASAP7_75t_R _21049_ (.A1(_12530_),
    .A2(_12688_),
    .B(_12311_),
    .Y(_12689_));
 AO21x1_ASAP7_75t_R _21050_ (.A1(_12210_),
    .A2(net577),
    .B(_12320_),
    .Y(_12690_));
 OA21x2_ASAP7_75t_R _21051_ (.A1(_12361_),
    .A2(_12252_),
    .B(_12383_),
    .Y(_12691_));
 OAI21x1_ASAP7_75t_R _21052_ (.A1(_12690_),
    .A2(_12691_),
    .B(_12272_),
    .Y(_12692_));
 OAI21x1_ASAP7_75t_R _21053_ (.A1(_12689_),
    .A2(_12692_),
    .B(_12323_),
    .Y(_12693_));
 AO21x1_ASAP7_75t_R _21054_ (.A1(_15838_),
    .A2(_12210_),
    .B(_12195_),
    .Y(_12694_));
 NAND2x1_ASAP7_75t_R _21055_ (.A(_12555_),
    .B(_12243_),
    .Y(_12695_));
 NOR2x1_ASAP7_75t_R _21056_ (.A(_12202_),
    .B(_12695_),
    .Y(_12696_));
 OAI21x1_ASAP7_75t_R _21057_ (.A1(_12694_),
    .A2(_12696_),
    .B(_12450_),
    .Y(_12697_));
 NAND2x1_ASAP7_75t_R _21058_ (.A(_12201_),
    .B(_12439_),
    .Y(_12698_));
 AOI21x1_ASAP7_75t_R _21059_ (.A1(_12307_),
    .A2(net10),
    .B(_12229_),
    .Y(_12699_));
 NAND3x1_ASAP7_75t_R _21060_ (.A(_12699_),
    .B(_12313_),
    .C(_12378_),
    .Y(_12700_));
 AOI21x1_ASAP7_75t_R _21061_ (.A1(_12698_),
    .A2(_12700_),
    .B(_12494_),
    .Y(_12701_));
 NOR2x1_ASAP7_75t_R _21062_ (.A(_12697_),
    .B(_12701_),
    .Y(_12702_));
 NOR2x1_ASAP7_75t_R _21063_ (.A(_12693_),
    .B(_12702_),
    .Y(_12703_));
 AO21x1_ASAP7_75t_R _21064_ (.A1(_12212_),
    .A2(_12383_),
    .B(_12384_),
    .Y(_12704_));
 OAI21x1_ASAP7_75t_R _21065_ (.A1(_12556_),
    .A2(_12704_),
    .B(_12272_),
    .Y(_12705_));
 INVx1_ASAP7_75t_R _21066_ (.A(_12648_),
    .Y(_12706_));
 AOI211x1_ASAP7_75t_R _21067_ (.A1(_12422_),
    .A2(_12354_),
    .B(_12706_),
    .C(_12494_),
    .Y(_12707_));
 OAI21x1_ASAP7_75t_R _21068_ (.A1(_12705_),
    .A2(_12707_),
    .B(_12226_),
    .Y(_12708_));
 OA21x2_ASAP7_75t_R _21069_ (.A1(_12519_),
    .A2(_12518_),
    .B(_12210_),
    .Y(_12709_));
 OAI21x1_ASAP7_75t_R _21070_ (.A1(_12709_),
    .A2(_12368_),
    .B(_12450_),
    .Y(_12710_));
 AO21x1_ASAP7_75t_R _21071_ (.A1(_12151_),
    .A2(_12149_),
    .B(_12472_),
    .Y(_12711_));
 AOI21x1_ASAP7_75t_R _21072_ (.A1(_12167_),
    .A2(_12711_),
    .B(_12230_),
    .Y(_12712_));
 OAI21x1_ASAP7_75t_R _21073_ (.A1(_12664_),
    .A2(_12288_),
    .B(_12365_),
    .Y(_12713_));
 NOR2x1_ASAP7_75t_R _21074_ (.A(_12712_),
    .B(_12713_),
    .Y(_12714_));
 NOR2x1_ASAP7_75t_R _21075_ (.A(_12710_),
    .B(_12714_),
    .Y(_12715_));
 OAI21x1_ASAP7_75t_R _21076_ (.A1(_12708_),
    .A2(_12715_),
    .B(_12284_),
    .Y(_12716_));
 OAI22x1_ASAP7_75t_R _21077_ (.A1(_12675_),
    .A2(_12687_),
    .B1(_12703_),
    .B2(_12716_),
    .Y(_00053_));
 NAND2x2_ASAP7_75t_R _21078_ (.A(_12243_),
    .B(_12290_),
    .Y(_12717_));
 AOI21x1_ASAP7_75t_R _21079_ (.A1(_12300_),
    .A2(_12717_),
    .B(_12346_),
    .Y(_12718_));
 AOI21x1_ASAP7_75t_R _21080_ (.A1(_12246_),
    .A2(_12411_),
    .B(_12365_),
    .Y(_12719_));
 OAI21x1_ASAP7_75t_R _21081_ (.A1(_12718_),
    .A2(_12719_),
    .B(_12369_),
    .Y(_12720_));
 OA21x2_ASAP7_75t_R _21082_ (.A1(_12352_),
    .A2(_12463_),
    .B(_12293_),
    .Y(_12721_));
 OAI21x1_ASAP7_75t_R _21083_ (.A1(_12327_),
    .A2(_12375_),
    .B(_12721_),
    .Y(_12722_));
 AOI21x1_ASAP7_75t_R _21084_ (.A1(_00518_),
    .A2(_12348_),
    .B(_12195_),
    .Y(_12723_));
 INVx1_ASAP7_75t_R _21085_ (.A(_12535_),
    .Y(_12724_));
 OAI21x1_ASAP7_75t_R _21086_ (.A1(_12724_),
    .A2(_12523_),
    .B(_12309_),
    .Y(_12725_));
 AOI21x1_ASAP7_75t_R _21087_ (.A1(_12723_),
    .A2(_12725_),
    .B(_12426_),
    .Y(_12726_));
 NAND2x1_ASAP7_75t_R _21088_ (.A(_12722_),
    .B(_12726_),
    .Y(_12727_));
 AOI21x1_ASAP7_75t_R _21089_ (.A1(_12720_),
    .A2(_12727_),
    .B(_12226_),
    .Y(_12728_));
 NOR2x1_ASAP7_75t_R _21090_ (.A(_12463_),
    .B(_12364_),
    .Y(_12729_));
 OA21x2_ASAP7_75t_R _21091_ (.A1(_12729_),
    .A2(_12496_),
    .B(_12352_),
    .Y(_12730_));
 AOI21x1_ASAP7_75t_R _21092_ (.A1(_12676_),
    .A2(_12591_),
    .B(_12426_),
    .Y(_12731_));
 OAI21x1_ASAP7_75t_R _21093_ (.A1(_12321_),
    .A2(_12730_),
    .B(_12731_),
    .Y(_12732_));
 NAND2x1_ASAP7_75t_R _21094_ (.A(net53),
    .B(_12422_),
    .Y(_12733_));
 NAND2x1_ASAP7_75t_R _21095_ (.A(_12327_),
    .B(_12555_),
    .Y(_12734_));
 NAND3x1_ASAP7_75t_R _21096_ (.A(_12733_),
    .B(_12561_),
    .C(_12734_),
    .Y(_12735_));
 AOI21x1_ASAP7_75t_R _21097_ (.A1(_12348_),
    .A2(_12415_),
    .B(_12334_),
    .Y(_12736_));
 OAI21x1_ASAP7_75t_R _21098_ (.A1(_12307_),
    .A2(_15838_),
    .B(net53),
    .Y(_12737_));
 NAND2x1_ASAP7_75t_R _21099_ (.A(_12309_),
    .B(_12737_),
    .Y(_12738_));
 AOI21x1_ASAP7_75t_R _21100_ (.A1(_12736_),
    .A2(_12738_),
    .B(_12303_),
    .Y(_12739_));
 NAND2x1_ASAP7_75t_R _21101_ (.A(_12735_),
    .B(_12739_),
    .Y(_12740_));
 AOI21x1_ASAP7_75t_R _21102_ (.A1(_12732_),
    .A2(_12740_),
    .B(_12323_),
    .Y(_12741_));
 OAI21x1_ASAP7_75t_R _21103_ (.A1(_12728_),
    .A2(_12741_),
    .B(_12391_),
    .Y(_12742_));
 AND2x2_ASAP7_75t_R _21104_ (.A(_12296_),
    .B(_12216_),
    .Y(_12743_));
 AO21x1_ASAP7_75t_R _21105_ (.A1(_12233_),
    .A2(_12232_),
    .B(_12472_),
    .Y(_12744_));
 AOI211x1_ASAP7_75t_R _21106_ (.A1(_12743_),
    .A2(_12744_),
    .B(_12669_),
    .C(_12236_),
    .Y(_12745_));
 NOR2x2_ASAP7_75t_R _21107_ (.A(_12364_),
    .B(_12664_),
    .Y(_12746_));
 INVx1_ASAP7_75t_R _21108_ (.A(_12746_),
    .Y(_12747_));
 AOI21x1_ASAP7_75t_R _21109_ (.A1(_15840_),
    .A2(net865),
    .B(_12307_),
    .Y(_12748_));
 OAI21x1_ASAP7_75t_R _21110_ (.A1(_12292_),
    .A2(_12748_),
    .B(_12348_),
    .Y(_12749_));
 AOI21x1_ASAP7_75t_R _21111_ (.A1(_12747_),
    .A2(_12749_),
    .B(_12384_),
    .Y(_12750_));
 OAI21x1_ASAP7_75t_R _21112_ (.A1(_12745_),
    .A2(_12750_),
    .B(_12369_),
    .Y(_12751_));
 AO21x1_ASAP7_75t_R _21113_ (.A1(_12431_),
    .A2(_12216_),
    .B(_12377_),
    .Y(_12752_));
 NOR2x1_ASAP7_75t_R _21114_ (.A(_12334_),
    .B(_12487_),
    .Y(_12753_));
 AOI21x1_ASAP7_75t_R _21115_ (.A1(_12752_),
    .A2(_12753_),
    .B(_12426_),
    .Y(_12754_));
 OAI21x1_ASAP7_75t_R _21116_ (.A1(_12361_),
    .A2(_12202_),
    .B(_12331_),
    .Y(_12755_));
 AO21x1_ASAP7_75t_R _21117_ (.A1(_01173_),
    .A2(_01171_),
    .B(_12207_),
    .Y(_12756_));
 NAND3x1_ASAP7_75t_R _21118_ (.A(_12755_),
    .B(_12320_),
    .C(_12756_),
    .Y(_12757_));
 AOI21x1_ASAP7_75t_R _21119_ (.A1(_12754_),
    .A2(_12757_),
    .B(_12237_),
    .Y(_12758_));
 NAND2x1_ASAP7_75t_R _21120_ (.A(_12751_),
    .B(_12758_),
    .Y(_12759_));
 OA21x2_ASAP7_75t_R _21121_ (.A1(_12313_),
    .A2(_12463_),
    .B(_12293_),
    .Y(_12760_));
 AO21x1_ASAP7_75t_R _21122_ (.A1(_12462_),
    .A2(_15838_),
    .B(_12555_),
    .Y(_12761_));
 AOI21x1_ASAP7_75t_R _21123_ (.A1(_12760_),
    .A2(_12761_),
    .B(_12303_),
    .Y(_12762_));
 AOI21x1_ASAP7_75t_R _21124_ (.A1(_12352_),
    .A2(_12353_),
    .B(_12293_),
    .Y(_12763_));
 AOI21x1_ASAP7_75t_R _21125_ (.A1(_12533_),
    .A2(_12711_),
    .B(_12207_),
    .Y(_12764_));
 NOR3x1_ASAP7_75t_R _21126_ (.A(_12229_),
    .B(_15840_),
    .C(_12153_),
    .Y(_12765_));
 NOR2x1_ASAP7_75t_R _21127_ (.A(_12764_),
    .B(_12765_),
    .Y(_12766_));
 NAND2x1_ASAP7_75t_R _21128_ (.A(_12763_),
    .B(_12766_),
    .Y(_12767_));
 AOI21x1_ASAP7_75t_R _21129_ (.A1(_12762_),
    .A2(_12767_),
    .B(_12225_),
    .Y(_12768_));
 AOI21x1_ASAP7_75t_R _21130_ (.A1(_12483_),
    .A2(_12482_),
    .B(_12563_),
    .Y(_12769_));
 AOI21x1_ASAP7_75t_R _21131_ (.A1(_12510_),
    .A2(_12651_),
    .B(_12195_),
    .Y(_12770_));
 OAI21x1_ASAP7_75t_R _21132_ (.A1(_15845_),
    .A2(_12354_),
    .B(_12699_),
    .Y(_12771_));
 AOI21x1_ASAP7_75t_R _21133_ (.A1(_12770_),
    .A2(_12771_),
    .B(_12426_),
    .Y(_12772_));
 OAI21x1_ASAP7_75t_R _21134_ (.A1(_12321_),
    .A2(_12769_),
    .B(_12772_),
    .Y(_12773_));
 AOI21x1_ASAP7_75t_R _21135_ (.A1(_12768_),
    .A2(_12773_),
    .B(_12391_),
    .Y(_12774_));
 NAND2x1_ASAP7_75t_R _21136_ (.A(_12759_),
    .B(_12774_),
    .Y(_12775_));
 NAND2x1_ASAP7_75t_R _21137_ (.A(_12742_),
    .B(_12775_),
    .Y(_00054_));
 AO21x1_ASAP7_75t_R _21138_ (.A1(_12377_),
    .A2(net53),
    .B(_12334_),
    .Y(_12776_));
 OR2x2_ASAP7_75t_R _21139_ (.A(_12776_),
    .B(_12629_),
    .Y(_12777_));
 NOR2x1_ASAP7_75t_R _21140_ (.A(_12344_),
    .B(_12695_),
    .Y(_12778_));
 AND2x2_ASAP7_75t_R _21141_ (.A(_12496_),
    .B(_12478_),
    .Y(_12779_));
 OAI21x1_ASAP7_75t_R _21142_ (.A1(_12778_),
    .A2(_12779_),
    .B(_12321_),
    .Y(_12780_));
 AOI21x1_ASAP7_75t_R _21143_ (.A1(_12777_),
    .A2(_12780_),
    .B(_12272_),
    .Y(_12781_));
 AOI211x1_ASAP7_75t_R _21144_ (.A1(_12465_),
    .A2(_12246_),
    .B(_12563_),
    .C(_12311_),
    .Y(_12782_));
 NOR2x1_ASAP7_75t_R _21145_ (.A(_12586_),
    .B(_12344_),
    .Y(_12783_));
 OAI21x1_ASAP7_75t_R _21146_ (.A1(_12230_),
    .A2(_12288_),
    .B(_12311_),
    .Y(_12784_));
 OAI21x1_ASAP7_75t_R _21147_ (.A1(_12784_),
    .A2(_12783_),
    .B(_12272_),
    .Y(_12785_));
 OAI21x1_ASAP7_75t_R _21148_ (.A1(_12782_),
    .A2(_12785_),
    .B(_12323_),
    .Y(_12786_));
 OAI21x1_ASAP7_75t_R _21149_ (.A1(_12781_),
    .A2(_12786_),
    .B(_12391_),
    .Y(_12787_));
 NAND3x1_ASAP7_75t_R _21150_ (.A(_12717_),
    .B(_12321_),
    .C(_12609_),
    .Y(_12788_));
 OAI21x1_ASAP7_75t_R _21151_ (.A1(_12249_),
    .A2(_12748_),
    .B(_12246_),
    .Y(_12789_));
 AO21x1_ASAP7_75t_R _21152_ (.A1(net10),
    .A2(_15845_),
    .B(_15840_),
    .Y(_12790_));
 AOI21x1_ASAP7_75t_R _21153_ (.A1(_12230_),
    .A2(_12790_),
    .B(_12494_),
    .Y(_12791_));
 AOI21x1_ASAP7_75t_R _21154_ (.A1(_12789_),
    .A2(_12791_),
    .B(_12272_),
    .Y(_12792_));
 OAI21x1_ASAP7_75t_R _21155_ (.A1(_12746_),
    .A2(_12504_),
    .B(_12321_),
    .Y(_12793_));
 NAND2x1_ASAP7_75t_R _21156_ (.A(_12412_),
    .B(_12336_),
    .Y(_12794_));
 AO21x1_ASAP7_75t_R _21157_ (.A1(_12794_),
    .A2(_12568_),
    .B(_12494_),
    .Y(_12795_));
 AOI21x1_ASAP7_75t_R _21158_ (.A1(_12793_),
    .A2(_12795_),
    .B(_12304_),
    .Y(_12796_));
 AOI211x1_ASAP7_75t_R _21159_ (.A1(_12788_),
    .A2(_12792_),
    .B(_12796_),
    .C(_12323_),
    .Y(_12797_));
 AO21x1_ASAP7_75t_R _21160_ (.A1(_12462_),
    .A2(_15838_),
    .B(_12348_),
    .Y(_12798_));
 NAND2x1_ASAP7_75t_R _21161_ (.A(_00517_),
    .B(_12463_),
    .Y(_12799_));
 AO21x1_ASAP7_75t_R _21162_ (.A1(_12253_),
    .A2(_12799_),
    .B(_12271_),
    .Y(_12800_));
 AO21x1_ASAP7_75t_R _21163_ (.A1(_12454_),
    .A2(_12798_),
    .B(_12800_),
    .Y(_12801_));
 NAND2x1_ASAP7_75t_R _21164_ (.A(_12555_),
    .B(_12382_),
    .Y(_12802_));
 AOI21x1_ASAP7_75t_R _21165_ (.A1(_12336_),
    .A2(_12328_),
    .B(_12320_),
    .Y(_12803_));
 OAI21x1_ASAP7_75t_R _21166_ (.A1(_12361_),
    .A2(_12802_),
    .B(_12803_),
    .Y(_12804_));
 NAND2x1_ASAP7_75t_R _21167_ (.A(_12335_),
    .B(_12383_),
    .Y(_12805_));
 OAI21x1_ASAP7_75t_R _21168_ (.A1(_01173_),
    .A2(_12377_),
    .B(_12334_),
    .Y(_12806_));
 NOR2x1_ASAP7_75t_R _21169_ (.A(_12217_),
    .B(_12806_),
    .Y(_12807_));
 AOI21x1_ASAP7_75t_R _21170_ (.A1(_12805_),
    .A2(_12807_),
    .B(_12450_),
    .Y(_12808_));
 AOI21x1_ASAP7_75t_R _21171_ (.A1(_12808_),
    .A2(_12804_),
    .B(_12226_),
    .Y(_12809_));
 AOI21x1_ASAP7_75t_R _21172_ (.A1(_12801_),
    .A2(_12809_),
    .B(_12391_),
    .Y(_12810_));
 AO21x1_ASAP7_75t_R _21173_ (.A1(_12382_),
    .A2(_15838_),
    .B(_12331_),
    .Y(_12811_));
 AND3x1_ASAP7_75t_R _21174_ (.A(_12811_),
    .B(_12311_),
    .C(_12548_),
    .Y(_12812_));
 OAI21x1_ASAP7_75t_R _21175_ (.A1(_12307_),
    .A2(_15838_),
    .B(_12330_),
    .Y(_12813_));
 INVx1_ASAP7_75t_R _21176_ (.A(_12683_),
    .Y(_12814_));
 OAI21x1_ASAP7_75t_R _21177_ (.A1(net560),
    .A2(_12814_),
    .B(_12348_),
    .Y(_12815_));
 OAI21x1_ASAP7_75t_R _21178_ (.A1(_12802_),
    .A2(_12813_),
    .B(_12815_),
    .Y(_12816_));
 AO21x1_ASAP7_75t_R _21179_ (.A1(_12816_),
    .A2(_12494_),
    .B(_12369_),
    .Y(_12817_));
 OA21x2_ASAP7_75t_R _21180_ (.A1(_12331_),
    .A2(_12165_),
    .B(_12293_),
    .Y(_12818_));
 AOI21x1_ASAP7_75t_R _21181_ (.A1(_12818_),
    .A2(_12755_),
    .B(_12450_),
    .Y(_12819_));
 NAND2x1_ASAP7_75t_R _21182_ (.A(_12348_),
    .B(_12813_),
    .Y(_12820_));
 INVx1_ASAP7_75t_R _21183_ (.A(_12253_),
    .Y(_12821_));
 NOR2x1_ASAP7_75t_R _21184_ (.A(_12487_),
    .B(_12821_),
    .Y(_12822_));
 NAND2x1_ASAP7_75t_R _21185_ (.A(_12820_),
    .B(_12822_),
    .Y(_12823_));
 AOI21x1_ASAP7_75t_R _21186_ (.A1(_12819_),
    .A2(_12823_),
    .B(_12237_),
    .Y(_12824_));
 OAI21x1_ASAP7_75t_R _21187_ (.A1(_12812_),
    .A2(_12817_),
    .B(_12824_),
    .Y(_12825_));
 NAND2x1_ASAP7_75t_R _21188_ (.A(_12825_),
    .B(_12810_),
    .Y(_12826_));
 OAI21x1_ASAP7_75t_R _21189_ (.A1(_12787_),
    .A2(_12797_),
    .B(_12826_),
    .Y(_00055_));
 AND2x2_ASAP7_75t_R _21190_ (.A(_10640_),
    .B(_00519_),
    .Y(_12827_));
 BUFx2_ASAP7_75t_R rebuffer204 (.A(_00756_),
    .Y(net657));
 BUFx6f_ASAP7_75t_R _21192_ (.A(_00763_),
    .Y(_12829_));
 XOR2x2_ASAP7_75t_R _21193_ (.A(_00756_),
    .B(_12829_),
    .Y(_12830_));
 BUFx6f_ASAP7_75t_R _21194_ (.A(_00821_),
    .Y(_12831_));
 XOR2x2_ASAP7_75t_R _21195_ (.A(_00789_),
    .B(_12831_),
    .Y(_12832_));
 XOR2x2_ASAP7_75t_R _21196_ (.A(_12832_),
    .B(_12830_),
    .Y(_12833_));
 BUFx6f_ASAP7_75t_R _21197_ (.A(_00788_),
    .Y(_12834_));
 XOR2x2_ASAP7_75t_R _21198_ (.A(_00795_),
    .B(_12834_),
    .Y(_12835_));
 BUFx6f_ASAP7_75t_R _21199_ (.A(_00853_),
    .Y(_12836_));
 INVx2_ASAP7_75t_R _21200_ (.A(_12836_),
    .Y(_12837_));
 XOR2x2_ASAP7_75t_R _21201_ (.A(_12837_),
    .B(_12835_),
    .Y(_12838_));
 XOR2x1_ASAP7_75t_R _21202_ (.A(_12838_),
    .Y(_12839_),
    .B(_12833_));
 NOR2x1_ASAP7_75t_R _21203_ (.A(_12095_),
    .B(_12839_),
    .Y(_12840_));
 INVx2_ASAP7_75t_R _21204_ (.A(_08191_),
    .Y(_12841_));
 OAI21x1_ASAP7_75t_R _21205_ (.A1(_12840_),
    .A2(_12827_),
    .B(_12841_),
    .Y(_12842_));
 NOR2x2_ASAP7_75t_R _21206_ (.A(_11356_),
    .B(_00519_),
    .Y(_12843_));
 XNOR2x1_ASAP7_75t_R _21207_ (.B(_12838_),
    .Y(_12844_),
    .A(_12833_));
 NOR2x1_ASAP7_75t_R _21208_ (.A(_12095_),
    .B(_12844_),
    .Y(_12845_));
 OAI21x1_ASAP7_75t_R _21209_ (.A1(_12843_),
    .A2(_12845_),
    .B(_08191_),
    .Y(_12846_));
 NAND2x2_ASAP7_75t_R _21210_ (.A(_12846_),
    .B(_12842_),
    .Y(_12847_));
 BUFx12f_ASAP7_75t_R _21211_ (.A(_12847_),
    .Y(_15855_));
 BUFx6f_ASAP7_75t_R _21212_ (.A(_00852_),
    .Y(_12848_));
 INVx2_ASAP7_75t_R _21213_ (.A(net664),
    .Y(_12849_));
 BUFx6f_ASAP7_75t_R _21214_ (.A(_00795_),
    .Y(_12850_));
 XOR2x2_ASAP7_75t_R _21215_ (.A(_12829_),
    .B(_12850_),
    .Y(_12851_));
 NAND2x1_ASAP7_75t_R _21216_ (.A(_12849_),
    .B(_12851_),
    .Y(_12852_));
 XNOR2x1_ASAP7_75t_R _21217_ (.B(_12850_),
    .Y(_12853_),
    .A(_12829_));
 NAND2x1_ASAP7_75t_R _21218_ (.A(net666),
    .B(_12853_),
    .Y(_12854_));
 XNOR2x1_ASAP7_75t_R _21219_ (.B(net911),
    .Y(_12855_),
    .A(_12834_));
 AOI21x1_ASAP7_75t_R _21220_ (.A1(_12852_),
    .A2(_12854_),
    .B(_12855_),
    .Y(_12856_));
 NAND2x1_ASAP7_75t_R _21221_ (.A(net664),
    .B(_12851_),
    .Y(_12857_));
 NAND2x1_ASAP7_75t_R _21222_ (.A(_12849_),
    .B(_12853_),
    .Y(_12858_));
 XOR2x2_ASAP7_75t_R _21223_ (.A(_12834_),
    .B(_00820_),
    .Y(_12859_));
 AOI21x1_ASAP7_75t_R _21224_ (.A1(_12857_),
    .A2(_12858_),
    .B(_12859_),
    .Y(_12860_));
 OAI21x1_ASAP7_75t_R _21225_ (.A1(_12856_),
    .A2(_12860_),
    .B(_11356_),
    .Y(_12861_));
 INVx2_ASAP7_75t_R _21226_ (.A(_01107_),
    .Y(_12862_));
 NOR2x2_ASAP7_75t_R _21227_ (.A(net621),
    .B(_00520_),
    .Y(_12863_));
 INVx3_ASAP7_75t_R _21228_ (.A(_12863_),
    .Y(_12864_));
 NAND3x2_ASAP7_75t_R _21229_ (.B(_12862_),
    .C(_12864_),
    .Y(_12865_),
    .A(_12861_));
 AO21x1_ASAP7_75t_R _21230_ (.A1(_12861_),
    .A2(_12864_),
    .B(_12862_),
    .Y(_12866_));
 NAND2x2_ASAP7_75t_R _21231_ (.A(_12866_),
    .B(_12865_),
    .Y(_12867_));
 BUFx12f_ASAP7_75t_R _21232_ (.A(_12867_),
    .Y(_15857_));
 BUFx6f_ASAP7_75t_R _21233_ (.A(_00790_),
    .Y(_12868_));
 INVx2_ASAP7_75t_R _21234_ (.A(_12868_),
    .Y(_12869_));
 BUFx6f_ASAP7_75t_R _21235_ (.A(_00757_),
    .Y(_12870_));
 XOR2x2_ASAP7_75t_R _21236_ (.A(_12870_),
    .B(_00789_),
    .Y(_12871_));
 NAND2x1_ASAP7_75t_R _21237_ (.A(_12869_),
    .B(_12871_),
    .Y(_12872_));
 XNOR2x2_ASAP7_75t_R _21238_ (.A(_00789_),
    .B(_12870_),
    .Y(_12873_));
 NAND2x1_ASAP7_75t_R _21239_ (.A(_12868_),
    .B(_12873_),
    .Y(_12874_));
 XNOR2x2_ASAP7_75t_R _21240_ (.A(_00822_),
    .B(_00854_),
    .Y(_12875_));
 AOI21x1_ASAP7_75t_R _21241_ (.A1(_12872_),
    .A2(_12874_),
    .B(_12875_),
    .Y(_12876_));
 NAND2x1_ASAP7_75t_R _21242_ (.A(_12868_),
    .B(_12871_),
    .Y(_12877_));
 NAND2x1_ASAP7_75t_R _21243_ (.A(_12869_),
    .B(_12873_),
    .Y(_12878_));
 BUFx6f_ASAP7_75t_R _21244_ (.A(_00822_),
    .Y(_12879_));
 BUFx6f_ASAP7_75t_R _21245_ (.A(_00854_),
    .Y(_12880_));
 XOR2x2_ASAP7_75t_R _21246_ (.A(_12879_),
    .B(_12880_),
    .Y(_12881_));
 AOI21x1_ASAP7_75t_R _21247_ (.A1(_12877_),
    .A2(_12878_),
    .B(_12881_),
    .Y(_12882_));
 OAI21x1_ASAP7_75t_R _21248_ (.A1(_12876_),
    .A2(_12882_),
    .B(net680),
    .Y(_12883_));
 NOR2x2_ASAP7_75t_R _21249_ (.A(net786),
    .B(_00522_),
    .Y(_12884_));
 INVx3_ASAP7_75t_R _21250_ (.A(_12884_),
    .Y(_12885_));
 NAND3x2_ASAP7_75t_R _21251_ (.B(_08198_),
    .C(_12883_),
    .Y(_12886_),
    .A(_12885_));
 AO21x1_ASAP7_75t_R _21252_ (.A1(_12883_),
    .A2(_12885_),
    .B(_08198_),
    .Y(_12887_));
 BUFx6f_ASAP7_75t_R _21253_ (.A(_12887_),
    .Y(_12888_));
 NAND2x2_ASAP7_75t_R _21254_ (.A(_12886_),
    .B(_12888_),
    .Y(_12889_));
 BUFx10_ASAP7_75t_R _21255_ (.A(_12889_),
    .Y(_12890_));
 BUFx12_ASAP7_75t_R _21256_ (.A(_12890_),
    .Y(_15865_));
 NAND3x2_ASAP7_75t_R _21257_ (.B(_01107_),
    .C(_12864_),
    .Y(_12891_),
    .A(_12861_));
 AO21x1_ASAP7_75t_R _21258_ (.A1(_12864_),
    .A2(_12861_),
    .B(_01107_),
    .Y(_12892_));
 NAND2x2_ASAP7_75t_R _21259_ (.A(_12892_),
    .B(_12891_),
    .Y(_12893_));
 BUFx12f_ASAP7_75t_R _21260_ (.A(_12893_),
    .Y(_15852_));
 INVx3_ASAP7_75t_R _21261_ (.A(_08198_),
    .Y(_12894_));
 NAND3x2_ASAP7_75t_R _21262_ (.B(_12894_),
    .C(_12885_),
    .Y(_12895_),
    .A(_12883_));
 AO21x1_ASAP7_75t_R _21263_ (.A1(_12883_),
    .A2(_12885_),
    .B(_12894_),
    .Y(_12896_));
 BUFx4f_ASAP7_75t_R _21264_ (.A(_12896_),
    .Y(_12897_));
 NAND2x2_ASAP7_75t_R _21265_ (.A(_12895_),
    .B(_12897_),
    .Y(_12898_));
 BUFx12_ASAP7_75t_R _21266_ (.A(_12898_),
    .Y(_12899_));
 BUFx10_ASAP7_75t_R _21267_ (.A(_12899_),
    .Y(_15862_));
 XOR2x2_ASAP7_75t_R _21268_ (.A(_00794_),
    .B(_00826_),
    .Y(_12900_));
 XOR2x1_ASAP7_75t_R _21269_ (.A(_12900_),
    .Y(_12901_),
    .B(_00858_));
 BUFx4f_ASAP7_75t_R _21270_ (.A(_00761_),
    .Y(_12902_));
 XNOR2x2_ASAP7_75t_R _21271_ (.A(_12902_),
    .B(_00793_),
    .Y(_12903_));
 XOR2x1_ASAP7_75t_R _21272_ (.A(_12901_),
    .Y(_12904_),
    .B(_12903_));
 NOR2x1_ASAP7_75t_R _21273_ (.A(_11450_),
    .B(_00692_),
    .Y(_12905_));
 AO21x1_ASAP7_75t_R _21274_ (.A1(_12904_),
    .A2(_10787_),
    .B(_12905_),
    .Y(_12906_));
 XNOR2x2_ASAP7_75t_R _21275_ (.A(_01114_),
    .B(_12906_),
    .Y(_12907_));
 BUFx10_ASAP7_75t_R _21276_ (.A(_12907_),
    .Y(_12908_));
 NOR2x2_ASAP7_75t_R _21277_ (.A(net769),
    .B(_12890_),
    .Y(_12909_));
 BUFx6f_ASAP7_75t_R _21278_ (.A(_00758_),
    .Y(_12910_));
 XOR2x2_ASAP7_75t_R _21279_ (.A(_12910_),
    .B(_12829_),
    .Y(_12911_));
 XNOR2x1_ASAP7_75t_R _21280_ (.B(_12911_),
    .Y(_12912_),
    .A(_00791_));
 BUFx6f_ASAP7_75t_R _21281_ (.A(_00823_),
    .Y(_12913_));
 XNOR2x2_ASAP7_75t_R _21282_ (.A(_12913_),
    .B(_00855_),
    .Y(_12914_));
 XOR2x2_ASAP7_75t_R _21283_ (.A(_12868_),
    .B(net72),
    .Y(_12915_));
 XOR2x1_ASAP7_75t_R _21284_ (.A(_12914_),
    .Y(_12916_),
    .B(_12915_));
 NOR2x1_ASAP7_75t_R _21285_ (.A(_12912_),
    .B(_12916_),
    .Y(_12917_));
 XOR2x1_ASAP7_75t_R _21286_ (.A(_12911_),
    .Y(_12918_),
    .B(_00791_));
 XOR2x2_ASAP7_75t_R _21287_ (.A(_12913_),
    .B(_00855_),
    .Y(_12919_));
 XOR2x1_ASAP7_75t_R _21288_ (.A(_12915_),
    .Y(_12920_),
    .B(_12919_));
 BUFx12f_ASAP7_75t_R _21289_ (.A(_10620_),
    .Y(_12921_));
 OAI21x1_ASAP7_75t_R _21290_ (.A1(_12918_),
    .A2(_12920_),
    .B(_12921_),
    .Y(_12922_));
 NAND2x1_ASAP7_75t_R _21291_ (.A(_00695_),
    .B(net849),
    .Y(_12923_));
 OAI21x1_ASAP7_75t_R _21292_ (.A1(_12917_),
    .A2(_12922_),
    .B(_12923_),
    .Y(_12924_));
 XOR2x2_ASAP7_75t_R _21293_ (.A(_12924_),
    .B(_10068_),
    .Y(_12925_));
 BUFx10_ASAP7_75t_R _21294_ (.A(_12925_),
    .Y(_12926_));
 BUFx6f_ASAP7_75t_R _21295_ (.A(_12926_),
    .Y(_12927_));
 XOR2x2_ASAP7_75t_R _21296_ (.A(_00759_),
    .B(net647),
    .Y(_12928_));
 XOR2x1_ASAP7_75t_R _21297_ (.A(_12928_),
    .Y(_12929_),
    .B(_00792_));
 XOR2x2_ASAP7_75t_R _21298_ (.A(_00791_),
    .B(_00795_),
    .Y(_12930_));
 XOR2x2_ASAP7_75t_R _21299_ (.A(_00824_),
    .B(_00856_),
    .Y(_12931_));
 XOR2x1_ASAP7_75t_R _21300_ (.A(_12930_),
    .Y(_12932_),
    .B(_12931_));
 OAI21x1_ASAP7_75t_R _21301_ (.A1(_12929_),
    .A2(_12932_),
    .B(net763),
    .Y(_12933_));
 AND2x2_ASAP7_75t_R _21302_ (.A(_12932_),
    .B(_12929_),
    .Y(_12934_));
 AND2x2_ASAP7_75t_R _21303_ (.A(net866),
    .B(_00694_),
    .Y(_12935_));
 INVx1_ASAP7_75t_R _21304_ (.A(_12935_),
    .Y(_12936_));
 OAI21x1_ASAP7_75t_R _21305_ (.A1(_12933_),
    .A2(_12934_),
    .B(_12936_),
    .Y(_12937_));
 XOR2x2_ASAP7_75t_R _21306_ (.A(_12937_),
    .B(_01111_),
    .Y(_12938_));
 BUFx6f_ASAP7_75t_R _21307_ (.A(_12938_),
    .Y(_12939_));
 BUFx4f_ASAP7_75t_R _21308_ (.A(_12939_),
    .Y(_12940_));
 AO21x1_ASAP7_75t_R _21309_ (.A1(_12909_),
    .A2(_12927_),
    .B(_12940_),
    .Y(_12941_));
 OAI21x1_ASAP7_75t_R _21310_ (.A1(_12827_),
    .A2(_12840_),
    .B(_08191_),
    .Y(_12942_));
 OAI21x1_ASAP7_75t_R _21311_ (.A1(_12845_),
    .A2(_12843_),
    .B(_12841_),
    .Y(_12943_));
 NAND2x2_ASAP7_75t_R _21312_ (.A(_12942_),
    .B(_12943_),
    .Y(_12944_));
 BUFx6f_ASAP7_75t_R _21313_ (.A(_12944_),
    .Y(_15853_));
 NOR2x2_ASAP7_75t_R _21314_ (.A(_15857_),
    .B(net34),
    .Y(_12945_));
 BUFx4f_ASAP7_75t_R _21315_ (.A(_01177_),
    .Y(_12946_));
 BUFx6f_ASAP7_75t_R _21316_ (.A(_12889_),
    .Y(_12947_));
 BUFx6f_ASAP7_75t_R _21317_ (.A(_12925_),
    .Y(_12948_));
 AOI21x1_ASAP7_75t_R _21318_ (.A1(_12946_),
    .A2(_12947_),
    .B(_12948_),
    .Y(_12949_));
 INVx1_ASAP7_75t_R _21319_ (.A(_12949_),
    .Y(_12950_));
 AOI21x1_ASAP7_75t_R _21320_ (.A1(_15862_),
    .A2(_12945_),
    .B(_12950_),
    .Y(_12951_));
 BUFx6f_ASAP7_75t_R _21321_ (.A(_00760_),
    .Y(_12952_));
 XNOR2x2_ASAP7_75t_R _21322_ (.A(_12952_),
    .B(_00792_),
    .Y(_12953_));
 XOR2x2_ASAP7_75t_R _21323_ (.A(_00793_),
    .B(_00825_),
    .Y(_12954_));
 BUFx6f_ASAP7_75t_R _21324_ (.A(_00857_),
    .Y(_12955_));
 INVx3_ASAP7_75t_R _21325_ (.A(_12955_),
    .Y(_12956_));
 XOR2x1_ASAP7_75t_R _21326_ (.A(_12954_),
    .Y(_12957_),
    .B(_12956_));
 NAND2x1_ASAP7_75t_R _21327_ (.A(_12953_),
    .B(_12957_),
    .Y(_12958_));
 XOR2x1_ASAP7_75t_R _21328_ (.A(_12952_),
    .Y(_12959_),
    .B(_00792_));
 XOR2x1_ASAP7_75t_R _21329_ (.A(_12954_),
    .Y(_12960_),
    .B(_12955_));
 NAND2x1_ASAP7_75t_R _21330_ (.A(_12959_),
    .B(_12960_),
    .Y(_12961_));
 AOI21x1_ASAP7_75t_R _21331_ (.A1(_12958_),
    .A2(_12961_),
    .B(_12160_),
    .Y(_12962_));
 INVx2_ASAP7_75t_R _21332_ (.A(_01112_),
    .Y(_12963_));
 NOR2x2_ASAP7_75t_R _21333_ (.A(net763),
    .B(_00693_),
    .Y(_12964_));
 NOR3x2_ASAP7_75t_R _21334_ (.B(_12963_),
    .C(_12964_),
    .Y(_12965_),
    .A(_12962_));
 OA21x2_ASAP7_75t_R _21335_ (.A1(_12962_),
    .A2(_12964_),
    .B(_12963_),
    .Y(_12966_));
 NOR2x2_ASAP7_75t_R _21336_ (.A(_12965_),
    .B(_12966_),
    .Y(_12967_));
 BUFx10_ASAP7_75t_R _21337_ (.A(_12967_),
    .Y(_12968_));
 OAI21x1_ASAP7_75t_R _21338_ (.A1(_12941_),
    .A2(_12951_),
    .B(_12968_),
    .Y(_12969_));
 INVx4_ASAP7_75t_R _21339_ (.A(_12938_),
    .Y(_12970_));
 BUFx6f_ASAP7_75t_R _21340_ (.A(_12970_),
    .Y(_12971_));
 BUFx10_ASAP7_75t_R _21341_ (.A(_12971_),
    .Y(_12972_));
 INVx2_ASAP7_75t_R _21342_ (.A(_00521_),
    .Y(_12973_));
 XOR2x2_ASAP7_75t_R _21343_ (.A(_12924_),
    .B(_01110_),
    .Y(_12974_));
 BUFx10_ASAP7_75t_R _21344_ (.A(_12974_),
    .Y(_12975_));
 AOI21x1_ASAP7_75t_R _21345_ (.A1(_12973_),
    .A2(_12947_),
    .B(_12975_),
    .Y(_12976_));
 INVx1_ASAP7_75t_R _21346_ (.A(_12976_),
    .Y(_12977_));
 AOI211x1_ASAP7_75t_R _21347_ (.A1(_12846_),
    .A2(_12842_),
    .B(_12947_),
    .C(_15857_),
    .Y(_12978_));
 BUFx6f_ASAP7_75t_R _21348_ (.A(_12975_),
    .Y(_12979_));
 NAND2x1_ASAP7_75t_R _21349_ (.A(_12979_),
    .B(_12909_),
    .Y(_12980_));
 OAI21x1_ASAP7_75t_R _21350_ (.A1(_12977_),
    .A2(_12978_),
    .B(_12980_),
    .Y(_12981_));
 NOR2x1_ASAP7_75t_R _21351_ (.A(_12972_),
    .B(_12981_),
    .Y(_12982_));
 AOI211x1_ASAP7_75t_R _21352_ (.A1(_12844_),
    .A2(_10786_),
    .B(_12827_),
    .C(_08191_),
    .Y(_12983_));
 AOI211x1_ASAP7_75t_R _21353_ (.A1(_12839_),
    .A2(_11451_),
    .B(_12843_),
    .C(_12841_),
    .Y(_12984_));
 OAI21x1_ASAP7_75t_R _21354_ (.A1(_12983_),
    .A2(_12984_),
    .B(_12898_),
    .Y(_12985_));
 BUFx10_ASAP7_75t_R _21355_ (.A(_12985_),
    .Y(_12986_));
 BUFx5_ASAP7_75t_R _21356_ (.A(_01176_),
    .Y(_12987_));
 AOI21x1_ASAP7_75t_R _21357_ (.A1(_12886_),
    .A2(_12888_),
    .B(_12987_),
    .Y(_12988_));
 AOI21x1_ASAP7_75t_R _21358_ (.A1(net661),
    .A2(_12899_),
    .B(_12988_),
    .Y(_12989_));
 BUFx6f_ASAP7_75t_R _21359_ (.A(_12974_),
    .Y(_12990_));
 BUFx6f_ASAP7_75t_R _21360_ (.A(_12990_),
    .Y(_12991_));
 AOI21x1_ASAP7_75t_R _21361_ (.A1(_12986_),
    .A2(_12989_),
    .B(_12991_),
    .Y(_12992_));
 BUFx6f_ASAP7_75t_R _21362_ (.A(_12925_),
    .Y(_12993_));
 BUFx6f_ASAP7_75t_R _21363_ (.A(_12993_),
    .Y(_12994_));
 INVx1_ASAP7_75t_R _21364_ (.A(_00523_),
    .Y(_12995_));
 AOI21x1_ASAP7_75t_R _21365_ (.A1(_12895_),
    .A2(_12897_),
    .B(_12995_),
    .Y(_12996_));
 AOI21x1_ASAP7_75t_R _21366_ (.A1(net659),
    .A2(_12947_),
    .B(_12996_),
    .Y(_12997_));
 BUFx6f_ASAP7_75t_R _21367_ (.A(_12948_),
    .Y(_12998_));
 AOI21x1_ASAP7_75t_R _21368_ (.A1(_12886_),
    .A2(_12888_),
    .B(net771),
    .Y(_12999_));
 BUFx6f_ASAP7_75t_R _21369_ (.A(_12939_),
    .Y(_13000_));
 AOI21x1_ASAP7_75t_R _21370_ (.A1(_12998_),
    .A2(_12999_),
    .B(_13000_),
    .Y(_13001_));
 OAI21x1_ASAP7_75t_R _21371_ (.A1(_12994_),
    .A2(_12997_),
    .B(_13001_),
    .Y(_13002_));
 OR2x2_ASAP7_75t_R _21372_ (.A(_01180_),
    .B(_12993_),
    .Y(_13003_));
 BUFx4f_ASAP7_75t_R _21373_ (.A(_12948_),
    .Y(_13004_));
 AOI21x1_ASAP7_75t_R _21374_ (.A1(_12886_),
    .A2(_12888_),
    .B(net455),
    .Y(_13005_));
 AOI21x1_ASAP7_75t_R _21375_ (.A1(_13004_),
    .A2(net66),
    .B(_12971_),
    .Y(_13006_));
 BUFx10_ASAP7_75t_R _21376_ (.A(_12967_),
    .Y(_13007_));
 AOI21x1_ASAP7_75t_R _21377_ (.A1(_13003_),
    .A2(_13006_),
    .B(_13007_),
    .Y(_13008_));
 OAI21x1_ASAP7_75t_R _21378_ (.A1(_12992_),
    .A2(_13002_),
    .B(_13008_),
    .Y(_13009_));
 OAI21x1_ASAP7_75t_R _21379_ (.A1(_12969_),
    .A2(_12982_),
    .B(_13009_),
    .Y(_13010_));
 BUFx6f_ASAP7_75t_R _21380_ (.A(_00827_),
    .Y(_13011_));
 XOR2x2_ASAP7_75t_R _21381_ (.A(net72),
    .B(net908),
    .Y(_13012_));
 BUFx6f_ASAP7_75t_R _21382_ (.A(_00725_),
    .Y(_13013_));
 XOR2x1_ASAP7_75t_R _21383_ (.A(_13012_),
    .Y(_13014_),
    .B(_13013_));
 XNOR2x2_ASAP7_75t_R _21384_ (.A(_00762_),
    .B(_00794_),
    .Y(_13015_));
 XOR2x1_ASAP7_75t_R _21385_ (.A(_13014_),
    .Y(_13016_),
    .B(_13015_));
 BUFx12f_ASAP7_75t_R _21386_ (.A(_10734_),
    .Y(_13017_));
 NOR2x1_ASAP7_75t_R _21387_ (.A(_13017_),
    .B(_00691_),
    .Y(_13018_));
 AO21x1_ASAP7_75t_R _21388_ (.A1(_13016_),
    .A2(_10831_),
    .B(_13018_),
    .Y(_13019_));
 XOR2x2_ASAP7_75t_R _21389_ (.A(_13019_),
    .B(_01115_),
    .Y(_13020_));
 CKINVDCx6p67_ASAP7_75t_R _21390_ (.A(_13020_),
    .Y(_13021_));
 OAI21x1_ASAP7_75t_R _21391_ (.A1(_12908_),
    .A2(_13010_),
    .B(_13021_),
    .Y(_13022_));
 NOR2x2_ASAP7_75t_R _21392_ (.A(net660),
    .B(_12898_),
    .Y(_13023_));
 NOR2x1_ASAP7_75t_R _21393_ (.A(_12926_),
    .B(_13023_),
    .Y(_13024_));
 AOI211x1_ASAP7_75t_R _21394_ (.A1(_12846_),
    .A2(_12842_),
    .B(_12889_),
    .C(net520),
    .Y(_13025_));
 INVx1_ASAP7_75t_R _21395_ (.A(_13025_),
    .Y(_13026_));
 AO21x1_ASAP7_75t_R _21396_ (.A1(_12988_),
    .A2(_12948_),
    .B(_12939_),
    .Y(_13027_));
 AOI21x1_ASAP7_75t_R _21397_ (.A1(_13024_),
    .A2(_13026_),
    .B(_13027_),
    .Y(_13028_));
 AOI21x1_ASAP7_75t_R _21398_ (.A1(_12895_),
    .A2(_12897_),
    .B(_12946_),
    .Y(_13029_));
 OA21x2_ASAP7_75t_R _21399_ (.A1(_12988_),
    .A2(_13029_),
    .B(_12926_),
    .Y(_13030_));
 NOR2x1_ASAP7_75t_R _21400_ (.A(_12869_),
    .B(_12871_),
    .Y(_13031_));
 NOR2x1_ASAP7_75t_R _21401_ (.A(_12868_),
    .B(_12873_),
    .Y(_13032_));
 OAI21x1_ASAP7_75t_R _21402_ (.A1(_13031_),
    .A2(_13032_),
    .B(_12881_),
    .Y(_13033_));
 NOR2x1_ASAP7_75t_R _21403_ (.A(_12868_),
    .B(_12871_),
    .Y(_13034_));
 NOR2x1_ASAP7_75t_R _21404_ (.A(_12869_),
    .B(_12873_),
    .Y(_13035_));
 OAI21x1_ASAP7_75t_R _21405_ (.A1(_13034_),
    .A2(_13035_),
    .B(_12875_),
    .Y(_13036_));
 AOI21x1_ASAP7_75t_R _21406_ (.A1(_13033_),
    .A2(_13036_),
    .B(_12160_),
    .Y(_13037_));
 NOR3x2_ASAP7_75t_R _21407_ (.B(_08198_),
    .C(_12884_),
    .Y(_13038_),
    .A(_13037_));
 OA21x2_ASAP7_75t_R _21408_ (.A1(_13037_),
    .A2(_12884_),
    .B(_08198_),
    .Y(_13039_));
 OAI21x1_ASAP7_75t_R _21409_ (.A1(_13038_),
    .A2(_13039_),
    .B(net454),
    .Y(_13040_));
 NAND2x2_ASAP7_75t_R _21410_ (.A(_12974_),
    .B(_13040_),
    .Y(_13041_));
 INVx2_ASAP7_75t_R _21411_ (.A(_13041_),
    .Y(_13042_));
 NOR3x1_ASAP7_75t_R _21412_ (.A(_13030_),
    .B(_13042_),
    .C(_12972_),
    .Y(_13043_));
 INVx4_ASAP7_75t_R _21413_ (.A(_12967_),
    .Y(_13044_));
 BUFx10_ASAP7_75t_R _21414_ (.A(_13044_),
    .Y(_13045_));
 OAI21x1_ASAP7_75t_R _21415_ (.A1(_13028_),
    .A2(_13043_),
    .B(_13045_),
    .Y(_13046_));
 AO21x1_ASAP7_75t_R _21416_ (.A1(_12888_),
    .A2(_12886_),
    .B(_00521_),
    .Y(_13047_));
 INVx1_ASAP7_75t_R _21417_ (.A(_13047_),
    .Y(_13048_));
 BUFx6f_ASAP7_75t_R _21418_ (.A(_12975_),
    .Y(_13049_));
 OAI21x1_ASAP7_75t_R _21419_ (.A1(_15857_),
    .A2(_12947_),
    .B(_13049_),
    .Y(_13050_));
 NAND2x2_ASAP7_75t_R _21420_ (.A(_12970_),
    .B(_12967_),
    .Y(_13051_));
 INVx2_ASAP7_75t_R _21421_ (.A(_13051_),
    .Y(_13052_));
 OAI21x1_ASAP7_75t_R _21422_ (.A1(_13048_),
    .A2(_13050_),
    .B(_13052_),
    .Y(_13053_));
 AOI21x1_ASAP7_75t_R _21423_ (.A1(_12899_),
    .A2(net662),
    .B(_12974_),
    .Y(_13054_));
 INVx2_ASAP7_75t_R _21424_ (.A(_13005_),
    .Y(_13055_));
 AND2x4_ASAP7_75t_R _21425_ (.A(_13054_),
    .B(_13055_),
    .Y(_13056_));
 NOR2x1_ASAP7_75t_R _21426_ (.A(_13053_),
    .B(_13056_),
    .Y(_13057_));
 AOI21x1_ASAP7_75t_R _21427_ (.A1(_12886_),
    .A2(_12888_),
    .B(_12995_),
    .Y(_13058_));
 INVx2_ASAP7_75t_R _21428_ (.A(_13058_),
    .Y(_13059_));
 INVx1_ASAP7_75t_R _21429_ (.A(_12909_),
    .Y(_13060_));
 BUFx6f_ASAP7_75t_R _21430_ (.A(_12975_),
    .Y(_13061_));
 AOI21x1_ASAP7_75t_R _21431_ (.A1(_13059_),
    .A2(_13060_),
    .B(_13061_),
    .Y(_13062_));
 AOI21x1_ASAP7_75t_R _21432_ (.A1(_12987_),
    .A2(_12899_),
    .B(_12948_),
    .Y(_13063_));
 NAND2x2_ASAP7_75t_R _21433_ (.A(_12938_),
    .B(_12967_),
    .Y(_13064_));
 NOR3x1_ASAP7_75t_R _21434_ (.A(_13062_),
    .B(_13063_),
    .C(_13064_),
    .Y(_13065_));
 NOR2x1_ASAP7_75t_R _21435_ (.A(_13057_),
    .B(_13065_),
    .Y(_13066_));
 CKINVDCx8_ASAP7_75t_R _21436_ (.A(_12907_),
    .Y(_13067_));
 BUFx10_ASAP7_75t_R _21437_ (.A(_13067_),
    .Y(_13068_));
 AOI21x1_ASAP7_75t_R _21438_ (.A1(_13046_),
    .A2(_13066_),
    .B(_13068_),
    .Y(_13069_));
 INVx1_ASAP7_75t_R _21439_ (.A(net769),
    .Y(_13070_));
 OA21x2_ASAP7_75t_R _21440_ (.A1(_12890_),
    .A2(_13070_),
    .B(_12948_),
    .Y(_13071_));
 NAND2x2_ASAP7_75t_R _21441_ (.A(_12890_),
    .B(net662),
    .Y(_13072_));
 AND2x2_ASAP7_75t_R _21442_ (.A(_13071_),
    .B(_13072_),
    .Y(_13073_));
 AO21x2_ASAP7_75t_R _21443_ (.A1(net518),
    .A2(_12890_),
    .B(_12948_),
    .Y(_13074_));
 BUFx6f_ASAP7_75t_R _21444_ (.A(_12970_),
    .Y(_13075_));
 OAI21x1_ASAP7_75t_R _21445_ (.A1(_13074_),
    .A2(_13025_),
    .B(_13075_),
    .Y(_13076_));
 NOR2x1_ASAP7_75t_R _21446_ (.A(_13073_),
    .B(_13076_),
    .Y(_13077_));
 INVx3_ASAP7_75t_R _21447_ (.A(_01178_),
    .Y(_13078_));
 NOR2x2_ASAP7_75t_R _21448_ (.A(_13078_),
    .B(_15865_),
    .Y(_13079_));
 BUFx6f_ASAP7_75t_R _21449_ (.A(_12939_),
    .Y(_13080_));
 OAI21x1_ASAP7_75t_R _21450_ (.A1(_13079_),
    .A2(_13074_),
    .B(_13080_),
    .Y(_13081_));
 NAND2x2_ASAP7_75t_R _21451_ (.A(_12993_),
    .B(_12986_),
    .Y(_13082_));
 AOI211x1_ASAP7_75t_R _21452_ (.A1(_12846_),
    .A2(_12842_),
    .B(_15862_),
    .C(_15857_),
    .Y(_13083_));
 NOR2x1_ASAP7_75t_R _21453_ (.A(_13082_),
    .B(_13083_),
    .Y(_13084_));
 OAI21x1_ASAP7_75t_R _21454_ (.A1(_13081_),
    .A2(_13084_),
    .B(_12908_),
    .Y(_13085_));
 OAI21x1_ASAP7_75t_R _21455_ (.A1(_13077_),
    .A2(_13085_),
    .B(_13045_),
    .Y(_13086_));
 BUFx10_ASAP7_75t_R _21456_ (.A(_13000_),
    .Y(_13087_));
 INVx3_ASAP7_75t_R _21457_ (.A(net454),
    .Y(_13088_));
 OAI21x1_ASAP7_75t_R _21458_ (.A1(_13038_),
    .A2(_13039_),
    .B(_13088_),
    .Y(_13089_));
 NAND2x2_ASAP7_75t_R _21459_ (.A(_12925_),
    .B(_13089_),
    .Y(_13090_));
 INVx2_ASAP7_75t_R _21460_ (.A(_13090_),
    .Y(_13091_));
 OA21x2_ASAP7_75t_R _21461_ (.A1(_12899_),
    .A2(_13088_),
    .B(_12975_),
    .Y(_13092_));
 AO21x1_ASAP7_75t_R _21462_ (.A1(_13091_),
    .A2(_13072_),
    .B(_13092_),
    .Y(_13093_));
 NAND2x1_ASAP7_75t_R _21463_ (.A(_12948_),
    .B(_12996_),
    .Y(_13094_));
 AND2x2_ASAP7_75t_R _21464_ (.A(_13094_),
    .B(_12970_),
    .Y(_13095_));
 INVx1_ASAP7_75t_R _21465_ (.A(_13095_),
    .Y(_13096_));
 BUFx10_ASAP7_75t_R _21466_ (.A(_12899_),
    .Y(_13097_));
 NOR2x2_ASAP7_75t_R _21467_ (.A(_00523_),
    .B(_13097_),
    .Y(_13098_));
 AO21x2_ASAP7_75t_R _21468_ (.A1(_12888_),
    .A2(_12886_),
    .B(_12973_),
    .Y(_13099_));
 OAI22x1_ASAP7_75t_R _21469_ (.A1(net691),
    .A2(_13098_),
    .B1(_12991_),
    .B2(_13099_),
    .Y(_13100_));
 OAI21x1_ASAP7_75t_R _21470_ (.A1(_13096_),
    .A2(_13100_),
    .B(_13067_),
    .Y(_13101_));
 AOI21x1_ASAP7_75t_R _21471_ (.A1(_13087_),
    .A2(_13093_),
    .B(_13101_),
    .Y(_13102_));
 NOR2x1_ASAP7_75t_R _21472_ (.A(_13086_),
    .B(_13102_),
    .Y(_13103_));
 AOI21x1_ASAP7_75t_R _21473_ (.A1(_12895_),
    .A2(_12897_),
    .B(_12973_),
    .Y(_13104_));
 OAI21x1_ASAP7_75t_R _21474_ (.A1(_13058_),
    .A2(_13104_),
    .B(_12979_),
    .Y(_13105_));
 NAND2x1_ASAP7_75t_R _21475_ (.A(_13075_),
    .B(_13105_),
    .Y(_13106_));
 INVx1_ASAP7_75t_R _21476_ (.A(_12842_),
    .Y(_13107_));
 INVx1_ASAP7_75t_R _21477_ (.A(_12846_),
    .Y(_13108_));
 OAI21x1_ASAP7_75t_R _21478_ (.A1(_13107_),
    .A2(_13108_),
    .B(net660),
    .Y(_13109_));
 INVx2_ASAP7_75t_R _21479_ (.A(_13109_),
    .Y(_13110_));
 NAND2x1_ASAP7_75t_R _21480_ (.A(_12926_),
    .B(_13040_),
    .Y(_13111_));
 AOI21x1_ASAP7_75t_R _21481_ (.A1(_15865_),
    .A2(_13110_),
    .B(_13111_),
    .Y(_13112_));
 OAI21x1_ASAP7_75t_R _21482_ (.A1(_13106_),
    .A2(_13112_),
    .B(_13067_),
    .Y(_13113_));
 NOR2x2_ASAP7_75t_R _21483_ (.A(net521),
    .B(_12899_),
    .Y(_13114_));
 OAI21x1_ASAP7_75t_R _21484_ (.A1(net660),
    .A2(_12944_),
    .B(_12990_),
    .Y(_13115_));
 OAI21x1_ASAP7_75t_R _21485_ (.A1(_13114_),
    .A2(_13115_),
    .B(_13080_),
    .Y(_13116_));
 NAND2x1_ASAP7_75t_R _21486_ (.A(_15852_),
    .B(_12944_),
    .Y(_13117_));
 NOR2x2_ASAP7_75t_R _21487_ (.A(net520),
    .B(_12889_),
    .Y(_13118_));
 NOR2x1_ASAP7_75t_R _21488_ (.A(_12975_),
    .B(_13118_),
    .Y(_13119_));
 NAND2x1_ASAP7_75t_R _21489_ (.A(_13117_),
    .B(_13119_),
    .Y(_13120_));
 INVx1_ASAP7_75t_R _21490_ (.A(_13120_),
    .Y(_13121_));
 NOR2x1_ASAP7_75t_R _21491_ (.A(_13116_),
    .B(_13121_),
    .Y(_13122_));
 NOR2x1_ASAP7_75t_R _21492_ (.A(_13113_),
    .B(_13122_),
    .Y(_13123_));
 NAND2x2_ASAP7_75t_R _21493_ (.A(net517),
    .B(_12899_),
    .Y(_13124_));
 AOI21x1_ASAP7_75t_R _21494_ (.A1(_15855_),
    .A2(_13023_),
    .B(_12990_),
    .Y(_13125_));
 NOR2x2_ASAP7_75t_R _21495_ (.A(_13078_),
    .B(_12899_),
    .Y(_13126_));
 OAI21x1_ASAP7_75t_R _21496_ (.A1(_13126_),
    .A2(_13041_),
    .B(_13087_),
    .Y(_13127_));
 AOI21x1_ASAP7_75t_R _21497_ (.A1(_13124_),
    .A2(_13125_),
    .B(_13127_),
    .Y(_13128_));
 OAI21x1_ASAP7_75t_R _21498_ (.A1(_15857_),
    .A2(_13097_),
    .B(_12993_),
    .Y(_13129_));
 NAND2x1_ASAP7_75t_R _21499_ (.A(_13075_),
    .B(_13129_),
    .Y(_13130_));
 INVx1_ASAP7_75t_R _21500_ (.A(_12987_),
    .Y(_13131_));
 OAI21x1_ASAP7_75t_R _21501_ (.A1(_13131_),
    .A2(_15865_),
    .B(_13061_),
    .Y(_13132_));
 AOI21x1_ASAP7_75t_R _21502_ (.A1(_15865_),
    .A2(_12945_),
    .B(_13132_),
    .Y(_13133_));
 OAI21x1_ASAP7_75t_R _21503_ (.A1(_13130_),
    .A2(_13133_),
    .B(_12908_),
    .Y(_13134_));
 OAI21x1_ASAP7_75t_R _21504_ (.A1(_13128_),
    .A2(_13134_),
    .B(_12968_),
    .Y(_13135_));
 OAI21x1_ASAP7_75t_R _21505_ (.A1(_13123_),
    .A2(_13135_),
    .B(_13020_),
    .Y(_13136_));
 OAI22x1_ASAP7_75t_R _21506_ (.A1(_13069_),
    .A2(_13022_),
    .B1(_13103_),
    .B2(_13136_),
    .Y(_00056_));
 OAI21x1_ASAP7_75t_R _21507_ (.A1(_13038_),
    .A2(_13039_),
    .B(_13131_),
    .Y(_13137_));
 INVx1_ASAP7_75t_R _21508_ (.A(_13137_),
    .Y(_13138_));
 AO21x1_ASAP7_75t_R _21509_ (.A1(_13138_),
    .A2(_12998_),
    .B(_12940_),
    .Y(_13139_));
 INVx2_ASAP7_75t_R _21510_ (.A(_13089_),
    .Y(_13140_));
 OAI21x1_ASAP7_75t_R _21511_ (.A1(_13097_),
    .A2(_13109_),
    .B(_13049_),
    .Y(_13141_));
 NOR2x1_ASAP7_75t_R _21512_ (.A(_13140_),
    .B(_13141_),
    .Y(_13142_));
 NOR2x1_ASAP7_75t_R _21513_ (.A(_13139_),
    .B(_13142_),
    .Y(_13143_));
 OAI21x1_ASAP7_75t_R _21514_ (.A1(net648),
    .A2(net34),
    .B(_15862_),
    .Y(_13144_));
 NOR2x1_ASAP7_75t_R _21515_ (.A(_12926_),
    .B(_13126_),
    .Y(_13145_));
 AOI21x1_ASAP7_75t_R _21516_ (.A1(_12986_),
    .A2(_13145_),
    .B(_12971_),
    .Y(_13146_));
 OA21x2_ASAP7_75t_R _21517_ (.A1(_12991_),
    .A2(_13144_),
    .B(_13146_),
    .Y(_13147_));
 OAI21x1_ASAP7_75t_R _21518_ (.A1(_13143_),
    .A2(_13147_),
    .B(_12968_),
    .Y(_13148_));
 INVx1_ASAP7_75t_R _21519_ (.A(_12988_),
    .Y(_13149_));
 BUFx6f_ASAP7_75t_R _21520_ (.A(_12970_),
    .Y(_13150_));
 AO21x1_ASAP7_75t_R _21521_ (.A1(_12997_),
    .A2(_12998_),
    .B(_13150_),
    .Y(_13151_));
 AO21x1_ASAP7_75t_R _21522_ (.A1(_13149_),
    .A2(_13042_),
    .B(_13151_),
    .Y(_13152_));
 NOR2x2_ASAP7_75t_R _21523_ (.A(_13005_),
    .B(_12975_),
    .Y(_13153_));
 NAND2x1_ASAP7_75t_R _21524_ (.A(_13124_),
    .B(_13153_),
    .Y(_13154_));
 NAND2x2_ASAP7_75t_R _21525_ (.A(_15857_),
    .B(net34),
    .Y(_13155_));
 NAND2x1_ASAP7_75t_R _21526_ (.A(_13155_),
    .B(_13024_),
    .Y(_13156_));
 NAND2x1_ASAP7_75t_R _21527_ (.A(_13154_),
    .B(_13156_),
    .Y(_13157_));
 AOI21x1_ASAP7_75t_R _21528_ (.A1(_12972_),
    .A2(_13157_),
    .B(_12968_),
    .Y(_13158_));
 AOI21x1_ASAP7_75t_R _21529_ (.A1(_13152_),
    .A2(_13158_),
    .B(_13068_),
    .Y(_13159_));
 NAND2x1_ASAP7_75t_R _21530_ (.A(_13148_),
    .B(_13159_),
    .Y(_13160_));
 NAND2x1_ASAP7_75t_R _21531_ (.A(_12890_),
    .B(_12975_),
    .Y(_13161_));
 AO21x2_ASAP7_75t_R _21532_ (.A1(net772),
    .A2(net648),
    .B(_13161_),
    .Y(_13162_));
 NAND2x1_ASAP7_75t_R _21533_ (.A(_13117_),
    .B(_13054_),
    .Y(_13163_));
 NAND2x1_ASAP7_75t_R _21534_ (.A(_13162_),
    .B(_13163_),
    .Y(_13164_));
 OAI21x1_ASAP7_75t_R _21535_ (.A1(_13138_),
    .A2(_13023_),
    .B(_12998_),
    .Y(_13165_));
 OAI21x1_ASAP7_75t_R _21536_ (.A1(_13140_),
    .A2(_13114_),
    .B(_13061_),
    .Y(_13166_));
 AOI21x1_ASAP7_75t_R _21537_ (.A1(_13165_),
    .A2(_13166_),
    .B(_13064_),
    .Y(_13167_));
 AOI21x1_ASAP7_75t_R _21538_ (.A1(_13052_),
    .A2(_13164_),
    .B(_13167_),
    .Y(_13168_));
 BUFx6f_ASAP7_75t_R _21539_ (.A(_12974_),
    .Y(_13169_));
 OA21x2_ASAP7_75t_R _21540_ (.A1(_13149_),
    .A2(_13169_),
    .B(_13000_),
    .Y(_13170_));
 INVx3_ASAP7_75t_R _21541_ (.A(_12985_),
    .Y(_13171_));
 AOI21x1_ASAP7_75t_R _21542_ (.A1(_13061_),
    .A2(_13072_),
    .B(_13171_),
    .Y(_13172_));
 AOI21x1_ASAP7_75t_R _21543_ (.A1(_13170_),
    .A2(_13172_),
    .B(_13007_),
    .Y(_13173_));
 AND2x2_ASAP7_75t_R _21544_ (.A(_12989_),
    .B(_12986_),
    .Y(_13174_));
 AOI21x1_ASAP7_75t_R _21545_ (.A1(_12895_),
    .A2(_12897_),
    .B(net580),
    .Y(_13175_));
 OAI21x1_ASAP7_75t_R _21546_ (.A1(_13175_),
    .A2(_13005_),
    .B(_12990_),
    .Y(_13176_));
 AND2x2_ASAP7_75t_R _21547_ (.A(_12971_),
    .B(_13176_),
    .Y(_13177_));
 OAI21x1_ASAP7_75t_R _21548_ (.A1(_12991_),
    .A2(_13174_),
    .B(_13177_),
    .Y(_13178_));
 NAND2x1_ASAP7_75t_R _21549_ (.A(_13173_),
    .B(_13178_),
    .Y(_13179_));
 NAND2x1_ASAP7_75t_R _21550_ (.A(_13168_),
    .B(_13179_),
    .Y(_13180_));
 AOI21x1_ASAP7_75t_R _21551_ (.A1(_13068_),
    .A2(_13180_),
    .B(_13020_),
    .Y(_13181_));
 NAND2x2_ASAP7_75t_R _21552_ (.A(_15862_),
    .B(_13049_),
    .Y(_13182_));
 INVx3_ASAP7_75t_R _21553_ (.A(_13064_),
    .Y(_13183_));
 OAI21x1_ASAP7_75t_R _21554_ (.A1(_13182_),
    .A2(_13110_),
    .B(_13183_),
    .Y(_13184_));
 INVx1_ASAP7_75t_R _21555_ (.A(_13162_),
    .Y(_13185_));
 AO21x1_ASAP7_75t_R _21556_ (.A1(net648),
    .A2(_13097_),
    .B(_12990_),
    .Y(_13186_));
 NOR2x1_ASAP7_75t_R _21557_ (.A(_13098_),
    .B(_13186_),
    .Y(_13187_));
 NOR3x1_ASAP7_75t_R _21558_ (.A(_13184_),
    .B(_13185_),
    .C(_13187_),
    .Y(_13188_));
 OAI21x1_ASAP7_75t_R _21559_ (.A1(_12983_),
    .A2(_12984_),
    .B(_12889_),
    .Y(_13189_));
 OAI21x1_ASAP7_75t_R _21560_ (.A1(_12965_),
    .A2(_12966_),
    .B(_12939_),
    .Y(_13190_));
 AOI21x1_ASAP7_75t_R _21561_ (.A1(_13189_),
    .A2(_13063_),
    .B(_13190_),
    .Y(_13191_));
 AO21x1_ASAP7_75t_R _21562_ (.A1(_13189_),
    .A2(_13124_),
    .B(_13049_),
    .Y(_13192_));
 NAND2x1_ASAP7_75t_R _21563_ (.A(_13191_),
    .B(_13192_),
    .Y(_13193_));
 OAI21x1_ASAP7_75t_R _21564_ (.A1(_15865_),
    .A2(_13109_),
    .B(_12976_),
    .Y(_13194_));
 NAND2x1_ASAP7_75t_R _21565_ (.A(_00525_),
    .B(_12990_),
    .Y(_13195_));
 OA21x2_ASAP7_75t_R _21566_ (.A1(_13195_),
    .A2(_12967_),
    .B(_12971_),
    .Y(_13196_));
 AOI21x1_ASAP7_75t_R _21567_ (.A1(_13194_),
    .A2(_13196_),
    .B(_12907_),
    .Y(_13197_));
 NAND2x1_ASAP7_75t_R _21568_ (.A(_13193_),
    .B(_13197_),
    .Y(_13198_));
 OAI21x1_ASAP7_75t_R _21569_ (.A1(_13188_),
    .A2(_13198_),
    .B(_13020_),
    .Y(_13199_));
 OAI21x1_ASAP7_75t_R _21570_ (.A1(net66),
    .A2(_12996_),
    .B(_13061_),
    .Y(_13200_));
 OAI21x1_ASAP7_75t_R _21571_ (.A1(_12909_),
    .A2(_13114_),
    .B(_12998_),
    .Y(_13201_));
 AOI21x1_ASAP7_75t_R _21572_ (.A1(_13200_),
    .A2(_13201_),
    .B(_13075_),
    .Y(_13202_));
 NAND2x2_ASAP7_75t_R _21573_ (.A(_13189_),
    .B(_13063_),
    .Y(_13203_));
 NOR2x2_ASAP7_75t_R _21574_ (.A(_15857_),
    .B(_12947_),
    .Y(_13204_));
 OAI21x1_ASAP7_75t_R _21575_ (.A1(_13058_),
    .A2(_13204_),
    .B(_12927_),
    .Y(_13205_));
 AOI21x1_ASAP7_75t_R _21576_ (.A1(_13203_),
    .A2(_13205_),
    .B(_13080_),
    .Y(_13206_));
 OAI21x1_ASAP7_75t_R _21577_ (.A1(_13202_),
    .A2(_13206_),
    .B(_12968_),
    .Y(_13207_));
 AOI21x1_ASAP7_75t_R _21578_ (.A1(net580),
    .A2(_13097_),
    .B(_12990_),
    .Y(_13208_));
 AO21x1_ASAP7_75t_R _21579_ (.A1(_12888_),
    .A2(_12886_),
    .B(_13070_),
    .Y(_13209_));
 AO21x1_ASAP7_75t_R _21580_ (.A1(_13208_),
    .A2(_13209_),
    .B(_13075_),
    .Y(_13210_));
 AOI21x1_ASAP7_75t_R _21581_ (.A1(net517),
    .A2(_12890_),
    .B(_12975_),
    .Y(_13211_));
 OAI21x1_ASAP7_75t_R _21582_ (.A1(_15865_),
    .A2(_13109_),
    .B(_13211_),
    .Y(_13212_));
 NOR2x1_ASAP7_75t_R _21583_ (.A(_13000_),
    .B(_13042_),
    .Y(_13213_));
 AOI21x1_ASAP7_75t_R _21584_ (.A1(_13212_),
    .A2(_13213_),
    .B(_13007_),
    .Y(_13214_));
 OAI21x1_ASAP7_75t_R _21585_ (.A1(_13142_),
    .A2(_13210_),
    .B(_13214_),
    .Y(_13215_));
 AOI21x1_ASAP7_75t_R _21586_ (.A1(_13207_),
    .A2(_13215_),
    .B(_13068_),
    .Y(_13216_));
 NOR2x1_ASAP7_75t_R _21587_ (.A(_13199_),
    .B(_13216_),
    .Y(_13217_));
 AOI21x1_ASAP7_75t_R _21588_ (.A1(_13160_),
    .A2(_13181_),
    .B(_13217_),
    .Y(_00057_));
 AND2x4_ASAP7_75t_R _21589_ (.A(_12987_),
    .B(_01175_),
    .Y(_13218_));
 INVx2_ASAP7_75t_R _21590_ (.A(_13218_),
    .Y(_13219_));
 AO21x2_ASAP7_75t_R _21591_ (.A1(_12897_),
    .A2(_12895_),
    .B(_13219_),
    .Y(_13220_));
 NAND2x1_ASAP7_75t_R _21592_ (.A(_13049_),
    .B(_13220_),
    .Y(_13221_));
 NOR2x2_ASAP7_75t_R _21593_ (.A(_13097_),
    .B(_13109_),
    .Y(_13222_));
 NOR2x1_ASAP7_75t_R _21594_ (.A(_13221_),
    .B(_13222_),
    .Y(_13223_));
 NAND2x1_ASAP7_75t_R _21595_ (.A(_13080_),
    .B(_13194_),
    .Y(_13224_));
 AO21x1_ASAP7_75t_R _21596_ (.A1(_13149_),
    .A2(_13089_),
    .B(_13004_),
    .Y(_13225_));
 AOI21x1_ASAP7_75t_R _21597_ (.A1(_13225_),
    .A2(_13095_),
    .B(_13044_),
    .Y(_13226_));
 OAI21x1_ASAP7_75t_R _21598_ (.A1(_13223_),
    .A2(_13224_),
    .B(_13226_),
    .Y(_13227_));
 NAND2x2_ASAP7_75t_R _21599_ (.A(net519),
    .B(_12890_),
    .Y(_13228_));
 OAI21x1_ASAP7_75t_R _21600_ (.A1(net34),
    .A2(_13228_),
    .B(_13004_),
    .Y(_13229_));
 NAND2x1_ASAP7_75t_R _21601_ (.A(_00526_),
    .B(_13169_),
    .Y(_13230_));
 NAND3x1_ASAP7_75t_R _21602_ (.A(_13229_),
    .B(_13150_),
    .C(_13230_),
    .Y(_13231_));
 OA21x2_ASAP7_75t_R _21603_ (.A1(_13049_),
    .A2(_01182_),
    .B(_13000_),
    .Y(_13232_));
 OAI21x1_ASAP7_75t_R _21604_ (.A1(net648),
    .A2(_13097_),
    .B(net772),
    .Y(_13233_));
 NAND2x1_ASAP7_75t_R _21605_ (.A(_12979_),
    .B(_13233_),
    .Y(_13234_));
 AOI21x1_ASAP7_75t_R _21606_ (.A1(_13232_),
    .A2(_13234_),
    .B(_13007_),
    .Y(_13235_));
 AOI21x1_ASAP7_75t_R _21607_ (.A1(_13231_),
    .A2(_13235_),
    .B(_12907_),
    .Y(_13236_));
 AOI21x1_ASAP7_75t_R _21608_ (.A1(_13227_),
    .A2(_13236_),
    .B(_13020_),
    .Y(_13237_));
 OA21x2_ASAP7_75t_R _21609_ (.A1(_01180_),
    .A2(_13169_),
    .B(_12970_),
    .Y(_13238_));
 NAND2x2_ASAP7_75t_R _21610_ (.A(net648),
    .B(_15855_),
    .Y(_13239_));
 OAI21x1_ASAP7_75t_R _21611_ (.A1(_15865_),
    .A2(_13239_),
    .B(_13092_),
    .Y(_13240_));
 AOI21x1_ASAP7_75t_R _21612_ (.A1(_13238_),
    .A2(_13240_),
    .B(_13044_),
    .Y(_13241_));
 AOI21x1_ASAP7_75t_R _21613_ (.A1(_12943_),
    .A2(_12942_),
    .B(_12898_),
    .Y(_13242_));
 AOI21x1_ASAP7_75t_R _21614_ (.A1(_13055_),
    .A2(_13054_),
    .B(_13150_),
    .Y(_13243_));
 OAI21x1_ASAP7_75t_R _21615_ (.A1(_13050_),
    .A2(_13242_),
    .B(_13243_),
    .Y(_13244_));
 AOI21x1_ASAP7_75t_R _21616_ (.A1(_13241_),
    .A2(_13244_),
    .B(_13067_),
    .Y(_13245_));
 INVx1_ASAP7_75t_R _21617_ (.A(_13104_),
    .Y(_13246_));
 NOR2x1_ASAP7_75t_R _21618_ (.A(_13004_),
    .B(_13005_),
    .Y(_13247_));
 AOI22x1_ASAP7_75t_R _21619_ (.A1(_13054_),
    .A2(_13059_),
    .B1(_13246_),
    .B2(_13247_),
    .Y(_13248_));
 NAND2x2_ASAP7_75t_R _21620_ (.A(_13097_),
    .B(net772),
    .Y(_13249_));
 AOI21x1_ASAP7_75t_R _21621_ (.A1(_15852_),
    .A2(_15853_),
    .B(_12926_),
    .Y(_13250_));
 AND2x2_ASAP7_75t_R _21622_ (.A(_12948_),
    .B(_00525_),
    .Y(_13251_));
 AOI21x1_ASAP7_75t_R _21623_ (.A1(_13249_),
    .A2(_13250_),
    .B(_13251_),
    .Y(_13252_));
 AOI21x1_ASAP7_75t_R _21624_ (.A1(_13075_),
    .A2(_13252_),
    .B(_13007_),
    .Y(_13253_));
 OAI21x1_ASAP7_75t_R _21625_ (.A1(_12972_),
    .A2(_13248_),
    .B(_13253_),
    .Y(_13254_));
 NAND2x1_ASAP7_75t_R _21626_ (.A(_13245_),
    .B(_13254_),
    .Y(_13255_));
 NAND2x1_ASAP7_75t_R _21627_ (.A(_13237_),
    .B(_13255_),
    .Y(_13256_));
 AOI21x1_ASAP7_75t_R _21628_ (.A1(_12987_),
    .A2(_12947_),
    .B(_12993_),
    .Y(_13257_));
 AO21x1_ASAP7_75t_R _21629_ (.A1(_12986_),
    .A2(_13257_),
    .B(_13030_),
    .Y(_13258_));
 INVx2_ASAP7_75t_R _21630_ (.A(_13029_),
    .Y(_13259_));
 NOR3x1_ASAP7_75t_R _21631_ (.A(_13037_),
    .B(_12894_),
    .C(_12884_),
    .Y(_13260_));
 OA21x2_ASAP7_75t_R _21632_ (.A1(_13037_),
    .A2(_12884_),
    .B(_12894_),
    .Y(_13261_));
 OAI21x1_ASAP7_75t_R _21633_ (.A1(_13260_),
    .A2(_13261_),
    .B(_13078_),
    .Y(_13262_));
 AO21x1_ASAP7_75t_R _21634_ (.A1(_13259_),
    .A2(_13262_),
    .B(_13049_),
    .Y(_13263_));
 AOI21x1_ASAP7_75t_R _21635_ (.A1(_13124_),
    .A2(_13257_),
    .B(_13150_),
    .Y(_13264_));
 AOI21x1_ASAP7_75t_R _21636_ (.A1(_13263_),
    .A2(_13264_),
    .B(_13007_),
    .Y(_13265_));
 OAI21x1_ASAP7_75t_R _21637_ (.A1(_13087_),
    .A2(_13258_),
    .B(_13265_),
    .Y(_13266_));
 AOI21x1_ASAP7_75t_R _21638_ (.A1(_12946_),
    .A2(_12947_),
    .B(_12975_),
    .Y(_13267_));
 NAND2x1_ASAP7_75t_R _21639_ (.A(_13124_),
    .B(_13267_),
    .Y(_13268_));
 AO21x2_ASAP7_75t_R _21640_ (.A1(_12888_),
    .A2(_12886_),
    .B(_13088_),
    .Y(_13269_));
 AO21x1_ASAP7_75t_R _21641_ (.A1(_13269_),
    .A2(net570),
    .B(_13004_),
    .Y(_13270_));
 AOI21x1_ASAP7_75t_R _21642_ (.A1(_13268_),
    .A2(_13270_),
    .B(_13080_),
    .Y(_13271_));
 NOR2x2_ASAP7_75t_R _21643_ (.A(_12926_),
    .B(_13242_),
    .Y(_13272_));
 OAI21x1_ASAP7_75t_R _21644_ (.A1(net581),
    .A2(_13097_),
    .B(_12993_),
    .Y(_13273_));
 OAI21x1_ASAP7_75t_R _21645_ (.A1(_13118_),
    .A2(_13273_),
    .B(_13000_),
    .Y(_13274_));
 AOI21x1_ASAP7_75t_R _21646_ (.A1(_13259_),
    .A2(_13272_),
    .B(_13274_),
    .Y(_13275_));
 OAI21x1_ASAP7_75t_R _21647_ (.A1(_13271_),
    .A2(_13275_),
    .B(_12968_),
    .Y(_13276_));
 AOI21x1_ASAP7_75t_R _21648_ (.A1(_13266_),
    .A2(_13276_),
    .B(_13068_),
    .Y(_13277_));
 NOR2x2_ASAP7_75t_R _21649_ (.A(_12948_),
    .B(_12988_),
    .Y(_13278_));
 INVx1_ASAP7_75t_R _21650_ (.A(_13278_),
    .Y(_13279_));
 NAND2x2_ASAP7_75t_R _21651_ (.A(net659),
    .B(_12899_),
    .Y(_13280_));
 NAND2x1_ASAP7_75t_R _21652_ (.A(_13280_),
    .B(_12986_),
    .Y(_13281_));
 OAI21x1_ASAP7_75t_R _21653_ (.A1(_13279_),
    .A2(_13281_),
    .B(_12971_),
    .Y(_13282_));
 NOR2x2_ASAP7_75t_R _21654_ (.A(_13056_),
    .B(_13282_),
    .Y(_13283_));
 AOI21x1_ASAP7_75t_R _21655_ (.A1(_13262_),
    .A2(_13137_),
    .B(_12990_),
    .Y(_13284_));
 AOI21x1_ASAP7_75t_R _21656_ (.A1(_12979_),
    .A2(_13233_),
    .B(_13284_),
    .Y(_13285_));
 BUFx6f_ASAP7_75t_R _21657_ (.A(_13044_),
    .Y(_13286_));
 OAI21x1_ASAP7_75t_R _21658_ (.A1(_13075_),
    .A2(_13285_),
    .B(_13286_),
    .Y(_13287_));
 NOR2x1_ASAP7_75t_R _21659_ (.A(_13287_),
    .B(_13283_),
    .Y(_13288_));
 NOR2x1_ASAP7_75t_R _21660_ (.A(_13051_),
    .B(_13125_),
    .Y(_13289_));
 OAI21x1_ASAP7_75t_R _21661_ (.A1(_13079_),
    .A2(_13141_),
    .B(_13289_),
    .Y(_13290_));
 OAI21x1_ASAP7_75t_R _21662_ (.A1(net770),
    .A2(_13097_),
    .B(_13169_),
    .Y(_13291_));
 OAI22x1_ASAP7_75t_R _21663_ (.A1(_13242_),
    .A2(_13090_),
    .B1(_13118_),
    .B2(_13291_),
    .Y(_13292_));
 AOI21x1_ASAP7_75t_R _21664_ (.A1(_13183_),
    .A2(_13292_),
    .B(_12907_),
    .Y(_13293_));
 NAND2x1_ASAP7_75t_R _21665_ (.A(_13290_),
    .B(_13293_),
    .Y(_13294_));
 NOR2x1_ASAP7_75t_R _21666_ (.A(_13288_),
    .B(_13294_),
    .Y(_13295_));
 OAI21x1_ASAP7_75t_R _21667_ (.A1(_13277_),
    .A2(_13295_),
    .B(_13020_),
    .Y(_13296_));
 NAND2x1_ASAP7_75t_R _21668_ (.A(_13296_),
    .B(_13256_),
    .Y(_00058_));
 NOR2x1_ASAP7_75t_R _21669_ (.A(_13104_),
    .B(_13114_),
    .Y(_13297_));
 NAND2x1_ASAP7_75t_R _21670_ (.A(_13297_),
    .B(_13272_),
    .Y(_13298_));
 AOI21x1_ASAP7_75t_R _21671_ (.A1(_13153_),
    .A2(_13144_),
    .B(_13080_),
    .Y(_13299_));
 NOR2x2_ASAP7_75t_R _21672_ (.A(_13114_),
    .B(_13115_),
    .Y(_13300_));
 INVx1_ASAP7_75t_R _21673_ (.A(_13300_),
    .Y(_13301_));
 INVx1_ASAP7_75t_R _21674_ (.A(_13099_),
    .Y(_13302_));
 OA21x2_ASAP7_75t_R _21675_ (.A1(_13111_),
    .A2(_13302_),
    .B(_12940_),
    .Y(_13303_));
 AOI22x1_ASAP7_75t_R _21676_ (.A1(_13298_),
    .A2(_13299_),
    .B1(_13301_),
    .B2(_13303_),
    .Y(_13304_));
 NOR2x1_ASAP7_75t_R _21677_ (.A(net659),
    .B(net772),
    .Y(_13305_));
 AO21x1_ASAP7_75t_R _21678_ (.A1(net659),
    .A2(_12890_),
    .B(_12939_),
    .Y(_13306_));
 NOR2x1_ASAP7_75t_R _21679_ (.A(_13305_),
    .B(_13306_),
    .Y(_13307_));
 AOI21x1_ASAP7_75t_R _21680_ (.A1(_13182_),
    .A2(_13307_),
    .B(_12967_),
    .Y(_13308_));
 AO21x1_ASAP7_75t_R _21681_ (.A1(_12946_),
    .A2(_12947_),
    .B(_13090_),
    .Y(_13309_));
 NAND2x1_ASAP7_75t_R _21682_ (.A(_13309_),
    .B(_13146_),
    .Y(_13310_));
 AOI21x1_ASAP7_75t_R _21683_ (.A1(_13308_),
    .A2(_13310_),
    .B(_13067_),
    .Y(_13311_));
 OAI21x1_ASAP7_75t_R _21684_ (.A1(_13045_),
    .A2(_13304_),
    .B(_13311_),
    .Y(_13312_));
 OAI21x1_ASAP7_75t_R _21685_ (.A1(_12988_),
    .A2(_13175_),
    .B(_12979_),
    .Y(_13313_));
 AOI21x1_ASAP7_75t_R _21686_ (.A1(_13189_),
    .A2(_13091_),
    .B(_13000_),
    .Y(_13314_));
 AOI21x1_ASAP7_75t_R _21687_ (.A1(_13313_),
    .A2(_13314_),
    .B(_13044_),
    .Y(_13315_));
 INVx1_ASAP7_75t_R _21688_ (.A(_12996_),
    .Y(_13316_));
 AND3x1_ASAP7_75t_R _21689_ (.A(_13269_),
    .B(_13169_),
    .C(_13316_),
    .Y(_13317_));
 NAND2x2_ASAP7_75t_R _21690_ (.A(net659),
    .B(_12890_),
    .Y(_13318_));
 AND3x1_ASAP7_75t_R _21691_ (.A(_13318_),
    .B(_13246_),
    .C(_12993_),
    .Y(_13319_));
 OAI21x1_ASAP7_75t_R _21692_ (.A1(_13317_),
    .A2(_13319_),
    .B(_13080_),
    .Y(_13320_));
 NAND2x1_ASAP7_75t_R _21693_ (.A(_13320_),
    .B(_13315_),
    .Y(_13321_));
 NOR2x1_ASAP7_75t_R _21694_ (.A(_12971_),
    .B(_13092_),
    .Y(_13322_));
 NAND3x1_ASAP7_75t_R _21695_ (.A(_13189_),
    .B(_13124_),
    .C(_12998_),
    .Y(_13323_));
 AOI21x1_ASAP7_75t_R _21696_ (.A1(_13322_),
    .A2(_13323_),
    .B(_13007_),
    .Y(_13324_));
 NAND2x1_ASAP7_75t_R _21697_ (.A(_13239_),
    .B(_13119_),
    .Y(_13325_));
 OA21x2_ASAP7_75t_R _21698_ (.A1(_13041_),
    .A2(_13242_),
    .B(_12971_),
    .Y(_13326_));
 NAND2x1_ASAP7_75t_R _21699_ (.A(_13325_),
    .B(_13326_),
    .Y(_13327_));
 AOI21x1_ASAP7_75t_R _21700_ (.A1(_13324_),
    .A2(_13327_),
    .B(_12908_),
    .Y(_13328_));
 AOI21x1_ASAP7_75t_R _21701_ (.A1(_13321_),
    .A2(_13328_),
    .B(_13020_),
    .Y(_13329_));
 NAND2x1_ASAP7_75t_R _21702_ (.A(_13312_),
    .B(_13329_),
    .Y(_13330_));
 AO21x1_ASAP7_75t_R _21703_ (.A1(_13228_),
    .A2(_13259_),
    .B(_13004_),
    .Y(_13331_));
 AO21x1_ASAP7_75t_R _21704_ (.A1(net570),
    .A2(_13262_),
    .B(_12979_),
    .Y(_13332_));
 AND3x1_ASAP7_75t_R _21705_ (.A(_13331_),
    .B(_13080_),
    .C(_13332_),
    .Y(_13333_));
 OA21x2_ASAP7_75t_R _21706_ (.A1(_12997_),
    .A2(_12998_),
    .B(_13150_),
    .Y(_13334_));
 AO21x1_ASAP7_75t_R _21707_ (.A1(_13334_),
    .A2(_13163_),
    .B(_13286_),
    .Y(_13335_));
 INVx1_ASAP7_75t_R _21708_ (.A(_13274_),
    .Y(_13336_));
 NAND2x1_ASAP7_75t_R _21709_ (.A(_13220_),
    .B(_12949_),
    .Y(_13337_));
 AOI21x1_ASAP7_75t_R _21710_ (.A1(_13337_),
    .A2(_13194_),
    .B(_13087_),
    .Y(_13338_));
 OAI21x1_ASAP7_75t_R _21711_ (.A1(_13336_),
    .A2(_13338_),
    .B(_13045_),
    .Y(_13339_));
 OAI21x1_ASAP7_75t_R _21712_ (.A1(_13333_),
    .A2(_13335_),
    .B(_13339_),
    .Y(_13340_));
 INVx1_ASAP7_75t_R _21713_ (.A(_12980_),
    .Y(_13341_));
 NOR2x1_ASAP7_75t_R _21714_ (.A(_13302_),
    .B(_13171_),
    .Y(_13342_));
 AO21x1_ASAP7_75t_R _21715_ (.A1(_13269_),
    .A2(_13049_),
    .B(_12967_),
    .Y(_13343_));
 AOI21x1_ASAP7_75t_R _21716_ (.A1(_12994_),
    .A2(_13342_),
    .B(_13343_),
    .Y(_13344_));
 OAI21x1_ASAP7_75t_R _21717_ (.A1(_13341_),
    .A2(_13344_),
    .B(_13087_),
    .Y(_13345_));
 NAND2x1_ASAP7_75t_R _21718_ (.A(_13040_),
    .B(_13211_),
    .Y(_13346_));
 INVx2_ASAP7_75t_R _21719_ (.A(_13126_),
    .Y(_13347_));
 NAND3x1_ASAP7_75t_R _21720_ (.A(_13347_),
    .B(_13220_),
    .C(_12979_),
    .Y(_13348_));
 NOR2x2_ASAP7_75t_R _21721_ (.A(_12939_),
    .B(_12967_),
    .Y(_13349_));
 INVx2_ASAP7_75t_R _21722_ (.A(_13349_),
    .Y(_13350_));
 AOI21x1_ASAP7_75t_R _21723_ (.A1(_13346_),
    .A2(_13348_),
    .B(_13350_),
    .Y(_13351_));
 NOR2x1_ASAP7_75t_R _21724_ (.A(_12993_),
    .B(_13259_),
    .Y(_13352_));
 AOI21x1_ASAP7_75t_R _21725_ (.A1(_13124_),
    .A2(_13267_),
    .B(_13352_),
    .Y(_13353_));
 NOR2x1_ASAP7_75t_R _21726_ (.A(_12990_),
    .B(_13040_),
    .Y(_13354_));
 AOI21x1_ASAP7_75t_R _21727_ (.A1(_13354_),
    .A2(_13183_),
    .B(_12907_),
    .Y(_13355_));
 OAI21x1_ASAP7_75t_R _21728_ (.A1(_13051_),
    .A2(_13353_),
    .B(_13355_),
    .Y(_13356_));
 NOR2x1_ASAP7_75t_R _21729_ (.A(_13351_),
    .B(_13356_),
    .Y(_13357_));
 AOI21x1_ASAP7_75t_R _21730_ (.A1(_13345_),
    .A2(_13357_),
    .B(_13021_),
    .Y(_13358_));
 OAI21x1_ASAP7_75t_R _21731_ (.A1(_13068_),
    .A2(_13340_),
    .B(_13358_),
    .Y(_13359_));
 NAND2x1_ASAP7_75t_R _21732_ (.A(_13330_),
    .B(_13359_),
    .Y(_00059_));
 AO21x1_ASAP7_75t_R _21733_ (.A1(_13208_),
    .A2(_13269_),
    .B(_12940_),
    .Y(_13360_));
 NOR2x1_ASAP7_75t_R _21734_ (.A(_12951_),
    .B(_13360_),
    .Y(_13361_));
 AOI21x1_ASAP7_75t_R _21735_ (.A1(_12991_),
    .A2(net66),
    .B(_13029_),
    .Y(_13362_));
 AO21x1_ASAP7_75t_R _21736_ (.A1(_13170_),
    .A2(_13362_),
    .B(_13286_),
    .Y(_13363_));
 AOI21x1_ASAP7_75t_R _21737_ (.A1(_13316_),
    .A2(_13072_),
    .B(_12994_),
    .Y(_13364_));
 OAI21x1_ASAP7_75t_R _21738_ (.A1(_12992_),
    .A2(_13364_),
    .B(_13349_),
    .Y(_13365_));
 OAI21x1_ASAP7_75t_R _21739_ (.A1(_13361_),
    .A2(_13363_),
    .B(_13365_),
    .Y(_13366_));
 NOR2x1_ASAP7_75t_R _21740_ (.A(_12927_),
    .B(_12978_),
    .Y(_13367_));
 AOI21x1_ASAP7_75t_R _21741_ (.A1(_13189_),
    .A2(_13367_),
    .B(_13284_),
    .Y(_13368_));
 OAI21x1_ASAP7_75t_R _21742_ (.A1(_13190_),
    .A2(_13368_),
    .B(_13068_),
    .Y(_13369_));
 OAI21x1_ASAP7_75t_R _21743_ (.A1(_13366_),
    .A2(_13369_),
    .B(_13021_),
    .Y(_13370_));
 NOR2x1_ASAP7_75t_R _21744_ (.A(_13150_),
    .B(_12909_),
    .Y(_13371_));
 AO21x1_ASAP7_75t_R _21745_ (.A1(_13371_),
    .A2(_12950_),
    .B(_13286_),
    .Y(_13372_));
 OAI21x1_ASAP7_75t_R _21746_ (.A1(_13098_),
    .A2(_13186_),
    .B(_13075_),
    .Y(_13373_));
 AO21x1_ASAP7_75t_R _21747_ (.A1(_12847_),
    .A2(_12947_),
    .B(_12926_),
    .Y(_13374_));
 NOR2x1_ASAP7_75t_R _21748_ (.A(_13204_),
    .B(_13374_),
    .Y(_13375_));
 NOR2x1_ASAP7_75t_R _21749_ (.A(_13373_),
    .B(_13375_),
    .Y(_13376_));
 OAI21x1_ASAP7_75t_R _21750_ (.A1(_13372_),
    .A2(_13376_),
    .B(_12908_),
    .Y(_13377_));
 AOI21x1_ASAP7_75t_R _21751_ (.A1(_13059_),
    .A2(_13249_),
    .B(_12927_),
    .Y(_13378_));
 NOR2x1_ASAP7_75t_R _21752_ (.A(_13110_),
    .B(_13082_),
    .Y(_13379_));
 OAI21x1_ASAP7_75t_R _21753_ (.A1(_13378_),
    .A2(_13379_),
    .B(_13087_),
    .Y(_13380_));
 AOI21x1_ASAP7_75t_R _21754_ (.A1(_13072_),
    .A2(_13155_),
    .B(_12994_),
    .Y(_13381_));
 INVx1_ASAP7_75t_R _21755_ (.A(_13192_),
    .Y(_13382_));
 OAI21x1_ASAP7_75t_R _21756_ (.A1(_13381_),
    .A2(_13382_),
    .B(_12972_),
    .Y(_13383_));
 AOI21x1_ASAP7_75t_R _21757_ (.A1(_13380_),
    .A2(_13383_),
    .B(_12968_),
    .Y(_13384_));
 NOR2x1_ASAP7_75t_R _21758_ (.A(_13377_),
    .B(_13384_),
    .Y(_13385_));
 NAND2x1_ASAP7_75t_R _21759_ (.A(_12979_),
    .B(_13005_),
    .Y(_13386_));
 INVx1_ASAP7_75t_R _21760_ (.A(_00527_),
    .Y(_13387_));
 AOI21x1_ASAP7_75t_R _21761_ (.A1(_13387_),
    .A2(_12994_),
    .B(_13051_),
    .Y(_13388_));
 AOI21x1_ASAP7_75t_R _21762_ (.A1(_13386_),
    .A2(_13388_),
    .B(_12907_),
    .Y(_13389_));
 OAI21x1_ASAP7_75t_R _21763_ (.A1(_13062_),
    .A2(_13300_),
    .B(_13349_),
    .Y(_13390_));
 NAND2x1_ASAP7_75t_R _21764_ (.A(_13389_),
    .B(_13390_),
    .Y(_13391_));
 OA211x2_ASAP7_75t_R _21765_ (.A1(_12946_),
    .A2(_15862_),
    .B(_13124_),
    .C(_12991_),
    .Y(_13392_));
 AOI21x1_ASAP7_75t_R _21766_ (.A1(_15862_),
    .A2(net34),
    .B(_12991_),
    .Y(_13393_));
 AO21x1_ASAP7_75t_R _21767_ (.A1(_13393_),
    .A2(_13109_),
    .B(_13190_),
    .Y(_13394_));
 NAND2x2_ASAP7_75t_R _21768_ (.A(_12986_),
    .B(_12949_),
    .Y(_13395_));
 INVx1_ASAP7_75t_R _21769_ (.A(_13395_),
    .Y(_13396_));
 OAI21x1_ASAP7_75t_R _21770_ (.A1(_15857_),
    .A2(net34),
    .B(_15862_),
    .Y(_13397_));
 NOR2x1_ASAP7_75t_R _21771_ (.A(_12991_),
    .B(_13397_),
    .Y(_13398_));
 OAI21x1_ASAP7_75t_R _21772_ (.A1(_13396_),
    .A2(_13398_),
    .B(_13183_),
    .Y(_13399_));
 OAI21x1_ASAP7_75t_R _21773_ (.A1(_13392_),
    .A2(_13394_),
    .B(_13399_),
    .Y(_13400_));
 OAI21x1_ASAP7_75t_R _21774_ (.A1(_13391_),
    .A2(_13400_),
    .B(_13020_),
    .Y(_13401_));
 AO21x1_ASAP7_75t_R _21775_ (.A1(_15862_),
    .A2(_12987_),
    .B(_13049_),
    .Y(_13402_));
 NOR2x1_ASAP7_75t_R _21776_ (.A(net66),
    .B(_13402_),
    .Y(_13403_));
 AOI21x1_ASAP7_75t_R _21777_ (.A1(_12927_),
    .A2(_13209_),
    .B(_13150_),
    .Y(_13404_));
 AOI21x1_ASAP7_75t_R _21778_ (.A1(_13404_),
    .A2(_13141_),
    .B(_13286_),
    .Y(_13405_));
 OA21x2_ASAP7_75t_R _21779_ (.A1(_13076_),
    .A2(_13403_),
    .B(_13405_),
    .Y(_13406_));
 AO21x1_ASAP7_75t_R _21780_ (.A1(_12926_),
    .A2(_12996_),
    .B(_12970_),
    .Y(_13407_));
 NOR2x1_ASAP7_75t_R _21781_ (.A(_12991_),
    .B(_13189_),
    .Y(_13408_));
 AOI211x1_ASAP7_75t_R _21782_ (.A1(_13063_),
    .A2(_13189_),
    .B(_13407_),
    .C(_13408_),
    .Y(_13409_));
 AO21x1_ASAP7_75t_R _21783_ (.A1(_13124_),
    .A2(_13262_),
    .B(_13061_),
    .Y(_13410_));
 AND2x2_ASAP7_75t_R _21784_ (.A(_13161_),
    .B(_12971_),
    .Y(_13411_));
 AO21x1_ASAP7_75t_R _21785_ (.A1(_13410_),
    .A2(_13411_),
    .B(_12968_),
    .Y(_13412_));
 OAI21x1_ASAP7_75t_R _21786_ (.A1(_13409_),
    .A2(_13412_),
    .B(_12908_),
    .Y(_13413_));
 NOR2x1_ASAP7_75t_R _21787_ (.A(_13406_),
    .B(_13413_),
    .Y(_13414_));
 OAI22x1_ASAP7_75t_R _21788_ (.A1(_13370_),
    .A2(_13385_),
    .B1(_13401_),
    .B2(_13414_),
    .Y(_00060_));
 OAI21x1_ASAP7_75t_R _21789_ (.A1(_13058_),
    .A2(net691),
    .B(_13273_),
    .Y(_13415_));
 AND2x2_ASAP7_75t_R _21790_ (.A(_13386_),
    .B(_13080_),
    .Y(_13416_));
 OAI21x1_ASAP7_75t_R _21791_ (.A1(_12999_),
    .A2(_13171_),
    .B(_12994_),
    .Y(_13417_));
 AOI221x1_ASAP7_75t_R _21792_ (.A1(_12972_),
    .A2(_13415_),
    .B1(_13416_),
    .B2(_13417_),
    .C(_12908_),
    .Y(_13418_));
 AND2x2_ASAP7_75t_R _21793_ (.A(_13111_),
    .B(_13150_),
    .Y(_13419_));
 AO21x1_ASAP7_75t_R _21794_ (.A1(_13331_),
    .A2(_13419_),
    .B(_13067_),
    .Y(_13420_));
 AND3x1_ASAP7_75t_R _21795_ (.A(_13162_),
    .B(_13087_),
    .C(_13402_),
    .Y(_13421_));
 OAI21x1_ASAP7_75t_R _21796_ (.A1(_13420_),
    .A2(_13421_),
    .B(_13045_),
    .Y(_13422_));
 OAI21x1_ASAP7_75t_R _21797_ (.A1(_13418_),
    .A2(_13422_),
    .B(_13021_),
    .Y(_13423_));
 NOR2x1_ASAP7_75t_R _21798_ (.A(_12927_),
    .B(net34),
    .Y(_13424_));
 OAI21x1_ASAP7_75t_R _21799_ (.A1(_13424_),
    .A2(_13379_),
    .B(_12972_),
    .Y(_13425_));
 OAI21x1_ASAP7_75t_R _21800_ (.A1(_13048_),
    .A2(_13025_),
    .B(_12991_),
    .Y(_13426_));
 OA21x2_ASAP7_75t_R _21801_ (.A1(_13110_),
    .A2(_13129_),
    .B(_12940_),
    .Y(_13427_));
 AOI21x1_ASAP7_75t_R _21802_ (.A1(_13426_),
    .A2(_13427_),
    .B(_12908_),
    .Y(_13428_));
 NAND2x1_ASAP7_75t_R _21803_ (.A(_13425_),
    .B(_13428_),
    .Y(_13429_));
 INVx1_ASAP7_75t_R _21804_ (.A(_12978_),
    .Y(_13430_));
 AO21x1_ASAP7_75t_R _21805_ (.A1(_13257_),
    .A2(_13219_),
    .B(_13075_),
    .Y(_13431_));
 AOI21x1_ASAP7_75t_R _21806_ (.A1(_13430_),
    .A2(_13267_),
    .B(_13431_),
    .Y(_13432_));
 AOI221x1_ASAP7_75t_R _21807_ (.A1(_13063_),
    .A2(_13347_),
    .B1(_13072_),
    .B2(_13071_),
    .C(_13087_),
    .Y(_13433_));
 OAI21x1_ASAP7_75t_R _21808_ (.A1(_13432_),
    .A2(_13433_),
    .B(_12908_),
    .Y(_13434_));
 AOI21x1_ASAP7_75t_R _21809_ (.A1(_13429_),
    .A2(_13434_),
    .B(_13045_),
    .Y(_13435_));
 INVx1_ASAP7_75t_R _21810_ (.A(_13145_),
    .Y(_13436_));
 AOI21x1_ASAP7_75t_R _21811_ (.A1(_13436_),
    .A2(_13170_),
    .B(_13286_),
    .Y(_13437_));
 AO21x1_ASAP7_75t_R _21812_ (.A1(_13169_),
    .A2(_13220_),
    .B(_12939_),
    .Y(_13438_));
 AO21x1_ASAP7_75t_R _21813_ (.A1(_13026_),
    .A2(_13125_),
    .B(_13438_),
    .Y(_13439_));
 NAND2x1_ASAP7_75t_R _21814_ (.A(_13439_),
    .B(_13437_),
    .Y(_13440_));
 NAND2x1_ASAP7_75t_R _21815_ (.A(_00521_),
    .B(_13061_),
    .Y(_13441_));
 OAI21x1_ASAP7_75t_R _21816_ (.A1(_15865_),
    .A2(_13109_),
    .B(_12927_),
    .Y(_13442_));
 AOI21x1_ASAP7_75t_R _21817_ (.A1(_13441_),
    .A2(_13442_),
    .B(_13350_),
    .Y(_13443_));
 AOI21x1_ASAP7_75t_R _21818_ (.A1(_13040_),
    .A2(_13262_),
    .B(_13049_),
    .Y(_13444_));
 AOI21x1_ASAP7_75t_R _21819_ (.A1(net570),
    .A2(_13099_),
    .B(_12993_),
    .Y(_13445_));
 INVx2_ASAP7_75t_R _21820_ (.A(_13190_),
    .Y(_13446_));
 OAI21x1_ASAP7_75t_R _21821_ (.A1(_13444_),
    .A2(_13445_),
    .B(_13446_),
    .Y(_13447_));
 NAND2x1_ASAP7_75t_R _21822_ (.A(_13067_),
    .B(_13447_),
    .Y(_13448_));
 NOR2x1_ASAP7_75t_R _21823_ (.A(_13443_),
    .B(_13448_),
    .Y(_13449_));
 AOI21x1_ASAP7_75t_R _21824_ (.A1(_13449_),
    .A2(_13440_),
    .B(_13021_),
    .Y(_13450_));
 AOI21x1_ASAP7_75t_R _21825_ (.A1(_12986_),
    .A2(_13267_),
    .B(_13150_),
    .Y(_13451_));
 OAI21x1_ASAP7_75t_R _21826_ (.A1(net691),
    .A2(_13083_),
    .B(_13451_),
    .Y(_13452_));
 OA21x2_ASAP7_75t_R _21827_ (.A1(net648),
    .A2(_13004_),
    .B(_12971_),
    .Y(_13453_));
 AOI21x1_ASAP7_75t_R _21828_ (.A1(_13453_),
    .A2(_13120_),
    .B(_13286_),
    .Y(_13454_));
 AOI21x1_ASAP7_75t_R _21829_ (.A1(_13452_),
    .A2(_13454_),
    .B(_13067_),
    .Y(_13455_));
 OA21x2_ASAP7_75t_R _21830_ (.A1(_13099_),
    .A2(_13004_),
    .B(_13000_),
    .Y(_13456_));
 NOR2x1_ASAP7_75t_R _21831_ (.A(_15857_),
    .B(_13169_),
    .Y(_13457_));
 OAI21x1_ASAP7_75t_R _21832_ (.A1(_13457_),
    .A2(_13054_),
    .B(_13347_),
    .Y(_13458_));
 AOI21x1_ASAP7_75t_R _21833_ (.A1(_13456_),
    .A2(_13458_),
    .B(_13007_),
    .Y(_13459_));
 NAND2x1_ASAP7_75t_R _21834_ (.A(_13004_),
    .B(_13118_),
    .Y(_13460_));
 NAND2x1_ASAP7_75t_R _21835_ (.A(_13460_),
    .B(_13028_),
    .Y(_13461_));
 NAND2x1_ASAP7_75t_R _21836_ (.A(_13459_),
    .B(_13461_),
    .Y(_13462_));
 NAND2x1_ASAP7_75t_R _21837_ (.A(_13455_),
    .B(_13462_),
    .Y(_13463_));
 NAND2x1_ASAP7_75t_R _21838_ (.A(_13463_),
    .B(_13450_),
    .Y(_13464_));
 OAI21x1_ASAP7_75t_R _21839_ (.A1(_13423_),
    .A2(_13435_),
    .B(_13464_),
    .Y(_00061_));
 OA21x2_ASAP7_75t_R _21840_ (.A1(_13029_),
    .A2(_12999_),
    .B(_12990_),
    .Y(_13465_));
 AO21x1_ASAP7_75t_R _21841_ (.A1(_13279_),
    .A2(_13460_),
    .B(_13465_),
    .Y(_13466_));
 AND2x2_ASAP7_75t_R _21842_ (.A(_13006_),
    .B(_13044_),
    .Y(_13467_));
 AO21x1_ASAP7_75t_R _21843_ (.A1(_13466_),
    .A2(_13467_),
    .B(_13068_),
    .Y(_13468_));
 NAND2x1_ASAP7_75t_R _21844_ (.A(_01181_),
    .B(_01179_),
    .Y(_13469_));
 AO21x1_ASAP7_75t_R _21845_ (.A1(_12993_),
    .A2(_13469_),
    .B(_12939_),
    .Y(_13470_));
 AO21x1_ASAP7_75t_R _21846_ (.A1(_13272_),
    .A2(_13239_),
    .B(_13470_),
    .Y(_13471_));
 OA21x2_ASAP7_75t_R _21847_ (.A1(_13465_),
    .A2(_13407_),
    .B(_12967_),
    .Y(_13472_));
 AND2x2_ASAP7_75t_R _21848_ (.A(_13471_),
    .B(_13472_),
    .Y(_13473_));
 AOI21x1_ASAP7_75t_R _21849_ (.A1(_12886_),
    .A2(_12888_),
    .B(_12946_),
    .Y(_13474_));
 OAI21x1_ASAP7_75t_R _21850_ (.A1(_13474_),
    .A2(_13175_),
    .B(_12998_),
    .Y(_13475_));
 NOR2x1_ASAP7_75t_R _21851_ (.A(_13023_),
    .B(_13242_),
    .Y(_13476_));
 AO21x1_ASAP7_75t_R _21852_ (.A1(_13476_),
    .A2(_13060_),
    .B(_12994_),
    .Y(_13477_));
 AOI21x1_ASAP7_75t_R _21853_ (.A1(_13475_),
    .A2(_13477_),
    .B(_13350_),
    .Y(_13478_));
 NOR3x2_ASAP7_75t_R _21854_ (.B(_13473_),
    .C(_13478_),
    .Y(_13479_),
    .A(_13468_));
 AO21x1_ASAP7_75t_R _21855_ (.A1(_13220_),
    .A2(_13153_),
    .B(_12940_),
    .Y(_13480_));
 AOI21x1_ASAP7_75t_R _21856_ (.A1(_13318_),
    .A2(_13367_),
    .B(_13480_),
    .Y(_13481_));
 AO21x1_ASAP7_75t_R _21857_ (.A1(_13280_),
    .A2(net772),
    .B(_12998_),
    .Y(_13482_));
 OA21x2_ASAP7_75t_R _21858_ (.A1(_13099_),
    .A2(_13061_),
    .B(_12940_),
    .Y(_13483_));
 AO21x1_ASAP7_75t_R _21859_ (.A1(_13482_),
    .A2(_13483_),
    .B(_12968_),
    .Y(_13484_));
 OAI21x1_ASAP7_75t_R _21860_ (.A1(_13484_),
    .A2(_13481_),
    .B(_13068_),
    .Y(_13485_));
 INVx1_ASAP7_75t_R _21861_ (.A(_13354_),
    .Y(_13486_));
 NAND2x1_ASAP7_75t_R _21862_ (.A(_13230_),
    .B(_13229_),
    .Y(_13487_));
 AOI21x1_ASAP7_75t_R _21863_ (.A1(_13486_),
    .A2(_13487_),
    .B(_12972_),
    .Y(_13488_));
 AO21x1_ASAP7_75t_R _21864_ (.A1(_13209_),
    .A2(_13091_),
    .B(_12940_),
    .Y(_13489_));
 NOR3x1_ASAP7_75t_R _21865_ (.A(_13083_),
    .B(_12927_),
    .C(_13171_),
    .Y(_13490_));
 OAI21x1_ASAP7_75t_R _21866_ (.A1(_13490_),
    .A2(_13489_),
    .B(_12968_),
    .Y(_13491_));
 NOR2x1_ASAP7_75t_R _21867_ (.A(_13488_),
    .B(_13491_),
    .Y(_13492_));
 OAI21x1_ASAP7_75t_R _21868_ (.A1(_13492_),
    .A2(_13485_),
    .B(_13021_),
    .Y(_13493_));
 AO21x1_ASAP7_75t_R _21869_ (.A1(_13114_),
    .A2(_12927_),
    .B(_13150_),
    .Y(_13494_));
 NOR2x1_ASAP7_75t_R _21870_ (.A(_13140_),
    .B(_13436_),
    .Y(_13495_));
 AOI21x1_ASAP7_75t_R _21871_ (.A1(_00528_),
    .A2(_13061_),
    .B(_13000_),
    .Y(_13496_));
 NAND2x1_ASAP7_75t_R _21872_ (.A(_12986_),
    .B(_13267_),
    .Y(_13497_));
 AOI21x1_ASAP7_75t_R _21873_ (.A1(_13496_),
    .A2(_13497_),
    .B(_13286_),
    .Y(_13498_));
 OAI21x1_ASAP7_75t_R _21874_ (.A1(_13494_),
    .A2(_13495_),
    .B(_13498_),
    .Y(_13499_));
 AO21x1_ASAP7_75t_R _21875_ (.A1(_13395_),
    .A2(_12977_),
    .B(_13190_),
    .Y(_13500_));
 AOI21x1_ASAP7_75t_R _21876_ (.A1(_13278_),
    .A2(_13397_),
    .B(_13080_),
    .Y(_13501_));
 AOI21x1_ASAP7_75t_R _21877_ (.A1(_13045_),
    .A2(_13501_),
    .B(_12907_),
    .Y(_13502_));
 NAND3x1_ASAP7_75t_R _21878_ (.A(_13499_),
    .B(_13500_),
    .C(_13502_),
    .Y(_13503_));
 OA21x2_ASAP7_75t_R _21879_ (.A1(_13250_),
    .A2(_13208_),
    .B(_13318_),
    .Y(_13504_));
 NOR2x1_ASAP7_75t_R _21880_ (.A(_13169_),
    .B(net772),
    .Y(_13505_));
 INVx1_ASAP7_75t_R _21881_ (.A(_13505_),
    .Y(_13506_));
 AOI21x1_ASAP7_75t_R _21882_ (.A1(_13506_),
    .A2(_13307_),
    .B(_13286_),
    .Y(_13507_));
 OAI21x1_ASAP7_75t_R _21883_ (.A1(_12972_),
    .A2(_13504_),
    .B(_13507_),
    .Y(_13508_));
 NAND2x1_ASAP7_75t_R _21884_ (.A(_13090_),
    .B(_13349_),
    .Y(_13509_));
 NOR2x1_ASAP7_75t_R _21885_ (.A(_13029_),
    .B(_13074_),
    .Y(_13510_));
 OAI21x1_ASAP7_75t_R _21886_ (.A1(_13509_),
    .A2(_13510_),
    .B(_12907_),
    .Y(_13511_));
 OAI21x1_ASAP7_75t_R _21887_ (.A1(_13211_),
    .A2(_13505_),
    .B(_13124_),
    .Y(_13512_));
 AOI21x1_ASAP7_75t_R _21888_ (.A1(_13374_),
    .A2(_13512_),
    .B(_13190_),
    .Y(_13513_));
 NOR2x1_ASAP7_75t_R _21889_ (.A(_13511_),
    .B(_13513_),
    .Y(_13514_));
 AOI21x1_ASAP7_75t_R _21890_ (.A1(_13508_),
    .A2(_13514_),
    .B(_13021_),
    .Y(_13515_));
 NAND2x1_ASAP7_75t_R _21891_ (.A(_13515_),
    .B(_13503_),
    .Y(_13516_));
 OAI21x1_ASAP7_75t_R _21892_ (.A1(_13493_),
    .A2(_13479_),
    .B(_13516_),
    .Y(_00062_));
 NOR2x1_ASAP7_75t_R _21893_ (.A(_13222_),
    .B(net639),
    .Y(_13517_));
 OAI21x1_ASAP7_75t_R _21894_ (.A1(_12994_),
    .A2(_12978_),
    .B(_13087_),
    .Y(_13518_));
 NOR2x1_ASAP7_75t_R _21895_ (.A(_13518_),
    .B(_13517_),
    .Y(_13519_));
 OA211x2_ASAP7_75t_R _21896_ (.A1(_13110_),
    .A2(_13182_),
    .B(_13486_),
    .C(_13075_),
    .Y(_13520_));
 OAI21x1_ASAP7_75t_R _21897_ (.A1(_13519_),
    .A2(_13520_),
    .B(_13045_),
    .Y(_13521_));
 OAI21x1_ASAP7_75t_R _21898_ (.A1(_13082_),
    .A2(_13222_),
    .B(_13007_),
    .Y(_13522_));
 AO21x1_ASAP7_75t_R _21899_ (.A1(_13250_),
    .A2(_13249_),
    .B(_12940_),
    .Y(_13523_));
 OAI21x1_ASAP7_75t_R _21900_ (.A1(_13522_),
    .A2(_13523_),
    .B(_13067_),
    .Y(_13524_));
 NAND2x2_ASAP7_75t_R _21901_ (.A(_15852_),
    .B(_12926_),
    .Y(_13525_));
 INVx1_ASAP7_75t_R _21902_ (.A(_13375_),
    .Y(_13526_));
 AOI21x1_ASAP7_75t_R _21903_ (.A1(_13525_),
    .A2(_13526_),
    .B(_13064_),
    .Y(_13527_));
 NOR2x1_ASAP7_75t_R _21904_ (.A(_13524_),
    .B(_13527_),
    .Y(_13528_));
 INVx1_ASAP7_75t_R _21905_ (.A(_13040_),
    .Y(_13529_));
 OAI21x1_ASAP7_75t_R _21906_ (.A1(_13529_),
    .A2(_13129_),
    .B(_13176_),
    .Y(_13530_));
 OAI21x1_ASAP7_75t_R _21907_ (.A1(_13050_),
    .A2(_13242_),
    .B(_13475_),
    .Y(_13531_));
 AOI22x1_ASAP7_75t_R _21908_ (.A1(_13530_),
    .A2(_13446_),
    .B1(_13531_),
    .B2(_13349_),
    .Y(_13532_));
 AOI21x1_ASAP7_75t_R _21909_ (.A1(_15865_),
    .A2(net34),
    .B(_12996_),
    .Y(_13533_));
 AOI21x1_ASAP7_75t_R _21910_ (.A1(_13228_),
    .A2(_13533_),
    .B(_12994_),
    .Y(_13534_));
 OAI21x1_ASAP7_75t_R _21911_ (.A1(_13129_),
    .A2(_12978_),
    .B(_13087_),
    .Y(_13535_));
 NOR2x1_ASAP7_75t_R _21912_ (.A(_12940_),
    .B(_13208_),
    .Y(_13536_));
 AOI21x1_ASAP7_75t_R _21913_ (.A1(_13395_),
    .A2(_13536_),
    .B(_13286_),
    .Y(_13537_));
 OAI21x1_ASAP7_75t_R _21914_ (.A1(_13534_),
    .A2(_13535_),
    .B(_13537_),
    .Y(_13538_));
 AOI21x1_ASAP7_75t_R _21915_ (.A1(_13532_),
    .A2(_13538_),
    .B(_13068_),
    .Y(_13539_));
 AOI21x1_ASAP7_75t_R _21916_ (.A1(_13521_),
    .A2(_13528_),
    .B(_13539_),
    .Y(_13540_));
 OAI21x1_ASAP7_75t_R _21917_ (.A1(_13169_),
    .A2(net772),
    .B(_12939_),
    .Y(_13541_));
 NOR2x1_ASAP7_75t_R _21918_ (.A(_15862_),
    .B(_13525_),
    .Y(_13542_));
 NOR2x1_ASAP7_75t_R _21919_ (.A(_13541_),
    .B(_13542_),
    .Y(_13543_));
 AO21x1_ASAP7_75t_R _21920_ (.A1(_13543_),
    .A2(_13337_),
    .B(_13045_),
    .Y(_13544_));
 AOI21x1_ASAP7_75t_R _21921_ (.A1(_13061_),
    .A2(_13242_),
    .B(_12996_),
    .Y(_13545_));
 AOI21x1_ASAP7_75t_R _21922_ (.A1(_13001_),
    .A2(_13545_),
    .B(_13007_),
    .Y(_13546_));
 INVx1_ASAP7_75t_R _21923_ (.A(_13272_),
    .Y(_13547_));
 OA21x2_ASAP7_75t_R _21924_ (.A1(_12979_),
    .A2(_12987_),
    .B(_13000_),
    .Y(_13548_));
 OAI21x1_ASAP7_75t_R _21925_ (.A1(_12945_),
    .A2(_13547_),
    .B(_13548_),
    .Y(_13549_));
 NAND2x1_ASAP7_75t_R _21926_ (.A(_13546_),
    .B(_13549_),
    .Y(_13550_));
 AOI21x1_ASAP7_75t_R _21927_ (.A1(net570),
    .A2(_13047_),
    .B(_12927_),
    .Y(_13551_));
 AOI21x1_ASAP7_75t_R _21928_ (.A1(_13211_),
    .A2(_13533_),
    .B(_13551_),
    .Y(_13552_));
 OAI21x1_ASAP7_75t_R _21929_ (.A1(_13051_),
    .A2(_13552_),
    .B(_12908_),
    .Y(_13553_));
 AOI21x1_ASAP7_75t_R _21930_ (.A1(_13544_),
    .A2(_13550_),
    .B(_13553_),
    .Y(_13554_));
 NAND2x1_ASAP7_75t_R _21931_ (.A(_12986_),
    .B(_13211_),
    .Y(_13555_));
 AO21x1_ASAP7_75t_R _21932_ (.A1(_13055_),
    .A2(_13040_),
    .B(_12998_),
    .Y(_13556_));
 AOI21x1_ASAP7_75t_R _21933_ (.A1(_13555_),
    .A2(_13556_),
    .B(_12972_),
    .Y(_13557_));
 AO21x1_ASAP7_75t_R _21934_ (.A1(_13269_),
    .A2(_13259_),
    .B(_12979_),
    .Y(_13558_));
 OA21x2_ASAP7_75t_R _21935_ (.A1(_01181_),
    .A2(_13004_),
    .B(_13044_),
    .Y(_13559_));
 AOI21x1_ASAP7_75t_R _21936_ (.A1(_13558_),
    .A2(_13559_),
    .B(_13446_),
    .Y(_13560_));
 OAI21x1_ASAP7_75t_R _21937_ (.A1(_13557_),
    .A2(_13560_),
    .B(_13067_),
    .Y(_13561_));
 OAI21x1_ASAP7_75t_R _21938_ (.A1(_13387_),
    .A2(_12994_),
    .B(_13001_),
    .Y(_13562_));
 NOR2x1_ASAP7_75t_R _21939_ (.A(_13169_),
    .B(_13280_),
    .Y(_13563_));
 NOR2x1_ASAP7_75t_R _21940_ (.A(_13541_),
    .B(_13563_),
    .Y(_13564_));
 NAND2x1_ASAP7_75t_R _21941_ (.A(_13203_),
    .B(_13564_),
    .Y(_13565_));
 AOI21x1_ASAP7_75t_R _21942_ (.A1(_13562_),
    .A2(_13565_),
    .B(_13045_),
    .Y(_13566_));
 NOR2x1_ASAP7_75t_R _21943_ (.A(_13566_),
    .B(_13561_),
    .Y(_13567_));
 OAI21x1_ASAP7_75t_R _21944_ (.A1(_13554_),
    .A2(_13567_),
    .B(_13021_),
    .Y(_13568_));
 OAI21x1_ASAP7_75t_R _21945_ (.A1(_13021_),
    .A2(_13540_),
    .B(_13568_),
    .Y(_00063_));
 INVx3_ASAP7_75t_R _21946_ (.A(_10676_),
    .Y(_13569_));
 XOR2x1_ASAP7_75t_R _21947_ (.A(_10623_),
    .Y(_13570_),
    .B(_13569_));
 XNOR2x2_ASAP7_75t_R _21948_ (.A(_00803_),
    .B(_00796_),
    .Y(_13571_));
 XOR2x2_ASAP7_75t_R _21949_ (.A(_00829_),
    .B(_10628_),
    .Y(_13572_));
 XOR2x1_ASAP7_75t_R _21950_ (.A(_13571_),
    .Y(_13573_),
    .B(_13572_));
 NOR2x1_ASAP7_75t_R _21951_ (.A(_13570_),
    .B(_13573_),
    .Y(_13574_));
 NOR2x1_ASAP7_75t_R _21952_ (.A(net49),
    .B(net726),
    .Y(_13575_));
 AND2x2_ASAP7_75t_R _21953_ (.A(net49),
    .B(_10653_),
    .Y(_13576_));
 OAI21x1_ASAP7_75t_R _21954_ (.A1(_13575_),
    .A2(_13576_),
    .B(_10676_),
    .Y(_13577_));
 INVx1_ASAP7_75t_R _21955_ (.A(_00764_),
    .Y(_13578_));
 NOR2x1_ASAP7_75t_R _21956_ (.A(net726),
    .B(_13578_),
    .Y(_13579_));
 INVx1_ASAP7_75t_R _21957_ (.A(_10653_),
    .Y(_13580_));
 NOR2x1_ASAP7_75t_R _21958_ (.A(net49),
    .B(_13580_),
    .Y(_13581_));
 OAI21x1_ASAP7_75t_R _21959_ (.A1(_13579_),
    .A2(_13581_),
    .B(_13569_),
    .Y(_13582_));
 NAND2x1_ASAP7_75t_R _21960_ (.A(_13577_),
    .B(_13582_),
    .Y(_13583_));
 XOR2x2_ASAP7_75t_R _21961_ (.A(_10826_),
    .B(_00796_),
    .Y(_13584_));
 XOR2x1_ASAP7_75t_R _21962_ (.A(_13584_),
    .Y(_13585_),
    .B(_13572_));
 OAI21x1_ASAP7_75t_R _21963_ (.A1(_13583_),
    .A2(_13585_),
    .B(_10665_),
    .Y(_13586_));
 NAND2x2_ASAP7_75t_R _21964_ (.A(_00529_),
    .B(_10639_),
    .Y(_13587_));
 OAI21x1_ASAP7_75t_R _21965_ (.A1(_13586_),
    .A2(_13574_),
    .B(_13587_),
    .Y(_13588_));
 XOR2x2_ASAP7_75t_R _21966_ (.A(_07969_),
    .B(net816),
    .Y(_15872_));
 NOR2x2_ASAP7_75t_R _21967_ (.A(_10620_),
    .B(_00530_),
    .Y(_13589_));
 NOR2x2_ASAP7_75t_R _21968_ (.A(_10634_),
    .B(_10825_),
    .Y(_13590_));
 AND2x2_ASAP7_75t_R _21969_ (.A(_10634_),
    .B(_10825_),
    .Y(_13591_));
 OAI21x1_ASAP7_75t_R _21970_ (.A1(_13590_),
    .A2(_13591_),
    .B(net671),
    .Y(_13592_));
 INVx1_ASAP7_75t_R _21971_ (.A(_13592_),
    .Y(_13593_));
 NOR3x1_ASAP7_75t_R _21972_ (.A(_13591_),
    .B(net671),
    .C(_13590_),
    .Y(_13594_));
 OAI21x1_ASAP7_75t_R _21973_ (.A1(_13593_),
    .A2(_13594_),
    .B(net678),
    .Y(_13595_));
 XOR2x1_ASAP7_75t_R _21974_ (.A(net25),
    .Y(_13596_),
    .B(_10825_));
 NAND2x2_ASAP7_75t_R _21975_ (.A(_10652_),
    .B(_13596_),
    .Y(_13597_));
 NAND3x1_ASAP7_75t_R _21976_ (.A(_13597_),
    .B(net724),
    .C(_13592_),
    .Y(_13598_));
 AOI21x1_ASAP7_75t_R _21977_ (.A1(_13595_),
    .A2(_13598_),
    .B(_10640_),
    .Y(_13599_));
 OAI21x1_ASAP7_75t_R _21978_ (.A1(_13589_),
    .A2(_13599_),
    .B(_07958_),
    .Y(_13600_));
 AOI21x1_ASAP7_75t_R _21979_ (.A1(_13592_),
    .A2(_13597_),
    .B(_13571_),
    .Y(_13601_));
 XOR2x1_ASAP7_75t_R _21980_ (.A(_10825_),
    .Y(_13602_),
    .B(net670));
 NAND2x1_ASAP7_75t_R _21981_ (.A(net25),
    .B(_13602_),
    .Y(_13603_));
 INVx1_ASAP7_75t_R _21982_ (.A(net25),
    .Y(_13604_));
 XNOR2x1_ASAP7_75t_R _21983_ (.B(net670),
    .Y(_13605_),
    .A(_10825_));
 NAND2x1_ASAP7_75t_R _21984_ (.A(_13604_),
    .B(_13605_),
    .Y(_13606_));
 AOI21x1_ASAP7_75t_R _21985_ (.A1(_13603_),
    .A2(_13606_),
    .B(net681),
    .Y(_13607_));
 OAI21x1_ASAP7_75t_R _21986_ (.A1(_13607_),
    .A2(_13601_),
    .B(_10621_),
    .Y(_13608_));
 INVx2_ASAP7_75t_R _21987_ (.A(_07958_),
    .Y(_13609_));
 INVx2_ASAP7_75t_R _21988_ (.A(_13589_),
    .Y(_13610_));
 NAND3x2_ASAP7_75t_R _21989_ (.B(_13609_),
    .C(_13610_),
    .Y(_13611_),
    .A(net819));
 NAND2x2_ASAP7_75t_R _21990_ (.A(_13611_),
    .B(_13600_),
    .Y(_13612_));
 BUFx12f_ASAP7_75t_R _21991_ (.A(_13612_),
    .Y(_15874_));
 NOR2x1_ASAP7_75t_R _21992_ (.A(_10741_),
    .B(_00532_),
    .Y(_13613_));
 INVx1_ASAP7_75t_R _21993_ (.A(_13613_),
    .Y(_13614_));
 INVx2_ASAP7_75t_R _21994_ (.A(_10711_),
    .Y(_13615_));
 NOR2x2_ASAP7_75t_R _21995_ (.A(_13615_),
    .B(_10683_),
    .Y(_13616_));
 NOR2x2_ASAP7_75t_R _21996_ (.A(_10711_),
    .B(_10687_),
    .Y(_13617_));
 OAI21x1_ASAP7_75t_R _21997_ (.A1(_13616_),
    .A2(_13617_),
    .B(net583),
    .Y(_13618_));
 INVx1_ASAP7_75t_R _21998_ (.A(_13618_),
    .Y(_13619_));
 NOR3x1_ASAP7_75t_R _21999_ (.A(_13617_),
    .B(_13616_),
    .C(net584),
    .Y(_13620_));
 OAI21x1_ASAP7_75t_R _22000_ (.A1(_13619_),
    .A2(_13620_),
    .B(net780),
    .Y(_13621_));
 INVx1_ASAP7_75t_R _22001_ (.A(_08002_),
    .Y(_13622_));
 AOI21x1_ASAP7_75t_R _22002_ (.A1(_13614_),
    .A2(_13621_),
    .B(_13622_),
    .Y(_13623_));
 BUFx6f_ASAP7_75t_R _22003_ (.A(_13623_),
    .Y(_13624_));
 NAND2x2_ASAP7_75t_R _22004_ (.A(_00532_),
    .B(net866),
    .Y(_13625_));
 NAND2x2_ASAP7_75t_R _22005_ (.A(_13615_),
    .B(_10683_),
    .Y(_13626_));
 INVx1_ASAP7_75t_R _22006_ (.A(net708),
    .Y(_13627_));
 NOR2x1_ASAP7_75t_R _22007_ (.A(_10681_),
    .B(_10682_),
    .Y(_13628_));
 AND2x2_ASAP7_75t_R _22008_ (.A(_10681_),
    .B(_10682_),
    .Y(_13629_));
 OAI21x1_ASAP7_75t_R _22009_ (.A1(_13628_),
    .A2(_13629_),
    .B(_10711_),
    .Y(_13630_));
 NAND3x2_ASAP7_75t_R _22010_ (.B(_13627_),
    .C(_13630_),
    .Y(_13631_),
    .A(_13626_));
 NAND3x2_ASAP7_75t_R _22011_ (.B(net780),
    .C(_13618_),
    .Y(_13632_),
    .A(_13631_));
 AOI21x1_ASAP7_75t_R _22012_ (.A1(_13625_),
    .A2(_13632_),
    .B(_08002_),
    .Y(_13633_));
 BUFx6f_ASAP7_75t_R _22013_ (.A(_13633_),
    .Y(_13634_));
 NOR2x2_ASAP7_75t_R _22014_ (.A(_13624_),
    .B(_13634_),
    .Y(_13635_));
 BUFx12f_ASAP7_75t_R _22015_ (.A(_13635_),
    .Y(_13636_));
 BUFx10_ASAP7_75t_R _22016_ (.A(_13636_),
    .Y(_15882_));
 OAI21x1_ASAP7_75t_R _22017_ (.A1(_13599_),
    .A2(_13589_),
    .B(_13609_),
    .Y(_13637_));
 NAND3x2_ASAP7_75t_R _22018_ (.B(_13608_),
    .C(_13610_),
    .Y(_13638_),
    .A(_07958_));
 NAND2x2_ASAP7_75t_R _22019_ (.A(_13637_),
    .B(_13638_),
    .Y(_13639_));
 BUFx6f_ASAP7_75t_R _22020_ (.A(_13639_),
    .Y(_15869_));
 AOI21x1_ASAP7_75t_R _22021_ (.A1(_13614_),
    .A2(_13621_),
    .B(_08002_),
    .Y(_13640_));
 BUFx6f_ASAP7_75t_R _22022_ (.A(_13640_),
    .Y(_13641_));
 AOI21x1_ASAP7_75t_R _22023_ (.A1(_13625_),
    .A2(_13632_),
    .B(_13622_),
    .Y(_13642_));
 NOR2x2_ASAP7_75t_R _22024_ (.A(_13642_),
    .B(_13641_),
    .Y(_13643_));
 BUFx16f_ASAP7_75t_R _22025_ (.A(_13643_),
    .Y(_13644_));
 BUFx12f_ASAP7_75t_R _22026_ (.A(_13644_),
    .Y(_15879_));
 NAND2x2_ASAP7_75t_R _22027_ (.A(net820),
    .B(_13635_),
    .Y(_13645_));
 NAND2x2_ASAP7_75t_R _22028_ (.A(net723),
    .B(net542),
    .Y(_13646_));
 NOR2x2_ASAP7_75t_R _22029_ (.A(net651),
    .B(_00715_),
    .Y(_13647_));
 NOR2x1_ASAP7_75t_R _22030_ (.A(_10674_),
    .B(_10825_),
    .Y(_13648_));
 AND2x2_ASAP7_75t_R _22031_ (.A(_10674_),
    .B(net726),
    .Y(_13649_));
 OAI21x1_ASAP7_75t_R _22032_ (.A1(_13648_),
    .A2(_13649_),
    .B(_00735_),
    .Y(_13650_));
 NOR2x1_ASAP7_75t_R _22033_ (.A(_10825_),
    .B(_10675_),
    .Y(_13651_));
 NOR2x1_ASAP7_75t_R _22034_ (.A(_10674_),
    .B(_13580_),
    .Y(_13652_));
 INVx1_ASAP7_75t_R _22035_ (.A(_00735_),
    .Y(_13653_));
 OAI21x1_ASAP7_75t_R _22036_ (.A1(_13651_),
    .A2(_13652_),
    .B(_13653_),
    .Y(_13654_));
 NAND2x1_ASAP7_75t_R _22037_ (.A(_13650_),
    .B(_13654_),
    .Y(_13655_));
 XOR2x2_ASAP7_75t_R _22038_ (.A(_10681_),
    .B(net58),
    .Y(_13656_));
 XOR2x1_ASAP7_75t_R _22039_ (.A(_10721_),
    .Y(_13657_),
    .B(_13656_));
 NAND2x1_ASAP7_75t_R _22040_ (.A(_13655_),
    .B(_13657_),
    .Y(_13658_));
 XOR2x1_ASAP7_75t_R _22041_ (.A(_10717_),
    .Y(_13659_),
    .B(_13653_));
 XOR2x1_ASAP7_75t_R _22042_ (.A(_10716_),
    .Y(_13660_),
    .B(_13656_));
 NAND2x1_ASAP7_75t_R _22043_ (.A(_13659_),
    .B(_13660_),
    .Y(_13661_));
 AOI21x1_ASAP7_75t_R _22044_ (.A1(_13658_),
    .A2(_13661_),
    .B(_11441_),
    .Y(_13662_));
 NOR2x1_ASAP7_75t_R _22045_ (.A(_13647_),
    .B(_13662_),
    .Y(_13663_));
 XOR2x2_ASAP7_75t_R _22046_ (.A(_13663_),
    .B(_07942_),
    .Y(_13664_));
 BUFx4f_ASAP7_75t_R _22047_ (.A(_13664_),
    .Y(_13665_));
 AO21x1_ASAP7_75t_R _22048_ (.A1(_13645_),
    .A2(_13646_),
    .B(_13665_),
    .Y(_13666_));
 NAND2x2_ASAP7_75t_R _22049_ (.A(_13664_),
    .B(_13646_),
    .Y(_13667_));
 NOR2x2_ASAP7_75t_R _22050_ (.A(net579),
    .B(_13644_),
    .Y(_13668_));
 AND2x2_ASAP7_75t_R _22051_ (.A(_11374_),
    .B(_00714_),
    .Y(_13669_));
 XOR2x2_ASAP7_75t_R _22052_ (.A(_10714_),
    .B(net58),
    .Y(_13670_));
 INVx2_ASAP7_75t_R _22053_ (.A(_00832_),
    .Y(_13671_));
 XOR2x1_ASAP7_75t_R _22054_ (.A(_13670_),
    .Y(_13672_),
    .B(_13671_));
 XOR2x2_ASAP7_75t_R _22055_ (.A(_10710_),
    .B(_10825_),
    .Y(_13673_));
 XOR2x2_ASAP7_75t_R _22056_ (.A(_10756_),
    .B(_00800_),
    .Y(_13674_));
 XOR2x1_ASAP7_75t_R _22057_ (.A(_13673_),
    .Y(_13675_),
    .B(_13674_));
 NAND2x1_ASAP7_75t_R _22058_ (.A(_13672_),
    .B(_13675_),
    .Y(_13676_));
 XOR2x2_ASAP7_75t_R _22059_ (.A(_13670_),
    .B(_00832_),
    .Y(_13677_));
 XOR2x1_ASAP7_75t_R _22060_ (.A(_10735_),
    .Y(_13678_),
    .B(_13674_));
 NAND2x1_ASAP7_75t_R _22061_ (.A(_13677_),
    .B(_13678_),
    .Y(_13679_));
 AOI21x1_ASAP7_75t_R _22062_ (.A1(_13676_),
    .A2(_13679_),
    .B(_12092_),
    .Y(_13680_));
 OAI21x1_ASAP7_75t_R _22063_ (.A1(_13669_),
    .A2(_13680_),
    .B(_01007_),
    .Y(_13681_));
 NOR2x1_ASAP7_75t_R _22064_ (.A(_10761_),
    .B(_00714_),
    .Y(_13682_));
 XOR2x1_ASAP7_75t_R _22065_ (.A(_13673_),
    .Y(_13683_),
    .B(_10756_));
 XOR2x1_ASAP7_75t_R _22066_ (.A(_10736_),
    .Y(_13684_),
    .B(_13670_));
 NAND2x1_ASAP7_75t_R _22067_ (.A(_13683_),
    .B(_13684_),
    .Y(_13685_));
 XNOR2x1_ASAP7_75t_R _22068_ (.B(_13673_),
    .Y(_13686_),
    .A(_10756_));
 XNOR2x1_ASAP7_75t_R _22069_ (.B(_13670_),
    .Y(_13687_),
    .A(_10736_));
 NAND2x1_ASAP7_75t_R _22070_ (.A(_13686_),
    .B(_13687_),
    .Y(_13688_));
 AOI21x1_ASAP7_75t_R _22071_ (.A1(_13685_),
    .A2(_13688_),
    .B(_11370_),
    .Y(_13689_));
 INVx1_ASAP7_75t_R _22072_ (.A(_01007_),
    .Y(_13690_));
 OAI21x1_ASAP7_75t_R _22073_ (.A1(_13682_),
    .A2(_13689_),
    .B(_13690_),
    .Y(_13691_));
 NAND2x2_ASAP7_75t_R _22074_ (.A(_13681_),
    .B(_13691_),
    .Y(_13692_));
 CKINVDCx6p67_ASAP7_75t_R _22075_ (.A(_13692_),
    .Y(_13693_));
 BUFx10_ASAP7_75t_R _22076_ (.A(_13693_),
    .Y(_13694_));
 OA21x2_ASAP7_75t_R _22077_ (.A1(_13667_),
    .A2(_13668_),
    .B(_13694_),
    .Y(_13695_));
 NAND2x1_ASAP7_75t_R _22078_ (.A(_13666_),
    .B(_13695_),
    .Y(_13696_));
 BUFx4f_ASAP7_75t_R _22079_ (.A(_13664_),
    .Y(_13697_));
 BUFx6f_ASAP7_75t_R _22080_ (.A(_13697_),
    .Y(_13698_));
 OAI21x1_ASAP7_75t_R _22081_ (.A1(_13641_),
    .A2(_13642_),
    .B(_00533_),
    .Y(_13699_));
 OAI21x1_ASAP7_75t_R _22082_ (.A1(_13624_),
    .A2(_13634_),
    .B(_00531_),
    .Y(_13700_));
 NAND2x1_ASAP7_75t_R _22083_ (.A(_13699_),
    .B(_13700_),
    .Y(_13701_));
 AOI21x1_ASAP7_75t_R _22084_ (.A1(_13698_),
    .A2(_13701_),
    .B(_13694_),
    .Y(_13702_));
 INVx1_ASAP7_75t_R _22085_ (.A(_07969_),
    .Y(_13703_));
 XOR2x2_ASAP7_75t_R _22086_ (.A(_13588_),
    .B(_13703_),
    .Y(_13704_));
 BUFx6f_ASAP7_75t_R _22087_ (.A(_13704_),
    .Y(_15870_));
 OAI21x1_ASAP7_75t_R _22088_ (.A1(net61),
    .A2(net60),
    .B(_15882_),
    .Y(_13705_));
 INVx3_ASAP7_75t_R _22089_ (.A(net469),
    .Y(_13706_));
 OAI21x1_ASAP7_75t_R _22090_ (.A1(_13624_),
    .A2(_13634_),
    .B(_13706_),
    .Y(_13707_));
 BUFx3_ASAP7_75t_R _22091_ (.A(_13707_),
    .Y(_13708_));
 AO21x1_ASAP7_75t_R _22092_ (.A1(_13705_),
    .A2(net67),
    .B(_13698_),
    .Y(_13709_));
 NOR2x1_ASAP7_75t_R _22093_ (.A(net641),
    .B(_00713_),
    .Y(_13710_));
 INVx1_ASAP7_75t_R _22094_ (.A(_13710_),
    .Y(_13711_));
 XNOR2x1_ASAP7_75t_R _22095_ (.B(_00768_),
    .Y(_13712_),
    .A(_10783_));
 XOR2x1_ASAP7_75t_R _22096_ (.A(_00800_),
    .Y(_13713_),
    .B(_00801_));
 INVx3_ASAP7_75t_R _22097_ (.A(_10758_),
    .Y(_13714_));
 XOR2x1_ASAP7_75t_R _22098_ (.A(_13713_),
    .Y(_13715_),
    .B(_13714_));
 NOR2x1_ASAP7_75t_R _22099_ (.A(_13712_),
    .B(_13715_),
    .Y(_13716_));
 AND2x2_ASAP7_75t_R _22100_ (.A(_13715_),
    .B(_13712_),
    .Y(_13717_));
 OAI21x1_ASAP7_75t_R _22101_ (.A1(_13716_),
    .A2(_13717_),
    .B(_11450_),
    .Y(_13718_));
 INVx1_ASAP7_75t_R _22102_ (.A(_01008_),
    .Y(_13719_));
 AOI21x1_ASAP7_75t_R _22103_ (.A1(_13711_),
    .A2(_13718_),
    .B(_13719_),
    .Y(_13720_));
 AND3x1_ASAP7_75t_R _22104_ (.A(_13718_),
    .B(_13719_),
    .C(_13711_),
    .Y(_13721_));
 NOR2x2_ASAP7_75t_R _22105_ (.A(_13720_),
    .B(_13721_),
    .Y(_13722_));
 BUFx10_ASAP7_75t_R _22106_ (.A(_13722_),
    .Y(_13723_));
 BUFx10_ASAP7_75t_R _22107_ (.A(_13723_),
    .Y(_13724_));
 AOI21x1_ASAP7_75t_R _22108_ (.A1(_13702_),
    .A2(_13709_),
    .B(_13724_),
    .Y(_13725_));
 NOR2x2_ASAP7_75t_R _22109_ (.A(net525),
    .B(net614),
    .Y(_13726_));
 INVx1_ASAP7_75t_R _22110_ (.A(_07942_),
    .Y(_13727_));
 OAI21x1_ASAP7_75t_R _22111_ (.A1(_13647_),
    .A2(_13662_),
    .B(_13727_),
    .Y(_13728_));
 NOR2x1_ASAP7_75t_R _22112_ (.A(_13655_),
    .B(_13657_),
    .Y(_13729_));
 NOR2x1_ASAP7_75t_R _22113_ (.A(_13659_),
    .B(_13660_),
    .Y(_13730_));
 OAI21x1_ASAP7_75t_R _22114_ (.A1(_13729_),
    .A2(_13730_),
    .B(_10761_),
    .Y(_13731_));
 INVx1_ASAP7_75t_R _22115_ (.A(_13647_),
    .Y(_13732_));
 NAND3x2_ASAP7_75t_R _22116_ (.B(_07942_),
    .C(_13732_),
    .Y(_13733_),
    .A(_13731_));
 NAND2x2_ASAP7_75t_R _22117_ (.A(_13728_),
    .B(_13733_),
    .Y(_13734_));
 BUFx6f_ASAP7_75t_R _22118_ (.A(_13734_),
    .Y(_13735_));
 BUFx6f_ASAP7_75t_R _22119_ (.A(_13735_),
    .Y(_13736_));
 NAND2x1_ASAP7_75t_R _22120_ (.A(net67),
    .B(_13736_),
    .Y(_13737_));
 OAI21x1_ASAP7_75t_R _22121_ (.A1(_13641_),
    .A2(_13642_),
    .B(net471),
    .Y(_13738_));
 BUFx6f_ASAP7_75t_R _22122_ (.A(_13664_),
    .Y(_13739_));
 BUFx6f_ASAP7_75t_R _22123_ (.A(_13692_),
    .Y(_13740_));
 AOI21x1_ASAP7_75t_R _22124_ (.A1(_13738_),
    .A2(_13739_),
    .B(_13740_),
    .Y(_13741_));
 OAI21x1_ASAP7_75t_R _22125_ (.A1(_13726_),
    .A2(_13737_),
    .B(_13741_),
    .Y(_13742_));
 BUFx6f_ASAP7_75t_R _22126_ (.A(_13735_),
    .Y(_13743_));
 AOI21x1_ASAP7_75t_R _22127_ (.A1(_13699_),
    .A2(net67),
    .B(_13743_),
    .Y(_13744_));
 OAI21x1_ASAP7_75t_R _22128_ (.A1(_13641_),
    .A2(_13642_),
    .B(_00531_),
    .Y(_13745_));
 BUFx6f_ASAP7_75t_R _22129_ (.A(_13745_),
    .Y(_13746_));
 OAI21x1_ASAP7_75t_R _22130_ (.A1(_13624_),
    .A2(_13634_),
    .B(_00533_),
    .Y(_13747_));
 BUFx6f_ASAP7_75t_R _22131_ (.A(_13664_),
    .Y(_13748_));
 BUFx6f_ASAP7_75t_R _22132_ (.A(_13748_),
    .Y(_13749_));
 AOI21x1_ASAP7_75t_R _22133_ (.A1(_13746_),
    .A2(_13747_),
    .B(_13749_),
    .Y(_13750_));
 BUFx6f_ASAP7_75t_R _22134_ (.A(_13692_),
    .Y(_13751_));
 BUFx10_ASAP7_75t_R _22135_ (.A(_13751_),
    .Y(_13752_));
 OAI21x1_ASAP7_75t_R _22136_ (.A1(_13744_),
    .A2(_13750_),
    .B(_13752_),
    .Y(_13753_));
 INVx4_ASAP7_75t_R _22137_ (.A(_13722_),
    .Y(_13754_));
 BUFx6f_ASAP7_75t_R _22138_ (.A(_13754_),
    .Y(_13755_));
 BUFx10_ASAP7_75t_R _22139_ (.A(_13755_),
    .Y(_13756_));
 AOI21x1_ASAP7_75t_R _22140_ (.A1(_13742_),
    .A2(_13753_),
    .B(_13756_),
    .Y(_13757_));
 XOR2x2_ASAP7_75t_R _22141_ (.A(_00802_),
    .B(_00834_),
    .Y(_13758_));
 XOR2x1_ASAP7_75t_R _22142_ (.A(_10755_),
    .Y(_13759_),
    .B(_00738_));
 XNOR2x1_ASAP7_75t_R _22143_ (.B(_13759_),
    .Y(_13760_),
    .A(_13758_));
 NOR2x1_ASAP7_75t_R _22144_ (.A(_10734_),
    .B(_00712_),
    .Y(_13761_));
 AO21x1_ASAP7_75t_R _22145_ (.A1(_13760_),
    .A2(_10829_),
    .B(_13761_),
    .Y(_13762_));
 XNOR2x2_ASAP7_75t_R _22146_ (.A(_01009_),
    .B(_13762_),
    .Y(_13763_));
 BUFx10_ASAP7_75t_R _22147_ (.A(_13763_),
    .Y(_13764_));
 AOI211x1_ASAP7_75t_R _22148_ (.A1(_13696_),
    .A2(_13725_),
    .B(_13757_),
    .C(_13764_),
    .Y(_13765_));
 INVx2_ASAP7_75t_R _22149_ (.A(_01186_),
    .Y(_13766_));
 NAND2x2_ASAP7_75t_R _22150_ (.A(_13766_),
    .B(_13644_),
    .Y(_13767_));
 AOI21x1_ASAP7_75t_R _22151_ (.A1(_13767_),
    .A2(_13645_),
    .B(_13743_),
    .Y(_13768_));
 AOI21x1_ASAP7_75t_R _22152_ (.A1(_13570_),
    .A2(net725),
    .B(_12161_),
    .Y(_13769_));
 INVx1_ASAP7_75t_R _22153_ (.A(_13574_),
    .Y(_13770_));
 NAND2x1_ASAP7_75t_R _22154_ (.A(_13769_),
    .B(_13770_),
    .Y(_13771_));
 AOI21x1_ASAP7_75t_R _22155_ (.A1(_13587_),
    .A2(_13771_),
    .B(_07969_),
    .Y(_13772_));
 NOR2x1_ASAP7_75t_R _22156_ (.A(_13703_),
    .B(_13588_),
    .Y(_13773_));
 OAI22x1_ASAP7_75t_R _22157_ (.A1(_13634_),
    .A2(_13624_),
    .B1(_13772_),
    .B2(_13773_),
    .Y(_13774_));
 OAI21x1_ASAP7_75t_R _22158_ (.A1(net63),
    .A2(_15874_),
    .B(_13636_),
    .Y(_13775_));
 AOI21x1_ASAP7_75t_R _22159_ (.A1(_13774_),
    .A2(_13775_),
    .B(_13749_),
    .Y(_13776_));
 BUFx6f_ASAP7_75t_R _22160_ (.A(_13693_),
    .Y(_13777_));
 BUFx10_ASAP7_75t_R _22161_ (.A(_13777_),
    .Y(_13778_));
 OAI21x1_ASAP7_75t_R _22162_ (.A1(_13768_),
    .A2(_13776_),
    .B(_13778_),
    .Y(_13779_));
 INVx1_ASAP7_75t_R _22163_ (.A(_01183_),
    .Y(_13780_));
 OAI21x1_ASAP7_75t_R _22164_ (.A1(_13624_),
    .A2(_13634_),
    .B(_13780_),
    .Y(_13781_));
 NAND2x2_ASAP7_75t_R _22165_ (.A(net525),
    .B(_13635_),
    .Y(_13782_));
 AOI21x1_ASAP7_75t_R _22166_ (.A1(_13781_),
    .A2(_13782_),
    .B(_13749_),
    .Y(_13783_));
 OAI21x1_ASAP7_75t_R _22167_ (.A1(net63),
    .A2(net62),
    .B(net614),
    .Y(_13784_));
 BUFx10_ASAP7_75t_R _22168_ (.A(_13734_),
    .Y(_13785_));
 AOI21x1_ASAP7_75t_R _22169_ (.A1(_13645_),
    .A2(_13784_),
    .B(_13785_),
    .Y(_13786_));
 OAI21x1_ASAP7_75t_R _22170_ (.A1(_13783_),
    .A2(_13786_),
    .B(_13752_),
    .Y(_13787_));
 AOI21x1_ASAP7_75t_R _22171_ (.A1(_13779_),
    .A2(_13787_),
    .B(_13756_),
    .Y(_13788_));
 NOR2x2_ASAP7_75t_R _22172_ (.A(_15874_),
    .B(_13644_),
    .Y(_13789_));
 BUFx10_ASAP7_75t_R _22173_ (.A(_13692_),
    .Y(_13790_));
 OAI21x1_ASAP7_75t_R _22174_ (.A1(_13698_),
    .A2(_13789_),
    .B(_13790_),
    .Y(_13791_));
 BUFx5_ASAP7_75t_R _22175_ (.A(_01184_),
    .Y(_13792_));
 INVx4_ASAP7_75t_R _22176_ (.A(_13792_),
    .Y(_13793_));
 NAND2x2_ASAP7_75t_R _22177_ (.A(_13793_),
    .B(net614),
    .Y(_13794_));
 AOI21x1_ASAP7_75t_R _22178_ (.A1(_13794_),
    .A2(_13775_),
    .B(_13743_),
    .Y(_13795_));
 BUFx10_ASAP7_75t_R _22179_ (.A(_13754_),
    .Y(_13796_));
 OAI21x1_ASAP7_75t_R _22180_ (.A1(_13791_),
    .A2(_13795_),
    .B(_13796_),
    .Y(_13797_));
 BUFx6f_ASAP7_75t_R _22181_ (.A(_13785_),
    .Y(_13798_));
 BUFx6f_ASAP7_75t_R _22182_ (.A(net614),
    .Y(_13799_));
 OAI21x1_ASAP7_75t_R _22183_ (.A1(net69),
    .A2(_13799_),
    .B(net60),
    .Y(_13800_));
 AOI21x1_ASAP7_75t_R _22184_ (.A1(_13798_),
    .A2(_13800_),
    .B(_13751_),
    .Y(_13801_));
 OAI21x1_ASAP7_75t_R _22185_ (.A1(_13641_),
    .A2(_13642_),
    .B(_13766_),
    .Y(_13802_));
 BUFx6f_ASAP7_75t_R _22186_ (.A(_13802_),
    .Y(_13803_));
 BUFx6f_ASAP7_75t_R _22187_ (.A(_13734_),
    .Y(_13804_));
 AO21x1_ASAP7_75t_R _22188_ (.A1(_13803_),
    .A2(_13708_),
    .B(_13804_),
    .Y(_13805_));
 AND2x2_ASAP7_75t_R _22189_ (.A(_13801_),
    .B(_13805_),
    .Y(_13806_));
 OAI21x1_ASAP7_75t_R _22190_ (.A1(_13806_),
    .A2(_13797_),
    .B(_13764_),
    .Y(_13807_));
 XOR2x1_ASAP7_75t_R _22191_ (.A(_00802_),
    .Y(_13808_),
    .B(net58));
 XOR2x1_ASAP7_75t_R _22192_ (.A(_13808_),
    .Y(_13809_),
    .B(_10823_));
 XOR2x1_ASAP7_75t_R _22193_ (.A(net50),
    .Y(_13810_),
    .B(_00770_));
 XOR2x1_ASAP7_75t_R _22194_ (.A(_13809_),
    .Y(_13811_),
    .B(_13810_));
 NOR2x1_ASAP7_75t_R _22195_ (.A(_13017_),
    .B(_00711_),
    .Y(_13812_));
 AO21x1_ASAP7_75t_R _22196_ (.A1(_13811_),
    .A2(_10831_),
    .B(_13812_),
    .Y(_13813_));
 XOR2x2_ASAP7_75t_R _22197_ (.A(_13813_),
    .B(_01010_),
    .Y(_13814_));
 OAI21x1_ASAP7_75t_R _22198_ (.A1(_13807_),
    .A2(_13788_),
    .B(_13814_),
    .Y(_13815_));
 OAI21x1_ASAP7_75t_R _22199_ (.A1(_13641_),
    .A2(_13642_),
    .B(_13706_),
    .Y(_13816_));
 INVx2_ASAP7_75t_R _22200_ (.A(_13816_),
    .Y(_13817_));
 AOI21x1_ASAP7_75t_R _22201_ (.A1(_13736_),
    .A2(_13817_),
    .B(_13751_),
    .Y(_13818_));
 INVx1_ASAP7_75t_R _22202_ (.A(_01188_),
    .Y(_13819_));
 BUFx6f_ASAP7_75t_R _22203_ (.A(_13748_),
    .Y(_13820_));
 NAND2x1_ASAP7_75t_R _22204_ (.A(_13819_),
    .B(_13820_),
    .Y(_13821_));
 AO21x1_ASAP7_75t_R _22205_ (.A1(_13818_),
    .A2(_13821_),
    .B(_13763_),
    .Y(_13822_));
 BUFx10_ASAP7_75t_R _22206_ (.A(_13664_),
    .Y(_13823_));
 OAI21x1_ASAP7_75t_R _22207_ (.A1(_13641_),
    .A2(_13642_),
    .B(_13793_),
    .Y(_13824_));
 INVx1_ASAP7_75t_R _22208_ (.A(_13824_),
    .Y(_13825_));
 AOI21x1_ASAP7_75t_R _22209_ (.A1(_13799_),
    .A2(_13646_),
    .B(_13825_),
    .Y(_13826_));
 NOR2x2_ASAP7_75t_R _22210_ (.A(_13826_),
    .B(_13823_),
    .Y(_13827_));
 OAI21x1_ASAP7_75t_R _22211_ (.A1(_15869_),
    .A2(_13799_),
    .B(_13747_),
    .Y(_13828_));
 INVx1_ASAP7_75t_R _22212_ (.A(_13828_),
    .Y(_13829_));
 OAI21x1_ASAP7_75t_R _22213_ (.A1(_13641_),
    .A2(_13642_),
    .B(_13780_),
    .Y(_13830_));
 INVx1_ASAP7_75t_R _22214_ (.A(_13830_),
    .Y(_13831_));
 BUFx6f_ASAP7_75t_R _22215_ (.A(_13693_),
    .Y(_13832_));
 AOI21x1_ASAP7_75t_R _22216_ (.A1(_13804_),
    .A2(_13831_),
    .B(_13832_),
    .Y(_13833_));
 OAI21x1_ASAP7_75t_R _22217_ (.A1(_13743_),
    .A2(_13829_),
    .B(_13833_),
    .Y(_13834_));
 NOR2x1_ASAP7_75t_R _22218_ (.A(_13834_),
    .B(_13827_),
    .Y(_13835_));
 OAI21x1_ASAP7_75t_R _22219_ (.A1(_13822_),
    .A2(_13835_),
    .B(_13724_),
    .Y(_13836_));
 OA21x2_ASAP7_75t_R _22220_ (.A1(_13748_),
    .A2(_13824_),
    .B(_13693_),
    .Y(_13837_));
 INVx2_ASAP7_75t_R _22221_ (.A(_01185_),
    .Y(_13838_));
 OAI21x1_ASAP7_75t_R _22222_ (.A1(_13624_),
    .A2(_13634_),
    .B(_13838_),
    .Y(_13839_));
 NOR2x2_ASAP7_75t_R _22223_ (.A(_13839_),
    .B(_13748_),
    .Y(_13840_));
 OAI21x1_ASAP7_75t_R _22224_ (.A1(_13624_),
    .A2(_13634_),
    .B(net470),
    .Y(_13841_));
 INVx2_ASAP7_75t_R _22225_ (.A(_13841_),
    .Y(_13842_));
 NOR2x2_ASAP7_75t_R _22226_ (.A(_13734_),
    .B(_13842_),
    .Y(_13843_));
 NOR2x1_ASAP7_75t_R _22227_ (.A(_13840_),
    .B(_13843_),
    .Y(_13844_));
 OAI21x1_ASAP7_75t_R _22228_ (.A1(_13824_),
    .A2(_13748_),
    .B(_13692_),
    .Y(_13845_));
 NOR2x1_ASAP7_75t_R _22229_ (.A(_13845_),
    .B(_13786_),
    .Y(_13846_));
 CKINVDCx8_ASAP7_75t_R _22230_ (.A(_13763_),
    .Y(_13847_));
 BUFx10_ASAP7_75t_R _22231_ (.A(_13847_),
    .Y(_13848_));
 AOI211x1_ASAP7_75t_R _22232_ (.A1(_13837_),
    .A2(_13844_),
    .B(_13846_),
    .C(_13848_),
    .Y(_13849_));
 INVx8_ASAP7_75t_R _22233_ (.A(_13814_),
    .Y(_13850_));
 OAI21x1_ASAP7_75t_R _22234_ (.A1(_13836_),
    .A2(_13849_),
    .B(_13850_),
    .Y(_13851_));
 OAI21x1_ASAP7_75t_R _22235_ (.A1(_13634_),
    .A2(_13624_),
    .B(net820),
    .Y(_13852_));
 AOI21x1_ASAP7_75t_R _22236_ (.A1(_13746_),
    .A2(_13852_),
    .B(_13736_),
    .Y(_13853_));
 OAI21x1_ASAP7_75t_R _22237_ (.A1(net61),
    .A2(_15882_),
    .B(net6),
    .Y(_13854_));
 NOR2x1_ASAP7_75t_R _22238_ (.A(_13749_),
    .B(_13854_),
    .Y(_13855_));
 BUFx6f_ASAP7_75t_R _22239_ (.A(_13740_),
    .Y(_13856_));
 OAI21x1_ASAP7_75t_R _22240_ (.A1(_13853_),
    .A2(_13855_),
    .B(_13856_),
    .Y(_13857_));
 AO21x1_ASAP7_75t_R _22241_ (.A1(_13781_),
    .A2(_13699_),
    .B(_13739_),
    .Y(_13858_));
 BUFx4f_ASAP7_75t_R _22242_ (.A(_13734_),
    .Y(_13859_));
 AOI21x1_ASAP7_75t_R _22243_ (.A1(_13792_),
    .A2(_15879_),
    .B(_13859_),
    .Y(_13860_));
 INVx1_ASAP7_75t_R _22244_ (.A(_13860_),
    .Y(_13861_));
 AO21x1_ASAP7_75t_R _22245_ (.A1(_13858_),
    .A2(_13861_),
    .B(_13856_),
    .Y(_13862_));
 AOI21x1_ASAP7_75t_R _22246_ (.A1(_13857_),
    .A2(_13862_),
    .B(_13847_),
    .Y(_13863_));
 OAI21x1_ASAP7_75t_R _22247_ (.A1(_13781_),
    .A2(_13785_),
    .B(_13693_),
    .Y(_13864_));
 OAI21x1_ASAP7_75t_R _22248_ (.A1(_15870_),
    .A2(_15874_),
    .B(_13799_),
    .Y(_13865_));
 AOI21x1_ASAP7_75t_R _22249_ (.A1(_13746_),
    .A2(_13865_),
    .B(_13749_),
    .Y(_13866_));
 OAI21x1_ASAP7_75t_R _22250_ (.A1(_13864_),
    .A2(_13866_),
    .B(_13847_),
    .Y(_13867_));
 NOR2x2_ASAP7_75t_R _22251_ (.A(net820),
    .B(net63),
    .Y(_13868_));
 NAND2x2_ASAP7_75t_R _22252_ (.A(_13644_),
    .B(_13868_),
    .Y(_13869_));
 AOI21x1_ASAP7_75t_R _22253_ (.A1(_01185_),
    .A2(_15882_),
    .B(_13735_),
    .Y(_13870_));
 NOR2x2_ASAP7_75t_R _22254_ (.A(_13781_),
    .B(_13664_),
    .Y(_13871_));
 AOI211x1_ASAP7_75t_R _22255_ (.A1(_13869_),
    .A2(_13870_),
    .B(_13871_),
    .C(_13694_),
    .Y(_13872_));
 OAI21x1_ASAP7_75t_R _22256_ (.A1(_13867_),
    .A2(_13872_),
    .B(_13756_),
    .Y(_13873_));
 NOR2x1_ASAP7_75t_R _22257_ (.A(_13863_),
    .B(_13873_),
    .Y(_13874_));
 OAI22x1_ASAP7_75t_R _22258_ (.A1(_13815_),
    .A2(_13765_),
    .B1(_13851_),
    .B2(_13874_),
    .Y(_00064_));
 NOR2x1_ASAP7_75t_R _22259_ (.A(net815),
    .B(_13636_),
    .Y(_13875_));
 OAI21x1_ASAP7_75t_R _22260_ (.A1(_13875_),
    .A2(_13817_),
    .B(_13739_),
    .Y(_13876_));
 NAND2x1_ASAP7_75t_R _22261_ (.A(_13751_),
    .B(_13876_),
    .Y(_13877_));
 BUFx6f_ASAP7_75t_R _22262_ (.A(_13664_),
    .Y(_13878_));
 NAND2x2_ASAP7_75t_R _22263_ (.A(_15872_),
    .B(_13635_),
    .Y(_13879_));
 NOR2x2_ASAP7_75t_R _22264_ (.A(net812),
    .B(_13635_),
    .Y(_13880_));
 AOI21x1_ASAP7_75t_R _22265_ (.A1(_13878_),
    .A2(_13879_),
    .B(_13880_),
    .Y(_13881_));
 AOI21x1_ASAP7_75t_R _22266_ (.A1(_13881_),
    .A2(_13837_),
    .B(_13755_),
    .Y(_13882_));
 OAI21x1_ASAP7_75t_R _22267_ (.A1(_13827_),
    .A2(_13877_),
    .B(_13882_),
    .Y(_13883_));
 NAND2x2_ASAP7_75t_R _22268_ (.A(net62),
    .B(_13636_),
    .Y(_13884_));
 AO21x1_ASAP7_75t_R _22269_ (.A1(_13884_),
    .A2(_13794_),
    .B(_13665_),
    .Y(_13885_));
 AOI21x1_ASAP7_75t_R _22270_ (.A1(_13884_),
    .A2(_13843_),
    .B(_13740_),
    .Y(_13886_));
 NAND2x1_ASAP7_75t_R _22271_ (.A(_13885_),
    .B(_13886_),
    .Y(_13887_));
 NOR2x2_ASAP7_75t_R _22272_ (.A(_15869_),
    .B(net540),
    .Y(_13888_));
 OAI21x1_ASAP7_75t_R _22273_ (.A1(_13888_),
    .A2(_13726_),
    .B(_13804_),
    .Y(_13889_));
 NOR2x2_ASAP7_75t_R _22274_ (.A(_13644_),
    .B(_13785_),
    .Y(_13890_));
 AOI21x1_ASAP7_75t_R _22275_ (.A1(_13646_),
    .A2(_13890_),
    .B(_13832_),
    .Y(_13891_));
 AOI21x1_ASAP7_75t_R _22276_ (.A1(_13889_),
    .A2(_13891_),
    .B(_13723_),
    .Y(_13892_));
 NAND2x1_ASAP7_75t_R _22277_ (.A(_13887_),
    .B(_13892_),
    .Y(_13893_));
 AOI21x1_ASAP7_75t_R _22278_ (.A1(_13883_),
    .A2(_13893_),
    .B(_13763_),
    .Y(_13894_));
 BUFx6f_ASAP7_75t_R _22279_ (.A(_13841_),
    .Y(_13895_));
 AO21x1_ASAP7_75t_R _22280_ (.A1(_13824_),
    .A2(net727),
    .B(_13859_),
    .Y(_13896_));
 INVx2_ASAP7_75t_R _22281_ (.A(_13747_),
    .Y(_13897_));
 BUFx10_ASAP7_75t_R _22282_ (.A(_13785_),
    .Y(_13898_));
 OAI21x1_ASAP7_75t_R _22283_ (.A1(_13897_),
    .A2(_13668_),
    .B(_13898_),
    .Y(_13899_));
 AOI21x1_ASAP7_75t_R _22284_ (.A1(_13896_),
    .A2(_13899_),
    .B(_13790_),
    .Y(_13900_));
 NOR2x2_ASAP7_75t_R _22285_ (.A(net578),
    .B(net63),
    .Y(_13901_));
 NOR2x2_ASAP7_75t_R _22286_ (.A(_15874_),
    .B(_13636_),
    .Y(_13902_));
 OAI21x1_ASAP7_75t_R _22287_ (.A1(_13901_),
    .A2(_13902_),
    .B(_13823_),
    .Y(_13903_));
 INVx3_ASAP7_75t_R _22288_ (.A(_13738_),
    .Y(_13904_));
 NOR2x2_ASAP7_75t_R _22289_ (.A(net579),
    .B(_13635_),
    .Y(_13905_));
 OAI21x1_ASAP7_75t_R _22290_ (.A1(_13904_),
    .A2(_13905_),
    .B(_13898_),
    .Y(_13906_));
 BUFx6f_ASAP7_75t_R _22291_ (.A(_13693_),
    .Y(_13907_));
 AOI21x1_ASAP7_75t_R _22292_ (.A1(_13903_),
    .A2(_13906_),
    .B(_13907_),
    .Y(_13908_));
 OAI21x1_ASAP7_75t_R _22293_ (.A1(_13900_),
    .A2(_13908_),
    .B(_13724_),
    .Y(_13909_));
 NAND2x2_ASAP7_75t_R _22294_ (.A(net62),
    .B(_13644_),
    .Y(_13910_));
 NAND2x2_ASAP7_75t_R _22295_ (.A(net526),
    .B(net614),
    .Y(_13911_));
 AO21x1_ASAP7_75t_R _22296_ (.A1(_13910_),
    .A2(_13911_),
    .B(_13665_),
    .Y(_13912_));
 AOI21x1_ASAP7_75t_R _22297_ (.A1(_01186_),
    .A2(_13636_),
    .B(_13785_),
    .Y(_13913_));
 AOI21x1_ASAP7_75t_R _22298_ (.A1(_13911_),
    .A2(_13913_),
    .B(_13740_),
    .Y(_13914_));
 NAND2x1_ASAP7_75t_R _22299_ (.A(_13912_),
    .B(_13914_),
    .Y(_13915_));
 NOR2x1_ASAP7_75t_R _22300_ (.A(_13792_),
    .B(_13636_),
    .Y(_13916_));
 AOI21x1_ASAP7_75t_R _22301_ (.A1(_13798_),
    .A2(_13916_),
    .B(_13832_),
    .Y(_13917_));
 AOI21x1_ASAP7_75t_R _22302_ (.A1(net69),
    .A2(_15874_),
    .B(_13799_),
    .Y(_13918_));
 OAI21x1_ASAP7_75t_R _22303_ (.A1(_13842_),
    .A2(_13918_),
    .B(_13739_),
    .Y(_13919_));
 AOI21x1_ASAP7_75t_R _22304_ (.A1(_13917_),
    .A2(_13919_),
    .B(_13723_),
    .Y(_13920_));
 NAND2x1_ASAP7_75t_R _22305_ (.A(_13915_),
    .B(_13920_),
    .Y(_13921_));
 AOI21x1_ASAP7_75t_R _22306_ (.A1(_13909_),
    .A2(_13921_),
    .B(_13848_),
    .Y(_13922_));
 OAI21x1_ASAP7_75t_R _22307_ (.A1(_13894_),
    .A2(_13922_),
    .B(_13850_),
    .Y(_13923_));
 AO21x1_ASAP7_75t_R _22308_ (.A1(_13784_),
    .A2(_13775_),
    .B(_13798_),
    .Y(_13924_));
 AO21x1_ASAP7_75t_R _22309_ (.A1(_13852_),
    .A2(_13699_),
    .B(_13878_),
    .Y(_13925_));
 BUFx6f_ASAP7_75t_R _22310_ (.A(_13722_),
    .Y(_13926_));
 AO21x1_ASAP7_75t_R _22311_ (.A1(_13924_),
    .A2(_13925_),
    .B(_13926_),
    .Y(_13927_));
 OAI21x1_ASAP7_75t_R _22312_ (.A1(_13726_),
    .A2(_13916_),
    .B(_13739_),
    .Y(_13928_));
 AOI21x1_ASAP7_75t_R _22313_ (.A1(_13910_),
    .A2(_13782_),
    .B(_13748_),
    .Y(_13929_));
 INVx1_ASAP7_75t_R _22314_ (.A(_13929_),
    .Y(_13930_));
 NAND2x1_ASAP7_75t_R _22315_ (.A(_13928_),
    .B(_13930_),
    .Y(_13931_));
 AOI21x1_ASAP7_75t_R _22316_ (.A1(_13724_),
    .A2(_13931_),
    .B(_13856_),
    .Y(_13932_));
 AO21x2_ASAP7_75t_R _22317_ (.A1(_13784_),
    .A2(_13746_),
    .B(_13748_),
    .Y(_13933_));
 INVx1_ASAP7_75t_R _22318_ (.A(_00535_),
    .Y(_13934_));
 NOR2x1_ASAP7_75t_R _22319_ (.A(_13934_),
    .B(_13859_),
    .Y(_13935_));
 AOI21x1_ASAP7_75t_R _22320_ (.A1(_13723_),
    .A2(_13935_),
    .B(_13907_),
    .Y(_13936_));
 AO21x1_ASAP7_75t_R _22321_ (.A1(_13933_),
    .A2(_13936_),
    .B(_13763_),
    .Y(_13937_));
 AOI21x1_ASAP7_75t_R _22322_ (.A1(_13927_),
    .A2(_13932_),
    .B(_13937_),
    .Y(_13938_));
 AO21x1_ASAP7_75t_R _22323_ (.A1(_13816_),
    .A2(_13747_),
    .B(_13804_),
    .Y(_13939_));
 INVx1_ASAP7_75t_R _22324_ (.A(_13781_),
    .Y(_13940_));
 OAI21x1_ASAP7_75t_R _22325_ (.A1(_13940_),
    .A2(_13668_),
    .B(_13898_),
    .Y(_13941_));
 AOI21x1_ASAP7_75t_R _22326_ (.A1(_13939_),
    .A2(_13941_),
    .B(_13790_),
    .Y(_13942_));
 INVx2_ASAP7_75t_R _22327_ (.A(_13699_),
    .Y(_13943_));
 OAI21x1_ASAP7_75t_R _22328_ (.A1(_13943_),
    .A2(_13902_),
    .B(_13898_),
    .Y(_13944_));
 AOI21x1_ASAP7_75t_R _22329_ (.A1(_13944_),
    .A2(_13928_),
    .B(_13694_),
    .Y(_13945_));
 OAI21x1_ASAP7_75t_R _22330_ (.A1(_13942_),
    .A2(_13945_),
    .B(_13796_),
    .Y(_13946_));
 OAI21x1_ASAP7_75t_R _22331_ (.A1(net814),
    .A2(_15882_),
    .B(_13830_),
    .Y(_13947_));
 AOI21x1_ASAP7_75t_R _22332_ (.A1(_13798_),
    .A2(_13947_),
    .B(_13751_),
    .Y(_13948_));
 AOI21x1_ASAP7_75t_R _22333_ (.A1(_13919_),
    .A2(_13948_),
    .B(_13755_),
    .Y(_13949_));
 NAND2x1_ASAP7_75t_R _22334_ (.A(_13799_),
    .B(_13901_),
    .Y(_13950_));
 AOI21x1_ASAP7_75t_R _22335_ (.A1(net60),
    .A2(_15882_),
    .B(_13665_),
    .Y(_13951_));
 AOI21x1_ASAP7_75t_R _22336_ (.A1(_13950_),
    .A2(_13951_),
    .B(_13843_),
    .Y(_13952_));
 NAND2x1_ASAP7_75t_R _22337_ (.A(_13790_),
    .B(_13952_),
    .Y(_13953_));
 NAND2x1_ASAP7_75t_R _22338_ (.A(_13949_),
    .B(_13953_),
    .Y(_13954_));
 AOI21x1_ASAP7_75t_R _22339_ (.A1(_13946_),
    .A2(_13954_),
    .B(_13848_),
    .Y(_13955_));
 OAI21x1_ASAP7_75t_R _22340_ (.A1(_13938_),
    .A2(_13955_),
    .B(_13814_),
    .Y(_13956_));
 NAND2x1_ASAP7_75t_R _22341_ (.A(_13923_),
    .B(_13956_),
    .Y(_00065_));
 AOI21x1_ASAP7_75t_R _22342_ (.A1(_13803_),
    .A2(_13794_),
    .B(_13820_),
    .Y(_13957_));
 BUFx6f_ASAP7_75t_R _22343_ (.A(_13785_),
    .Y(_13958_));
 AOI21x1_ASAP7_75t_R _22344_ (.A1(_15874_),
    .A2(_15882_),
    .B(net61),
    .Y(_13959_));
 NOR2x1_ASAP7_75t_R _22345_ (.A(_13958_),
    .B(_13959_),
    .Y(_13960_));
 OAI21x1_ASAP7_75t_R _22346_ (.A1(_13957_),
    .A2(_13960_),
    .B(_13778_),
    .Y(_13961_));
 AOI21x1_ASAP7_75t_R _22347_ (.A1(net6),
    .A2(_13774_),
    .B(_13698_),
    .Y(_13962_));
 AOI21x1_ASAP7_75t_R _22348_ (.A1(net813),
    .A2(_13865_),
    .B(_13743_),
    .Y(_13963_));
 OAI21x1_ASAP7_75t_R _22349_ (.A1(_13962_),
    .A2(_13963_),
    .B(_13752_),
    .Y(_13964_));
 AOI21x1_ASAP7_75t_R _22350_ (.A1(_13961_),
    .A2(_13964_),
    .B(_13756_),
    .Y(_13965_));
 NAND3x1_ASAP7_75t_R _22351_ (.A(_13852_),
    .B(_13749_),
    .C(_13830_),
    .Y(_13966_));
 AO21x1_ASAP7_75t_R _22352_ (.A1(_13879_),
    .A2(net727),
    .B(_13665_),
    .Y(_13967_));
 AOI21x1_ASAP7_75t_R _22353_ (.A1(_13966_),
    .A2(_13967_),
    .B(_13752_),
    .Y(_13968_));
 AOI21x1_ASAP7_75t_R _22354_ (.A1(_13767_),
    .A2(_13705_),
    .B(_13743_),
    .Y(_13969_));
 OAI21x1_ASAP7_75t_R _22355_ (.A1(_15879_),
    .A2(_13646_),
    .B(_13898_),
    .Y(_13970_));
 NAND2x1_ASAP7_75t_R _22356_ (.A(_13790_),
    .B(_13970_),
    .Y(_13971_));
 OAI21x1_ASAP7_75t_R _22357_ (.A1(_13969_),
    .A2(_13971_),
    .B(_13796_),
    .Y(_13972_));
 OAI21x1_ASAP7_75t_R _22358_ (.A1(_13968_),
    .A2(_13972_),
    .B(_13848_),
    .Y(_13973_));
 OAI21x1_ASAP7_75t_R _22359_ (.A1(_13965_),
    .A2(_13973_),
    .B(_13814_),
    .Y(_13974_));
 AOI21x1_ASAP7_75t_R _22360_ (.A1(_13738_),
    .A2(net67),
    .B(_13736_),
    .Y(_13975_));
 OAI21x1_ASAP7_75t_R _22361_ (.A1(_13641_),
    .A2(_13642_),
    .B(_13838_),
    .Y(_13976_));
 AOI21x1_ASAP7_75t_R _22362_ (.A1(_13976_),
    .A2(_13852_),
    .B(_13748_),
    .Y(_13977_));
 OAI21x1_ASAP7_75t_R _22363_ (.A1(_13975_),
    .A2(_13977_),
    .B(_13856_),
    .Y(_13978_));
 AOI21x1_ASAP7_75t_R _22364_ (.A1(_13803_),
    .A2(_13852_),
    .B(_13749_),
    .Y(_13979_));
 AOI21x1_ASAP7_75t_R _22365_ (.A1(_13839_),
    .A2(_13782_),
    .B(_13736_),
    .Y(_13980_));
 OAI21x1_ASAP7_75t_R _22366_ (.A1(_13979_),
    .A2(_13980_),
    .B(_13694_),
    .Y(_13981_));
 AOI21x1_ASAP7_75t_R _22367_ (.A1(_13978_),
    .A2(_13981_),
    .B(_13724_),
    .Y(_13982_));
 AOI21x1_ASAP7_75t_R _22368_ (.A1(_13839_),
    .A2(_13803_),
    .B(_13820_),
    .Y(_13983_));
 AOI21x1_ASAP7_75t_R _22369_ (.A1(net813),
    .A2(_13852_),
    .B(_13736_),
    .Y(_13984_));
 OAI21x1_ASAP7_75t_R _22370_ (.A1(_13983_),
    .A2(_13984_),
    .B(_13694_),
    .Y(_13985_));
 AOI21x1_ASAP7_75t_R _22371_ (.A1(net813),
    .A2(_13839_),
    .B(_13820_),
    .Y(_13986_));
 AOI21x1_ASAP7_75t_R _22372_ (.A1(net813),
    .A2(_13774_),
    .B(_13736_),
    .Y(_13987_));
 OAI21x1_ASAP7_75t_R _22373_ (.A1(_13986_),
    .A2(_13987_),
    .B(_13856_),
    .Y(_13988_));
 AOI21x1_ASAP7_75t_R _22374_ (.A1(_13985_),
    .A2(_13988_),
    .B(_13796_),
    .Y(_13989_));
 NOR3x1_ASAP7_75t_R _22375_ (.A(_13982_),
    .B(_13989_),
    .C(_13848_),
    .Y(_13990_));
 NAND2x1_ASAP7_75t_R _22376_ (.A(_13699_),
    .B(_13774_),
    .Y(_13991_));
 AOI21x1_ASAP7_75t_R _22377_ (.A1(net6),
    .A2(_13700_),
    .B(_13736_),
    .Y(_13992_));
 AOI21x1_ASAP7_75t_R _22378_ (.A1(_13743_),
    .A2(_13991_),
    .B(_13992_),
    .Y(_13993_));
 AOI21x1_ASAP7_75t_R _22379_ (.A1(_13778_),
    .A2(_13993_),
    .B(_13847_),
    .Y(_13994_));
 OAI21x1_ASAP7_75t_R _22380_ (.A1(_13888_),
    .A2(_13726_),
    .B(_13878_),
    .Y(_13995_));
 AO21x1_ASAP7_75t_R _22381_ (.A1(_13733_),
    .A2(_13728_),
    .B(_13934_),
    .Y(_13996_));
 NAND3x1_ASAP7_75t_R _22382_ (.A(_13995_),
    .B(_13752_),
    .C(_13996_),
    .Y(_13997_));
 AND3x1_ASAP7_75t_R _22383_ (.A(_13733_),
    .B(_00536_),
    .C(_13728_),
    .Y(_13998_));
 AOI21x1_ASAP7_75t_R _22384_ (.A1(_13636_),
    .A2(_13868_),
    .B(_13748_),
    .Y(_13999_));
 OAI21x1_ASAP7_75t_R _22385_ (.A1(_13998_),
    .A2(_13999_),
    .B(_13752_),
    .Y(_14000_));
 NOR2x1_ASAP7_75t_R _22386_ (.A(_01190_),
    .B(_13749_),
    .Y(_14001_));
 OAI21x1_ASAP7_75t_R _22387_ (.A1(_14001_),
    .A2(_13960_),
    .B(_13778_),
    .Y(_14002_));
 AOI21x1_ASAP7_75t_R _22388_ (.A1(_14000_),
    .A2(_14002_),
    .B(_13764_),
    .Y(_14003_));
 AOI211x1_ASAP7_75t_R _22389_ (.A1(_13994_),
    .A2(_13997_),
    .B(_14003_),
    .C(_13756_),
    .Y(_14004_));
 AO21x1_ASAP7_75t_R _22390_ (.A1(_13958_),
    .A2(_13819_),
    .B(_13777_),
    .Y(_14005_));
 AOI21x1_ASAP7_75t_R _22391_ (.A1(net6),
    .A2(_13865_),
    .B(_13743_),
    .Y(_14006_));
 OAI21x1_ASAP7_75t_R _22392_ (.A1(_14005_),
    .A2(_14006_),
    .B(_13763_),
    .Y(_14007_));
 OAI21x1_ASAP7_75t_R _22393_ (.A1(_13905_),
    .A2(_13726_),
    .B(_13823_),
    .Y(_14008_));
 INVx1_ASAP7_75t_R _22394_ (.A(_14008_),
    .Y(_14009_));
 OAI21x1_ASAP7_75t_R _22395_ (.A1(_13749_),
    .A2(_13854_),
    .B(_13694_),
    .Y(_14010_));
 NOR2x1_ASAP7_75t_R _22396_ (.A(_14009_),
    .B(_14010_),
    .Y(_14011_));
 OAI21x1_ASAP7_75t_R _22397_ (.A1(_14007_),
    .A2(_14011_),
    .B(_13756_),
    .Y(_14012_));
 AND2x2_ASAP7_75t_R _22398_ (.A(_01183_),
    .B(_13792_),
    .Y(_14013_));
 INVx1_ASAP7_75t_R _22399_ (.A(_14013_),
    .Y(_14014_));
 OAI21x1_ASAP7_75t_R _22400_ (.A1(_13624_),
    .A2(_13634_),
    .B(_14014_),
    .Y(_14015_));
 INVx1_ASAP7_75t_R _22401_ (.A(_14015_),
    .Y(_14016_));
 NAND2x2_ASAP7_75t_R _22402_ (.A(_15874_),
    .B(net541),
    .Y(_14017_));
 AOI221x1_ASAP7_75t_R _22403_ (.A1(_13698_),
    .A2(_14016_),
    .B1(_14017_),
    .B2(_13890_),
    .C(_13856_),
    .Y(_14018_));
 AO21x1_ASAP7_75t_R _22404_ (.A1(_13897_),
    .A2(_13958_),
    .B(_13907_),
    .Y(_14019_));
 INVx2_ASAP7_75t_R _22405_ (.A(_13707_),
    .Y(_14020_));
 OA21x2_ASAP7_75t_R _22406_ (.A1(_13825_),
    .A2(_14020_),
    .B(_13820_),
    .Y(_14021_));
 OAI21x1_ASAP7_75t_R _22407_ (.A1(_14019_),
    .A2(_14021_),
    .B(_13847_),
    .Y(_14022_));
 AOI21x1_ASAP7_75t_R _22408_ (.A1(_13933_),
    .A2(_14018_),
    .B(_14022_),
    .Y(_14023_));
 OAI21x1_ASAP7_75t_R _22409_ (.A1(_14012_),
    .A2(_14023_),
    .B(_13850_),
    .Y(_14024_));
 OAI22x1_ASAP7_75t_R _22410_ (.A1(_13990_),
    .A2(_13974_),
    .B1(_14004_),
    .B2(_14024_),
    .Y(_00066_));
 NAND2x1_ASAP7_75t_R _22411_ (.A(_15879_),
    .B(_13739_),
    .Y(_14025_));
 NOR2x2_ASAP7_75t_R _22412_ (.A(_15874_),
    .B(net69),
    .Y(_14026_));
 OAI21x1_ASAP7_75t_R _22413_ (.A1(_15869_),
    .A2(_13644_),
    .B(_13692_),
    .Y(_14027_));
 NOR2x2_ASAP7_75t_R _22414_ (.A(_14026_),
    .B(_14027_),
    .Y(_14028_));
 AOI21x1_ASAP7_75t_R _22415_ (.A1(_14025_),
    .A2(_14028_),
    .B(_13754_),
    .Y(_14029_));
 AO21x1_ASAP7_75t_R _22416_ (.A1(_13976_),
    .A2(_13895_),
    .B(_13665_),
    .Y(_14030_));
 NAND2x1_ASAP7_75t_R _22417_ (.A(_14030_),
    .B(_13914_),
    .Y(_14031_));
 AOI21x1_ASAP7_75t_R _22418_ (.A1(_14029_),
    .A2(_14031_),
    .B(_13847_),
    .Y(_14032_));
 AND3x1_ASAP7_75t_R _22419_ (.A(_13785_),
    .B(_13745_),
    .C(net727),
    .Y(_14033_));
 OAI21x1_ASAP7_75t_R _22420_ (.A1(_13668_),
    .A2(_13667_),
    .B(_13832_),
    .Y(_14034_));
 NOR2x1_ASAP7_75t_R _22421_ (.A(_14033_),
    .B(_14034_),
    .Y(_14035_));
 AO21x1_ASAP7_75t_R _22422_ (.A1(_13775_),
    .A2(_13700_),
    .B(_13859_),
    .Y(_14036_));
 AO21x1_ASAP7_75t_R _22423_ (.A1(_13784_),
    .A2(_13816_),
    .B(_13697_),
    .Y(_14037_));
 AOI21x1_ASAP7_75t_R _22424_ (.A1(_14036_),
    .A2(_14037_),
    .B(_13907_),
    .Y(_14038_));
 OAI21x1_ASAP7_75t_R _22425_ (.A1(_14035_),
    .A2(_14038_),
    .B(_13796_),
    .Y(_14039_));
 NAND2x1_ASAP7_75t_R _22426_ (.A(_14032_),
    .B(_14039_),
    .Y(_14040_));
 OAI21x1_ASAP7_75t_R _22427_ (.A1(_14026_),
    .A2(_13668_),
    .B(_13798_),
    .Y(_14041_));
 AOI21x1_ASAP7_75t_R _22428_ (.A1(_13782_),
    .A2(_13843_),
    .B(_13832_),
    .Y(_14042_));
 NAND2x1_ASAP7_75t_R _22429_ (.A(_14042_),
    .B(_14041_),
    .Y(_14043_));
 AO21x1_ASAP7_75t_R _22430_ (.A1(_13879_),
    .A2(_13852_),
    .B(_13697_),
    .Y(_14044_));
 AOI21x1_ASAP7_75t_R _22431_ (.A1(_13741_),
    .A2(_14044_),
    .B(_13755_),
    .Y(_14045_));
 AOI21x1_ASAP7_75t_R _22432_ (.A1(_14045_),
    .A2(_14043_),
    .B(_13763_),
    .Y(_14046_));
 AO21x1_ASAP7_75t_R _22433_ (.A1(_13738_),
    .A2(_13747_),
    .B(_13859_),
    .Y(_14047_));
 AO21x1_ASAP7_75t_R _22434_ (.A1(_13645_),
    .A2(_13700_),
    .B(_13697_),
    .Y(_14048_));
 AOI21x1_ASAP7_75t_R _22435_ (.A1(_14047_),
    .A2(_14048_),
    .B(_13790_),
    .Y(_14049_));
 AO21x1_ASAP7_75t_R _22436_ (.A1(_13767_),
    .A2(_13824_),
    .B(_13859_),
    .Y(_14050_));
 AOI21x1_ASAP7_75t_R _22437_ (.A1(_14050_),
    .A2(_13967_),
    .B(_13907_),
    .Y(_14051_));
 OAI21x1_ASAP7_75t_R _22438_ (.A1(_14049_),
    .A2(_14051_),
    .B(_13796_),
    .Y(_14052_));
 AOI21x1_ASAP7_75t_R _22439_ (.A1(_14052_),
    .A2(_14046_),
    .B(_13814_),
    .Y(_14053_));
 NAND2x1_ASAP7_75t_R _22440_ (.A(_14053_),
    .B(_14040_),
    .Y(_14054_));
 INVx2_ASAP7_75t_R _22441_ (.A(_13976_),
    .Y(_14055_));
 OAI21x1_ASAP7_75t_R _22442_ (.A1(_14055_),
    .A2(_14016_),
    .B(_13739_),
    .Y(_14056_));
 NAND2x1_ASAP7_75t_R _22443_ (.A(_14056_),
    .B(_13933_),
    .Y(_14057_));
 NAND2x1_ASAP7_75t_R _22444_ (.A(_13802_),
    .B(_13735_),
    .Y(_14058_));
 OAI21x1_ASAP7_75t_R _22445_ (.A1(_13905_),
    .A2(_14058_),
    .B(_13832_),
    .Y(_14059_));
 NAND2x1_ASAP7_75t_R _22446_ (.A(_13723_),
    .B(_14059_),
    .Y(_14060_));
 AOI21x1_ASAP7_75t_R _22447_ (.A1(_13856_),
    .A2(_14057_),
    .B(_14060_),
    .Y(_14061_));
 AOI21x1_ASAP7_75t_R _22448_ (.A1(_13878_),
    .A2(_13828_),
    .B(_13832_),
    .Y(_14062_));
 NAND2x1_ASAP7_75t_R _22449_ (.A(_13889_),
    .B(_14062_),
    .Y(_14063_));
 INVx3_ASAP7_75t_R _22450_ (.A(_13839_),
    .Y(_14064_));
 OAI21x1_ASAP7_75t_R _22451_ (.A1(_14064_),
    .A2(_13789_),
    .B(_13697_),
    .Y(_14065_));
 AO21x1_ASAP7_75t_R _22452_ (.A1(_13708_),
    .A2(_13803_),
    .B(_13665_),
    .Y(_14066_));
 NAND3x1_ASAP7_75t_R _22453_ (.A(_14066_),
    .B(_14065_),
    .C(_13907_),
    .Y(_14067_));
 AOI21x1_ASAP7_75t_R _22454_ (.A1(_14063_),
    .A2(_14067_),
    .B(_13926_),
    .Y(_14068_));
 OAI21x1_ASAP7_75t_R _22455_ (.A1(_14061_),
    .A2(_14068_),
    .B(_13764_),
    .Y(_14069_));
 AOI21x1_ASAP7_75t_R _22456_ (.A1(_13878_),
    .A2(_14064_),
    .B(_13722_),
    .Y(_14070_));
 INVx1_ASAP7_75t_R _22457_ (.A(_13977_),
    .Y(_14071_));
 AOI21x1_ASAP7_75t_R _22458_ (.A1(_14070_),
    .A2(_14071_),
    .B(_13907_),
    .Y(_14072_));
 OAI21x1_ASAP7_75t_R _22459_ (.A1(_14020_),
    .A2(_13668_),
    .B(_13804_),
    .Y(_14073_));
 AO21x1_ASAP7_75t_R _22460_ (.A1(_13803_),
    .A2(_14015_),
    .B(_13735_),
    .Y(_14074_));
 NAND3x1_ASAP7_75t_R _22461_ (.A(_14073_),
    .B(_14074_),
    .C(_13723_),
    .Y(_14075_));
 AOI21x1_ASAP7_75t_R _22462_ (.A1(_14072_),
    .A2(_14075_),
    .B(_13763_),
    .Y(_14076_));
 NOR2x1_ASAP7_75t_R _22463_ (.A(net727),
    .B(_13665_),
    .Y(_14077_));
 AO22x1_ASAP7_75t_R _22464_ (.A1(_13823_),
    .A2(_13940_),
    .B1(_14077_),
    .B2(_13754_),
    .Y(_14078_));
 NAND2x1_ASAP7_75t_R _22465_ (.A(_13878_),
    .B(_13904_),
    .Y(_14079_));
 AO21x1_ASAP7_75t_R _22466_ (.A1(_13911_),
    .A2(_13746_),
    .B(_13697_),
    .Y(_14080_));
 AOI21x1_ASAP7_75t_R _22467_ (.A1(_14079_),
    .A2(_14080_),
    .B(_13755_),
    .Y(_14081_));
 OAI21x1_ASAP7_75t_R _22468_ (.A1(_14078_),
    .A2(_14081_),
    .B(_13778_),
    .Y(_14082_));
 AOI21x1_ASAP7_75t_R _22469_ (.A1(_14076_),
    .A2(_14082_),
    .B(_13850_),
    .Y(_14083_));
 NAND2x1_ASAP7_75t_R _22470_ (.A(_14069_),
    .B(_14083_),
    .Y(_14084_));
 NAND2x1_ASAP7_75t_R _22471_ (.A(_14084_),
    .B(_14054_),
    .Y(_00067_));
 AOI21x1_ASAP7_75t_R _22472_ (.A1(_13879_),
    .A2(_13865_),
    .B(_13743_),
    .Y(_14085_));
 OAI21x1_ASAP7_75t_R _22473_ (.A1(_13957_),
    .A2(_14085_),
    .B(_13778_),
    .Y(_14086_));
 BUFx6f_ASAP7_75t_R _22474_ (.A(_13664_),
    .Y(_14087_));
 OA21x2_ASAP7_75t_R _22475_ (.A1(_13726_),
    .A2(_13897_),
    .B(_14087_),
    .Y(_14088_));
 OAI21x1_ASAP7_75t_R _22476_ (.A1(_14088_),
    .A2(_13827_),
    .B(_13752_),
    .Y(_14089_));
 AOI21x1_ASAP7_75t_R _22477_ (.A1(_14086_),
    .A2(_14089_),
    .B(_13756_),
    .Y(_14090_));
 NOR2x2_ASAP7_75t_R _22478_ (.A(_13816_),
    .B(_13785_),
    .Y(_14091_));
 NOR2x1_ASAP7_75t_R _22479_ (.A(_14064_),
    .B(_14091_),
    .Y(_14092_));
 AO21x1_ASAP7_75t_R _22480_ (.A1(_14092_),
    .A2(_13837_),
    .B(_13926_),
    .Y(_14093_));
 AO21x2_ASAP7_75t_R _22481_ (.A1(net815),
    .A2(_13799_),
    .B(_13748_),
    .Y(_14094_));
 NOR2x1_ASAP7_75t_R _22482_ (.A(_13904_),
    .B(_14094_),
    .Y(_14095_));
 AO21x1_ASAP7_75t_R _22483_ (.A1(_13869_),
    .A2(_13870_),
    .B(_13777_),
    .Y(_14096_));
 NOR2x1_ASAP7_75t_R _22484_ (.A(_14095_),
    .B(_14096_),
    .Y(_14097_));
 OAI21x1_ASAP7_75t_R _22485_ (.A1(_14097_),
    .A2(_14093_),
    .B(_13848_),
    .Y(_14098_));
 NOR2x1_ASAP7_75t_R _22486_ (.A(_14090_),
    .B(_14098_),
    .Y(_14099_));
 OAI21x1_ASAP7_75t_R _22487_ (.A1(_13838_),
    .A2(_15879_),
    .B(_13823_),
    .Y(_14100_));
 NOR2x1_ASAP7_75t_R _22488_ (.A(_13751_),
    .B(_13940_),
    .Y(_14101_));
 AO21x1_ASAP7_75t_R _22489_ (.A1(_14100_),
    .A2(_14101_),
    .B(_13926_),
    .Y(_14102_));
 AOI21x1_ASAP7_75t_R _22490_ (.A1(_13852_),
    .A2(_13782_),
    .B(_13798_),
    .Y(_14103_));
 OAI21x1_ASAP7_75t_R _22491_ (.A1(net539),
    .A2(_15879_),
    .B(_13898_),
    .Y(_14104_));
 OAI21x1_ASAP7_75t_R _22492_ (.A1(_13902_),
    .A2(_14104_),
    .B(_13790_),
    .Y(_14105_));
 NOR2x1_ASAP7_75t_R _22493_ (.A(_14103_),
    .B(_14105_),
    .Y(_14106_));
 OAI21x1_ASAP7_75t_R _22494_ (.A1(_14102_),
    .A2(_14106_),
    .B(_13764_),
    .Y(_14107_));
 AOI21x1_ASAP7_75t_R _22495_ (.A1(_13699_),
    .A2(_13774_),
    .B(_13743_),
    .Y(_14108_));
 AOI21x1_ASAP7_75t_R _22496_ (.A1(_13646_),
    .A2(_13782_),
    .B(_13698_),
    .Y(_14109_));
 OAI21x1_ASAP7_75t_R _22497_ (.A1(_14108_),
    .A2(_14109_),
    .B(_13778_),
    .Y(_14110_));
 INVx1_ASAP7_75t_R _22498_ (.A(_13995_),
    .Y(_14111_));
 OAI21x1_ASAP7_75t_R _22499_ (.A1(_13929_),
    .A2(_14111_),
    .B(_13752_),
    .Y(_14112_));
 AOI21x1_ASAP7_75t_R _22500_ (.A1(_14110_),
    .A2(_14112_),
    .B(_13756_),
    .Y(_14113_));
 OAI21x1_ASAP7_75t_R _22501_ (.A1(_14107_),
    .A2(_14113_),
    .B(_13850_),
    .Y(_14114_));
 AOI21x1_ASAP7_75t_R _22502_ (.A1(_13803_),
    .A2(_13910_),
    .B(_13698_),
    .Y(_14115_));
 AO21x1_ASAP7_75t_R _22503_ (.A1(_13820_),
    .A2(_15882_),
    .B(_13907_),
    .Y(_14116_));
 OAI21x1_ASAP7_75t_R _22504_ (.A1(_14115_),
    .A2(_14116_),
    .B(_13724_),
    .Y(_14117_));
 OAI21x1_ASAP7_75t_R _22505_ (.A1(_13747_),
    .A2(_13749_),
    .B(_13907_),
    .Y(_14118_));
 NOR2x2_ASAP7_75t_R _22506_ (.A(_13664_),
    .B(_13782_),
    .Y(_14119_));
 AOI211x1_ASAP7_75t_R _22507_ (.A1(_13860_),
    .A2(_13782_),
    .B(_14118_),
    .C(_14119_),
    .Y(_14120_));
 OAI21x1_ASAP7_75t_R _22508_ (.A1(_14117_),
    .A2(_14120_),
    .B(_13764_),
    .Y(_14121_));
 NOR2x1_ASAP7_75t_R _22509_ (.A(_13778_),
    .B(_13786_),
    .Y(_14122_));
 AO21x1_ASAP7_75t_R _22510_ (.A1(_13794_),
    .A2(_13738_),
    .B(_13698_),
    .Y(_14123_));
 OA21x2_ASAP7_75t_R _22511_ (.A1(_14017_),
    .A2(_15879_),
    .B(_13820_),
    .Y(_14124_));
 NAND2x1_ASAP7_75t_R _22512_ (.A(_01183_),
    .B(_13636_),
    .Y(_14125_));
 AO21x1_ASAP7_75t_R _22513_ (.A1(_14125_),
    .A2(_13958_),
    .B(_13751_),
    .Y(_14126_));
 OAI21x1_ASAP7_75t_R _22514_ (.A1(_14124_),
    .A2(_14126_),
    .B(_13796_),
    .Y(_14127_));
 AOI21x1_ASAP7_75t_R _22515_ (.A1(_14122_),
    .A2(_14123_),
    .B(_14127_),
    .Y(_14128_));
 OAI21x1_ASAP7_75t_R _22516_ (.A1(_14121_),
    .A2(_14128_),
    .B(_13814_),
    .Y(_14129_));
 OAI21x1_ASAP7_75t_R _22517_ (.A1(_00537_),
    .A2(_14087_),
    .B(_13751_),
    .Y(_14130_));
 OA21x2_ASAP7_75t_R _22518_ (.A1(_14130_),
    .A2(_14091_),
    .B(_13755_),
    .Y(_14131_));
 NOR2x1_ASAP7_75t_R _22519_ (.A(_14087_),
    .B(_13865_),
    .Y(_14132_));
 NOR2x1_ASAP7_75t_R _22520_ (.A(net61),
    .B(_13636_),
    .Y(_14133_));
 OAI21x1_ASAP7_75t_R _22521_ (.A1(_14055_),
    .A2(_14133_),
    .B(_13823_),
    .Y(_14134_));
 INVx1_ASAP7_75t_R _22522_ (.A(_14134_),
    .Y(_14135_));
 OAI21x1_ASAP7_75t_R _22523_ (.A1(_14132_),
    .A2(_14135_),
    .B(_13778_),
    .Y(_14136_));
 NAND2x1_ASAP7_75t_R _22524_ (.A(_14131_),
    .B(_14136_),
    .Y(_14137_));
 NOR2x2_ASAP7_75t_R _22525_ (.A(_13693_),
    .B(_13871_),
    .Y(_14138_));
 INVx1_ASAP7_75t_R _22526_ (.A(_14138_),
    .Y(_14139_));
 NAND2x1_ASAP7_75t_R _22527_ (.A(_13798_),
    .B(_13943_),
    .Y(_14140_));
 OAI21x1_ASAP7_75t_R _22528_ (.A1(_13668_),
    .A2(_13667_),
    .B(_14140_),
    .Y(_14141_));
 NOR2x1_ASAP7_75t_R _22529_ (.A(_14139_),
    .B(_14141_),
    .Y(_14142_));
 OA21x2_ASAP7_75t_R _22530_ (.A1(_13880_),
    .A2(_13901_),
    .B(_13735_),
    .Y(_14143_));
 OAI21x1_ASAP7_75t_R _22531_ (.A1(_13905_),
    .A2(_14100_),
    .B(_13694_),
    .Y(_14144_));
 NOR2x1_ASAP7_75t_R _22532_ (.A(_14143_),
    .B(_14144_),
    .Y(_14145_));
 OAI21x1_ASAP7_75t_R _22533_ (.A1(_14142_),
    .A2(_14145_),
    .B(_13724_),
    .Y(_14146_));
 AOI21x1_ASAP7_75t_R _22534_ (.A1(_14137_),
    .A2(_14146_),
    .B(_13764_),
    .Y(_14147_));
 OAI22x1_ASAP7_75t_R _22535_ (.A1(_14099_),
    .A2(_14114_),
    .B1(_14129_),
    .B2(_14147_),
    .Y(_00068_));
 NAND2x1_ASAP7_75t_R _22536_ (.A(_14013_),
    .B(_13799_),
    .Y(_14148_));
 AO21x1_ASAP7_75t_R _22537_ (.A1(_14148_),
    .A2(_14087_),
    .B(_13777_),
    .Y(_14149_));
 AND2x2_ASAP7_75t_R _22538_ (.A(_13999_),
    .B(_13950_),
    .Y(_14150_));
 INVx1_ASAP7_75t_R _22539_ (.A(_13913_),
    .Y(_14151_));
 AOI21x1_ASAP7_75t_R _22540_ (.A1(_14151_),
    .A2(_13837_),
    .B(_13723_),
    .Y(_14152_));
 OAI21x1_ASAP7_75t_R _22541_ (.A1(_14149_),
    .A2(_14150_),
    .B(_14152_),
    .Y(_14153_));
 INVx1_ASAP7_75t_R _22542_ (.A(_00531_),
    .Y(_14154_));
 OA21x2_ASAP7_75t_R _22543_ (.A1(_13735_),
    .A2(_14154_),
    .B(_13692_),
    .Y(_14155_));
 AO21x1_ASAP7_75t_R _22544_ (.A1(_13901_),
    .A2(_13799_),
    .B(_13697_),
    .Y(_14156_));
 AOI21x1_ASAP7_75t_R _22545_ (.A1(_14155_),
    .A2(_14156_),
    .B(_13754_),
    .Y(_14157_));
 AO21x1_ASAP7_75t_R _22546_ (.A1(_13895_),
    .A2(_13803_),
    .B(_13665_),
    .Y(_14158_));
 AO21x1_ASAP7_75t_R _22547_ (.A1(_13746_),
    .A2(_13708_),
    .B(_13735_),
    .Y(_14159_));
 NAND3x1_ASAP7_75t_R _22548_ (.A(_14158_),
    .B(_14159_),
    .C(_13907_),
    .Y(_14160_));
 AOI21x1_ASAP7_75t_R _22549_ (.A1(_14157_),
    .A2(_14160_),
    .B(_13763_),
    .Y(_14161_));
 AOI21x1_ASAP7_75t_R _22550_ (.A1(_14153_),
    .A2(_14161_),
    .B(_13850_),
    .Y(_14162_));
 NAND2x1_ASAP7_75t_R _22551_ (.A(_13804_),
    .B(_13905_),
    .Y(_14163_));
 AND2x2_ASAP7_75t_R _22552_ (.A(_13846_),
    .B(_14163_),
    .Y(_14164_));
 AO21x1_ASAP7_75t_R _22553_ (.A1(_13784_),
    .A2(_13803_),
    .B(_13878_),
    .Y(_14165_));
 OA21x2_ASAP7_75t_R _22554_ (.A1(_13804_),
    .A2(_13746_),
    .B(_13832_),
    .Y(_14166_));
 AO21x1_ASAP7_75t_R _22555_ (.A1(_14165_),
    .A2(_14166_),
    .B(_13796_),
    .Y(_14167_));
 OA21x2_ASAP7_75t_R _22556_ (.A1(_13735_),
    .A2(net60),
    .B(_13692_),
    .Y(_14168_));
 AOI21x1_ASAP7_75t_R _22557_ (.A1(_14168_),
    .A2(_13666_),
    .B(_13723_),
    .Y(_14169_));
 AO21x1_ASAP7_75t_R _22558_ (.A1(_13775_),
    .A2(_13708_),
    .B(_13859_),
    .Y(_14170_));
 OA21x2_ASAP7_75t_R _22559_ (.A1(_13838_),
    .A2(_13644_),
    .B(_13734_),
    .Y(_14171_));
 AOI21x1_ASAP7_75t_R _22560_ (.A1(_13911_),
    .A2(_14171_),
    .B(_13740_),
    .Y(_14172_));
 NAND2x1_ASAP7_75t_R _22561_ (.A(_14170_),
    .B(_14172_),
    .Y(_14173_));
 AOI21x1_ASAP7_75t_R _22562_ (.A1(_14169_),
    .A2(_14173_),
    .B(_13847_),
    .Y(_14174_));
 OAI21x1_ASAP7_75t_R _22563_ (.A1(_14164_),
    .A2(_14167_),
    .B(_14174_),
    .Y(_14175_));
 NAND2x1_ASAP7_75t_R _22564_ (.A(_14162_),
    .B(_14175_),
    .Y(_14176_));
 NAND2x1_ASAP7_75t_R _22565_ (.A(_13792_),
    .B(_13644_),
    .Y(_14177_));
 AOI21x1_ASAP7_75t_R _22566_ (.A1(_13798_),
    .A2(_14177_),
    .B(_13740_),
    .Y(_14178_));
 OAI21x1_ASAP7_75t_R _22567_ (.A1(_13736_),
    .A2(_13775_),
    .B(_14178_),
    .Y(_14179_));
 AO21x1_ASAP7_75t_R _22568_ (.A1(_13785_),
    .A2(_13895_),
    .B(_13693_),
    .Y(_14180_));
 INVx1_ASAP7_75t_R _22569_ (.A(_14180_),
    .Y(_14181_));
 AOI21x1_ASAP7_75t_R _22570_ (.A1(_14065_),
    .A2(_14181_),
    .B(_13754_),
    .Y(_14182_));
 AOI21x1_ASAP7_75t_R _22571_ (.A1(_14179_),
    .A2(_14182_),
    .B(_13847_),
    .Y(_14183_));
 NAND2x1_ASAP7_75t_R _22572_ (.A(_13869_),
    .B(_14171_),
    .Y(_14184_));
 AOI21x1_ASAP7_75t_R _22573_ (.A1(_13793_),
    .A2(_13878_),
    .B(_13864_),
    .Y(_14185_));
 AOI21x1_ASAP7_75t_R _22574_ (.A1(_14184_),
    .A2(_14185_),
    .B(_13723_),
    .Y(_14186_));
 NAND2x1_ASAP7_75t_R _22575_ (.A(_14177_),
    .B(_13913_),
    .Y(_14187_));
 INVx1_ASAP7_75t_R _22576_ (.A(_14119_),
    .Y(_14188_));
 NAND3x1_ASAP7_75t_R _22577_ (.A(_14187_),
    .B(_14138_),
    .C(_14188_),
    .Y(_14189_));
 NAND2x1_ASAP7_75t_R _22578_ (.A(_14186_),
    .B(_14189_),
    .Y(_14190_));
 AOI21x1_ASAP7_75t_R _22579_ (.A1(_14183_),
    .A2(_14190_),
    .B(_13814_),
    .Y(_14191_));
 AO21x1_ASAP7_75t_R _22580_ (.A1(_13665_),
    .A2(net61),
    .B(_13693_),
    .Y(_14192_));
 NOR2x1_ASAP7_75t_R _22581_ (.A(_14192_),
    .B(_14143_),
    .Y(_14193_));
 AO21x1_ASAP7_75t_R _22582_ (.A1(_13884_),
    .A2(_14017_),
    .B(_13697_),
    .Y(_14194_));
 AO21x1_ASAP7_75t_R _22583_ (.A1(_13784_),
    .A2(_13746_),
    .B(_13859_),
    .Y(_14195_));
 AOI21x1_ASAP7_75t_R _22584_ (.A1(_14194_),
    .A2(_14195_),
    .B(_13790_),
    .Y(_14196_));
 OAI21x1_ASAP7_75t_R _22585_ (.A1(_14193_),
    .A2(_14196_),
    .B(_13796_),
    .Y(_14197_));
 NAND2x1_ASAP7_75t_R _22586_ (.A(_13830_),
    .B(_13911_),
    .Y(_14198_));
 AOI21x1_ASAP7_75t_R _22587_ (.A1(_13798_),
    .A2(_14198_),
    .B(_14091_),
    .Y(_14199_));
 INVx1_ASAP7_75t_R _22588_ (.A(_13843_),
    .Y(_14200_));
 AOI21x1_ASAP7_75t_R _22589_ (.A1(_13735_),
    .A2(_13803_),
    .B(_13693_),
    .Y(_14201_));
 OAI21x1_ASAP7_75t_R _22590_ (.A1(_13943_),
    .A2(_14200_),
    .B(_14201_),
    .Y(_14202_));
 OAI21x1_ASAP7_75t_R _22591_ (.A1(_13790_),
    .A2(_14199_),
    .B(_14202_),
    .Y(_14203_));
 AOI21x1_ASAP7_75t_R _22592_ (.A1(_13926_),
    .A2(_14203_),
    .B(_13763_),
    .Y(_14204_));
 NAND2x1_ASAP7_75t_R _22593_ (.A(_14197_),
    .B(_14204_),
    .Y(_14205_));
 NAND2x1_ASAP7_75t_R _22594_ (.A(_14191_),
    .B(_14205_),
    .Y(_14206_));
 NAND2x1_ASAP7_75t_R _22595_ (.A(_14176_),
    .B(_14206_),
    .Y(_00069_));
 AOI21x1_ASAP7_75t_R _22596_ (.A1(_13781_),
    .A2(_13705_),
    .B(_13736_),
    .Y(_14207_));
 OAI21x1_ASAP7_75t_R _22597_ (.A1(_14055_),
    .A2(_13875_),
    .B(_13898_),
    .Y(_14208_));
 INVx1_ASAP7_75t_R _22598_ (.A(_14208_),
    .Y(_14209_));
 OAI21x1_ASAP7_75t_R _22599_ (.A1(_14207_),
    .A2(_14209_),
    .B(_13856_),
    .Y(_14210_));
 NOR2x1_ASAP7_75t_R _22600_ (.A(_14013_),
    .B(_13799_),
    .Y(_14211_));
 OA21x2_ASAP7_75t_R _22601_ (.A1(_14211_),
    .A2(_14064_),
    .B(_14087_),
    .Y(_14212_));
 OA21x2_ASAP7_75t_R _22602_ (.A1(_13904_),
    .A2(_13902_),
    .B(_13958_),
    .Y(_14213_));
 OAI21x1_ASAP7_75t_R _22603_ (.A1(_14212_),
    .A2(_14213_),
    .B(_13778_),
    .Y(_14214_));
 AOI21x1_ASAP7_75t_R _22604_ (.A1(_14214_),
    .A2(_14210_),
    .B(_13756_),
    .Y(_14215_));
 OA21x2_ASAP7_75t_R _22605_ (.A1(_14064_),
    .A2(_13831_),
    .B(_14087_),
    .Y(_14216_));
 NAND2x1_ASAP7_75t_R _22606_ (.A(_01187_),
    .B(_01189_),
    .Y(_14217_));
 AOI21x1_ASAP7_75t_R _22607_ (.A1(_13958_),
    .A2(_14217_),
    .B(_13777_),
    .Y(_14218_));
 OAI21x1_ASAP7_75t_R _22608_ (.A1(_13901_),
    .A2(_13880_),
    .B(_13823_),
    .Y(_14219_));
 AOI21x1_ASAP7_75t_R _22609_ (.A1(_14218_),
    .A2(_14219_),
    .B(_13926_),
    .Y(_14220_));
 OA21x2_ASAP7_75t_R _22610_ (.A1(_14118_),
    .A2(_14216_),
    .B(_14220_),
    .Y(_14221_));
 NOR3x1_ASAP7_75t_R _22611_ (.A(_14215_),
    .B(_13848_),
    .C(_14221_),
    .Y(_14222_));
 NOR2x1_ASAP7_75t_R _22612_ (.A(_15879_),
    .B(_13646_),
    .Y(_14223_));
 NAND2x1_ASAP7_75t_R _22613_ (.A(_14087_),
    .B(_13911_),
    .Y(_14224_));
 NAND2x1_ASAP7_75t_R _22614_ (.A(_13898_),
    .B(_14125_),
    .Y(_14225_));
 OAI21x1_ASAP7_75t_R _22615_ (.A1(_14223_),
    .A2(_14224_),
    .B(_14225_),
    .Y(_14226_));
 OA21x2_ASAP7_75t_R _22616_ (.A1(_13697_),
    .A2(_13708_),
    .B(_13740_),
    .Y(_14227_));
 INVx1_ASAP7_75t_R _22617_ (.A(_13998_),
    .Y(_14228_));
 OAI21x1_ASAP7_75t_R _22618_ (.A1(net727),
    .A2(_14087_),
    .B(_13777_),
    .Y(_14229_));
 AOI21x1_ASAP7_75t_R _22619_ (.A1(_14228_),
    .A2(_13970_),
    .B(_14229_),
    .Y(_14230_));
 AOI21x1_ASAP7_75t_R _22620_ (.A1(_14226_),
    .A2(_14227_),
    .B(_14230_),
    .Y(_14231_));
 NOR2x1_ASAP7_75t_R _22621_ (.A(_13668_),
    .B(_13667_),
    .Y(_14232_));
 AO21x1_ASAP7_75t_R _22622_ (.A1(_13738_),
    .A2(_14015_),
    .B(_13739_),
    .Y(_14233_));
 AOI21x1_ASAP7_75t_R _22623_ (.A1(net60),
    .A2(_13890_),
    .B(_13777_),
    .Y(_14234_));
 NAND2x1_ASAP7_75t_R _22624_ (.A(_14233_),
    .B(_14234_),
    .Y(_14235_));
 OAI21x1_ASAP7_75t_R _22625_ (.A1(net61),
    .A2(_13905_),
    .B(_13820_),
    .Y(_14236_));
 OA21x2_ASAP7_75t_R _22626_ (.A1(_13739_),
    .A2(_13746_),
    .B(_13832_),
    .Y(_14237_));
 AOI21x1_ASAP7_75t_R _22627_ (.A1(_14236_),
    .A2(_14237_),
    .B(_13796_),
    .Y(_14238_));
 OAI21x1_ASAP7_75t_R _22628_ (.A1(_14232_),
    .A2(_14235_),
    .B(_14238_),
    .Y(_14239_));
 OAI21x1_ASAP7_75t_R _22629_ (.A1(_13724_),
    .A2(_14231_),
    .B(_14239_),
    .Y(_14240_));
 OAI21x1_ASAP7_75t_R _22630_ (.A1(_13764_),
    .A2(_14240_),
    .B(_13850_),
    .Y(_14241_));
 NAND2x1_ASAP7_75t_R _22631_ (.A(_13878_),
    .B(_13879_),
    .Y(_14242_));
 NAND2x1_ASAP7_75t_R _22632_ (.A(_14242_),
    .B(_13801_),
    .Y(_14243_));
 AOI21x1_ASAP7_75t_R _22633_ (.A1(_14065_),
    .A2(_14227_),
    .B(_13755_),
    .Y(_14244_));
 NAND2x1_ASAP7_75t_R _22634_ (.A(_14244_),
    .B(_14243_),
    .Y(_14245_));
 OAI21x1_ASAP7_75t_R _22635_ (.A1(net69),
    .A2(_15874_),
    .B(_13820_),
    .Y(_14246_));
 AOI21x1_ASAP7_75t_R _22636_ (.A1(_14246_),
    .A2(_14094_),
    .B(_13668_),
    .Y(_14247_));
 NAND2x1_ASAP7_75t_R _22637_ (.A(net61),
    .B(_13958_),
    .Y(_14248_));
 AOI21x1_ASAP7_75t_R _22638_ (.A1(_14248_),
    .A2(_14028_),
    .B(_13926_),
    .Y(_14249_));
 OAI21x1_ASAP7_75t_R _22639_ (.A1(_13752_),
    .A2(_14247_),
    .B(_14249_),
    .Y(_14250_));
 AOI21x1_ASAP7_75t_R _22640_ (.A1(_14245_),
    .A2(_14250_),
    .B(_13848_),
    .Y(_14251_));
 NOR2x1_ASAP7_75t_R _22641_ (.A(_14020_),
    .B(_14151_),
    .Y(_14252_));
 AO21x1_ASAP7_75t_R _22642_ (.A1(_13668_),
    .A2(_13958_),
    .B(_13751_),
    .Y(_14253_));
 AOI21x1_ASAP7_75t_R _22643_ (.A1(_00538_),
    .A2(_13820_),
    .B(_13777_),
    .Y(_14254_));
 OAI21x1_ASAP7_75t_R _22644_ (.A1(_14055_),
    .A2(_14133_),
    .B(_13958_),
    .Y(_14255_));
 AOI21x1_ASAP7_75t_R _22645_ (.A1(_14254_),
    .A2(_14255_),
    .B(_13926_),
    .Y(_14256_));
 OAI21x1_ASAP7_75t_R _22646_ (.A1(_14252_),
    .A2(_14253_),
    .B(_14256_),
    .Y(_14257_));
 AOI21x1_ASAP7_75t_R _22647_ (.A1(_13698_),
    .A2(_13826_),
    .B(_13694_),
    .Y(_14258_));
 AO21x1_ASAP7_75t_R _22648_ (.A1(_14154_),
    .A2(_15882_),
    .B(_13878_),
    .Y(_14259_));
 AOI21x1_ASAP7_75t_R _22649_ (.A1(_14259_),
    .A2(_14134_),
    .B(_13856_),
    .Y(_14260_));
 OAI21x1_ASAP7_75t_R _22650_ (.A1(_14258_),
    .A2(_14260_),
    .B(_13724_),
    .Y(_14261_));
 AOI21x1_ASAP7_75t_R _22651_ (.A1(_14257_),
    .A2(_14261_),
    .B(_13764_),
    .Y(_14262_));
 OAI21x1_ASAP7_75t_R _22652_ (.A1(_14251_),
    .A2(_14262_),
    .B(_13814_),
    .Y(_14263_));
 OAI21x1_ASAP7_75t_R _22653_ (.A1(_14241_),
    .A2(_14222_),
    .B(_14263_),
    .Y(_00070_));
 AND3x1_ASAP7_75t_R _22654_ (.A(_14134_),
    .B(_14094_),
    .C(_13856_),
    .Y(_14264_));
 NAND2x1_ASAP7_75t_R _22655_ (.A(_13747_),
    .B(_13705_),
    .Y(_14265_));
 AOI211x1_ASAP7_75t_R _22656_ (.A1(_13698_),
    .A2(_14265_),
    .B(_14253_),
    .C(_14132_),
    .Y(_14266_));
 OAI21x1_ASAP7_75t_R _22657_ (.A1(_14264_),
    .A2(_14266_),
    .B(_13756_),
    .Y(_14267_));
 AOI21x1_ASAP7_75t_R _22658_ (.A1(_13876_),
    .A2(_14073_),
    .B(_13790_),
    .Y(_14268_));
 AOI21x1_ASAP7_75t_R _22659_ (.A1(_14208_),
    .A2(_14008_),
    .B(_13694_),
    .Y(_14269_));
 NOR2x1_ASAP7_75t_R _22660_ (.A(_14269_),
    .B(_14268_),
    .Y(_14270_));
 AOI21x1_ASAP7_75t_R _22661_ (.A1(_13724_),
    .A2(_14270_),
    .B(_13848_),
    .Y(_14271_));
 OAI21x1_ASAP7_75t_R _22662_ (.A1(_15882_),
    .A2(_13646_),
    .B(_13823_),
    .Y(_14272_));
 OAI21x1_ASAP7_75t_R _22663_ (.A1(_15879_),
    .A2(_14017_),
    .B(_13798_),
    .Y(_14273_));
 OAI21x1_ASAP7_75t_R _22664_ (.A1(net67),
    .A2(_13823_),
    .B(_13777_),
    .Y(_14274_));
 AOI21x1_ASAP7_75t_R _22665_ (.A1(_14272_),
    .A2(_14273_),
    .B(_14274_),
    .Y(_14275_));
 AOI21x1_ASAP7_75t_R _22666_ (.A1(_15879_),
    .A2(_14017_),
    .B(_13898_),
    .Y(_14276_));
 OAI21x1_ASAP7_75t_R _22667_ (.A1(_14276_),
    .A2(_14180_),
    .B(_13723_),
    .Y(_14277_));
 OAI21x1_ASAP7_75t_R _22668_ (.A1(_14275_),
    .A2(_14277_),
    .B(_13847_),
    .Y(_14278_));
 OAI21x1_ASAP7_75t_R _22669_ (.A1(_13880_),
    .A2(_14273_),
    .B(_13995_),
    .Y(_14279_));
 AO21x1_ASAP7_75t_R _22670_ (.A1(_13859_),
    .A2(net60),
    .B(_13740_),
    .Y(_14280_));
 OAI21x1_ASAP7_75t_R _22671_ (.A1(_14280_),
    .A2(_14103_),
    .B(_13755_),
    .Y(_14281_));
 AOI21x1_ASAP7_75t_R _22672_ (.A1(_13752_),
    .A2(_14279_),
    .B(_14281_),
    .Y(_14282_));
 NOR2x1_ASAP7_75t_R _22673_ (.A(_14282_),
    .B(_14278_),
    .Y(_14283_));
 AOI21x1_ASAP7_75t_R _22674_ (.A1(_14267_),
    .A2(_14271_),
    .B(_14283_),
    .Y(_14284_));
 AOI21x1_ASAP7_75t_R _22675_ (.A1(net61),
    .A2(_13804_),
    .B(_13740_),
    .Y(_14285_));
 NAND2x1_ASAP7_75t_R _22676_ (.A(_14285_),
    .B(_14163_),
    .Y(_14286_));
 INVx1_ASAP7_75t_R _22677_ (.A(_13928_),
    .Y(_14287_));
 NAND2x1_ASAP7_75t_R _22678_ (.A(_00537_),
    .B(_14087_),
    .Y(_14288_));
 AOI21x1_ASAP7_75t_R _22679_ (.A1(_14288_),
    .A2(_13833_),
    .B(_13926_),
    .Y(_14289_));
 OAI21x1_ASAP7_75t_R _22680_ (.A1(_14286_),
    .A2(_14287_),
    .B(_14289_),
    .Y(_14290_));
 NAND2x1_ASAP7_75t_R _22681_ (.A(_13895_),
    .B(_13816_),
    .Y(_14291_));
 AOI21x1_ASAP7_75t_R _22682_ (.A1(_13823_),
    .A2(_14291_),
    .B(_13751_),
    .Y(_14292_));
 AO21x1_ASAP7_75t_R _22683_ (.A1(_13645_),
    .A2(_13774_),
    .B(_13739_),
    .Y(_14293_));
 NAND2x1_ASAP7_75t_R _22684_ (.A(_14292_),
    .B(_14293_),
    .Y(_14294_));
 NAND2x1_ASAP7_75t_R _22685_ (.A(_13898_),
    .B(_13904_),
    .Y(_14295_));
 OAI21x1_ASAP7_75t_R _22686_ (.A1(_01189_),
    .A2(_13859_),
    .B(_13740_),
    .Y(_14296_));
 NOR2x1_ASAP7_75t_R _22687_ (.A(_13840_),
    .B(_14296_),
    .Y(_14297_));
 AOI21x1_ASAP7_75t_R _22688_ (.A1(_14295_),
    .A2(_14297_),
    .B(_13755_),
    .Y(_14298_));
 NAND2x1_ASAP7_75t_R _22689_ (.A(_14294_),
    .B(_14298_),
    .Y(_14299_));
 AOI21x1_ASAP7_75t_R _22690_ (.A1(_14290_),
    .A2(_14299_),
    .B(_13764_),
    .Y(_14300_));
 OA21x2_ASAP7_75t_R _22691_ (.A1(_13697_),
    .A2(_13792_),
    .B(_13832_),
    .Y(_14301_));
 AOI21x1_ASAP7_75t_R _22692_ (.A1(_14219_),
    .A2(_14301_),
    .B(_13755_),
    .Y(_14302_));
 OA21x2_ASAP7_75t_R _22693_ (.A1(_13782_),
    .A2(_13804_),
    .B(_13747_),
    .Y(_14303_));
 NAND2x1_ASAP7_75t_R _22694_ (.A(_13833_),
    .B(_14303_),
    .Y(_14304_));
 NAND2x1_ASAP7_75t_R _22695_ (.A(_14302_),
    .B(_14304_),
    .Y(_14305_));
 NAND2x1_ASAP7_75t_R _22696_ (.A(_13804_),
    .B(_13789_),
    .Y(_14306_));
 NAND3x1_ASAP7_75t_R _22697_ (.A(_14056_),
    .B(_14306_),
    .C(_14285_),
    .Y(_14307_));
 NAND2x1_ASAP7_75t_R _22698_ (.A(_13746_),
    .B(_13895_),
    .Y(_14308_));
 AOI21x1_ASAP7_75t_R _22699_ (.A1(_14087_),
    .A2(_14308_),
    .B(_13777_),
    .Y(_14309_));
 OAI21x1_ASAP7_75t_R _22700_ (.A1(_13897_),
    .A2(_13918_),
    .B(_13958_),
    .Y(_14310_));
 AOI21x1_ASAP7_75t_R _22701_ (.A1(_14309_),
    .A2(_14310_),
    .B(_13926_),
    .Y(_14311_));
 NAND2x1_ASAP7_75t_R _22702_ (.A(_14307_),
    .B(_14311_),
    .Y(_14312_));
 AOI21x1_ASAP7_75t_R _22703_ (.A1(_14305_),
    .A2(_14312_),
    .B(_13848_),
    .Y(_14313_));
 OAI21x1_ASAP7_75t_R _22704_ (.A1(_14300_),
    .A2(_14313_),
    .B(_13850_),
    .Y(_14314_));
 OAI21x1_ASAP7_75t_R _22705_ (.A1(_14284_),
    .A2(_13850_),
    .B(_14314_),
    .Y(_00071_));
 INVx2_ASAP7_75t_R _22706_ (.A(net789),
    .Y(_14315_));
 XOR2x1_ASAP7_75t_R _22707_ (.A(_14315_),
    .Y(_14316_),
    .B(_11359_));
 XNOR2x2_ASAP7_75t_R _22708_ (.A(_11539_),
    .B(_11388_),
    .Y(_14317_));
 XOR2x2_ASAP7_75t_R _22709_ (.A(_11360_),
    .B(_11365_),
    .Y(_14318_));
 XOR2x1_ASAP7_75t_R _22710_ (.A(_14317_),
    .Y(_14319_),
    .B(_14318_));
 NOR2x1_ASAP7_75t_R _22711_ (.A(_14319_),
    .B(_14316_),
    .Y(_14320_));
 XOR2x1_ASAP7_75t_R _22712_ (.A(_11359_),
    .Y(_14321_),
    .B(net789));
 XOR2x2_ASAP7_75t_R _22713_ (.A(_11388_),
    .B(_11539_),
    .Y(_14322_));
 XOR2x1_ASAP7_75t_R _22714_ (.A(_14318_),
    .Y(_14323_),
    .B(_14322_));
 OAI21x1_ASAP7_75t_R _22715_ (.A1(_14321_),
    .A2(_14323_),
    .B(_10742_),
    .Y(_14324_));
 NAND2x1_ASAP7_75t_R _22716_ (.A(_00539_),
    .B(_11373_),
    .Y(_14325_));
 OAI21x1_ASAP7_75t_R _22717_ (.A1(_14320_),
    .A2(_14324_),
    .B(_14325_),
    .Y(_14326_));
 XOR2x2_ASAP7_75t_R _22718_ (.A(_07970_),
    .B(_14326_),
    .Y(_15889_));
 NOR2x2_ASAP7_75t_R _22719_ (.A(net767),
    .B(_00540_),
    .Y(_14327_));
 XOR2x1_ASAP7_75t_R _22720_ (.A(_11362_),
    .Y(_14328_),
    .B(_11383_));
 NAND2x1_ASAP7_75t_R _22721_ (.A(_11382_),
    .B(_14328_),
    .Y(_14329_));
 XNOR2x1_ASAP7_75t_R _22722_ (.B(_11383_),
    .Y(_14330_),
    .A(_11362_));
 NAND2x1_ASAP7_75t_R _22723_ (.A(net776),
    .B(_14330_),
    .Y(_14331_));
 AOI21x1_ASAP7_75t_R _22724_ (.A1(_14329_),
    .A2(_14331_),
    .B(_14317_),
    .Y(_14332_));
 XOR2x1_ASAP7_75t_R _22725_ (.A(_11383_),
    .Y(_14333_),
    .B(net776));
 NAND2x1_ASAP7_75t_R _22726_ (.A(net19),
    .B(_14333_),
    .Y(_14334_));
 INVx1_ASAP7_75t_R _22727_ (.A(net19),
    .Y(_14335_));
 XNOR2x1_ASAP7_75t_R _22728_ (.B(net776),
    .Y(_14336_),
    .A(_11383_));
 NAND2x1_ASAP7_75t_R _22729_ (.A(_14335_),
    .B(_14336_),
    .Y(_14337_));
 AOI21x1_ASAP7_75t_R _22730_ (.A1(_14334_),
    .A2(_14337_),
    .B(net696),
    .Y(_14338_));
 OAI21x1_ASAP7_75t_R _22731_ (.A1(_14332_),
    .A2(_14338_),
    .B(_10723_),
    .Y(_14339_));
 INVx2_ASAP7_75t_R _22732_ (.A(_14339_),
    .Y(_14340_));
 OAI21x1_ASAP7_75t_R _22733_ (.A1(_14327_),
    .A2(_14340_),
    .B(_07960_),
    .Y(_14341_));
 INVx2_ASAP7_75t_R _22734_ (.A(_07960_),
    .Y(_14342_));
 INVx2_ASAP7_75t_R _22735_ (.A(_14327_),
    .Y(_14343_));
 NAND3x2_ASAP7_75t_R _22736_ (.B(_14342_),
    .C(_14343_),
    .Y(_14344_),
    .A(net632));
 NAND2x2_ASAP7_75t_R _22737_ (.A(_14344_),
    .B(_14341_),
    .Y(_14345_));
 BUFx12f_ASAP7_75t_R _22738_ (.A(_14345_),
    .Y(_15891_));
 NOR2x1_ASAP7_75t_R _22739_ (.A(net680),
    .B(_00542_),
    .Y(_14346_));
 INVx2_ASAP7_75t_R _22740_ (.A(_14346_),
    .Y(_14347_));
 INVx2_ASAP7_75t_R _22741_ (.A(_11433_),
    .Y(_14348_));
 NOR2x2_ASAP7_75t_R _22742_ (.A(_14348_),
    .B(_11415_),
    .Y(_14349_));
 NOR2x2_ASAP7_75t_R _22743_ (.A(_11433_),
    .B(_11411_),
    .Y(_14350_));
 OAI21x1_ASAP7_75t_R _22744_ (.A1(_14349_),
    .A2(_14350_),
    .B(_11366_),
    .Y(_14351_));
 INVx1_ASAP7_75t_R _22745_ (.A(_14351_),
    .Y(_14352_));
 NOR3x1_ASAP7_75t_R _22746_ (.A(_14350_),
    .B(_14349_),
    .C(_11366_),
    .Y(_14353_));
 OAI21x1_ASAP7_75t_R _22747_ (.A1(_14352_),
    .A2(_14353_),
    .B(_10742_),
    .Y(_14354_));
 INVx2_ASAP7_75t_R _22748_ (.A(_08004_),
    .Y(_14355_));
 AOI21x1_ASAP7_75t_R _22749_ (.A1(_14347_),
    .A2(_14354_),
    .B(_14355_),
    .Y(_14356_));
 NAND2x2_ASAP7_75t_R _22750_ (.A(_00542_),
    .B(_10643_),
    .Y(_14357_));
 NAND2x2_ASAP7_75t_R _22751_ (.A(_14348_),
    .B(_11415_),
    .Y(_14358_));
 INVx1_ASAP7_75t_R _22752_ (.A(_11366_),
    .Y(_14359_));
 NOR2x1_ASAP7_75t_R _22753_ (.A(_11409_),
    .B(_11410_),
    .Y(_14360_));
 AND2x2_ASAP7_75t_R _22754_ (.A(_11409_),
    .B(_11410_),
    .Y(_14361_));
 OAI21x1_ASAP7_75t_R _22755_ (.A1(_14360_),
    .A2(_14361_),
    .B(_11433_),
    .Y(_14362_));
 NAND3x2_ASAP7_75t_R _22756_ (.B(_14359_),
    .C(_14362_),
    .Y(_14363_),
    .A(_14358_));
 NAND3x2_ASAP7_75t_R _22757_ (.B(_10742_),
    .C(_14351_),
    .Y(_14364_),
    .A(_14363_));
 AOI21x1_ASAP7_75t_R _22758_ (.A1(_14357_),
    .A2(_14364_),
    .B(_08004_),
    .Y(_14365_));
 NOR2x2_ASAP7_75t_R _22759_ (.A(_14365_),
    .B(_14356_),
    .Y(_14366_));
 BUFx12_ASAP7_75t_R _22760_ (.A(_14366_),
    .Y(_15899_));
 OAI21x1_ASAP7_75t_R _22761_ (.A1(_14327_),
    .A2(_14340_),
    .B(_14342_),
    .Y(_14367_));
 NAND3x2_ASAP7_75t_R _22762_ (.B(_07960_),
    .C(_14343_),
    .Y(_14368_),
    .A(_14339_));
 NAND2x2_ASAP7_75t_R _22763_ (.A(_14368_),
    .B(_14367_),
    .Y(_14369_));
 BUFx12f_ASAP7_75t_R _22764_ (.A(_14369_),
    .Y(_15886_));
 AOI21x1_ASAP7_75t_R _22765_ (.A1(_14347_),
    .A2(_14354_),
    .B(_08004_),
    .Y(_14370_));
 AOI21x1_ASAP7_75t_R _22766_ (.A1(_14357_),
    .A2(_14364_),
    .B(_14355_),
    .Y(_14371_));
 NOR2x2_ASAP7_75t_R _22767_ (.A(_14370_),
    .B(_14371_),
    .Y(_14372_));
 BUFx12f_ASAP7_75t_R _22768_ (.A(_14372_),
    .Y(_14373_));
 BUFx12_ASAP7_75t_R _22769_ (.A(_14373_),
    .Y(_15896_));
 XOR2x1_ASAP7_75t_R _22770_ (.A(_11436_),
    .Y(_14374_),
    .B(_00743_));
 XOR2x2_ASAP7_75t_R _22771_ (.A(_11409_),
    .B(net698),
    .Y(_14375_));
 XOR2x1_ASAP7_75t_R _22772_ (.A(_11437_),
    .Y(_14376_),
    .B(_14375_));
 NOR2x1_ASAP7_75t_R _22773_ (.A(_14374_),
    .B(_14376_),
    .Y(_14377_));
 XNOR2x1_ASAP7_75t_R _22774_ (.B(_11436_),
    .Y(_14378_),
    .A(_00743_));
 XNOR2x1_ASAP7_75t_R _22775_ (.B(_14375_),
    .Y(_14379_),
    .A(_11437_));
 NOR2x1_ASAP7_75t_R _22776_ (.A(_14378_),
    .B(_14379_),
    .Y(_14380_));
 OAI21x1_ASAP7_75t_R _22777_ (.A1(_14377_),
    .A2(_14380_),
    .B(net867),
    .Y(_14381_));
 NOR2x1_ASAP7_75t_R _22778_ (.A(_10742_),
    .B(_00655_),
    .Y(_14382_));
 INVx3_ASAP7_75t_R _22779_ (.A(_14382_),
    .Y(_14383_));
 NAND3x2_ASAP7_75t_R _22780_ (.B(_01037_),
    .C(_14383_),
    .Y(_14384_),
    .A(_14381_));
 AO21x2_ASAP7_75t_R _22781_ (.A1(_14381_),
    .A2(_14383_),
    .B(_01037_),
    .Y(_14385_));
 NAND2x2_ASAP7_75t_R _22782_ (.A(_14384_),
    .B(_14385_),
    .Y(_14386_));
 BUFx6f_ASAP7_75t_R _22783_ (.A(_14386_),
    .Y(_14387_));
 AOI21x1_ASAP7_75t_R _22784_ (.A1(net703),
    .A2(_15899_),
    .B(_14387_),
    .Y(_14388_));
 BUFx12f_ASAP7_75t_R _22785_ (.A(_14372_),
    .Y(_14389_));
 XNOR2x2_ASAP7_75t_R _22786_ (.A(_07970_),
    .B(_14326_),
    .Y(_14390_));
 NOR2x2_ASAP7_75t_R _22787_ (.A(_14369_),
    .B(net695),
    .Y(_14391_));
 NAND2x2_ASAP7_75t_R _22788_ (.A(_14389_),
    .B(_14391_),
    .Y(_14392_));
 INVx3_ASAP7_75t_R _22789_ (.A(_01192_),
    .Y(_14393_));
 OAI21x1_ASAP7_75t_R _22790_ (.A1(_14370_),
    .A2(_14371_),
    .B(_14393_),
    .Y(_14394_));
 BUFx10_ASAP7_75t_R _22791_ (.A(_14394_),
    .Y(_14395_));
 NAND3x2_ASAP7_75t_R _22792_ (.B(_08297_),
    .C(_14383_),
    .Y(_14396_),
    .A(_14381_));
 AO21x2_ASAP7_75t_R _22793_ (.A1(_14381_),
    .A2(_14383_),
    .B(_08297_),
    .Y(_14397_));
 NAND2x2_ASAP7_75t_R _22794_ (.A(_14396_),
    .B(_14397_),
    .Y(_14398_));
 BUFx6f_ASAP7_75t_R _22795_ (.A(_14398_),
    .Y(_14399_));
 XOR2x1_ASAP7_75t_R _22796_ (.A(_00744_),
    .Y(_14400_),
    .B(_00808_));
 XOR2x1_ASAP7_75t_R _22797_ (.A(_11465_),
    .Y(_14401_),
    .B(_14400_));
 XOR2x1_ASAP7_75t_R _22798_ (.A(_00807_),
    .Y(_14402_),
    .B(net28));
 XOR2x2_ASAP7_75t_R _22799_ (.A(_14402_),
    .B(_00840_),
    .Y(_14403_));
 XOR2x1_ASAP7_75t_R _22800_ (.A(_14401_),
    .Y(_14404_),
    .B(_14403_));
 AND2x2_ASAP7_75t_R _22801_ (.A(_12095_),
    .B(_00654_),
    .Y(_14405_));
 AOI21x1_ASAP7_75t_R _22802_ (.A1(_10787_),
    .A2(_14404_),
    .B(_14405_),
    .Y(_14406_));
 XOR2x2_ASAP7_75t_R _22803_ (.A(_14406_),
    .B(_01039_),
    .Y(_14407_));
 OAI21x1_ASAP7_75t_R _22804_ (.A1(_14395_),
    .A2(_14399_),
    .B(_14407_),
    .Y(_14408_));
 AOI21x1_ASAP7_75t_R _22805_ (.A1(_14388_),
    .A2(_14392_),
    .B(_14408_),
    .Y(_14409_));
 BUFx12_ASAP7_75t_R _22806_ (.A(_14398_),
    .Y(_14410_));
 BUFx6f_ASAP7_75t_R _22807_ (.A(_14410_),
    .Y(_14411_));
 OAI21x1_ASAP7_75t_R _22808_ (.A1(_14356_),
    .A2(_14365_),
    .B(net464),
    .Y(_14412_));
 BUFx6f_ASAP7_75t_R _22809_ (.A(_14407_),
    .Y(_14413_));
 AO21x1_ASAP7_75t_R _22810_ (.A1(_14411_),
    .A2(net54),
    .B(_14413_),
    .Y(_14414_));
 INVx3_ASAP7_75t_R _22811_ (.A(_01193_),
    .Y(_14415_));
 NAND2x2_ASAP7_75t_R _22812_ (.A(_14415_),
    .B(_14373_),
    .Y(_14416_));
 BUFx6f_ASAP7_75t_R _22813_ (.A(_14410_),
    .Y(_14417_));
 AOI21x1_ASAP7_75t_R _22814_ (.A1(_14395_),
    .A2(_14416_),
    .B(_14417_),
    .Y(_14418_));
 NOR2x1_ASAP7_75t_R _22815_ (.A(_11450_),
    .B(_00653_),
    .Y(_14419_));
 XOR2x1_ASAP7_75t_R _22816_ (.A(_00808_),
    .Y(_14420_),
    .B(_00809_));
 XOR2x1_ASAP7_75t_R _22817_ (.A(_14420_),
    .Y(_14421_),
    .B(_11485_));
 XNOR2x1_ASAP7_75t_R _22818_ (.B(_00776_),
    .Y(_14422_),
    .A(_00745_));
 AND2x2_ASAP7_75t_R _22819_ (.A(_14421_),
    .B(_14422_),
    .Y(_14423_));
 NOR2x1_ASAP7_75t_R _22820_ (.A(_14422_),
    .B(_14421_),
    .Y(_14424_));
 OA21x2_ASAP7_75t_R _22821_ (.A1(_14423_),
    .A2(_14424_),
    .B(_10761_),
    .Y(_14425_));
 NOR2x1_ASAP7_75t_R _22822_ (.A(_14419_),
    .B(_14425_),
    .Y(_14426_));
 XOR2x2_ASAP7_75t_R _22823_ (.A(_14426_),
    .B(_01040_),
    .Y(_14427_));
 INVx6_ASAP7_75t_R _22824_ (.A(_14427_),
    .Y(_14428_));
 BUFx6f_ASAP7_75t_R _22825_ (.A(_14428_),
    .Y(_14429_));
 OAI21x1_ASAP7_75t_R _22826_ (.A1(_14414_),
    .A2(_14418_),
    .B(_14429_),
    .Y(_14430_));
 NOR2x1_ASAP7_75t_R _22827_ (.A(_14409_),
    .B(_14430_),
    .Y(_14431_));
 INVx2_ASAP7_75t_R _22828_ (.A(_01191_),
    .Y(_14432_));
 NAND2x2_ASAP7_75t_R _22829_ (.A(_14432_),
    .B(_14373_),
    .Y(_14433_));
 INVx2_ASAP7_75t_R _22830_ (.A(_14370_),
    .Y(_14434_));
 INVx2_ASAP7_75t_R _22831_ (.A(_14371_),
    .Y(_14435_));
 INVx1_ASAP7_75t_R _22832_ (.A(_00543_),
    .Y(_14436_));
 AOI21x1_ASAP7_75t_R _22833_ (.A1(_14434_),
    .A2(_14435_),
    .B(_14436_),
    .Y(_14437_));
 INVx1_ASAP7_75t_R _22834_ (.A(_14437_),
    .Y(_14438_));
 BUFx6f_ASAP7_75t_R _22835_ (.A(_14410_),
    .Y(_14439_));
 AOI21x1_ASAP7_75t_R _22836_ (.A1(_14433_),
    .A2(_14438_),
    .B(_14439_),
    .Y(_14440_));
 INVx1_ASAP7_75t_R _22837_ (.A(_14356_),
    .Y(_14441_));
 NAND3x1_ASAP7_75t_R _22838_ (.A(_14354_),
    .B(_14355_),
    .C(_14347_),
    .Y(_14442_));
 AOI21x1_ASAP7_75t_R _22839_ (.A1(_14441_),
    .A2(_14442_),
    .B(_14393_),
    .Y(_14443_));
 INVx1_ASAP7_75t_R _22840_ (.A(_14443_),
    .Y(_14444_));
 BUFx4f_ASAP7_75t_R _22841_ (.A(_14407_),
    .Y(_14445_));
 AO21x1_ASAP7_75t_R _22842_ (.A1(_14444_),
    .A2(_14417_),
    .B(_14445_),
    .Y(_14446_));
 BUFx10_ASAP7_75t_R _22843_ (.A(_14427_),
    .Y(_14447_));
 OAI21x1_ASAP7_75t_R _22844_ (.A1(_14440_),
    .A2(_14446_),
    .B(_14447_),
    .Y(_14448_));
 NOR2x2_ASAP7_75t_R _22845_ (.A(_15886_),
    .B(net706),
    .Y(_14449_));
 INVx2_ASAP7_75t_R _22846_ (.A(_00541_),
    .Y(_14450_));
 NOR2x2_ASAP7_75t_R _22847_ (.A(_14450_),
    .B(_14389_),
    .Y(_14451_));
 OA21x2_ASAP7_75t_R _22848_ (.A1(_14449_),
    .A2(_14451_),
    .B(_14411_),
    .Y(_14452_));
 BUFx12f_ASAP7_75t_R _22849_ (.A(_14366_),
    .Y(_14453_));
 OAI21x1_ASAP7_75t_R _22850_ (.A1(_14370_),
    .A2(_14371_),
    .B(net465),
    .Y(_14454_));
 OAI21x1_ASAP7_75t_R _22851_ (.A1(net721),
    .A2(_14453_),
    .B(_14454_),
    .Y(_14455_));
 BUFx4f_ASAP7_75t_R _22852_ (.A(_14386_),
    .Y(_14456_));
 XOR2x2_ASAP7_75t_R _22853_ (.A(_14406_),
    .B(_07992_),
    .Y(_14457_));
 BUFx4f_ASAP7_75t_R _22854_ (.A(_14457_),
    .Y(_14458_));
 AO21x1_ASAP7_75t_R _22855_ (.A1(_14455_),
    .A2(_14456_),
    .B(_14458_),
    .Y(_14459_));
 NOR2x1_ASAP7_75t_R _22856_ (.A(_14452_),
    .B(_14459_),
    .Y(_14460_));
 XOR2x2_ASAP7_75t_R _22857_ (.A(_00810_),
    .B(_00842_),
    .Y(_14461_));
 XOR2x1_ASAP7_75t_R _22858_ (.A(_11487_),
    .Y(_14462_),
    .B(_00746_));
 XNOR2x1_ASAP7_75t_R _22859_ (.B(_14462_),
    .Y(_14463_),
    .A(_14461_));
 NOR2x1_ASAP7_75t_R _22860_ (.A(_10786_),
    .B(_00652_),
    .Y(_14464_));
 AO21x1_ASAP7_75t_R _22861_ (.A1(_14463_),
    .A2(_13017_),
    .B(_14464_),
    .Y(_14465_));
 XOR2x2_ASAP7_75t_R _22862_ (.A(_14465_),
    .B(_01041_),
    .Y(_14466_));
 CKINVDCx5p33_ASAP7_75t_R _22863_ (.A(_14466_),
    .Y(_14467_));
 BUFx10_ASAP7_75t_R _22864_ (.A(_14467_),
    .Y(_14468_));
 OAI21x1_ASAP7_75t_R _22865_ (.A1(_14448_),
    .A2(_14460_),
    .B(_14468_),
    .Y(_14469_));
 XOR2x1_ASAP7_75t_R _22866_ (.A(_00810_),
    .Y(_14470_),
    .B(net28));
 XOR2x1_ASAP7_75t_R _22867_ (.A(_14470_),
    .Y(_14471_),
    .B(_11537_));
 XOR2x1_ASAP7_75t_R _22868_ (.A(_11363_),
    .Y(_14472_),
    .B(_00778_));
 XOR2x1_ASAP7_75t_R _22869_ (.A(_14471_),
    .Y(_14473_),
    .B(_14472_));
 NOR2x1_ASAP7_75t_R _22870_ (.A(_13017_),
    .B(_00651_),
    .Y(_14474_));
 AO21x1_ASAP7_75t_R _22871_ (.A1(_14473_),
    .A2(_10831_),
    .B(_14474_),
    .Y(_14475_));
 XOR2x2_ASAP7_75t_R _22872_ (.A(_14475_),
    .B(_01042_),
    .Y(_14476_));
 CKINVDCx6p67_ASAP7_75t_R _22873_ (.A(_14476_),
    .Y(_14477_));
 OAI21x1_ASAP7_75t_R _22874_ (.A1(_14431_),
    .A2(_14469_),
    .B(_14477_),
    .Y(_14478_));
 BUFx10_ASAP7_75t_R _22875_ (.A(_14413_),
    .Y(_14479_));
 NOR2x2_ASAP7_75t_R _22876_ (.A(net760),
    .B(net692),
    .Y(_14480_));
 NAND2x2_ASAP7_75t_R _22877_ (.A(_14389_),
    .B(_14480_),
    .Y(_14481_));
 AOI21x1_ASAP7_75t_R _22878_ (.A1(_14434_),
    .A2(_14435_),
    .B(_14415_),
    .Y(_14482_));
 NOR2x2_ASAP7_75t_R _22879_ (.A(_14386_),
    .B(_14482_),
    .Y(_14483_));
 BUFx6f_ASAP7_75t_R _22880_ (.A(_14386_),
    .Y(_14484_));
 BUFx6f_ASAP7_75t_R _22881_ (.A(_14484_),
    .Y(_14485_));
 NOR2x2_ASAP7_75t_R _22882_ (.A(_01191_),
    .B(net706),
    .Y(_14486_));
 AOI22x1_ASAP7_75t_R _22883_ (.A1(_14481_),
    .A2(_14483_),
    .B1(_14485_),
    .B2(_14486_),
    .Y(_14487_));
 BUFx6f_ASAP7_75t_R _22884_ (.A(_14410_),
    .Y(_14488_));
 AO21x1_ASAP7_75t_R _22885_ (.A1(_14486_),
    .A2(_14488_),
    .B(_14413_),
    .Y(_14489_));
 NAND2x2_ASAP7_75t_R _22886_ (.A(_15886_),
    .B(net720),
    .Y(_14490_));
 NOR2x1_ASAP7_75t_R _22887_ (.A(_15899_),
    .B(_14490_),
    .Y(_14491_));
 NAND2x2_ASAP7_75t_R _22888_ (.A(_14450_),
    .B(_14453_),
    .Y(_14492_));
 NAND2x2_ASAP7_75t_R _22889_ (.A(_14484_),
    .B(_14492_),
    .Y(_14493_));
 NOR2x1_ASAP7_75t_R _22890_ (.A(_14491_),
    .B(_14493_),
    .Y(_14494_));
 BUFx6f_ASAP7_75t_R _22891_ (.A(_14427_),
    .Y(_14495_));
 OAI21x1_ASAP7_75t_R _22892_ (.A1(_14489_),
    .A2(_14494_),
    .B(_14495_),
    .Y(_14496_));
 AOI21x1_ASAP7_75t_R _22893_ (.A1(_14479_),
    .A2(_14487_),
    .B(_14496_),
    .Y(_14497_));
 BUFx4f_ASAP7_75t_R _22894_ (.A(_14398_),
    .Y(_14498_));
 INVx3_ASAP7_75t_R _22895_ (.A(net464),
    .Y(_14499_));
 OAI21x1_ASAP7_75t_R _22896_ (.A1(_14370_),
    .A2(_14371_),
    .B(_14499_),
    .Y(_14500_));
 BUFx6f_ASAP7_75t_R _22897_ (.A(_14457_),
    .Y(_14501_));
 OA21x2_ASAP7_75t_R _22898_ (.A1(_14500_),
    .A2(_14498_),
    .B(_14501_),
    .Y(_14502_));
 AO21x1_ASAP7_75t_R _22899_ (.A1(_14397_),
    .A2(_14396_),
    .B(_01196_),
    .Y(_14503_));
 AO21x1_ASAP7_75t_R _22900_ (.A1(_14503_),
    .A2(_14502_),
    .B(_14495_),
    .Y(_14504_));
 NAND2x2_ASAP7_75t_R _22901_ (.A(_01191_),
    .B(net630),
    .Y(_14505_));
 NAND2x2_ASAP7_75t_R _22902_ (.A(_14505_),
    .B(_15899_),
    .Y(_14506_));
 OAI21x1_ASAP7_75t_R _22903_ (.A1(net760),
    .A2(_14390_),
    .B(_14373_),
    .Y(_14507_));
 NAND2x1_ASAP7_75t_R _22904_ (.A(_14506_),
    .B(_14507_),
    .Y(_14508_));
 OAI21x1_ASAP7_75t_R _22905_ (.A1(_14356_),
    .A2(_14365_),
    .B(_00543_),
    .Y(_14509_));
 NAND2x2_ASAP7_75t_R _22906_ (.A(net760),
    .B(_14366_),
    .Y(_14510_));
 AOI21x1_ASAP7_75t_R _22907_ (.A1(_14509_),
    .A2(_14510_),
    .B(_14456_),
    .Y(_14511_));
 BUFx6f_ASAP7_75t_R _22908_ (.A(_14501_),
    .Y(_14512_));
 AOI211x1_ASAP7_75t_R _22909_ (.A1(_14508_),
    .A2(_14485_),
    .B(_14511_),
    .C(_14512_),
    .Y(_14513_));
 BUFx10_ASAP7_75t_R _22910_ (.A(_14466_),
    .Y(_14514_));
 OAI21x1_ASAP7_75t_R _22911_ (.A1(_14513_),
    .A2(_14504_),
    .B(_14514_),
    .Y(_14515_));
 NOR2x1_ASAP7_75t_R _22912_ (.A(_14515_),
    .B(_14497_),
    .Y(_14516_));
 NOR2x2_ASAP7_75t_R _22913_ (.A(_15889_),
    .B(_14389_),
    .Y(_14517_));
 BUFx6f_ASAP7_75t_R _22914_ (.A(_14386_),
    .Y(_14518_));
 OA21x2_ASAP7_75t_R _22915_ (.A1(_14486_),
    .A2(_14517_),
    .B(_14518_),
    .Y(_14519_));
 NAND2x2_ASAP7_75t_R _22916_ (.A(_15891_),
    .B(net720),
    .Y(_14520_));
 NOR2x2_ASAP7_75t_R _22917_ (.A(_14453_),
    .B(_14520_),
    .Y(_14521_));
 NAND2x2_ASAP7_75t_R _22918_ (.A(net703),
    .B(net706),
    .Y(_14522_));
 NAND2x1_ASAP7_75t_R _22919_ (.A(_14498_),
    .B(_14522_),
    .Y(_14523_));
 OAI21x1_ASAP7_75t_R _22920_ (.A1(_14521_),
    .A2(_14523_),
    .B(_14445_),
    .Y(_14524_));
 NOR2x1_ASAP7_75t_R _22921_ (.A(_14519_),
    .B(_14524_),
    .Y(_14525_));
 NAND2x2_ASAP7_75t_R _22922_ (.A(net719),
    .B(_14373_),
    .Y(_14526_));
 OAI21x1_ASAP7_75t_R _22923_ (.A1(_15891_),
    .A2(_14390_),
    .B(_14453_),
    .Y(_14527_));
 BUFx6f_ASAP7_75t_R _22924_ (.A(_14399_),
    .Y(_14528_));
 AOI21x1_ASAP7_75t_R _22925_ (.A1(_14526_),
    .A2(_14527_),
    .B(_14528_),
    .Y(_14529_));
 NOR2x2_ASAP7_75t_R _22926_ (.A(_15891_),
    .B(_15896_),
    .Y(_14530_));
 INVx5_ASAP7_75t_R _22927_ (.A(_01194_),
    .Y(_14531_));
 BUFx6f_ASAP7_75t_R _22928_ (.A(_14410_),
    .Y(_14532_));
 OAI21x1_ASAP7_75t_R _22929_ (.A1(_14531_),
    .A2(_15899_),
    .B(_14532_),
    .Y(_14533_));
 BUFx10_ASAP7_75t_R _22930_ (.A(_14457_),
    .Y(_14534_));
 OAI21x1_ASAP7_75t_R _22931_ (.A1(_14530_),
    .A2(_14533_),
    .B(_14534_),
    .Y(_14535_));
 OAI21x1_ASAP7_75t_R _22932_ (.A1(_14529_),
    .A2(_14535_),
    .B(_14429_),
    .Y(_14536_));
 NOR2x1_ASAP7_75t_R _22933_ (.A(_14525_),
    .B(_14536_),
    .Y(_14537_));
 NAND2x2_ASAP7_75t_R _22934_ (.A(_14393_),
    .B(_14373_),
    .Y(_14538_));
 AOI21x1_ASAP7_75t_R _22935_ (.A1(_14538_),
    .A2(_14527_),
    .B(_14485_),
    .Y(_14539_));
 AO21x1_ASAP7_75t_R _22936_ (.A1(_14522_),
    .A2(_14456_),
    .B(_14458_),
    .Y(_14540_));
 OAI21x1_ASAP7_75t_R _22937_ (.A1(_14539_),
    .A2(_14540_),
    .B(_14447_),
    .Y(_14541_));
 BUFx6f_ASAP7_75t_R _22938_ (.A(_14390_),
    .Y(_15887_));
 AO21x1_ASAP7_75t_R _22939_ (.A1(_15899_),
    .A2(net56),
    .B(_15891_),
    .Y(_14542_));
 AOI21x1_ASAP7_75t_R _22940_ (.A1(_14434_),
    .A2(_14435_),
    .B(_14531_),
    .Y(_14543_));
 NAND2x2_ASAP7_75t_R _22941_ (.A(_14412_),
    .B(_14398_),
    .Y(_14544_));
 OAI21x1_ASAP7_75t_R _22942_ (.A1(_14543_),
    .A2(_14544_),
    .B(_14534_),
    .Y(_14545_));
 AOI21x1_ASAP7_75t_R _22943_ (.A1(_14485_),
    .A2(_14542_),
    .B(_14545_),
    .Y(_14546_));
 OAI21x1_ASAP7_75t_R _22944_ (.A1(_14541_),
    .A2(_14546_),
    .B(_14468_),
    .Y(_14547_));
 OAI21x1_ASAP7_75t_R _22945_ (.A1(_14537_),
    .A2(_14547_),
    .B(_14476_),
    .Y(_14548_));
 NOR2x2_ASAP7_75t_R _22946_ (.A(net575),
    .B(_15896_),
    .Y(_14549_));
 NOR2x1_ASAP7_75t_R _22947_ (.A(_14549_),
    .B(_14544_),
    .Y(_14550_));
 INVx1_ASAP7_75t_R _22948_ (.A(_14509_),
    .Y(_14551_));
 BUFx6f_ASAP7_75t_R _22949_ (.A(_14386_),
    .Y(_14552_));
 OA21x2_ASAP7_75t_R _22950_ (.A1(_14451_),
    .A2(_14551_),
    .B(_14552_),
    .Y(_14553_));
 BUFx6f_ASAP7_75t_R _22951_ (.A(_14407_),
    .Y(_14554_));
 BUFx10_ASAP7_75t_R _22952_ (.A(_14554_),
    .Y(_14555_));
 OAI21x1_ASAP7_75t_R _22953_ (.A1(_14550_),
    .A2(_14553_),
    .B(_14555_),
    .Y(_14556_));
 NOR2x2_ASAP7_75t_R _22954_ (.A(_14454_),
    .B(_14518_),
    .Y(_14557_));
 NOR2x2_ASAP7_75t_R _22955_ (.A(_15887_),
    .B(_14389_),
    .Y(_14558_));
 OAI21x1_ASAP7_75t_R _22956_ (.A1(_14356_),
    .A2(_14365_),
    .B(_14499_),
    .Y(_14559_));
 INVx2_ASAP7_75t_R _22957_ (.A(_14559_),
    .Y(_14560_));
 OA21x2_ASAP7_75t_R _22958_ (.A1(_14558_),
    .A2(_14560_),
    .B(_14456_),
    .Y(_14561_));
 OAI21x1_ASAP7_75t_R _22959_ (.A1(_14557_),
    .A2(_14561_),
    .B(_14512_),
    .Y(_14562_));
 BUFx10_ASAP7_75t_R _22960_ (.A(_14427_),
    .Y(_14563_));
 BUFx6f_ASAP7_75t_R _22961_ (.A(_14563_),
    .Y(_14564_));
 AOI21x1_ASAP7_75t_R _22962_ (.A1(_14556_),
    .A2(_14562_),
    .B(_14564_),
    .Y(_14565_));
 AND3x1_ASAP7_75t_R _22963_ (.A(_14510_),
    .B(_14498_),
    .C(_14490_),
    .Y(_14566_));
 NOR2x2_ASAP7_75t_R _22964_ (.A(_15886_),
    .B(_14373_),
    .Y(_14567_));
 BUFx6f_ASAP7_75t_R _22965_ (.A(_14386_),
    .Y(_14568_));
 OAI21x1_ASAP7_75t_R _22966_ (.A1(_14480_),
    .A2(_14567_),
    .B(_14568_),
    .Y(_14569_));
 NAND2x1_ASAP7_75t_R _22967_ (.A(_14458_),
    .B(_14569_),
    .Y(_14570_));
 NOR2x1_ASAP7_75t_R _22968_ (.A(_14566_),
    .B(_14570_),
    .Y(_14571_));
 OAI21x1_ASAP7_75t_R _22969_ (.A1(net699),
    .A2(_14390_),
    .B(_14366_),
    .Y(_14572_));
 AOI21x1_ASAP7_75t_R _22970_ (.A1(net55),
    .A2(_14572_),
    .B(_14528_),
    .Y(_14573_));
 OA21x2_ASAP7_75t_R _22971_ (.A1(_14365_),
    .A2(_14356_),
    .B(_00541_),
    .Y(_14574_));
 OAI21x1_ASAP7_75t_R _22972_ (.A1(_14437_),
    .A2(_14574_),
    .B(_14488_),
    .Y(_14575_));
 NAND2x1_ASAP7_75t_R _22973_ (.A(_14445_),
    .B(_14575_),
    .Y(_14576_));
 OAI21x1_ASAP7_75t_R _22974_ (.A1(_14573_),
    .A2(_14576_),
    .B(_14495_),
    .Y(_14577_));
 BUFx10_ASAP7_75t_R _22975_ (.A(_14466_),
    .Y(_14578_));
 OAI21x1_ASAP7_75t_R _22976_ (.A1(_14571_),
    .A2(_14577_),
    .B(_14578_),
    .Y(_14579_));
 NOR2x1_ASAP7_75t_R _22977_ (.A(_14565_),
    .B(_14579_),
    .Y(_14580_));
 OAI22x1_ASAP7_75t_R _22978_ (.A1(_14516_),
    .A2(_14478_),
    .B1(_14548_),
    .B2(_14580_),
    .Y(_00072_));
 OAI21x1_ASAP7_75t_R _22979_ (.A1(net703),
    .A2(net56),
    .B(_14389_),
    .Y(_14581_));
 AO21x1_ASAP7_75t_R _22980_ (.A1(_14581_),
    .A2(_14527_),
    .B(_14518_),
    .Y(_14582_));
 NAND2x2_ASAP7_75t_R _22981_ (.A(_15891_),
    .B(_14373_),
    .Y(_14583_));
 AO21x1_ASAP7_75t_R _22982_ (.A1(_14438_),
    .A2(_14583_),
    .B(_14532_),
    .Y(_14584_));
 AO21x1_ASAP7_75t_R _22983_ (.A1(_14582_),
    .A2(_14584_),
    .B(_14429_),
    .Y(_14585_));
 NOR2x1_ASAP7_75t_R _22984_ (.A(_01192_),
    .B(_14453_),
    .Y(_14586_));
 OAI21x1_ASAP7_75t_R _22985_ (.A1(_14558_),
    .A2(_14586_),
    .B(_14532_),
    .Y(_14587_));
 NAND2x2_ASAP7_75t_R _22986_ (.A(net699),
    .B(_14373_),
    .Y(_14588_));
 NAND2x2_ASAP7_75t_R _22987_ (.A(_15887_),
    .B(net706),
    .Y(_14589_));
 AO21x1_ASAP7_75t_R _22988_ (.A1(_14588_),
    .A2(_14589_),
    .B(_14399_),
    .Y(_14590_));
 NAND2x1_ASAP7_75t_R _22989_ (.A(_14587_),
    .B(_14590_),
    .Y(_14591_));
 AOI21x1_ASAP7_75t_R _22990_ (.A1(_14429_),
    .A2(_14591_),
    .B(_14555_),
    .Y(_14592_));
 NOR2x2_ASAP7_75t_R _22991_ (.A(_14521_),
    .B(_14493_),
    .Y(_14593_));
 AND3x1_ASAP7_75t_R _22992_ (.A(_14385_),
    .B(_14384_),
    .C(_00545_),
    .Y(_14594_));
 AO21x1_ASAP7_75t_R _22993_ (.A1(_14428_),
    .A2(_14594_),
    .B(_14458_),
    .Y(_14595_));
 OAI21x1_ASAP7_75t_R _22994_ (.A1(_14593_),
    .A2(_14595_),
    .B(_14514_),
    .Y(_14596_));
 AOI21x1_ASAP7_75t_R _22995_ (.A1(_14585_),
    .A2(_14592_),
    .B(_14596_),
    .Y(_14597_));
 OAI21x1_ASAP7_75t_R _22996_ (.A1(_14370_),
    .A2(_14371_),
    .B(_14432_),
    .Y(_14598_));
 OAI21x1_ASAP7_75t_R _22997_ (.A1(_14356_),
    .A2(_14365_),
    .B(_14531_),
    .Y(_14599_));
 NAND2x1_ASAP7_75t_R _22998_ (.A(_14598_),
    .B(_14599_),
    .Y(_14600_));
 AOI21x1_ASAP7_75t_R _22999_ (.A1(_14568_),
    .A2(_14600_),
    .B(_14554_),
    .Y(_14601_));
 AO21x1_ASAP7_75t_R _23000_ (.A1(_14572_),
    .A2(_14412_),
    .B(_14387_),
    .Y(_14602_));
 NAND2x1_ASAP7_75t_R _23001_ (.A(_14601_),
    .B(_14602_),
    .Y(_14603_));
 INVx2_ASAP7_75t_R _23002_ (.A(_14412_),
    .Y(_14604_));
 NOR2x1_ASAP7_75t_R _23003_ (.A(_14387_),
    .B(_14604_),
    .Y(_14605_));
 NOR2x1_ASAP7_75t_R _23004_ (.A(_14501_),
    .B(_14605_),
    .Y(_14606_));
 AOI21x1_ASAP7_75t_R _23005_ (.A1(_15889_),
    .A2(_15891_),
    .B(_14453_),
    .Y(_14607_));
 OAI21x1_ASAP7_75t_R _23006_ (.A1(_14567_),
    .A2(_14607_),
    .B(_14552_),
    .Y(_14608_));
 AOI21x1_ASAP7_75t_R _23007_ (.A1(_14606_),
    .A2(_14608_),
    .B(_14563_),
    .Y(_14609_));
 NAND2x1_ASAP7_75t_R _23008_ (.A(_14603_),
    .B(_14609_),
    .Y(_14610_));
 AO21x1_ASAP7_75t_R _23009_ (.A1(_14500_),
    .A2(_14509_),
    .B(_14568_),
    .Y(_14611_));
 OAI21x1_ASAP7_75t_R _23010_ (.A1(_14567_),
    .A2(_14486_),
    .B(_14552_),
    .Y(_14612_));
 BUFx6f_ASAP7_75t_R _23011_ (.A(_14407_),
    .Y(_14613_));
 AOI21x1_ASAP7_75t_R _23012_ (.A1(_14611_),
    .A2(_14612_),
    .B(_14613_),
    .Y(_14614_));
 NOR2x2_ASAP7_75t_R _23013_ (.A(_15891_),
    .B(_14453_),
    .Y(_14615_));
 OAI21x1_ASAP7_75t_R _23014_ (.A1(_14437_),
    .A2(_14615_),
    .B(_14552_),
    .Y(_14616_));
 AOI21x1_ASAP7_75t_R _23015_ (.A1(_14616_),
    .A2(_14587_),
    .B(_14534_),
    .Y(_14617_));
 OAI21x1_ASAP7_75t_R _23016_ (.A1(_14614_),
    .A2(_14617_),
    .B(_14447_),
    .Y(_14618_));
 AOI21x1_ASAP7_75t_R _23017_ (.A1(_14610_),
    .A2(_14618_),
    .B(_14514_),
    .Y(_14619_));
 OAI21x1_ASAP7_75t_R _23018_ (.A1(_14597_),
    .A2(_14619_),
    .B(_14476_),
    .Y(_14620_));
 AO21x1_ASAP7_75t_R _23019_ (.A1(_14510_),
    .A2(_14559_),
    .B(_14484_),
    .Y(_14621_));
 NOR2x2_ASAP7_75t_R _23020_ (.A(_14410_),
    .B(_14443_),
    .Y(_14622_));
 AOI21x1_ASAP7_75t_R _23021_ (.A1(_14510_),
    .A2(_14622_),
    .B(_14554_),
    .Y(_14623_));
 NAND2x1_ASAP7_75t_R _23022_ (.A(_14621_),
    .B(_14623_),
    .Y(_14624_));
 NAND2x1_ASAP7_75t_R _23023_ (.A(_15891_),
    .B(_15887_),
    .Y(_14625_));
 NAND2x2_ASAP7_75t_R _23024_ (.A(net718),
    .B(net706),
    .Y(_14626_));
 AOI21x1_ASAP7_75t_R _23025_ (.A1(_14625_),
    .A2(_14626_),
    .B(_14410_),
    .Y(_14627_));
 INVx1_ASAP7_75t_R _23026_ (.A(_14627_),
    .Y(_14628_));
 NOR2x1_ASAP7_75t_R _23027_ (.A(_15896_),
    .B(_14387_),
    .Y(_14629_));
 AOI21x1_ASAP7_75t_R _23028_ (.A1(_14490_),
    .A2(_14629_),
    .B(_14501_),
    .Y(_14630_));
 AOI21x1_ASAP7_75t_R _23029_ (.A1(_14628_),
    .A2(_14630_),
    .B(_14428_),
    .Y(_14631_));
 NAND2x1_ASAP7_75t_R _23030_ (.A(_14624_),
    .B(_14631_),
    .Y(_14632_));
 NAND2x1_ASAP7_75t_R _23031_ (.A(_14599_),
    .B(_14500_),
    .Y(_14633_));
 AOI21x1_ASAP7_75t_R _23032_ (.A1(_14532_),
    .A2(_14633_),
    .B(_14501_),
    .Y(_14634_));
 AOI21x1_ASAP7_75t_R _23033_ (.A1(_14394_),
    .A2(_14507_),
    .B(_14410_),
    .Y(_14635_));
 INVx1_ASAP7_75t_R _23034_ (.A(_14635_),
    .Y(_14636_));
 NAND2x1_ASAP7_75t_R _23035_ (.A(_14636_),
    .B(_14634_),
    .Y(_14637_));
 NAND2x2_ASAP7_75t_R _23036_ (.A(net693),
    .B(_14373_),
    .Y(_14638_));
 BUFx6f_ASAP7_75t_R _23037_ (.A(_14638_),
    .Y(_14639_));
 AO21x1_ASAP7_75t_R _23038_ (.A1(_14639_),
    .A2(_14395_),
    .B(_14498_),
    .Y(_14640_));
 NOR2x2_ASAP7_75t_R _23039_ (.A(_14453_),
    .B(_14386_),
    .Y(_14641_));
 OAI21x1_ASAP7_75t_R _23040_ (.A1(net720),
    .A2(_14387_),
    .B(_14457_),
    .Y(_14642_));
 NOR2x1_ASAP7_75t_R _23041_ (.A(_14641_),
    .B(_14642_),
    .Y(_14643_));
 AOI21x1_ASAP7_75t_R _23042_ (.A1(_14640_),
    .A2(_14643_),
    .B(_14563_),
    .Y(_14644_));
 NAND2x1_ASAP7_75t_R _23043_ (.A(_14637_),
    .B(_14644_),
    .Y(_14645_));
 AOI21x1_ASAP7_75t_R _23044_ (.A1(_14632_),
    .A2(_14645_),
    .B(_14467_),
    .Y(_14646_));
 AO21x1_ASAP7_75t_R _23045_ (.A1(_14395_),
    .A2(_14412_),
    .B(_14568_),
    .Y(_14647_));
 OAI21x1_ASAP7_75t_R _23046_ (.A1(_14551_),
    .A2(_14567_),
    .B(_14552_),
    .Y(_14648_));
 AOI21x1_ASAP7_75t_R _23047_ (.A1(_14647_),
    .A2(_14648_),
    .B(_14613_),
    .Y(_14649_));
 OAI21x1_ASAP7_75t_R _23048_ (.A1(_14391_),
    .A2(_14615_),
    .B(_14411_),
    .Y(_14650_));
 INVx3_ASAP7_75t_R _23049_ (.A(_14454_),
    .Y(_14651_));
 OAI21x1_ASAP7_75t_R _23050_ (.A1(_14651_),
    .A2(_14449_),
    .B(_14552_),
    .Y(_14652_));
 AOI21x1_ASAP7_75t_R _23051_ (.A1(_14650_),
    .A2(_14652_),
    .B(_14534_),
    .Y(_14653_));
 BUFx10_ASAP7_75t_R _23052_ (.A(_14428_),
    .Y(_14654_));
 OAI21x1_ASAP7_75t_R _23053_ (.A1(_14649_),
    .A2(_14653_),
    .B(_14654_),
    .Y(_14655_));
 OA21x2_ASAP7_75t_R _23054_ (.A1(_14538_),
    .A2(_14399_),
    .B(_14407_),
    .Y(_14656_));
 NAND2x1_ASAP7_75t_R _23055_ (.A(_14656_),
    .B(_14602_),
    .Y(_14657_));
 NAND2x1_ASAP7_75t_R _23056_ (.A(_14518_),
    .B(_14607_),
    .Y(_14658_));
 NOR2x2_ASAP7_75t_R _23057_ (.A(_14387_),
    .B(_14543_),
    .Y(_14659_));
 AOI21x1_ASAP7_75t_R _23058_ (.A1(_14639_),
    .A2(_14659_),
    .B(_14413_),
    .Y(_14660_));
 AOI21x1_ASAP7_75t_R _23059_ (.A1(_14658_),
    .A2(_14660_),
    .B(_14428_),
    .Y(_14661_));
 NAND2x1_ASAP7_75t_R _23060_ (.A(_14657_),
    .B(_14661_),
    .Y(_14662_));
 AOI21x1_ASAP7_75t_R _23061_ (.A1(_14655_),
    .A2(_14662_),
    .B(_14514_),
    .Y(_14663_));
 OAI21x1_ASAP7_75t_R _23062_ (.A1(_14646_),
    .A2(_14663_),
    .B(_14477_),
    .Y(_14664_));
 NAND2x1_ASAP7_75t_R _23063_ (.A(_14620_),
    .B(_14664_),
    .Y(_00073_));
 NAND2x2_ASAP7_75t_R _23064_ (.A(_14531_),
    .B(net706),
    .Y(_14665_));
 AOI21x1_ASAP7_75t_R _23065_ (.A1(_14665_),
    .A2(_14538_),
    .B(_14498_),
    .Y(_14666_));
 INVx1_ASAP7_75t_R _23066_ (.A(_14666_),
    .Y(_14667_));
 OAI21x1_ASAP7_75t_R _23067_ (.A1(net56),
    .A2(_14567_),
    .B(_14411_),
    .Y(_14668_));
 AO21x1_ASAP7_75t_R _23068_ (.A1(_14667_),
    .A2(_14668_),
    .B(_14613_),
    .Y(_14669_));
 NAND3x2_ASAP7_75t_R _23069_ (.B(_14411_),
    .C(_14395_),
    .Y(_14670_),
    .A(_14507_));
 BUFx6f_ASAP7_75t_R _23070_ (.A(_14387_),
    .Y(_14671_));
 NAND2x1_ASAP7_75t_R _23071_ (.A(_14671_),
    .B(_14455_),
    .Y(_14672_));
 NAND3x1_ASAP7_75t_R _23072_ (.A(_14670_),
    .B(_14555_),
    .C(_14672_),
    .Y(_14673_));
 AOI21x1_ASAP7_75t_R _23073_ (.A1(_14669_),
    .A2(_14673_),
    .B(_14564_),
    .Y(_14674_));
 NAND2x1_ASAP7_75t_R _23074_ (.A(_14599_),
    .B(_14572_),
    .Y(_14675_));
 BUFx6f_ASAP7_75t_R _23075_ (.A(_14399_),
    .Y(_14676_));
 OAI21x1_ASAP7_75t_R _23076_ (.A1(_15896_),
    .A2(_14490_),
    .B(_14518_),
    .Y(_14677_));
 INVx1_ASAP7_75t_R _23077_ (.A(_14677_),
    .Y(_14678_));
 AOI211x1_ASAP7_75t_R _23078_ (.A1(_14675_),
    .A2(_14676_),
    .B(_14678_),
    .C(_14512_),
    .Y(_14679_));
 AOI21x1_ASAP7_75t_R _23079_ (.A1(net54),
    .A2(_14626_),
    .B(_14488_),
    .Y(_14680_));
 NAND2x1_ASAP7_75t_R _23080_ (.A(_01191_),
    .B(_15899_),
    .Y(_14681_));
 AOI21x1_ASAP7_75t_R _23081_ (.A1(_14588_),
    .A2(_14681_),
    .B(_14552_),
    .Y(_14682_));
 OAI21x1_ASAP7_75t_R _23082_ (.A1(_14680_),
    .A2(_14682_),
    .B(_14534_),
    .Y(_14683_));
 NAND2x1_ASAP7_75t_R _23083_ (.A(_14495_),
    .B(_14683_),
    .Y(_14684_));
 OAI21x1_ASAP7_75t_R _23084_ (.A1(_14679_),
    .A2(_14684_),
    .B(_14578_),
    .Y(_14685_));
 OAI21x1_ASAP7_75t_R _23085_ (.A1(_14674_),
    .A2(_14685_),
    .B(_14476_),
    .Y(_14686_));
 NAND2x2_ASAP7_75t_R _23086_ (.A(_14415_),
    .B(_15899_),
    .Y(_14687_));
 AOI21x1_ASAP7_75t_R _23087_ (.A1(_14583_),
    .A2(_14687_),
    .B(_14439_),
    .Y(_14688_));
 INVx2_ASAP7_75t_R _23088_ (.A(_14500_),
    .Y(_14689_));
 NOR2x1_ASAP7_75t_R _23089_ (.A(_14689_),
    .B(_14544_),
    .Y(_14690_));
 OAI21x1_ASAP7_75t_R _23090_ (.A1(_14688_),
    .A2(_14690_),
    .B(_14555_),
    .Y(_14691_));
 NOR2x2_ASAP7_75t_R _23091_ (.A(net707),
    .B(_14453_),
    .Y(_14692_));
 OA21x2_ASAP7_75t_R _23092_ (.A1(_14692_),
    .A2(_14517_),
    .B(_14417_),
    .Y(_14693_));
 NOR2x1_ASAP7_75t_R _23093_ (.A(_01194_),
    .B(_14389_),
    .Y(_14694_));
 OA21x2_ASAP7_75t_R _23094_ (.A1(_14449_),
    .A2(_14694_),
    .B(_14456_),
    .Y(_14695_));
 BUFx10_ASAP7_75t_R _23095_ (.A(_14501_),
    .Y(_14696_));
 OAI21x1_ASAP7_75t_R _23096_ (.A1(_14693_),
    .A2(_14695_),
    .B(_14696_),
    .Y(_14697_));
 AOI21x1_ASAP7_75t_R _23097_ (.A1(_14691_),
    .A2(_14697_),
    .B(_14654_),
    .Y(_14698_));
 AOI21x1_ASAP7_75t_R _23098_ (.A1(_14395_),
    .A2(_14526_),
    .B(_14671_),
    .Y(_14699_));
 OAI21x1_ASAP7_75t_R _23099_ (.A1(_14418_),
    .A2(_14699_),
    .B(_14613_),
    .Y(_14700_));
 AOI21x1_ASAP7_75t_R _23100_ (.A1(_14395_),
    .A2(_14583_),
    .B(_14671_),
    .Y(_14701_));
 AOI21x1_ASAP7_75t_R _23101_ (.A1(_14416_),
    .A2(_14665_),
    .B(_14528_),
    .Y(_14702_));
 OAI21x1_ASAP7_75t_R _23102_ (.A1(_14701_),
    .A2(_14702_),
    .B(_14512_),
    .Y(_14703_));
 AOI21x1_ASAP7_75t_R _23103_ (.A1(_14700_),
    .A2(_14703_),
    .B(_14447_),
    .Y(_14704_));
 NOR3x1_ASAP7_75t_R _23104_ (.A(_14698_),
    .B(_14578_),
    .C(_14704_),
    .Y(_14705_));
 NAND2x2_ASAP7_75t_R _23105_ (.A(_14505_),
    .B(_14389_),
    .Y(_14706_));
 AOI21x1_ASAP7_75t_R _23106_ (.A1(_14706_),
    .A2(_14572_),
    .B(_14485_),
    .Y(_14707_));
 NOR2x2_ASAP7_75t_R _23107_ (.A(net759),
    .B(_14389_),
    .Y(_14708_));
 NOR2x1_ASAP7_75t_R _23108_ (.A(_14399_),
    .B(_14708_),
    .Y(_14709_));
 AO21x1_ASAP7_75t_R _23109_ (.A1(_14709_),
    .A2(_14392_),
    .B(_14445_),
    .Y(_14710_));
 AO21x1_ASAP7_75t_R _23110_ (.A1(_14395_),
    .A2(_14559_),
    .B(_14568_),
    .Y(_14711_));
 OA21x2_ASAP7_75t_R _23111_ (.A1(_14498_),
    .A2(_14509_),
    .B(_14554_),
    .Y(_14712_));
 AOI21x1_ASAP7_75t_R _23112_ (.A1(_14711_),
    .A2(_14712_),
    .B(_14429_),
    .Y(_14713_));
 OAI21x1_ASAP7_75t_R _23113_ (.A1(_14707_),
    .A2(_14710_),
    .B(_14713_),
    .Y(_14714_));
 OA21x2_ASAP7_75t_R _23114_ (.A1(_14498_),
    .A2(_01198_),
    .B(_14501_),
    .Y(_14715_));
 AOI21x1_ASAP7_75t_R _23115_ (.A1(_14668_),
    .A2(_14715_),
    .B(_14563_),
    .Y(_14716_));
 NAND2x1_ASAP7_75t_R _23116_ (.A(_00546_),
    .B(_14498_),
    .Y(_14717_));
 NAND3x1_ASAP7_75t_R _23117_ (.A(_14677_),
    .B(_14613_),
    .C(_14717_),
    .Y(_14718_));
 AOI21x1_ASAP7_75t_R _23118_ (.A1(_14716_),
    .A2(_14718_),
    .B(_14467_),
    .Y(_14719_));
 AOI21x1_ASAP7_75t_R _23119_ (.A1(_14714_),
    .A2(_14719_),
    .B(_14476_),
    .Y(_14720_));
 AO21x1_ASAP7_75t_R _23120_ (.A1(_14583_),
    .A2(_14626_),
    .B(_14484_),
    .Y(_14721_));
 AOI21x1_ASAP7_75t_R _23121_ (.A1(_14518_),
    .A2(_14455_),
    .B(_14554_),
    .Y(_14722_));
 NAND2x1_ASAP7_75t_R _23122_ (.A(_14721_),
    .B(_14722_),
    .Y(_14723_));
 OA21x2_ASAP7_75t_R _23123_ (.A1(_14399_),
    .A2(_01196_),
    .B(_14554_),
    .Y(_14724_));
 NOR2x1_ASAP7_75t_R _23124_ (.A(_14651_),
    .B(_14387_),
    .Y(_14725_));
 NAND2x1_ASAP7_75t_R _23125_ (.A(_14481_),
    .B(_14725_),
    .Y(_14726_));
 AOI21x1_ASAP7_75t_R _23126_ (.A1(_14724_),
    .A2(_14726_),
    .B(_14428_),
    .Y(_14727_));
 AOI21x1_ASAP7_75t_R _23127_ (.A1(_14727_),
    .A2(_14723_),
    .B(_14514_),
    .Y(_14728_));
 AOI21x1_ASAP7_75t_R _23128_ (.A1(_14625_),
    .A2(_14626_),
    .B(_14484_),
    .Y(_14729_));
 AND3x1_ASAP7_75t_R _23129_ (.A(_14397_),
    .B(_14396_),
    .C(_00545_),
    .Y(_14730_));
 OA21x2_ASAP7_75t_R _23130_ (.A1(_14729_),
    .A2(_14730_),
    .B(_14445_),
    .Y(_14731_));
 NAND2x2_ASAP7_75t_R _23131_ (.A(net758),
    .B(_14389_),
    .Y(_14732_));
 AO21x1_ASAP7_75t_R _23132_ (.A1(_14732_),
    .A2(_14500_),
    .B(_14568_),
    .Y(_14733_));
 AO21x1_ASAP7_75t_R _23133_ (.A1(_14438_),
    .A2(_14526_),
    .B(_14532_),
    .Y(_14734_));
 AOI21x1_ASAP7_75t_R _23134_ (.A1(_14733_),
    .A2(_14734_),
    .B(_14613_),
    .Y(_14735_));
 OAI21x1_ASAP7_75t_R _23135_ (.A1(_14731_),
    .A2(_14735_),
    .B(_14654_),
    .Y(_14736_));
 NAND2x1_ASAP7_75t_R _23136_ (.A(_14728_),
    .B(_14736_),
    .Y(_14737_));
 NAND2x1_ASAP7_75t_R _23137_ (.A(_14720_),
    .B(_14737_),
    .Y(_14738_));
 OAI21x1_ASAP7_75t_R _23138_ (.A1(_14686_),
    .A2(_14705_),
    .B(_14738_),
    .Y(_00074_));
 NAND2x1_ASAP7_75t_R _23139_ (.A(_14395_),
    .B(_14599_),
    .Y(_14739_));
 AOI211x1_ASAP7_75t_R _23140_ (.A1(_14676_),
    .A2(_14739_),
    .B(_14680_),
    .C(_14429_),
    .Y(_14740_));
 NOR2x1_ASAP7_75t_R _23141_ (.A(_14517_),
    .B(_14544_),
    .Y(_14741_));
 NAND2x1_ASAP7_75t_R _23142_ (.A(_14490_),
    .B(_14583_),
    .Y(_14742_));
 OAI21x1_ASAP7_75t_R _23143_ (.A1(_14528_),
    .A2(_14742_),
    .B(_14428_),
    .Y(_14743_));
 OAI21x1_ASAP7_75t_R _23144_ (.A1(_14741_),
    .A2(_14743_),
    .B(_14555_),
    .Y(_14744_));
 NOR2x1_ASAP7_75t_R _23145_ (.A(_14740_),
    .B(_14744_),
    .Y(_14745_));
 AO21x1_ASAP7_75t_R _23146_ (.A1(_14411_),
    .A2(_14454_),
    .B(_14563_),
    .Y(_14746_));
 AND3x1_ASAP7_75t_R _23147_ (.A(_14588_),
    .B(_14589_),
    .C(_14518_),
    .Y(_14747_));
 OAI21x1_ASAP7_75t_R _23148_ (.A1(_14746_),
    .A2(_14747_),
    .B(_14696_),
    .Y(_14748_));
 NAND2x1_ASAP7_75t_R _23149_ (.A(_15896_),
    .B(_14532_),
    .Y(_14749_));
 OAI21x1_ASAP7_75t_R _23150_ (.A1(_14436_),
    .A2(_14749_),
    .B(_14563_),
    .Y(_14750_));
 AOI21x1_ASAP7_75t_R _23151_ (.A1(_14510_),
    .A2(_14732_),
    .B(_14417_),
    .Y(_14751_));
 NOR3x1_ASAP7_75t_R _23152_ (.A(_14750_),
    .B(_14557_),
    .C(_14751_),
    .Y(_14752_));
 OAI21x1_ASAP7_75t_R _23153_ (.A1(_14748_),
    .A2(_14752_),
    .B(_14578_),
    .Y(_14753_));
 NOR2x1_ASAP7_75t_R _23154_ (.A(_14745_),
    .B(_14753_),
    .Y(_14754_));
 BUFx6f_ASAP7_75t_R _23155_ (.A(_14484_),
    .Y(_14755_));
 AOI21x1_ASAP7_75t_R _23156_ (.A1(_14490_),
    .A2(_14510_),
    .B(_14755_),
    .Y(_14756_));
 NAND2x2_ASAP7_75t_R _23157_ (.A(net759),
    .B(_14453_),
    .Y(_14757_));
 AOI21x1_ASAP7_75t_R _23158_ (.A1(net54),
    .A2(_14757_),
    .B(_14528_),
    .Y(_14758_));
 OAI21x1_ASAP7_75t_R _23159_ (.A1(_14756_),
    .A2(_14758_),
    .B(_14696_),
    .Y(_14759_));
 AOI21x1_ASAP7_75t_R _23160_ (.A1(_14732_),
    .A2(_14527_),
    .B(_14755_),
    .Y(_14760_));
 AOI21x1_ASAP7_75t_R _23161_ (.A1(_14500_),
    .A2(_14581_),
    .B(_14676_),
    .Y(_14761_));
 OAI21x1_ASAP7_75t_R _23162_ (.A1(_14760_),
    .A2(_14761_),
    .B(_14479_),
    .Y(_14762_));
 AOI21x1_ASAP7_75t_R _23163_ (.A1(_14759_),
    .A2(_14762_),
    .B(_14654_),
    .Y(_14763_));
 NAND2x2_ASAP7_75t_R _23164_ (.A(net703),
    .B(net56),
    .Y(_14764_));
 NAND3x2_ASAP7_75t_R _23165_ (.B(_14764_),
    .C(_14413_),
    .Y(_14765_),
    .A(_14510_));
 OAI21x1_ASAP7_75t_R _23166_ (.A1(_14641_),
    .A2(_14765_),
    .B(_14654_),
    .Y(_14766_));
 INVx3_ASAP7_75t_R _23167_ (.A(_14638_),
    .Y(_14767_));
 OAI21x1_ASAP7_75t_R _23168_ (.A1(_14531_),
    .A2(_15896_),
    .B(_14532_),
    .Y(_14768_));
 OAI21x1_ASAP7_75t_R _23169_ (.A1(_14767_),
    .A2(_14768_),
    .B(_14534_),
    .Y(_14769_));
 NOR2x2_ASAP7_75t_R _23170_ (.A(_14398_),
    .B(_14482_),
    .Y(_14770_));
 AND2x2_ASAP7_75t_R _23171_ (.A(_14770_),
    .B(net55),
    .Y(_14771_));
 NOR2x1_ASAP7_75t_R _23172_ (.A(_14769_),
    .B(_14771_),
    .Y(_14772_));
 OAI21x1_ASAP7_75t_R _23173_ (.A1(_14766_),
    .A2(_14772_),
    .B(_14468_),
    .Y(_14773_));
 OAI21x1_ASAP7_75t_R _23174_ (.A1(_14763_),
    .A2(_14773_),
    .B(_14477_),
    .Y(_14774_));
 NAND3x1_ASAP7_75t_R _23175_ (.A(_14583_),
    .B(_14665_),
    .C(_14671_),
    .Y(_14775_));
 AOI21x1_ASAP7_75t_R _23176_ (.A1(_14512_),
    .A2(_14775_),
    .B(_14495_),
    .Y(_14776_));
 AOI21x1_ASAP7_75t_R _23177_ (.A1(_14687_),
    .A2(_14706_),
    .B(_14671_),
    .Y(_14777_));
 OAI21x1_ASAP7_75t_R _23178_ (.A1(_14777_),
    .A2(_14593_),
    .B(_14479_),
    .Y(_14778_));
 NAND2x1_ASAP7_75t_R _23179_ (.A(_14776_),
    .B(_14778_),
    .Y(_14779_));
 AOI21x1_ASAP7_75t_R _23180_ (.A1(net55),
    .A2(_14665_),
    .B(_14528_),
    .Y(_14780_));
 AOI21x1_ASAP7_75t_R _23181_ (.A1(_14522_),
    .A2(_14416_),
    .B(_14387_),
    .Y(_14781_));
 OAI21x1_ASAP7_75t_R _23182_ (.A1(_14780_),
    .A2(_14781_),
    .B(_14696_),
    .Y(_14782_));
 OAI21x1_ASAP7_75t_R _23183_ (.A1(_14511_),
    .A2(_14627_),
    .B(_14555_),
    .Y(_14783_));
 NAND3x1_ASAP7_75t_R _23184_ (.A(_14782_),
    .B(_14783_),
    .C(_14447_),
    .Y(_14784_));
 AOI21x1_ASAP7_75t_R _23185_ (.A1(_14779_),
    .A2(_14784_),
    .B(_14578_),
    .Y(_14785_));
 NOR2x2_ASAP7_75t_R _23186_ (.A(_14412_),
    .B(_14399_),
    .Y(_14786_));
 AOI22x1_ASAP7_75t_R _23187_ (.A1(_14786_),
    .A2(_14495_),
    .B1(_14676_),
    .B2(_14486_),
    .Y(_14787_));
 AOI21x1_ASAP7_75t_R _23188_ (.A1(_14639_),
    .A2(_14757_),
    .B(_14676_),
    .Y(_14788_));
 OAI21x1_ASAP7_75t_R _23189_ (.A1(_14557_),
    .A2(_14788_),
    .B(_14654_),
    .Y(_14789_));
 AOI21x1_ASAP7_75t_R _23190_ (.A1(_14787_),
    .A2(_14789_),
    .B(_14479_),
    .Y(_14790_));
 OAI21x1_ASAP7_75t_R _23191_ (.A1(_14485_),
    .A2(_14416_),
    .B(_14563_),
    .Y(_14791_));
 OAI21x1_ASAP7_75t_R _23192_ (.A1(_14688_),
    .A2(_14791_),
    .B(_14479_),
    .Y(_14792_));
 AOI21x1_ASAP7_75t_R _23193_ (.A1(_14665_),
    .A2(_14706_),
    .B(_14755_),
    .Y(_14793_));
 OAI21x1_ASAP7_75t_R _23194_ (.A1(_15891_),
    .A2(_15896_),
    .B(net54),
    .Y(_14794_));
 OAI21x1_ASAP7_75t_R _23195_ (.A1(_14676_),
    .A2(_14794_),
    .B(_14428_),
    .Y(_14795_));
 NOR2x1_ASAP7_75t_R _23196_ (.A(_14793_),
    .B(_14795_),
    .Y(_14796_));
 OAI21x1_ASAP7_75t_R _23197_ (.A1(_14792_),
    .A2(_14796_),
    .B(_14578_),
    .Y(_14797_));
 OAI21x1_ASAP7_75t_R _23198_ (.A1(_14790_),
    .A2(_14797_),
    .B(_14476_),
    .Y(_14798_));
 OAI22x1_ASAP7_75t_R _23199_ (.A1(_14754_),
    .A2(_14774_),
    .B1(_14785_),
    .B2(_14798_),
    .Y(_00075_));
 NOR2x1_ASAP7_75t_R _23200_ (.A(_14413_),
    .B(_14486_),
    .Y(_14799_));
 INVx1_ASAP7_75t_R _23201_ (.A(_14483_),
    .Y(_14800_));
 AO21x1_ASAP7_75t_R _23202_ (.A1(_14799_),
    .A2(_14800_),
    .B(_14429_),
    .Y(_14801_));
 AND3x1_ASAP7_75t_R _23203_ (.A(_14588_),
    .B(_14626_),
    .C(_14532_),
    .Y(_14802_));
 NAND2x1_ASAP7_75t_R _23204_ (.A(_14518_),
    .B(_14588_),
    .Y(_14803_));
 OAI21x1_ASAP7_75t_R _23205_ (.A1(_14549_),
    .A2(_14803_),
    .B(_14613_),
    .Y(_14804_));
 NOR2x1_ASAP7_75t_R _23206_ (.A(_14802_),
    .B(_14804_),
    .Y(_14805_));
 OAI21x1_ASAP7_75t_R _23207_ (.A1(_14801_),
    .A2(_14805_),
    .B(_14468_),
    .Y(_14806_));
 NAND2x1_ASAP7_75t_R _23208_ (.A(_14520_),
    .B(_14639_),
    .Y(_14807_));
 NOR2x1_ASAP7_75t_R _23209_ (.A(_14439_),
    .B(_14807_),
    .Y(_14808_));
 NAND2x1_ASAP7_75t_R _23210_ (.A(_14532_),
    .B(_14639_),
    .Y(_14809_));
 NOR2x1_ASAP7_75t_R _23211_ (.A(_14549_),
    .B(_14809_),
    .Y(_14810_));
 OAI21x1_ASAP7_75t_R _23212_ (.A1(_14808_),
    .A2(_14810_),
    .B(_14696_),
    .Y(_14811_));
 INVx1_ASAP7_75t_R _23213_ (.A(_14729_),
    .Y(_14812_));
 AO21x1_ASAP7_75t_R _23214_ (.A1(_14590_),
    .A2(_14812_),
    .B(_14534_),
    .Y(_14813_));
 AOI21x1_ASAP7_75t_R _23215_ (.A1(_14811_),
    .A2(_14813_),
    .B(_14564_),
    .Y(_14814_));
 NOR2x1_ASAP7_75t_R _23216_ (.A(_14806_),
    .B(_14814_),
    .Y(_14815_));
 AOI21x1_ASAP7_75t_R _23217_ (.A1(_14626_),
    .A2(_14507_),
    .B(_14755_),
    .Y(_14816_));
 OAI21x1_ASAP7_75t_R _23218_ (.A1(_14666_),
    .A2(_14816_),
    .B(_14696_),
    .Y(_14817_));
 AOI21x1_ASAP7_75t_R _23219_ (.A1(_14509_),
    .A2(_14626_),
    .B(_14755_),
    .Y(_14818_));
 OAI21x1_ASAP7_75t_R _23220_ (.A1(_14818_),
    .A2(_14635_),
    .B(_14479_),
    .Y(_14819_));
 AOI21x1_ASAP7_75t_R _23221_ (.A1(_14817_),
    .A2(_14819_),
    .B(_14564_),
    .Y(_14820_));
 OAI21x1_ASAP7_75t_R _23222_ (.A1(_14395_),
    .A2(_14399_),
    .B(_14457_),
    .Y(_14821_));
 NAND2x2_ASAP7_75t_R _23223_ (.A(_14410_),
    .B(_14689_),
    .Y(_14822_));
 NAND2x1_ASAP7_75t_R _23224_ (.A(_14416_),
    .B(_14822_),
    .Y(_14823_));
 OAI21x1_ASAP7_75t_R _23225_ (.A1(_14821_),
    .A2(_14823_),
    .B(_14447_),
    .Y(_14824_));
 AOI21x1_ASAP7_75t_R _23226_ (.A1(_14500_),
    .A2(_14599_),
    .B(_14528_),
    .Y(_14825_));
 AOI211x1_ASAP7_75t_R _23227_ (.A1(_14481_),
    .A2(_14483_),
    .B(_14825_),
    .C(_14512_),
    .Y(_14826_));
 OAI21x1_ASAP7_75t_R _23228_ (.A1(_14826_),
    .A2(_14824_),
    .B(_14578_),
    .Y(_14827_));
 OAI21x1_ASAP7_75t_R _23229_ (.A1(_14820_),
    .A2(_14827_),
    .B(_14477_),
    .Y(_14828_));
 OAI21x1_ASAP7_75t_R _23230_ (.A1(_14439_),
    .A2(_14507_),
    .B(_14534_),
    .Y(_14829_));
 NOR2x2_ASAP7_75t_R _23231_ (.A(_14767_),
    .B(_14800_),
    .Y(_14830_));
 NOR2x1_ASAP7_75t_R _23232_ (.A(_14829_),
    .B(_14830_),
    .Y(_14831_));
 AO21x1_ASAP7_75t_R _23233_ (.A1(_14385_),
    .A2(_14384_),
    .B(_00547_),
    .Y(_14832_));
 AO21x1_ASAP7_75t_R _23234_ (.A1(_14832_),
    .A2(_14822_),
    .B(_14501_),
    .Y(_14833_));
 NAND2x1_ASAP7_75t_R _23235_ (.A(_14495_),
    .B(_14833_),
    .Y(_14834_));
 OAI21x1_ASAP7_75t_R _23236_ (.A1(_14834_),
    .A2(_14831_),
    .B(_14578_),
    .Y(_14835_));
 OAI21x1_ASAP7_75t_R _23237_ (.A1(_14440_),
    .A2(_14566_),
    .B(_14479_),
    .Y(_14836_));
 AO21x1_ASAP7_75t_R _23238_ (.A1(_14639_),
    .A2(_14520_),
    .B(_14488_),
    .Y(_14837_));
 NAND2x1_ASAP7_75t_R _23239_ (.A(_14583_),
    .B(_14483_),
    .Y(_14838_));
 AO21x1_ASAP7_75t_R _23240_ (.A1(_14837_),
    .A2(_14838_),
    .B(_14613_),
    .Y(_14839_));
 AOI21x1_ASAP7_75t_R _23241_ (.A1(_14836_),
    .A2(_14839_),
    .B(_14564_),
    .Y(_14840_));
 NOR2x1_ASAP7_75t_R _23242_ (.A(_14840_),
    .B(_14835_),
    .Y(_14841_));
 AO21x1_ASAP7_75t_R _23243_ (.A1(_14411_),
    .A2(_15899_),
    .B(_14458_),
    .Y(_14842_));
 AOI21x1_ASAP7_75t_R _23244_ (.A1(_14588_),
    .A2(_14665_),
    .B(_14676_),
    .Y(_14843_));
 OAI21x1_ASAP7_75t_R _23245_ (.A1(_14842_),
    .A2(_14843_),
    .B(_14429_),
    .Y(_14844_));
 NOR2x1_ASAP7_75t_R _23246_ (.A(_14671_),
    .B(_14443_),
    .Y(_14845_));
 OAI21x1_ASAP7_75t_R _23247_ (.A1(_14509_),
    .A2(_14439_),
    .B(_14534_),
    .Y(_14846_));
 NOR2x1_ASAP7_75t_R _23248_ (.A(_14439_),
    .B(_14589_),
    .Y(_14847_));
 AOI211x1_ASAP7_75t_R _23249_ (.A1(_14845_),
    .A2(_14589_),
    .B(_14846_),
    .C(_14847_),
    .Y(_14848_));
 OAI21x1_ASAP7_75t_R _23250_ (.A1(_14844_),
    .A2(_14848_),
    .B(_14468_),
    .Y(_14849_));
 INVx1_ASAP7_75t_R _23251_ (.A(_14524_),
    .Y(_14850_));
 NAND2x1_ASAP7_75t_R _23252_ (.A(_14500_),
    .B(_14622_),
    .Y(_14851_));
 OA21x2_ASAP7_75t_R _23253_ (.A1(_14520_),
    .A2(_15896_),
    .B(_14417_),
    .Y(_14852_));
 AO21x1_ASAP7_75t_R _23254_ (.A1(_14681_),
    .A2(_14456_),
    .B(_14445_),
    .Y(_14853_));
 OAI21x1_ASAP7_75t_R _23255_ (.A1(_14852_),
    .A2(_14853_),
    .B(_14447_),
    .Y(_14854_));
 AOI21x1_ASAP7_75t_R _23256_ (.A1(_14850_),
    .A2(_14851_),
    .B(_14854_),
    .Y(_14855_));
 OAI21x1_ASAP7_75t_R _23257_ (.A1(_14849_),
    .A2(_14855_),
    .B(_14476_),
    .Y(_14856_));
 OAI22x1_ASAP7_75t_R _23258_ (.A1(_14828_),
    .A2(_14815_),
    .B1(_14841_),
    .B2(_14856_),
    .Y(_00076_));
 AOI211x1_ASAP7_75t_R _23259_ (.A1(_14444_),
    .A2(_14659_),
    .B(_14519_),
    .C(_14512_),
    .Y(_14857_));
 AO21x1_ASAP7_75t_R _23260_ (.A1(_14433_),
    .A2(_01192_),
    .B(_14484_),
    .Y(_14858_));
 NAND2x1_ASAP7_75t_R _23261_ (.A(_14770_),
    .B(_14481_),
    .Y(_14859_));
 NAND2x1_ASAP7_75t_R _23262_ (.A(_14858_),
    .B(_14859_),
    .Y(_14860_));
 OAI21x1_ASAP7_75t_R _23263_ (.A1(_14555_),
    .A2(_14860_),
    .B(_14467_),
    .Y(_14861_));
 NOR2x1_ASAP7_75t_R _23264_ (.A(_14857_),
    .B(_14861_),
    .Y(_14862_));
 AO21x1_ASAP7_75t_R _23265_ (.A1(_14392_),
    .A2(_14492_),
    .B(_14456_),
    .Y(_14863_));
 NAND2x1_ASAP7_75t_R _23266_ (.A(_14484_),
    .B(_14522_),
    .Y(_14864_));
 OA21x2_ASAP7_75t_R _23267_ (.A1(_14864_),
    .A2(_14391_),
    .B(_14458_),
    .Y(_14865_));
 AO21x1_ASAP7_75t_R _23268_ (.A1(_14498_),
    .A2(net56),
    .B(_14457_),
    .Y(_14866_));
 AOI21x1_ASAP7_75t_R _23269_ (.A1(_14755_),
    .A2(_14807_),
    .B(_14866_),
    .Y(_14867_));
 AOI21x1_ASAP7_75t_R _23270_ (.A1(_14863_),
    .A2(_14865_),
    .B(_14867_),
    .Y(_14868_));
 OAI21x1_ASAP7_75t_R _23271_ (.A1(_14468_),
    .A2(_14868_),
    .B(_14564_),
    .Y(_14869_));
 NOR2x1_ASAP7_75t_R _23272_ (.A(_14862_),
    .B(_14869_),
    .Y(_14870_));
 AO21x1_ASAP7_75t_R _23273_ (.A1(_14639_),
    .A2(_14598_),
    .B(_14498_),
    .Y(_14871_));
 AOI21x1_ASAP7_75t_R _23274_ (.A1(_14822_),
    .A2(_14871_),
    .B(_14445_),
    .Y(_14872_));
 NOR2x1_ASAP7_75t_R _23275_ (.A(_14437_),
    .B(_14544_),
    .Y(_14873_));
 AO21x1_ASAP7_75t_R _23276_ (.A1(_14665_),
    .A2(_14568_),
    .B(_14457_),
    .Y(_14874_));
 OAI21x1_ASAP7_75t_R _23277_ (.A1(_14873_),
    .A2(_14874_),
    .B(_14514_),
    .Y(_14875_));
 NOR2x1_ASAP7_75t_R _23278_ (.A(_14875_),
    .B(_14872_),
    .Y(_14876_));
 OA21x2_ASAP7_75t_R _23279_ (.A1(_14604_),
    .A2(_14399_),
    .B(_14554_),
    .Y(_14877_));
 INVx1_ASAP7_75t_R _23280_ (.A(_14781_),
    .Y(_14878_));
 NAND2x1_ASAP7_75t_R _23281_ (.A(_14877_),
    .B(_14878_),
    .Y(_14879_));
 NOR2x1_ASAP7_75t_R _23282_ (.A(_14413_),
    .B(_14622_),
    .Y(_14880_));
 OAI21x1_ASAP7_75t_R _23283_ (.A1(_14485_),
    .A2(_14527_),
    .B(_14880_),
    .Y(_14881_));
 AOI21x1_ASAP7_75t_R _23284_ (.A1(_14879_),
    .A2(_14881_),
    .B(_14514_),
    .Y(_14882_));
 OAI21x1_ASAP7_75t_R _23285_ (.A1(_14882_),
    .A2(_14876_),
    .B(_14654_),
    .Y(_14883_));
 NAND2x1_ASAP7_75t_R _23286_ (.A(_14477_),
    .B(_14883_),
    .Y(_14884_));
 AO21x1_ASAP7_75t_R _23287_ (.A1(_14581_),
    .A2(_14527_),
    .B(_14488_),
    .Y(_14885_));
 AO21x1_ASAP7_75t_R _23288_ (.A1(_14442_),
    .A2(_14441_),
    .B(_14505_),
    .Y(_14886_));
 AOI21x1_ASAP7_75t_R _23289_ (.A1(_14417_),
    .A2(_14886_),
    .B(_14458_),
    .Y(_14887_));
 OAI21x1_ASAP7_75t_R _23290_ (.A1(_14659_),
    .A2(_14821_),
    .B(_14563_),
    .Y(_14888_));
 AO21x1_ASAP7_75t_R _23291_ (.A1(_14885_),
    .A2(_14887_),
    .B(_14888_),
    .Y(_14889_));
 OA21x2_ASAP7_75t_R _23292_ (.A1(_14484_),
    .A2(_14450_),
    .B(_14554_),
    .Y(_14890_));
 AO21x1_ASAP7_75t_R _23293_ (.A1(_14391_),
    .A2(_15896_),
    .B(_14532_),
    .Y(_14891_));
 AOI21x1_ASAP7_75t_R _23294_ (.A1(_14890_),
    .A2(_14891_),
    .B(_14563_),
    .Y(_14892_));
 NAND2x1_ASAP7_75t_R _23295_ (.A(_14492_),
    .B(_14605_),
    .Y(_14893_));
 NAND2x1_ASAP7_75t_R _23296_ (.A(_14559_),
    .B(_14387_),
    .Y(_14894_));
 OA21x2_ASAP7_75t_R _23297_ (.A1(_14894_),
    .A2(_14543_),
    .B(_14457_),
    .Y(_14895_));
 NAND2x1_ASAP7_75t_R _23298_ (.A(_14893_),
    .B(_14895_),
    .Y(_14896_));
 AOI21x1_ASAP7_75t_R _23299_ (.A1(_14892_),
    .A2(_14896_),
    .B(_14467_),
    .Y(_14897_));
 NAND2x1_ASAP7_75t_R _23300_ (.A(_14889_),
    .B(_14897_),
    .Y(_14898_));
 OAI21x1_ASAP7_75t_R _23301_ (.A1(_14694_),
    .A2(_14607_),
    .B(_14552_),
    .Y(_14899_));
 OA21x2_ASAP7_75t_R _23302_ (.A1(_14757_),
    .A2(_14484_),
    .B(_14457_),
    .Y(_14900_));
 AOI21x1_ASAP7_75t_R _23303_ (.A1(_14899_),
    .A2(_14900_),
    .B(_14563_),
    .Y(_14901_));
 NAND2x1_ASAP7_75t_R _23304_ (.A(_14568_),
    .B(_14449_),
    .Y(_14902_));
 NAND2x1_ASAP7_75t_R _23305_ (.A(_14902_),
    .B(_14409_),
    .Y(_14903_));
 NAND2x1_ASAP7_75t_R _23306_ (.A(_14901_),
    .B(_14903_),
    .Y(_14904_));
 OA21x2_ASAP7_75t_R _23307_ (.A1(_14568_),
    .A2(net703),
    .B(_14554_),
    .Y(_14905_));
 AOI21x1_ASAP7_75t_R _23308_ (.A1(_14569_),
    .A2(_14905_),
    .B(_14429_),
    .Y(_14906_));
 AOI21x1_ASAP7_75t_R _23309_ (.A1(_14639_),
    .A2(_14770_),
    .B(_14413_),
    .Y(_14907_));
 AO21x1_ASAP7_75t_R _23310_ (.A1(_14527_),
    .A2(_14559_),
    .B(_14518_),
    .Y(_14908_));
 NAND2x1_ASAP7_75t_R _23311_ (.A(_14907_),
    .B(_14908_),
    .Y(_14909_));
 AOI21x1_ASAP7_75t_R _23312_ (.A1(_14906_),
    .A2(_14909_),
    .B(_14514_),
    .Y(_14910_));
 AOI21x1_ASAP7_75t_R _23313_ (.A1(_14904_),
    .A2(_14910_),
    .B(_14477_),
    .Y(_14911_));
 NAND2x1_ASAP7_75t_R _23314_ (.A(_14898_),
    .B(_14911_),
    .Y(_14912_));
 OAI21x1_ASAP7_75t_R _23315_ (.A1(_14870_),
    .A2(_14884_),
    .B(_14912_),
    .Y(_00077_));
 AOI21x1_ASAP7_75t_R _23316_ (.A1(_14599_),
    .A2(_14687_),
    .B(_14417_),
    .Y(_14913_));
 AOI21x1_ASAP7_75t_R _23317_ (.A1(_14433_),
    .A2(_14572_),
    .B(_14755_),
    .Y(_14914_));
 OAI21x1_ASAP7_75t_R _23318_ (.A1(_14913_),
    .A2(_14914_),
    .B(_14479_),
    .Y(_14915_));
 AOI21x1_ASAP7_75t_R _23319_ (.A1(_14416_),
    .A2(_14506_),
    .B(_14755_),
    .Y(_14916_));
 OA21x2_ASAP7_75t_R _23320_ (.A1(_14615_),
    .A2(_14651_),
    .B(_14671_),
    .Y(_14917_));
 OAI21x1_ASAP7_75t_R _23321_ (.A1(_14916_),
    .A2(_14917_),
    .B(_14696_),
    .Y(_14918_));
 AOI21x1_ASAP7_75t_R _23322_ (.A1(_14915_),
    .A2(_14918_),
    .B(_14564_),
    .Y(_14919_));
 AOI21x1_ASAP7_75t_R _23323_ (.A1(_14520_),
    .A2(_14639_),
    .B(_14671_),
    .Y(_14920_));
 AOI21x1_ASAP7_75t_R _23324_ (.A1(_01197_),
    .A2(_01195_),
    .B(_14439_),
    .Y(_14921_));
 NOR3x1_ASAP7_75t_R _23325_ (.A(_14920_),
    .B(_14921_),
    .C(_14512_),
    .Y(_14922_));
 INVx1_ASAP7_75t_R _23326_ (.A(_14598_),
    .Y(_14923_));
 OA21x2_ASAP7_75t_R _23327_ (.A1(_14692_),
    .A2(_14923_),
    .B(_14439_),
    .Y(_14924_));
 OAI21x1_ASAP7_75t_R _23328_ (.A1(_14846_),
    .A2(_14924_),
    .B(_14447_),
    .Y(_14925_));
 OAI21x1_ASAP7_75t_R _23329_ (.A1(_14922_),
    .A2(_14925_),
    .B(_14468_),
    .Y(_14926_));
 OAI21x1_ASAP7_75t_R _23330_ (.A1(_14919_),
    .A2(_14926_),
    .B(_14477_),
    .Y(_14927_));
 AOI21x1_ASAP7_75t_R _23331_ (.A1(_14526_),
    .A2(_14527_),
    .B(_14671_),
    .Y(_14928_));
 OA21x2_ASAP7_75t_R _23332_ (.A1(_14923_),
    .A2(_14604_),
    .B(_14552_),
    .Y(_14929_));
 OAI21x1_ASAP7_75t_R _23333_ (.A1(_14928_),
    .A2(_14929_),
    .B(_14555_),
    .Y(_14930_));
 AO21x1_ASAP7_75t_R _23334_ (.A1(_14604_),
    .A2(_14518_),
    .B(_14554_),
    .Y(_14931_));
 AO21x1_ASAP7_75t_R _23335_ (.A1(_14677_),
    .A2(_14717_),
    .B(_14931_),
    .Y(_14932_));
 AOI21x1_ASAP7_75t_R _23336_ (.A1(_14930_),
    .A2(_14932_),
    .B(_14654_),
    .Y(_14933_));
 AO21x1_ASAP7_75t_R _23337_ (.A1(_14451_),
    .A2(_14552_),
    .B(_14413_),
    .Y(_14934_));
 OA21x2_ASAP7_75t_R _23338_ (.A1(_14449_),
    .A2(net56),
    .B(_14411_),
    .Y(_14935_));
 OAI21x1_ASAP7_75t_R _23339_ (.A1(_14934_),
    .A2(_14935_),
    .B(_14429_),
    .Y(_14936_));
 NAND2x1_ASAP7_75t_R _23340_ (.A(_14522_),
    .B(_14507_),
    .Y(_14937_));
 AOI21x1_ASAP7_75t_R _23341_ (.A1(_14454_),
    .A2(_14706_),
    .B(_14439_),
    .Y(_14938_));
 AOI211x1_ASAP7_75t_R _23342_ (.A1(_14937_),
    .A2(_14676_),
    .B(_14938_),
    .C(_14512_),
    .Y(_14939_));
 OAI21x1_ASAP7_75t_R _23343_ (.A1(_14936_),
    .A2(_14939_),
    .B(_14514_),
    .Y(_14940_));
 NOR2x1_ASAP7_75t_R _23344_ (.A(_14933_),
    .B(_14940_),
    .Y(_14941_));
 AOI21x1_ASAP7_75t_R _23345_ (.A1(_14555_),
    .A2(_14670_),
    .B(_14467_),
    .Y(_14942_));
 OAI21x1_ASAP7_75t_R _23346_ (.A1(_14709_),
    .A2(_14830_),
    .B(_14696_),
    .Y(_14943_));
 NAND2x1_ASAP7_75t_R _23347_ (.A(_14942_),
    .B(_14943_),
    .Y(_14944_));
 AO21x1_ASAP7_75t_R _23348_ (.A1(_14560_),
    .A2(_14456_),
    .B(_14458_),
    .Y(_14945_));
 NOR2x1_ASAP7_75t_R _23349_ (.A(_14781_),
    .B(_14945_),
    .Y(_14946_));
 AOI211x1_ASAP7_75t_R _23350_ (.A1(_14542_),
    .A2(_14485_),
    .B(_14642_),
    .C(_14641_),
    .Y(_14947_));
 OAI21x1_ASAP7_75t_R _23351_ (.A1(_14946_),
    .A2(_14947_),
    .B(_14468_),
    .Y(_14948_));
 AOI21x1_ASAP7_75t_R _23352_ (.A1(_14944_),
    .A2(_14948_),
    .B(_14564_),
    .Y(_14949_));
 AO21x1_ASAP7_75t_R _23353_ (.A1(_14488_),
    .A2(_00548_),
    .B(_14501_),
    .Y(_14950_));
 AOI21x1_ASAP7_75t_R _23354_ (.A1(_14639_),
    .A2(_14770_),
    .B(_14950_),
    .Y(_14951_));
 NOR2x1_ASAP7_75t_R _23355_ (.A(_14560_),
    .B(_14768_),
    .Y(_14952_));
 AO21x1_ASAP7_75t_R _23356_ (.A1(_14567_),
    .A2(_14456_),
    .B(_14413_),
    .Y(_14953_));
 OAI21x1_ASAP7_75t_R _23357_ (.A1(_14952_),
    .A2(_14953_),
    .B(_14514_),
    .Y(_14954_));
 NOR2x1_ASAP7_75t_R _23358_ (.A(_14951_),
    .B(_14954_),
    .Y(_14955_));
 NOR2x2_ASAP7_75t_R _23359_ (.A(net720),
    .B(_14410_),
    .Y(_14956_));
 OAI21x1_ASAP7_75t_R _23360_ (.A1(_14956_),
    .A2(_14765_),
    .B(_14467_),
    .Y(_14957_));
 OAI21x1_ASAP7_75t_R _23361_ (.A1(_14531_),
    .A2(_15899_),
    .B(_14568_),
    .Y(_14958_));
 NAND2x1_ASAP7_75t_R _23362_ (.A(_14488_),
    .B(_14764_),
    .Y(_14959_));
 NAND2x1_ASAP7_75t_R _23363_ (.A(_14958_),
    .B(_14959_),
    .Y(_14960_));
 AOI21x1_ASAP7_75t_R _23364_ (.A1(_14510_),
    .A2(_14960_),
    .B(_14479_),
    .Y(_14961_));
 OAI21x1_ASAP7_75t_R _23365_ (.A1(_14957_),
    .A2(_14961_),
    .B(_14564_),
    .Y(_14962_));
 OAI21x1_ASAP7_75t_R _23366_ (.A1(_14955_),
    .A2(_14962_),
    .B(_14476_),
    .Y(_14963_));
 OAI22x1_ASAP7_75t_R _23367_ (.A1(_14927_),
    .A2(_14941_),
    .B1(_14949_),
    .B2(_14963_),
    .Y(_00078_));
 NOR2x1_ASAP7_75t_R _23368_ (.A(net703),
    .B(_14528_),
    .Y(_14964_));
 AOI21x1_ASAP7_75t_R _23369_ (.A1(_14588_),
    .A2(_14626_),
    .B(_14755_),
    .Y(_14965_));
 OAI21x1_ASAP7_75t_R _23370_ (.A1(_14964_),
    .A2(_14965_),
    .B(_14696_),
    .Y(_14966_));
 AOI21x1_ASAP7_75t_R _23371_ (.A1(_14526_),
    .A2(_14572_),
    .B(_14676_),
    .Y(_14967_));
 OAI21x1_ASAP7_75t_R _23372_ (.A1(_14729_),
    .A2(_14967_),
    .B(_14479_),
    .Y(_14968_));
 AOI21x1_ASAP7_75t_R _23373_ (.A1(_14966_),
    .A2(_14968_),
    .B(_14654_),
    .Y(_14969_));
 AOI21x1_ASAP7_75t_R _23374_ (.A1(net54),
    .A2(_14572_),
    .B(_14528_),
    .Y(_14970_));
 OAI21x1_ASAP7_75t_R _23375_ (.A1(_14755_),
    .A2(_14491_),
    .B(_14534_),
    .Y(_14971_));
 NOR2x1_ASAP7_75t_R _23376_ (.A(_14970_),
    .B(_14971_),
    .Y(_14972_));
 NOR2x1_ASAP7_75t_R _23377_ (.A(_14458_),
    .B(_14786_),
    .Y(_14973_));
 NAND2x1_ASAP7_75t_R _23378_ (.A(_14417_),
    .B(_14607_),
    .Y(_14974_));
 AO21x1_ASAP7_75t_R _23379_ (.A1(_14973_),
    .A2(_14974_),
    .B(_14495_),
    .Y(_14975_));
 OAI21x1_ASAP7_75t_R _23380_ (.A1(_14972_),
    .A2(_14975_),
    .B(_14578_),
    .Y(_14976_));
 OAI21x1_ASAP7_75t_R _23381_ (.A1(_14969_),
    .A2(_14976_),
    .B(_14476_),
    .Y(_14977_));
 NOR2x1_ASAP7_75t_R _23382_ (.A(_14439_),
    .B(_14794_),
    .Y(_14978_));
 NOR2x1_ASAP7_75t_R _23383_ (.A(_14651_),
    .B(_14533_),
    .Y(_14979_));
 OAI21x1_ASAP7_75t_R _23384_ (.A1(_14978_),
    .A2(_14979_),
    .B(_14512_),
    .Y(_14980_));
 OA21x2_ASAP7_75t_R _23385_ (.A1(_14449_),
    .A2(_14558_),
    .B(_14411_),
    .Y(_14981_));
 OAI21x1_ASAP7_75t_R _23386_ (.A1(_14913_),
    .A2(_14981_),
    .B(_14555_),
    .Y(_14982_));
 AOI21x1_ASAP7_75t_R _23387_ (.A1(_14980_),
    .A2(_14982_),
    .B(_14447_),
    .Y(_14983_));
 NAND2x1_ASAP7_75t_R _23388_ (.A(_14445_),
    .B(_14958_),
    .Y(_14984_));
 OAI21x1_ASAP7_75t_R _23389_ (.A1(_14984_),
    .A2(_14830_),
    .B(_14495_),
    .Y(_14985_));
 NOR2x1_ASAP7_75t_R _23390_ (.A(_14417_),
    .B(_14530_),
    .Y(_14986_));
 AOI21x1_ASAP7_75t_R _23391_ (.A1(_14509_),
    .A2(_14572_),
    .B(_14671_),
    .Y(_14987_));
 AOI211x1_ASAP7_75t_R _23392_ (.A1(_14986_),
    .A2(_14481_),
    .B(_14987_),
    .C(_14613_),
    .Y(_14988_));
 OAI21x1_ASAP7_75t_R _23393_ (.A1(_14985_),
    .A2(_14988_),
    .B(_14468_),
    .Y(_14989_));
 NOR2x1_ASAP7_75t_R _23394_ (.A(_14983_),
    .B(_14989_),
    .Y(_14990_));
 NOR2x1_ASAP7_75t_R _23395_ (.A(_14651_),
    .B(_14692_),
    .Y(_14991_));
 AO21x1_ASAP7_75t_R _23396_ (.A1(_14488_),
    .A2(_01197_),
    .B(_14501_),
    .Y(_14992_));
 AO21x1_ASAP7_75t_R _23397_ (.A1(_14485_),
    .A2(_14991_),
    .B(_14992_),
    .Y(_14993_));
 AND3x1_ASAP7_75t_R _23398_ (.A(_14488_),
    .B(_14454_),
    .C(net55),
    .Y(_14994_));
 NOR2x1_ASAP7_75t_R _23399_ (.A(_14767_),
    .B(_14864_),
    .Y(_14995_));
 OAI21x1_ASAP7_75t_R _23400_ (.A1(_14994_),
    .A2(_14995_),
    .B(_14696_),
    .Y(_14996_));
 AOI21x1_ASAP7_75t_R _23401_ (.A1(_14993_),
    .A2(_14996_),
    .B(_14564_),
    .Y(_14997_));
 NOR2x2_ASAP7_75t_R _23402_ (.A(_14598_),
    .B(_14411_),
    .Y(_14998_));
 AO21x1_ASAP7_75t_R _23403_ (.A1(_14417_),
    .A2(_00547_),
    .B(_14458_),
    .Y(_14999_));
 OAI21x1_ASAP7_75t_R _23404_ (.A1(_14998_),
    .A2(_14999_),
    .B(_14495_),
    .Y(_15000_));
 INVx1_ASAP7_75t_R _23405_ (.A(_14587_),
    .Y(_15001_));
 NOR2x2_ASAP7_75t_R _23406_ (.A(_14407_),
    .B(_14956_),
    .Y(_15002_));
 NAND2x1_ASAP7_75t_R _23407_ (.A(_14902_),
    .B(_15002_),
    .Y(_15003_));
 NOR2x1_ASAP7_75t_R _23408_ (.A(_15001_),
    .B(_15003_),
    .Y(_15004_));
 OAI21x1_ASAP7_75t_R _23409_ (.A1(_15000_),
    .A2(_15004_),
    .B(_14578_),
    .Y(_15005_));
 NOR2x1_ASAP7_75t_R _23410_ (.A(_14997_),
    .B(_15005_),
    .Y(_15006_));
 NAND2x1_ASAP7_75t_R _23411_ (.A(_14509_),
    .B(_14445_),
    .Y(_15007_));
 AOI211x1_ASAP7_75t_R _23412_ (.A1(_14517_),
    .A2(_14676_),
    .B(_15007_),
    .C(_14998_),
    .Y(_15008_));
 AO21x1_ASAP7_75t_R _23413_ (.A1(_14456_),
    .A2(_14393_),
    .B(_14445_),
    .Y(_15009_));
 OAI21x1_ASAP7_75t_R _23414_ (.A1(_15009_),
    .A2(_14920_),
    .B(_14654_),
    .Y(_15010_));
 OAI21x1_ASAP7_75t_R _23415_ (.A1(_15008_),
    .A2(_15010_),
    .B(_14468_),
    .Y(_15011_));
 AOI21x1_ASAP7_75t_R _23416_ (.A1(_14485_),
    .A2(_14530_),
    .B(_14777_),
    .Y(_15012_));
 AOI21x1_ASAP7_75t_R _23417_ (.A1(_14509_),
    .A2(_14572_),
    .B(_14528_),
    .Y(_15013_));
 NAND2x1_ASAP7_75t_R _23418_ (.A(net55),
    .B(_14488_),
    .Y(_15014_));
 OAI21x1_ASAP7_75t_R _23419_ (.A1(_14708_),
    .A2(_15014_),
    .B(_14613_),
    .Y(_15015_));
 OAI21x1_ASAP7_75t_R _23420_ (.A1(_15013_),
    .A2(_15015_),
    .B(_14447_),
    .Y(_15016_));
 AOI21x1_ASAP7_75t_R _23421_ (.A1(_15002_),
    .A2(_15012_),
    .B(_15016_),
    .Y(_15017_));
 OAI21x1_ASAP7_75t_R _23422_ (.A1(_15011_),
    .A2(_15017_),
    .B(_14477_),
    .Y(_15018_));
 OAI22x1_ASAP7_75t_R _23423_ (.A1(_14977_),
    .A2(_14990_),
    .B1(_15006_),
    .B2(_15018_),
    .Y(_00079_));
 INVx2_ASAP7_75t_R _23424_ (.A(_12127_),
    .Y(_15019_));
 XOR2x2_ASAP7_75t_R _23425_ (.A(_15019_),
    .B(_12081_),
    .Y(_15020_));
 XNOR2x2_ASAP7_75t_R _23426_ (.A(_00819_),
    .B(_00812_),
    .Y(_15021_));
 XOR2x2_ASAP7_75t_R _23427_ (.A(_12082_),
    .B(_12087_),
    .Y(_15022_));
 XOR2x1_ASAP7_75t_R _23428_ (.A(_15021_),
    .Y(_15023_),
    .B(_15022_));
 NOR2x1_ASAP7_75t_R _23429_ (.A(_15023_),
    .B(_15020_),
    .Y(_15024_));
 NOR2x1_ASAP7_75t_R _23430_ (.A(net20),
    .B(_12108_),
    .Y(_15025_));
 AND2x2_ASAP7_75t_R _23431_ (.A(net20),
    .B(_12080_),
    .Y(_15026_));
 OAI21x1_ASAP7_75t_R _23432_ (.A1(_15026_),
    .A2(_15025_),
    .B(_12127_),
    .Y(_15027_));
 INVx1_ASAP7_75t_R _23433_ (.A(net20),
    .Y(_15028_));
 NOR2x1_ASAP7_75t_R _23434_ (.A(_12108_),
    .B(_15028_),
    .Y(_15029_));
 INVx1_ASAP7_75t_R _23435_ (.A(_12080_),
    .Y(_15030_));
 NOR2x1_ASAP7_75t_R _23436_ (.A(net20),
    .B(_15030_),
    .Y(_15031_));
 OAI21x1_ASAP7_75t_R _23437_ (.A1(_15031_),
    .A2(_15029_),
    .B(_15019_),
    .Y(_15032_));
 NAND2x2_ASAP7_75t_R _23438_ (.A(_15032_),
    .B(_15027_),
    .Y(_15033_));
 XOR2x2_ASAP7_75t_R _23439_ (.A(_00812_),
    .B(_00819_),
    .Y(_15034_));
 XOR2x1_ASAP7_75t_R _23440_ (.A(_15034_),
    .Y(_15035_),
    .B(_15022_));
 OAI21x1_ASAP7_75t_R _23441_ (.A1(_15035_),
    .A2(_15033_),
    .B(_10723_),
    .Y(_15036_));
 NAND2x2_ASAP7_75t_R _23442_ (.A(_00549_),
    .B(_11373_),
    .Y(_15037_));
 OAI21x1_ASAP7_75t_R _23443_ (.A1(_15024_),
    .A2(_15036_),
    .B(_15037_),
    .Y(_15038_));
 XOR2x2_ASAP7_75t_R _23444_ (.A(_15038_),
    .B(_07972_),
    .Y(_15039_));
 BUFx12f_ASAP7_75t_R _23445_ (.A(_15039_),
    .Y(_15906_));
 NOR2x2_ASAP7_75t_R _23446_ (.A(_10668_),
    .B(_00550_),
    .Y(_15040_));
 NOR2x2_ASAP7_75t_R _23447_ (.A(net38),
    .B(_12108_),
    .Y(_15041_));
 AND2x4_ASAP7_75t_R _23448_ (.A(net921),
    .B(_12108_),
    .Y(_15042_));
 OAI21x1_ASAP7_75t_R _23449_ (.A1(_15042_),
    .A2(_15041_),
    .B(_12104_),
    .Y(_15043_));
 INVx1_ASAP7_75t_R _23450_ (.A(_15043_),
    .Y(_15044_));
 NOR3x1_ASAP7_75t_R _23451_ (.A(_15042_),
    .B(_12104_),
    .C(_15041_),
    .Y(_15045_));
 OAI21x1_ASAP7_75t_R _23452_ (.A1(_15044_),
    .A2(_15045_),
    .B(_15034_),
    .Y(_15046_));
 XOR2x1_ASAP7_75t_R _23453_ (.A(net921),
    .Y(_15047_),
    .B(_12108_));
 NAND2x2_ASAP7_75t_R _23454_ (.A(_12105_),
    .B(_15047_),
    .Y(_15048_));
 NAND3x1_ASAP7_75t_R _23455_ (.A(_15048_),
    .B(_15021_),
    .C(_15043_),
    .Y(_15049_));
 AOI21x1_ASAP7_75t_R _23456_ (.A1(_15046_),
    .A2(_15049_),
    .B(_12160_),
    .Y(_15050_));
 OAI21x1_ASAP7_75t_R _23457_ (.A1(_15040_),
    .A2(_15050_),
    .B(_07961_),
    .Y(_15051_));
 AOI21x1_ASAP7_75t_R _23458_ (.A1(_15043_),
    .A2(_15048_),
    .B(_15021_),
    .Y(_15052_));
 XOR2x1_ASAP7_75t_R _23459_ (.A(_12108_),
    .Y(_15053_),
    .B(_12104_));
 NAND2x1_ASAP7_75t_R _23460_ (.A(net38),
    .B(_15053_),
    .Y(_15054_));
 INVx1_ASAP7_75t_R _23461_ (.A(net38),
    .Y(_15055_));
 XNOR2x1_ASAP7_75t_R _23462_ (.B(_12104_),
    .Y(_15056_),
    .A(_12108_));
 NAND2x1_ASAP7_75t_R _23463_ (.A(_15055_),
    .B(_15056_),
    .Y(_15057_));
 AOI21x1_ASAP7_75t_R _23464_ (.A1(_15054_),
    .A2(_15057_),
    .B(net903),
    .Y(_15058_));
 OAI21x1_ASAP7_75t_R _23465_ (.A1(_15058_),
    .A2(_15052_),
    .B(_10763_),
    .Y(_15059_));
 INVx2_ASAP7_75t_R _23466_ (.A(_07961_),
    .Y(_15060_));
 INVx2_ASAP7_75t_R _23467_ (.A(_15040_),
    .Y(_15061_));
 NAND3x2_ASAP7_75t_R _23468_ (.B(_15060_),
    .C(_15061_),
    .Y(_15062_),
    .A(_15059_));
 NAND2x2_ASAP7_75t_R _23469_ (.A(_15051_),
    .B(_15062_),
    .Y(_15063_));
 BUFx10_ASAP7_75t_R _23470_ (.A(_15063_),
    .Y(_15908_));
 NOR2x1_ASAP7_75t_R _23471_ (.A(net668),
    .B(_00552_),
    .Y(_15064_));
 INVx1_ASAP7_75t_R _23472_ (.A(_15064_),
    .Y(_15065_));
 INVx2_ASAP7_75t_R _23473_ (.A(_12169_),
    .Y(_15066_));
 NOR2x2_ASAP7_75t_R _23474_ (.A(_15066_),
    .B(_12138_),
    .Y(_15067_));
 NOR2x2_ASAP7_75t_R _23475_ (.A(_12169_),
    .B(_12134_),
    .Y(_15068_));
 OAI21x1_ASAP7_75t_R _23476_ (.A1(_15067_),
    .A2(_15068_),
    .B(net610),
    .Y(_15069_));
 INVx1_ASAP7_75t_R _23477_ (.A(_15069_),
    .Y(_15070_));
 NOR3x1_ASAP7_75t_R _23478_ (.A(_15068_),
    .B(_15067_),
    .C(net609),
    .Y(_15071_));
 OAI21x1_ASAP7_75t_R _23479_ (.A1(_15070_),
    .A2(_15071_),
    .B(net767),
    .Y(_15072_));
 AOI21x1_ASAP7_75t_R _23480_ (.A1(_15065_),
    .A2(_15072_),
    .B(_08293_),
    .Y(_15073_));
 BUFx6f_ASAP7_75t_R _23481_ (.A(_15073_),
    .Y(_15074_));
 NAND2x1_ASAP7_75t_R _23482_ (.A(_00552_),
    .B(_10639_),
    .Y(_15075_));
 NAND2x2_ASAP7_75t_R _23483_ (.A(_15066_),
    .B(_12138_),
    .Y(_15076_));
 INVx1_ASAP7_75t_R _23484_ (.A(net608),
    .Y(_15077_));
 NOR2x1_ASAP7_75t_R _23485_ (.A(_12132_),
    .B(_12133_),
    .Y(_15078_));
 AND2x2_ASAP7_75t_R _23486_ (.A(_12132_),
    .B(_12133_),
    .Y(_15079_));
 OAI21x1_ASAP7_75t_R _23487_ (.A1(_15078_),
    .A2(_15079_),
    .B(_12169_),
    .Y(_15080_));
 NAND3x2_ASAP7_75t_R _23488_ (.B(_15077_),
    .C(_15080_),
    .Y(_15081_),
    .A(_15076_));
 NAND3x2_ASAP7_75t_R _23489_ (.B(_10620_),
    .C(_15069_),
    .Y(_15082_),
    .A(_15081_));
 AOI21x1_ASAP7_75t_R _23490_ (.A1(_15075_),
    .A2(_15082_),
    .B(_08007_),
    .Y(_15083_));
 NOR2x2_ASAP7_75t_R _23491_ (.A(_15083_),
    .B(_15074_),
    .Y(_15084_));
 BUFx12f_ASAP7_75t_R _23492_ (.A(_15084_),
    .Y(_15085_));
 BUFx10_ASAP7_75t_R _23493_ (.A(_15085_),
    .Y(_15916_));
 OAI21x1_ASAP7_75t_R _23494_ (.A1(_15040_),
    .A2(_15050_),
    .B(_15060_),
    .Y(_15086_));
 NAND3x2_ASAP7_75t_R _23495_ (.B(_07961_),
    .C(_15061_),
    .Y(_15087_),
    .A(_15059_));
 NAND2x2_ASAP7_75t_R _23496_ (.A(_15087_),
    .B(_15086_),
    .Y(_15088_));
 BUFx12_ASAP7_75t_R _23497_ (.A(_15088_),
    .Y(_15903_));
 AOI21x1_ASAP7_75t_R _23498_ (.A1(_15065_),
    .A2(_15072_),
    .B(_08007_),
    .Y(_15089_));
 BUFx6f_ASAP7_75t_R _23499_ (.A(_15089_),
    .Y(_15090_));
 AOI21x1_ASAP7_75t_R _23500_ (.A1(_15075_),
    .A2(_15082_),
    .B(_08293_),
    .Y(_15091_));
 NOR2x2_ASAP7_75t_R _23501_ (.A(_15090_),
    .B(_15091_),
    .Y(_15092_));
 BUFx12f_ASAP7_75t_R _23502_ (.A(_15092_),
    .Y(_15913_));
 INVx3_ASAP7_75t_R _23503_ (.A(_01201_),
    .Y(_15093_));
 BUFx10_ASAP7_75t_R _23504_ (.A(_15092_),
    .Y(_15094_));
 INVx1_ASAP7_75t_R _23505_ (.A(_00751_),
    .Y(_15095_));
 XOR2x1_ASAP7_75t_R _23506_ (.A(_12173_),
    .Y(_15096_),
    .B(_15095_));
 XOR2x2_ASAP7_75t_R _23507_ (.A(_12132_),
    .B(_00819_),
    .Y(_15097_));
 XOR2x1_ASAP7_75t_R _23508_ (.A(_12172_),
    .Y(_15098_),
    .B(_15097_));
 NOR2x1_ASAP7_75t_R _23509_ (.A(_15096_),
    .B(_15098_),
    .Y(_15099_));
 XOR2x1_ASAP7_75t_R _23510_ (.A(_12173_),
    .Y(_15100_),
    .B(_00751_));
 XNOR2x1_ASAP7_75t_R _23511_ (.B(_12172_),
    .Y(_15101_),
    .A(_15097_));
 NOR2x1_ASAP7_75t_R _23512_ (.A(_15100_),
    .B(_15101_),
    .Y(_15102_));
 OAI21x1_ASAP7_75t_R _23513_ (.A1(_15099_),
    .A2(_15102_),
    .B(net621),
    .Y(_15103_));
 INVx2_ASAP7_75t_R _23514_ (.A(_01069_),
    .Y(_15104_));
 NOR2x2_ASAP7_75t_R _23515_ (.A(net650),
    .B(_00678_),
    .Y(_15105_));
 INVx3_ASAP7_75t_R _23516_ (.A(_15105_),
    .Y(_15106_));
 NAND3x2_ASAP7_75t_R _23517_ (.B(_15104_),
    .C(_15106_),
    .Y(_15107_),
    .A(_15103_));
 AO21x1_ASAP7_75t_R _23518_ (.A1(_15103_),
    .A2(_15106_),
    .B(_15104_),
    .Y(_15108_));
 NAND2x2_ASAP7_75t_R _23519_ (.A(_15107_),
    .B(_15108_),
    .Y(_15109_));
 BUFx6f_ASAP7_75t_R _23520_ (.A(_15109_),
    .Y(_15110_));
 OAI21x1_ASAP7_75t_R _23521_ (.A1(_15093_),
    .A2(_15094_),
    .B(_15110_),
    .Y(_15111_));
 NAND2x2_ASAP7_75t_R _23522_ (.A(net840),
    .B(_15039_),
    .Y(_15112_));
 NOR2x2_ASAP7_75t_R _23523_ (.A(_15916_),
    .B(_15112_),
    .Y(_15113_));
 NOR2x1_ASAP7_75t_R _23524_ (.A(_15111_),
    .B(_15113_),
    .Y(_15114_));
 NOR2x2_ASAP7_75t_R _23525_ (.A(net868),
    .B(_15085_),
    .Y(_15115_));
 INVx1_ASAP7_75t_R _23526_ (.A(_15103_),
    .Y(_15116_));
 OAI21x1_ASAP7_75t_R _23527_ (.A1(_15105_),
    .A2(_15116_),
    .B(_15104_),
    .Y(_15117_));
 NAND3x2_ASAP7_75t_R _23528_ (.B(_01069_),
    .C(_15106_),
    .Y(_15118_),
    .A(_15103_));
 NAND2x2_ASAP7_75t_R _23529_ (.A(_15117_),
    .B(_15118_),
    .Y(_15119_));
 BUFx12_ASAP7_75t_R _23530_ (.A(_15119_),
    .Y(_15120_));
 BUFx6f_ASAP7_75t_R _23531_ (.A(_15120_),
    .Y(_15121_));
 AND2x2_ASAP7_75t_R _23532_ (.A(_11370_),
    .B(_00677_),
    .Y(_15122_));
 XOR2x2_ASAP7_75t_R _23533_ (.A(_12187_),
    .B(_00752_),
    .Y(_15123_));
 XOR2x2_ASAP7_75t_R _23534_ (.A(_00815_),
    .B(net40),
    .Y(_15124_));
 XOR2x2_ASAP7_75t_R _23535_ (.A(_12188_),
    .B(_15124_),
    .Y(_15125_));
 XOR2x1_ASAP7_75t_R _23536_ (.A(_15123_),
    .Y(_15126_),
    .B(_15125_));
 NOR2x1_ASAP7_75t_R _23537_ (.A(_12092_),
    .B(_15126_),
    .Y(_15127_));
 INVx1_ASAP7_75t_R _23538_ (.A(_07994_),
    .Y(_15128_));
 OAI21x1_ASAP7_75t_R _23539_ (.A1(_15122_),
    .A2(_15127_),
    .B(_15128_),
    .Y(_15129_));
 NOR2x2_ASAP7_75t_R _23540_ (.A(_11450_),
    .B(_00677_),
    .Y(_15130_));
 XNOR2x1_ASAP7_75t_R _23541_ (.B(_15123_),
    .Y(_15131_),
    .A(_15125_));
 NOR2x1_ASAP7_75t_R _23542_ (.A(_12092_),
    .B(_15131_),
    .Y(_15132_));
 OAI21x1_ASAP7_75t_R _23543_ (.A1(_15130_),
    .A2(_15132_),
    .B(_07994_),
    .Y(_15133_));
 NAND2x2_ASAP7_75t_R _23544_ (.A(_15129_),
    .B(_15133_),
    .Y(_15134_));
 BUFx6f_ASAP7_75t_R _23545_ (.A(_15134_),
    .Y(_15135_));
 AO21x1_ASAP7_75t_R _23546_ (.A1(_15115_),
    .A2(_15121_),
    .B(_15135_),
    .Y(_15136_));
 NOR2x1_ASAP7_75t_R _23547_ (.A(_15114_),
    .B(_15136_),
    .Y(_15137_));
 OAI21x1_ASAP7_75t_R _23548_ (.A1(_15090_),
    .A2(_15091_),
    .B(_00551_),
    .Y(_15138_));
 INVx1_ASAP7_75t_R _23549_ (.A(_07972_),
    .Y(_15139_));
 XOR2x2_ASAP7_75t_R _23550_ (.A(_15038_),
    .B(_15139_),
    .Y(_15140_));
 OAI21x1_ASAP7_75t_R _23551_ (.A1(_15140_),
    .A2(_15063_),
    .B(_15092_),
    .Y(_15141_));
 BUFx6f_ASAP7_75t_R _23552_ (.A(_15110_),
    .Y(_15142_));
 AOI21x1_ASAP7_75t_R _23553_ (.A1(_15138_),
    .A2(_15141_),
    .B(_15142_),
    .Y(_15143_));
 BUFx6f_ASAP7_75t_R _23554_ (.A(_15109_),
    .Y(_15144_));
 BUFx6f_ASAP7_75t_R _23555_ (.A(_15144_),
    .Y(_15145_));
 OAI21x1_ASAP7_75t_R _23556_ (.A1(_15122_),
    .A2(_15127_),
    .B(_07994_),
    .Y(_15146_));
 OAI21x1_ASAP7_75t_R _23557_ (.A1(_15130_),
    .A2(_15132_),
    .B(_15128_),
    .Y(_15147_));
 NAND2x2_ASAP7_75t_R _23558_ (.A(_15146_),
    .B(_15147_),
    .Y(_15148_));
 BUFx6f_ASAP7_75t_R _23559_ (.A(_15148_),
    .Y(_15149_));
 AO21x1_ASAP7_75t_R _23560_ (.A1(_15115_),
    .A2(_15145_),
    .B(_15149_),
    .Y(_15150_));
 XOR2x2_ASAP7_75t_R _23561_ (.A(_00818_),
    .B(_00850_),
    .Y(_15151_));
 XOR2x1_ASAP7_75t_R _23562_ (.A(_12258_),
    .Y(_15152_),
    .B(_00754_));
 XNOR2x1_ASAP7_75t_R _23563_ (.B(_15152_),
    .Y(_15153_),
    .A(_15151_));
 NOR2x1_ASAP7_75t_R _23564_ (.A(_10734_),
    .B(_00675_),
    .Y(_15154_));
 AO21x1_ASAP7_75t_R _23565_ (.A1(_15153_),
    .A2(_10829_),
    .B(_15154_),
    .Y(_15155_));
 XOR2x2_ASAP7_75t_R _23566_ (.A(_15155_),
    .B(_01073_),
    .Y(_15156_));
 BUFx10_ASAP7_75t_R _23567_ (.A(_15156_),
    .Y(_15157_));
 OAI21x1_ASAP7_75t_R _23568_ (.A1(_15143_),
    .A2(_15150_),
    .B(_15157_),
    .Y(_15158_));
 XNOR2x1_ASAP7_75t_R _23569_ (.B(_00784_),
    .Y(_15159_),
    .A(_00753_));
 INVx1_ASAP7_75t_R _23570_ (.A(_15159_),
    .Y(_15160_));
 XOR2x2_ASAP7_75t_R _23571_ (.A(_00816_),
    .B(_00817_),
    .Y(_15161_));
 XOR2x1_ASAP7_75t_R _23572_ (.A(_15161_),
    .Y(_15162_),
    .B(_12259_));
 NOR2x1_ASAP7_75t_R _23573_ (.A(_15160_),
    .B(_15162_),
    .Y(_15163_));
 XOR2x1_ASAP7_75t_R _23574_ (.A(_15161_),
    .Y(_15164_),
    .B(_12260_));
 NOR2x1_ASAP7_75t_R _23575_ (.A(_15159_),
    .B(_15164_),
    .Y(_15165_));
 OAI21x1_ASAP7_75t_R _23576_ (.A1(_15163_),
    .A2(_15165_),
    .B(_10742_),
    .Y(_15166_));
 NOR2x1_ASAP7_75t_R _23577_ (.A(net780),
    .B(_00676_),
    .Y(_15167_));
 INVx1_ASAP7_75t_R _23578_ (.A(_15167_),
    .Y(_15168_));
 AND2x2_ASAP7_75t_R _23579_ (.A(_15166_),
    .B(_15168_),
    .Y(_15169_));
 XNOR2x2_ASAP7_75t_R _23580_ (.A(_07984_),
    .B(_15169_),
    .Y(_15170_));
 INVx2_ASAP7_75t_R _23581_ (.A(_15170_),
    .Y(_15171_));
 BUFx10_ASAP7_75t_R _23582_ (.A(_15171_),
    .Y(_15172_));
 BUFx10_ASAP7_75t_R _23583_ (.A(_15172_),
    .Y(_15173_));
 OAI21x1_ASAP7_75t_R _23584_ (.A1(_15137_),
    .A2(_15158_),
    .B(_15173_),
    .Y(_15174_));
 INVx1_ASAP7_75t_R _23585_ (.A(_15074_),
    .Y(_15175_));
 INVx1_ASAP7_75t_R _23586_ (.A(_15083_),
    .Y(_15176_));
 INVx3_ASAP7_75t_R _23587_ (.A(_01200_),
    .Y(_15177_));
 AOI21x1_ASAP7_75t_R _23588_ (.A1(_15175_),
    .A2(_15176_),
    .B(_15177_),
    .Y(_15178_));
 NOR2x2_ASAP7_75t_R _23589_ (.A(_15120_),
    .B(_15178_),
    .Y(_15179_));
 INVx1_ASAP7_75t_R _23590_ (.A(_15090_),
    .Y(_15180_));
 INVx1_ASAP7_75t_R _23591_ (.A(_15091_),
    .Y(_15181_));
 INVx1_ASAP7_75t_R _23592_ (.A(_00553_),
    .Y(_15182_));
 AOI21x1_ASAP7_75t_R _23593_ (.A1(_15180_),
    .A2(_15181_),
    .B(_15182_),
    .Y(_15183_));
 BUFx6f_ASAP7_75t_R _23594_ (.A(_15119_),
    .Y(_15184_));
 BUFx6f_ASAP7_75t_R _23595_ (.A(_15184_),
    .Y(_15185_));
 OA21x2_ASAP7_75t_R _23596_ (.A1(_15115_),
    .A2(_15183_),
    .B(_15185_),
    .Y(_15186_));
 BUFx10_ASAP7_75t_R _23597_ (.A(_15135_),
    .Y(_15187_));
 OAI21x1_ASAP7_75t_R _23598_ (.A1(_15179_),
    .A2(_15186_),
    .B(_15187_),
    .Y(_15188_));
 BUFx6f_ASAP7_75t_R _23599_ (.A(_15140_),
    .Y(_15904_));
 INVx3_ASAP7_75t_R _23600_ (.A(net477),
    .Y(_15189_));
 OAI21x1_ASAP7_75t_R _23601_ (.A1(_15090_),
    .A2(_15091_),
    .B(_15189_),
    .Y(_15190_));
 OAI21x1_ASAP7_75t_R _23602_ (.A1(net9),
    .A2(_15916_),
    .B(net5),
    .Y(_15191_));
 NOR2x1_ASAP7_75t_R _23603_ (.A(_15142_),
    .B(_15191_),
    .Y(_15192_));
 NOR2x2_ASAP7_75t_R _23604_ (.A(net904),
    .B(_15085_),
    .Y(_15193_));
 INVx3_ASAP7_75t_R _23605_ (.A(_15138_),
    .Y(_15194_));
 OA21x2_ASAP7_75t_R _23606_ (.A1(_15193_),
    .A2(_15194_),
    .B(_15145_),
    .Y(_15195_));
 BUFx10_ASAP7_75t_R _23607_ (.A(_15149_),
    .Y(_15196_));
 OAI21x1_ASAP7_75t_R _23608_ (.A1(_15192_),
    .A2(_15195_),
    .B(_15196_),
    .Y(_15197_));
 BUFx10_ASAP7_75t_R _23609_ (.A(_15156_),
    .Y(_15198_));
 AOI21x1_ASAP7_75t_R _23610_ (.A1(_15188_),
    .A2(_15197_),
    .B(_15198_),
    .Y(_15199_));
 NAND2x2_ASAP7_75t_R _23611_ (.A(_15063_),
    .B(_15906_),
    .Y(_15200_));
 NOR2x2_ASAP7_75t_R _23612_ (.A(_15085_),
    .B(_15200_),
    .Y(_15201_));
 OAI21x1_ASAP7_75t_R _23613_ (.A1(_15090_),
    .A2(_15091_),
    .B(_15088_),
    .Y(_15202_));
 NAND2x2_ASAP7_75t_R _23614_ (.A(_15110_),
    .B(_15202_),
    .Y(_15203_));
 BUFx10_ASAP7_75t_R _23615_ (.A(_15120_),
    .Y(_15204_));
 OAI21x1_ASAP7_75t_R _23616_ (.A1(_15090_),
    .A2(_15091_),
    .B(_15177_),
    .Y(_15205_));
 INVx1_ASAP7_75t_R _23617_ (.A(_15205_),
    .Y(_15206_));
 BUFx6f_ASAP7_75t_R _23618_ (.A(_15134_),
    .Y(_15207_));
 AOI21x1_ASAP7_75t_R _23619_ (.A1(_15204_),
    .A2(_15206_),
    .B(_15207_),
    .Y(_15208_));
 OAI21x1_ASAP7_75t_R _23620_ (.A1(_15201_),
    .A2(_15203_),
    .B(_15208_),
    .Y(_15209_));
 BUFx6f_ASAP7_75t_R _23621_ (.A(_15109_),
    .Y(_15210_));
 OAI21x1_ASAP7_75t_R _23622_ (.A1(_15074_),
    .A2(_15083_),
    .B(net478),
    .Y(_15211_));
 BUFx6f_ASAP7_75t_R _23623_ (.A(_15211_),
    .Y(_15212_));
 BUFx6f_ASAP7_75t_R _23624_ (.A(_15148_),
    .Y(_15213_));
 AOI21x1_ASAP7_75t_R _23625_ (.A1(_15210_),
    .A2(net900),
    .B(_15213_),
    .Y(_15214_));
 OAI21x1_ASAP7_75t_R _23626_ (.A1(_15074_),
    .A2(_15083_),
    .B(_15093_),
    .Y(_15215_));
 INVx2_ASAP7_75t_R _23627_ (.A(_15215_),
    .Y(_15216_));
 OAI21x1_ASAP7_75t_R _23628_ (.A1(_15206_),
    .A2(_15216_),
    .B(_15185_),
    .Y(_15217_));
 AOI21x1_ASAP7_75t_R _23629_ (.A1(_15214_),
    .A2(_15217_),
    .B(_15157_),
    .Y(_15218_));
 AOI21x1_ASAP7_75t_R _23630_ (.A1(_15209_),
    .A2(_15218_),
    .B(_15172_),
    .Y(_15219_));
 BUFx6f_ASAP7_75t_R _23631_ (.A(_15205_),
    .Y(_15220_));
 AOI21x1_ASAP7_75t_R _23632_ (.A1(_15220_),
    .A2(_15141_),
    .B(_15210_),
    .Y(_15221_));
 BUFx6f_ASAP7_75t_R _23633_ (.A(_15120_),
    .Y(_15222_));
 NOR2x2_ASAP7_75t_R _23634_ (.A(net869),
    .B(_15092_),
    .Y(_15223_));
 AOI21x1_ASAP7_75t_R _23635_ (.A1(_15222_),
    .A2(_15223_),
    .B(_15207_),
    .Y(_15224_));
 OAI21x1_ASAP7_75t_R _23636_ (.A1(_15074_),
    .A2(_15083_),
    .B(_00553_),
    .Y(_15225_));
 INVx2_ASAP7_75t_R _23637_ (.A(_15225_),
    .Y(_15226_));
 NOR2x2_ASAP7_75t_R _23638_ (.A(net841),
    .B(_15092_),
    .Y(_15227_));
 OAI21x1_ASAP7_75t_R _23639_ (.A1(_15226_),
    .A2(_15227_),
    .B(_15210_),
    .Y(_15228_));
 NAND2x1_ASAP7_75t_R _23640_ (.A(_15224_),
    .B(_15228_),
    .Y(_15229_));
 AO21x1_ASAP7_75t_R _23641_ (.A1(_15108_),
    .A2(_15107_),
    .B(_01204_),
    .Y(_15230_));
 INVx2_ASAP7_75t_R _23642_ (.A(_15190_),
    .Y(_15231_));
 AOI21x1_ASAP7_75t_R _23643_ (.A1(_15222_),
    .A2(_15231_),
    .B(_15148_),
    .Y(_15232_));
 CKINVDCx8_ASAP7_75t_R _23644_ (.A(_15156_),
    .Y(_15233_));
 AOI21x1_ASAP7_75t_R _23645_ (.A1(_15230_),
    .A2(_15232_),
    .B(_15233_),
    .Y(_15234_));
 OAI21x1_ASAP7_75t_R _23646_ (.A1(_15221_),
    .A2(_15229_),
    .B(_15234_),
    .Y(_15235_));
 NAND2x1_ASAP7_75t_R _23647_ (.A(_15219_),
    .B(_15235_),
    .Y(_15236_));
 OAI21x1_ASAP7_75t_R _23648_ (.A1(_15174_),
    .A2(_15199_),
    .B(_15236_),
    .Y(_15237_));
 XOR2x1_ASAP7_75t_R _23649_ (.A(_00818_),
    .Y(_15238_),
    .B(net40));
 XOR2x1_ASAP7_75t_R _23650_ (.A(_15238_),
    .Y(_15239_),
    .B(_12276_));
 XOR2x1_ASAP7_75t_R _23651_ (.A(_12085_),
    .Y(_15240_),
    .B(_00786_));
 XOR2x1_ASAP7_75t_R _23652_ (.A(_15239_),
    .Y(_15241_),
    .B(_15240_));
 NOR2x1_ASAP7_75t_R _23653_ (.A(_13017_),
    .B(_00674_),
    .Y(_15242_));
 AO21x1_ASAP7_75t_R _23654_ (.A1(_15241_),
    .A2(_10830_),
    .B(_15242_),
    .Y(_15243_));
 XOR2x2_ASAP7_75t_R _23655_ (.A(_15243_),
    .B(_01074_),
    .Y(_15244_));
 INVx8_ASAP7_75t_R _23656_ (.A(_15244_),
    .Y(_15245_));
 OAI21x1_ASAP7_75t_R _23657_ (.A1(_15906_),
    .A2(_15913_),
    .B(net904),
    .Y(_15246_));
 NAND2x2_ASAP7_75t_R _23658_ (.A(_15204_),
    .B(_15246_),
    .Y(_15247_));
 NAND2x1_ASAP7_75t_R _23659_ (.A(_15212_),
    .B(_15110_),
    .Y(_15248_));
 BUFx4f_ASAP7_75t_R _23660_ (.A(_01202_),
    .Y(_15249_));
 INVx2_ASAP7_75t_R _23661_ (.A(_15249_),
    .Y(_15250_));
 NOR2x2_ASAP7_75t_R _23662_ (.A(_15250_),
    .B(_15094_),
    .Y(_15251_));
 BUFx6f_ASAP7_75t_R _23663_ (.A(_15207_),
    .Y(_15252_));
 OA21x2_ASAP7_75t_R _23664_ (.A1(_15248_),
    .A2(_15251_),
    .B(_15252_),
    .Y(_15253_));
 NAND2x2_ASAP7_75t_R _23665_ (.A(_15177_),
    .B(_15092_),
    .Y(_15254_));
 OAI21x1_ASAP7_75t_R _23666_ (.A1(net39),
    .A2(_15908_),
    .B(_15085_),
    .Y(_15255_));
 BUFx6f_ASAP7_75t_R _23667_ (.A(_15184_),
    .Y(_15256_));
 AOI21x1_ASAP7_75t_R _23668_ (.A1(_15254_),
    .A2(_15255_),
    .B(_15256_),
    .Y(_15257_));
 BUFx6f_ASAP7_75t_R _23669_ (.A(_15134_),
    .Y(_15258_));
 AO21x1_ASAP7_75t_R _23670_ (.A1(_15202_),
    .A2(_15121_),
    .B(_15258_),
    .Y(_15259_));
 BUFx10_ASAP7_75t_R _23671_ (.A(_15172_),
    .Y(_15260_));
 OAI21x1_ASAP7_75t_R _23672_ (.A1(_15257_),
    .A2(_15259_),
    .B(_15260_),
    .Y(_15261_));
 AOI21x1_ASAP7_75t_R _23673_ (.A1(_15247_),
    .A2(_15253_),
    .B(_15261_),
    .Y(_15262_));
 NAND2x1_ASAP7_75t_R _23674_ (.A(_15033_),
    .B(_15035_),
    .Y(_15263_));
 AOI21x1_ASAP7_75t_R _23675_ (.A1(_15020_),
    .A2(net870),
    .B(_12161_),
    .Y(_15264_));
 NAND2x1_ASAP7_75t_R _23676_ (.A(_15263_),
    .B(_15264_),
    .Y(_15265_));
 AOI21x1_ASAP7_75t_R _23677_ (.A1(_15037_),
    .A2(_15265_),
    .B(_07972_),
    .Y(_15266_));
 NOR2x1_ASAP7_75t_R _23678_ (.A(_15139_),
    .B(_15038_),
    .Y(_15267_));
 OAI22x1_ASAP7_75t_R _23679_ (.A1(_15083_),
    .A2(_15074_),
    .B1(_15266_),
    .B2(_15267_),
    .Y(_15268_));
 AOI21x1_ASAP7_75t_R _23680_ (.A1(_15268_),
    .A2(_15255_),
    .B(_15142_),
    .Y(_15269_));
 NAND2x2_ASAP7_75t_R _23681_ (.A(_15063_),
    .B(net843),
    .Y(_15270_));
 NOR2x2_ASAP7_75t_R _23682_ (.A(_15249_),
    .B(_15085_),
    .Y(_15271_));
 INVx1_ASAP7_75t_R _23683_ (.A(_15271_),
    .Y(_15272_));
 BUFx4f_ASAP7_75t_R _23684_ (.A(_15120_),
    .Y(_15273_));
 BUFx6f_ASAP7_75t_R _23685_ (.A(_15273_),
    .Y(_15274_));
 AOI21x1_ASAP7_75t_R _23686_ (.A1(_15270_),
    .A2(_15272_),
    .B(_15274_),
    .Y(_15275_));
 OAI21x1_ASAP7_75t_R _23687_ (.A1(_15269_),
    .A2(_15275_),
    .B(_15187_),
    .Y(_15276_));
 NOR2x2_ASAP7_75t_R _23688_ (.A(_15201_),
    .B(_15203_),
    .Y(_15277_));
 NOR2x1_ASAP7_75t_R _23689_ (.A(_15906_),
    .B(_15913_),
    .Y(_15278_));
 OA21x2_ASAP7_75t_R _23690_ (.A1(_15115_),
    .A2(_15278_),
    .B(_15121_),
    .Y(_15279_));
 OAI21x1_ASAP7_75t_R _23691_ (.A1(_15277_),
    .A2(_15279_),
    .B(_15196_),
    .Y(_15280_));
 AOI21x1_ASAP7_75t_R _23692_ (.A1(_15276_),
    .A2(_15280_),
    .B(_15173_),
    .Y(_15281_));
 BUFx10_ASAP7_75t_R _23693_ (.A(_15233_),
    .Y(_15282_));
 OAI21x1_ASAP7_75t_R _23694_ (.A1(_15262_),
    .A2(_15281_),
    .B(_15282_),
    .Y(_15283_));
 OAI21x1_ASAP7_75t_R _23695_ (.A1(_15074_),
    .A2(_15083_),
    .B(_15189_),
    .Y(_15284_));
 INVx1_ASAP7_75t_R _23696_ (.A(_15284_),
    .Y(_15285_));
 BUFx4f_ASAP7_75t_R _23697_ (.A(_15144_),
    .Y(_15286_));
 OA21x2_ASAP7_75t_R _23698_ (.A1(_15285_),
    .A2(_15183_),
    .B(_15286_),
    .Y(_15287_));
 OA21x2_ASAP7_75t_R _23699_ (.A1(_15226_),
    .A2(_15194_),
    .B(_15121_),
    .Y(_15288_));
 OAI21x1_ASAP7_75t_R _23700_ (.A1(_15287_),
    .A2(_15288_),
    .B(_15196_),
    .Y(_15289_));
 BUFx6f_ASAP7_75t_R _23701_ (.A(_15109_),
    .Y(_15290_));
 OAI21x1_ASAP7_75t_R _23702_ (.A1(_15090_),
    .A2(_15091_),
    .B(net479),
    .Y(_15291_));
 AOI21x1_ASAP7_75t_R _23703_ (.A1(_15290_),
    .A2(_15291_),
    .B(_15213_),
    .Y(_15292_));
 NAND2x2_ASAP7_75t_R _23704_ (.A(_15039_),
    .B(net842),
    .Y(_15293_));
 NAND2x2_ASAP7_75t_R _23705_ (.A(_15284_),
    .B(_15120_),
    .Y(_15294_));
 INVx2_ASAP7_75t_R _23706_ (.A(_15294_),
    .Y(_15295_));
 NAND2x1_ASAP7_75t_R _23707_ (.A(_15293_),
    .B(_15295_),
    .Y(_15296_));
 AOI21x1_ASAP7_75t_R _23708_ (.A1(_15292_),
    .A2(_15296_),
    .B(_15260_),
    .Y(_15297_));
 AOI21x1_ASAP7_75t_R _23709_ (.A1(_15297_),
    .A2(_15289_),
    .B(_15282_),
    .Y(_15298_));
 AOI21x1_ASAP7_75t_R _23710_ (.A1(_15112_),
    .A2(_15270_),
    .B(_15286_),
    .Y(_15299_));
 OAI21x1_ASAP7_75t_R _23711_ (.A1(net9),
    .A2(_15908_),
    .B(_15144_),
    .Y(_15300_));
 OAI21x1_ASAP7_75t_R _23712_ (.A1(_15227_),
    .A2(_15300_),
    .B(_15207_),
    .Y(_15301_));
 NOR2x1_ASAP7_75t_R _23713_ (.A(_15299_),
    .B(_15301_),
    .Y(_15302_));
 OAI21x1_ASAP7_75t_R _23714_ (.A1(net39),
    .A2(net841),
    .B(_15085_),
    .Y(_15303_));
 BUFx6f_ASAP7_75t_R _23715_ (.A(_15110_),
    .Y(_15304_));
 AOI21x1_ASAP7_75t_R _23716_ (.A1(net558),
    .A2(_15303_),
    .B(_15304_),
    .Y(_15305_));
 OA21x2_ASAP7_75t_R _23717_ (.A1(_15083_),
    .A2(_15074_),
    .B(_00551_),
    .Y(_15306_));
 OAI21x1_ASAP7_75t_R _23718_ (.A1(_15183_),
    .A2(_15306_),
    .B(_15210_),
    .Y(_15307_));
 NAND2x1_ASAP7_75t_R _23719_ (.A(_15149_),
    .B(_15307_),
    .Y(_15308_));
 NOR2x1_ASAP7_75t_R _23720_ (.A(_15305_),
    .B(_15308_),
    .Y(_15309_));
 OAI21x1_ASAP7_75t_R _23721_ (.A1(_15302_),
    .A2(_15309_),
    .B(_15173_),
    .Y(_15310_));
 AOI21x1_ASAP7_75t_R _23722_ (.A1(_15310_),
    .A2(_15298_),
    .B(_15245_),
    .Y(_15311_));
 AOI22x1_ASAP7_75t_R _23723_ (.A1(_15237_),
    .A2(_15245_),
    .B1(_15311_),
    .B2(_15283_),
    .Y(_00080_));
 AO21x1_ASAP7_75t_R _23724_ (.A1(_15225_),
    .A2(_15190_),
    .B(_15273_),
    .Y(_15312_));
 OAI21x1_ASAP7_75t_R _23725_ (.A1(_15227_),
    .A2(_15115_),
    .B(_15204_),
    .Y(_15313_));
 AOI21x1_ASAP7_75t_R _23726_ (.A1(_15312_),
    .A2(_15313_),
    .B(_15149_),
    .Y(_15314_));
 NOR2x2_ASAP7_75t_R _23727_ (.A(_15908_),
    .B(_15085_),
    .Y(_15315_));
 OAI21x1_ASAP7_75t_R _23728_ (.A1(_15183_),
    .A2(_15315_),
    .B(_15204_),
    .Y(_15316_));
 NAND2x2_ASAP7_75t_R _23729_ (.A(net567),
    .B(net843),
    .Y(_15317_));
 BUFx6f_ASAP7_75t_R _23730_ (.A(_15317_),
    .Y(_15318_));
 NAND2x1_ASAP7_75t_R _23731_ (.A(_15318_),
    .B(_15179_),
    .Y(_15319_));
 AOI21x1_ASAP7_75t_R _23732_ (.A1(_15316_),
    .A2(_15319_),
    .B(_15258_),
    .Y(_15320_));
 OAI21x1_ASAP7_75t_R _23733_ (.A1(_15314_),
    .A2(_15320_),
    .B(_15172_),
    .Y(_15321_));
 BUFx6f_ASAP7_75t_R _23734_ (.A(_15213_),
    .Y(_15322_));
 INVx2_ASAP7_75t_R _23735_ (.A(net869),
    .Y(_15323_));
 NOR2x2_ASAP7_75t_R _23736_ (.A(_15323_),
    .B(_15913_),
    .Y(_15324_));
 AOI21x1_ASAP7_75t_R _23737_ (.A1(_15249_),
    .A2(_15094_),
    .B(_15144_),
    .Y(_15325_));
 INVx1_ASAP7_75t_R _23738_ (.A(_15325_),
    .Y(_15326_));
 INVx3_ASAP7_75t_R _23739_ (.A(_15211_),
    .Y(_15327_));
 AOI21x1_ASAP7_75t_R _23740_ (.A1(_15906_),
    .A2(_15908_),
    .B(_15094_),
    .Y(_15328_));
 OAI21x1_ASAP7_75t_R _23741_ (.A1(_15327_),
    .A2(_15328_),
    .B(_15290_),
    .Y(_15329_));
 OAI21x1_ASAP7_75t_R _23742_ (.A1(_15324_),
    .A2(_15326_),
    .B(_15329_),
    .Y(_15330_));
 NOR2x2_ASAP7_75t_R _23743_ (.A(_15120_),
    .B(_15327_),
    .Y(_15331_));
 NOR2x1_ASAP7_75t_R _23744_ (.A(_15207_),
    .B(_15331_),
    .Y(_15332_));
 AOI21x1_ASAP7_75t_R _23745_ (.A1(_15906_),
    .A2(_15908_),
    .B(_15085_),
    .Y(_15333_));
 BUFx6f_ASAP7_75t_R _23746_ (.A(_15120_),
    .Y(_15334_));
 OAI21x1_ASAP7_75t_R _23747_ (.A1(_15227_),
    .A2(_15333_),
    .B(_15334_),
    .Y(_15335_));
 AOI21x1_ASAP7_75t_R _23748_ (.A1(_15332_),
    .A2(_15335_),
    .B(_15172_),
    .Y(_15336_));
 OAI21x1_ASAP7_75t_R _23749_ (.A1(_15322_),
    .A2(_15330_),
    .B(_15336_),
    .Y(_15337_));
 AOI21x1_ASAP7_75t_R _23750_ (.A1(_15321_),
    .A2(_15337_),
    .B(_15157_),
    .Y(_15338_));
 INVx1_ASAP7_75t_R _23751_ (.A(_15183_),
    .Y(_15339_));
 OAI21x1_ASAP7_75t_R _23752_ (.A1(_15083_),
    .A2(_15074_),
    .B(_15063_),
    .Y(_15340_));
 AO21x1_ASAP7_75t_R _23753_ (.A1(_15339_),
    .A2(_15340_),
    .B(_15110_),
    .Y(_15341_));
 OAI21x1_ASAP7_75t_R _23754_ (.A1(net39),
    .A2(_15903_),
    .B(_15092_),
    .Y(_15342_));
 AO21x1_ASAP7_75t_R _23755_ (.A1(_15342_),
    .A2(_15255_),
    .B(_15273_),
    .Y(_15343_));
 AOI21x1_ASAP7_75t_R _23756_ (.A1(_15341_),
    .A2(_15343_),
    .B(_15149_),
    .Y(_15344_));
 BUFx6f_ASAP7_75t_R _23757_ (.A(_15134_),
    .Y(_15345_));
 OAI21x1_ASAP7_75t_R _23758_ (.A1(_15194_),
    .A2(_15333_),
    .B(_15204_),
    .Y(_15346_));
 NAND2x1_ASAP7_75t_R _23759_ (.A(_00555_),
    .B(_15144_),
    .Y(_15347_));
 AO21x1_ASAP7_75t_R _23760_ (.A1(_15347_),
    .A2(_15148_),
    .B(_15171_),
    .Y(_15348_));
 OAI21x1_ASAP7_75t_R _23761_ (.A1(_15345_),
    .A2(_15346_),
    .B(_15348_),
    .Y(_15349_));
 NAND2x2_ASAP7_75t_R _23762_ (.A(_15903_),
    .B(_15092_),
    .Y(_15350_));
 BUFx4f_ASAP7_75t_R _23763_ (.A(_15109_),
    .Y(_15351_));
 AO21x1_ASAP7_75t_R _23764_ (.A1(_15350_),
    .A2(_15317_),
    .B(_15351_),
    .Y(_15352_));
 AND3x1_ASAP7_75t_R _23765_ (.A(_15166_),
    .B(_07984_),
    .C(_15168_),
    .Y(_15353_));
 NOR2x1_ASAP7_75t_R _23766_ (.A(_07984_),
    .B(_15169_),
    .Y(_15354_));
 OAI21x1_ASAP7_75t_R _23767_ (.A1(_15353_),
    .A2(_15354_),
    .B(_15134_),
    .Y(_15355_));
 AOI21x1_ASAP7_75t_R _23768_ (.A1(_15318_),
    .A2(_15179_),
    .B(_15355_),
    .Y(_15356_));
 AOI21x1_ASAP7_75t_R _23769_ (.A1(_15352_),
    .A2(_15356_),
    .B(_15233_),
    .Y(_15357_));
 OAI21x1_ASAP7_75t_R _23770_ (.A1(_15344_),
    .A2(_15349_),
    .B(_15357_),
    .Y(_15358_));
 NAND2x1_ASAP7_75t_R _23771_ (.A(_15244_),
    .B(_15358_),
    .Y(_15359_));
 NOR2x1_ASAP7_75t_R _23772_ (.A(_15338_),
    .B(_15359_),
    .Y(_15360_));
 AND2x2_ASAP7_75t_R _23773_ (.A(_15141_),
    .B(_15205_),
    .Y(_15361_));
 NAND2x2_ASAP7_75t_R _23774_ (.A(_15249_),
    .B(_15094_),
    .Y(_15362_));
 INVx2_ASAP7_75t_R _23775_ (.A(_15291_),
    .Y(_15363_));
 NOR2x2_ASAP7_75t_R _23776_ (.A(_15363_),
    .B(_15120_),
    .Y(_15364_));
 AOI21x1_ASAP7_75t_R _23777_ (.A1(_15364_),
    .A2(_15362_),
    .B(_15207_),
    .Y(_15365_));
 OAI21x1_ASAP7_75t_R _23778_ (.A1(_15145_),
    .A2(_15361_),
    .B(_15365_),
    .Y(_15366_));
 OA21x2_ASAP7_75t_R _23779_ (.A1(_15144_),
    .A2(_15220_),
    .B(_15134_),
    .Y(_15367_));
 NOR2x2_ASAP7_75t_R _23780_ (.A(net39),
    .B(_15092_),
    .Y(_15368_));
 NOR2x2_ASAP7_75t_R _23781_ (.A(_15039_),
    .B(net842),
    .Y(_15369_));
 INVx2_ASAP7_75t_R _23782_ (.A(_15369_),
    .Y(_15370_));
 OA21x2_ASAP7_75t_R _23783_ (.A1(_15368_),
    .A2(_15184_),
    .B(_15370_),
    .Y(_15371_));
 AOI21x1_ASAP7_75t_R _23784_ (.A1(_15367_),
    .A2(_15371_),
    .B(_15172_),
    .Y(_15372_));
 NAND2x1_ASAP7_75t_R _23785_ (.A(_15372_),
    .B(_15366_),
    .Y(_15373_));
 OAI21x1_ASAP7_75t_R _23786_ (.A1(net904),
    .A2(_15094_),
    .B(_15284_),
    .Y(_15374_));
 NAND2x1_ASAP7_75t_R _23787_ (.A(_15374_),
    .B(_15290_),
    .Y(_15375_));
 NOR2x2_ASAP7_75t_R _23788_ (.A(_15144_),
    .B(_15178_),
    .Y(_15376_));
 AOI21x1_ASAP7_75t_R _23789_ (.A1(_15270_),
    .A2(_15376_),
    .B(_15213_),
    .Y(_15377_));
 NAND2x1_ASAP7_75t_R _23790_ (.A(_15377_),
    .B(_15375_),
    .Y(_15378_));
 NOR2x1_ASAP7_75t_R _23791_ (.A(_15903_),
    .B(_15906_),
    .Y(_15379_));
 OAI21x1_ASAP7_75t_R _23792_ (.A1(_15379_),
    .A2(_15368_),
    .B(_15204_),
    .Y(_15380_));
 NOR2x2_ASAP7_75t_R _23793_ (.A(_15094_),
    .B(_15184_),
    .Y(_15381_));
 AOI21x1_ASAP7_75t_R _23794_ (.A1(_15112_),
    .A2(_15381_),
    .B(_15135_),
    .Y(_15382_));
 AOI21x1_ASAP7_75t_R _23795_ (.A1(_15380_),
    .A2(_15382_),
    .B(_15170_),
    .Y(_15383_));
 AOI21x1_ASAP7_75t_R _23796_ (.A1(_15383_),
    .A2(_15378_),
    .B(_15233_),
    .Y(_15384_));
 NAND2x1_ASAP7_75t_R _23797_ (.A(_15373_),
    .B(_15384_),
    .Y(_15385_));
 AO21x1_ASAP7_75t_R _23798_ (.A1(_15220_),
    .A2(_15212_),
    .B(_15273_),
    .Y(_15386_));
 AO21x1_ASAP7_75t_R _23799_ (.A1(_15270_),
    .A2(_15225_),
    .B(_15351_),
    .Y(_15387_));
 AOI21x1_ASAP7_75t_R _23800_ (.A1(_15386_),
    .A2(_15387_),
    .B(_15149_),
    .Y(_15388_));
 AO21x1_ASAP7_75t_R _23801_ (.A1(_15340_),
    .A2(_15291_),
    .B(_15351_),
    .Y(_15389_));
 AO21x1_ASAP7_75t_R _23802_ (.A1(_15350_),
    .A2(_15200_),
    .B(_15222_),
    .Y(_15390_));
 AOI21x1_ASAP7_75t_R _23803_ (.A1(_15389_),
    .A2(_15390_),
    .B(_15345_),
    .Y(_15391_));
 BUFx6f_ASAP7_75t_R _23804_ (.A(_15170_),
    .Y(_15392_));
 OAI21x1_ASAP7_75t_R _23805_ (.A1(_15388_),
    .A2(_15391_),
    .B(_15392_),
    .Y(_15393_));
 NAND2x1_ASAP7_75t_R _23806_ (.A(_15204_),
    .B(_15333_),
    .Y(_15394_));
 AOI21x1_ASAP7_75t_R _23807_ (.A1(_15249_),
    .A2(_15085_),
    .B(_15184_),
    .Y(_15395_));
 AOI21x1_ASAP7_75t_R _23808_ (.A1(_15370_),
    .A2(_15395_),
    .B(_15213_),
    .Y(_15396_));
 NAND2x1_ASAP7_75t_R _23809_ (.A(_15394_),
    .B(_15396_),
    .Y(_15397_));
 OA21x2_ASAP7_75t_R _23810_ (.A1(_15254_),
    .A2(_15351_),
    .B(_15148_),
    .Y(_15398_));
 AOI21x1_ASAP7_75t_R _23811_ (.A1(_15329_),
    .A2(_15398_),
    .B(_15170_),
    .Y(_15399_));
 AOI21x1_ASAP7_75t_R _23812_ (.A1(_15397_),
    .A2(_15399_),
    .B(_15157_),
    .Y(_15400_));
 NAND2x1_ASAP7_75t_R _23813_ (.A(_15393_),
    .B(_15400_),
    .Y(_15401_));
 AOI21x1_ASAP7_75t_R _23814_ (.A1(_15385_),
    .A2(_15401_),
    .B(_15244_),
    .Y(_15402_));
 NOR2x2_ASAP7_75t_R _23815_ (.A(_15402_),
    .B(_15360_),
    .Y(_00081_));
 AOI21x1_ASAP7_75t_R _23816_ (.A1(net5),
    .A2(_15268_),
    .B(_15142_),
    .Y(_15403_));
 AOI21x1_ASAP7_75t_R _23817_ (.A1(_15220_),
    .A2(_15141_),
    .B(_15274_),
    .Y(_15404_));
 OAI21x1_ASAP7_75t_R _23818_ (.A1(_15403_),
    .A2(_15404_),
    .B(_15196_),
    .Y(_15405_));
 AOI21x1_ASAP7_75t_R _23819_ (.A1(_15908_),
    .A2(_15916_),
    .B(net9),
    .Y(_15406_));
 NOR2x2_ASAP7_75t_R _23820_ (.A(_15121_),
    .B(_15406_),
    .Y(_15407_));
 OAI21x1_ASAP7_75t_R _23821_ (.A1(_15177_),
    .A2(_15916_),
    .B(_15222_),
    .Y(_15408_));
 NOR2x1_ASAP7_75t_R _23822_ (.A(_15251_),
    .B(_15408_),
    .Y(_15409_));
 OAI21x1_ASAP7_75t_R _23823_ (.A1(_15407_),
    .A2(_15409_),
    .B(_15187_),
    .Y(_15410_));
 AOI21x1_ASAP7_75t_R _23824_ (.A1(_15405_),
    .A2(_15410_),
    .B(_15173_),
    .Y(_15411_));
 NAND2x1_ASAP7_75t_R _23825_ (.A(_15318_),
    .B(_15295_),
    .Y(_15412_));
 BUFx6f_ASAP7_75t_R _23826_ (.A(_15340_),
    .Y(_15413_));
 AOI21x1_ASAP7_75t_R _23827_ (.A1(_15323_),
    .A2(_15916_),
    .B(_15334_),
    .Y(_15414_));
 NAND2x1_ASAP7_75t_R _23828_ (.A(_15413_),
    .B(_15414_),
    .Y(_15415_));
 AOI21x1_ASAP7_75t_R _23829_ (.A1(_15415_),
    .A2(_15412_),
    .B(_15196_),
    .Y(_15416_));
 AOI21x1_ASAP7_75t_R _23830_ (.A1(_15303_),
    .A2(_15272_),
    .B(_15274_),
    .Y(_15417_));
 BUFx6f_ASAP7_75t_R _23831_ (.A(_15148_),
    .Y(_15418_));
 OAI21x1_ASAP7_75t_R _23832_ (.A1(_15913_),
    .A2(_15112_),
    .B(_15185_),
    .Y(_15419_));
 NAND2x1_ASAP7_75t_R _23833_ (.A(_15418_),
    .B(_15419_),
    .Y(_15420_));
 OAI21x1_ASAP7_75t_R _23834_ (.A1(_15417_),
    .A2(_15420_),
    .B(_15260_),
    .Y(_15421_));
 OAI21x1_ASAP7_75t_R _23835_ (.A1(_15421_),
    .A2(_15416_),
    .B(_15198_),
    .Y(_15422_));
 OAI21x1_ASAP7_75t_R _23836_ (.A1(_15422_),
    .A2(_15411_),
    .B(_15244_),
    .Y(_15423_));
 AOI21x1_ASAP7_75t_R _23837_ (.A1(_15291_),
    .A2(_15284_),
    .B(_15256_),
    .Y(_15424_));
 OAI21x1_ASAP7_75t_R _23838_ (.A1(_15090_),
    .A2(_15091_),
    .B(_15093_),
    .Y(_15425_));
 AOI21x1_ASAP7_75t_R _23839_ (.A1(_15425_),
    .A2(_15340_),
    .B(_15110_),
    .Y(_15426_));
 OAI21x1_ASAP7_75t_R _23840_ (.A1(_15424_),
    .A2(_15426_),
    .B(_15322_),
    .Y(_15427_));
 OAI21x1_ASAP7_75t_R _23841_ (.A1(_15090_),
    .A2(_15091_),
    .B(_15250_),
    .Y(_15428_));
 AOI21x1_ASAP7_75t_R _23842_ (.A1(_15428_),
    .A2(_15413_),
    .B(_15304_),
    .Y(_15429_));
 AOI21x1_ASAP7_75t_R _23843_ (.A1(_15215_),
    .A2(_15318_),
    .B(_15256_),
    .Y(_15430_));
 OAI21x1_ASAP7_75t_R _23844_ (.A1(_15429_),
    .A2(_15430_),
    .B(_15252_),
    .Y(_15431_));
 BUFx10_ASAP7_75t_R _23845_ (.A(_15170_),
    .Y(_15432_));
 AOI21x1_ASAP7_75t_R _23846_ (.A1(_15427_),
    .A2(_15431_),
    .B(_15432_),
    .Y(_15433_));
 AOI21x1_ASAP7_75t_R _23847_ (.A1(_15215_),
    .A2(_15428_),
    .B(_15145_),
    .Y(_15434_));
 AOI21x1_ASAP7_75t_R _23848_ (.A1(_15220_),
    .A2(_15413_),
    .B(_15121_),
    .Y(_15435_));
 OAI21x1_ASAP7_75t_R _23849_ (.A1(_15434_),
    .A2(_15435_),
    .B(_15252_),
    .Y(_15436_));
 AOI21x1_ASAP7_75t_R _23850_ (.A1(_15220_),
    .A2(_15215_),
    .B(_15145_),
    .Y(_15437_));
 AOI21x1_ASAP7_75t_R _23851_ (.A1(_15220_),
    .A2(_15268_),
    .B(_15256_),
    .Y(_15438_));
 OAI21x1_ASAP7_75t_R _23852_ (.A1(_15437_),
    .A2(_15438_),
    .B(_15322_),
    .Y(_15439_));
 AOI21x1_ASAP7_75t_R _23853_ (.A1(_15436_),
    .A2(_15439_),
    .B(_15260_),
    .Y(_15440_));
 NOR3x1_ASAP7_75t_R _23854_ (.A(_15433_),
    .B(_15440_),
    .C(_15198_),
    .Y(_15441_));
 NAND2x1_ASAP7_75t_R _23855_ (.A(_00551_),
    .B(_15092_),
    .Y(_15442_));
 AND3x1_ASAP7_75t_R _23856_ (.A(_15442_),
    .B(_15304_),
    .C(net5),
    .Y(_15443_));
 AND3x1_ASAP7_75t_R _23857_ (.A(_15339_),
    .B(_15268_),
    .C(_15256_),
    .Y(_15444_));
 OAI21x1_ASAP7_75t_R _23858_ (.A1(_15443_),
    .A2(_15444_),
    .B(_15187_),
    .Y(_15445_));
 NAND2x1_ASAP7_75t_R _23859_ (.A(_00555_),
    .B(_15274_),
    .Y(_15446_));
 NAND2x2_ASAP7_75t_R _23860_ (.A(net904),
    .B(_15904_),
    .Y(_15447_));
 AOI21x1_ASAP7_75t_R _23861_ (.A1(_15906_),
    .A2(_15094_),
    .B(_15120_),
    .Y(_15448_));
 AOI21x1_ASAP7_75t_R _23862_ (.A1(_15447_),
    .A2(_15448_),
    .B(_15207_),
    .Y(_15449_));
 AOI21x1_ASAP7_75t_R _23863_ (.A1(_15446_),
    .A2(_15449_),
    .B(_15198_),
    .Y(_15450_));
 AND3x2_ASAP7_75t_R _23864_ (.A(_15118_),
    .B(_15117_),
    .C(_00556_),
    .Y(_15451_));
 NOR2x2_ASAP7_75t_R _23865_ (.A(_15063_),
    .B(net569),
    .Y(_15452_));
 AOI21x1_ASAP7_75t_R _23866_ (.A1(_15916_),
    .A2(_15452_),
    .B(_15304_),
    .Y(_15453_));
 OAI21x1_ASAP7_75t_R _23867_ (.A1(_15451_),
    .A2(_15453_),
    .B(_15196_),
    .Y(_15454_));
 NOR2x1_ASAP7_75t_R _23868_ (.A(_01206_),
    .B(_15304_),
    .Y(_15455_));
 OAI21x1_ASAP7_75t_R _23869_ (.A1(_15455_),
    .A2(_15407_),
    .B(_15187_),
    .Y(_15456_));
 AOI21x1_ASAP7_75t_R _23870_ (.A1(_15454_),
    .A2(_15456_),
    .B(_15282_),
    .Y(_15457_));
 AOI211x1_ASAP7_75t_R _23871_ (.A1(_15445_),
    .A2(_15450_),
    .B(_15457_),
    .C(_15173_),
    .Y(_15458_));
 OAI21x1_ASAP7_75t_R _23872_ (.A1(_01204_),
    .A2(_15142_),
    .B(_15418_),
    .Y(_15459_));
 AOI21x1_ASAP7_75t_R _23873_ (.A1(net5),
    .A2(_15141_),
    .B(_15274_),
    .Y(_15460_));
 OAI21x1_ASAP7_75t_R _23874_ (.A1(_15459_),
    .A2(_15460_),
    .B(_15282_),
    .Y(_15461_));
 OAI21x1_ASAP7_75t_R _23875_ (.A1(_15304_),
    .A2(_15191_),
    .B(_15345_),
    .Y(_15462_));
 NAND2x2_ASAP7_75t_R _23876_ (.A(_15109_),
    .B(_15317_),
    .Y(_15463_));
 NOR2x1_ASAP7_75t_R _23877_ (.A(_15315_),
    .B(_15463_),
    .Y(_15464_));
 NOR2x1_ASAP7_75t_R _23878_ (.A(_15462_),
    .B(_15464_),
    .Y(_15465_));
 OAI21x1_ASAP7_75t_R _23879_ (.A1(_15461_),
    .A2(_15465_),
    .B(_15173_),
    .Y(_15466_));
 AND2x2_ASAP7_75t_R _23880_ (.A(_01199_),
    .B(_01200_),
    .Y(_15467_));
 INVx1_ASAP7_75t_R _23881_ (.A(_15467_),
    .Y(_15468_));
 OAI21x1_ASAP7_75t_R _23882_ (.A1(_15074_),
    .A2(_15083_),
    .B(_15468_),
    .Y(_15469_));
 AO21x1_ASAP7_75t_R _23883_ (.A1(_15303_),
    .A2(_15469_),
    .B(_15274_),
    .Y(_15470_));
 AND2x2_ASAP7_75t_R _23884_ (.A(_15346_),
    .B(_15345_),
    .Y(_15471_));
 OA21x2_ASAP7_75t_R _23885_ (.A1(_15290_),
    .A2(_15225_),
    .B(_15213_),
    .Y(_15472_));
 AO21x1_ASAP7_75t_R _23886_ (.A1(_15220_),
    .A2(_15284_),
    .B(_15334_),
    .Y(_15473_));
 AO21x1_ASAP7_75t_R _23887_ (.A1(_15472_),
    .A2(_15473_),
    .B(_15233_),
    .Y(_15474_));
 AOI21x1_ASAP7_75t_R _23888_ (.A1(_15470_),
    .A2(_15471_),
    .B(_15474_),
    .Y(_15475_));
 OAI21x1_ASAP7_75t_R _23889_ (.A1(_15466_),
    .A2(_15475_),
    .B(_15245_),
    .Y(_15476_));
 OAI22x1_ASAP7_75t_R _23890_ (.A1(_15423_),
    .A2(_15441_),
    .B1(_15458_),
    .B2(_15476_),
    .Y(_00082_));
 AO21x1_ASAP7_75t_R _23891_ (.A1(_15228_),
    .A2(_15380_),
    .B(_15252_),
    .Y(_15477_));
 AOI21x1_ASAP7_75t_R _23892_ (.A1(_15215_),
    .A2(_15202_),
    .B(_15222_),
    .Y(_15478_));
 INVx1_ASAP7_75t_R _23893_ (.A(_15478_),
    .Y(_15479_));
 AO21x1_ASAP7_75t_R _23894_ (.A1(_15284_),
    .A2(_15428_),
    .B(_15290_),
    .Y(_15480_));
 AO21x1_ASAP7_75t_R _23895_ (.A1(_15479_),
    .A2(_15480_),
    .B(_15322_),
    .Y(_15481_));
 AOI21x1_ASAP7_75t_R _23896_ (.A1(_15477_),
    .A2(_15481_),
    .B(_15432_),
    .Y(_15482_));
 AO21x1_ASAP7_75t_R _23897_ (.A1(_15425_),
    .A2(_15469_),
    .B(_15273_),
    .Y(_15483_));
 NAND2x1_ASAP7_75t_R _23898_ (.A(_15483_),
    .B(_15346_),
    .Y(_15484_));
 AND2x2_ASAP7_75t_R _23899_ (.A(_15273_),
    .B(_15428_),
    .Y(_15485_));
 AOI21x1_ASAP7_75t_R _23900_ (.A1(_15413_),
    .A2(_15485_),
    .B(_15418_),
    .Y(_15486_));
 AOI21x1_ASAP7_75t_R _23901_ (.A1(_15322_),
    .A2(_15484_),
    .B(_15486_),
    .Y(_15487_));
 OAI21x1_ASAP7_75t_R _23902_ (.A1(_15173_),
    .A2(_15487_),
    .B(_15282_),
    .Y(_15488_));
 NAND2x2_ASAP7_75t_R _23903_ (.A(_15184_),
    .B(_15327_),
    .Y(_15489_));
 INVx1_ASAP7_75t_R _23904_ (.A(_15115_),
    .Y(_15490_));
 OAI22x1_ASAP7_75t_R _23905_ (.A1(_15489_),
    .A2(_15170_),
    .B1(_15256_),
    .B2(_15490_),
    .Y(_15491_));
 NAND2x1_ASAP7_75t_R _23906_ (.A(_15290_),
    .B(_15363_),
    .Y(_15492_));
 OAI21x1_ASAP7_75t_R _23907_ (.A1(_15194_),
    .A2(_15369_),
    .B(_15185_),
    .Y(_15493_));
 AOI21x1_ASAP7_75t_R _23908_ (.A1(_15492_),
    .A2(_15493_),
    .B(_15172_),
    .Y(_15494_));
 OAI21x1_ASAP7_75t_R _23909_ (.A1(_15491_),
    .A2(_15494_),
    .B(_15252_),
    .Y(_15495_));
 AO21x1_ASAP7_75t_R _23910_ (.A1(_15428_),
    .A2(_15469_),
    .B(_15222_),
    .Y(_15496_));
 AOI21x1_ASAP7_75t_R _23911_ (.A1(_15334_),
    .A2(_15374_),
    .B(_15171_),
    .Y(_15497_));
 NAND2x1_ASAP7_75t_R _23912_ (.A(_15496_),
    .B(_15497_),
    .Y(_15498_));
 AOI21x1_ASAP7_75t_R _23913_ (.A1(_15210_),
    .A2(_15216_),
    .B(_15170_),
    .Y(_15499_));
 INVx1_ASAP7_75t_R _23914_ (.A(_15426_),
    .Y(_15500_));
 AOI21x1_ASAP7_75t_R _23915_ (.A1(_15499_),
    .A2(_15500_),
    .B(_15345_),
    .Y(_15501_));
 AOI21x1_ASAP7_75t_R _23916_ (.A1(_15498_),
    .A2(_15501_),
    .B(_15233_),
    .Y(_15502_));
 AOI21x1_ASAP7_75t_R _23917_ (.A1(_15495_),
    .A2(_15502_),
    .B(_15245_),
    .Y(_15503_));
 OAI21x1_ASAP7_75t_R _23918_ (.A1(_15482_),
    .A2(_15488_),
    .B(_15503_),
    .Y(_15504_));
 NAND2x1_ASAP7_75t_R _23919_ (.A(_15442_),
    .B(_15270_),
    .Y(_15505_));
 NOR2x1_ASAP7_75t_R _23920_ (.A(_15286_),
    .B(_15505_),
    .Y(_15506_));
 AO21x1_ASAP7_75t_R _23921_ (.A1(_15225_),
    .A2(_15364_),
    .B(_15506_),
    .Y(_15507_));
 OA21x2_ASAP7_75t_R _23922_ (.A1(_15271_),
    .A2(_15206_),
    .B(_15286_),
    .Y(_15508_));
 AO21x1_ASAP7_75t_R _23923_ (.A1(_15318_),
    .A2(_15295_),
    .B(_15135_),
    .Y(_15509_));
 OAI21x1_ASAP7_75t_R _23924_ (.A1(_15508_),
    .A2(_15509_),
    .B(_15157_),
    .Y(_15510_));
 AOI21x1_ASAP7_75t_R _23925_ (.A1(_15187_),
    .A2(_15507_),
    .B(_15510_),
    .Y(_15511_));
 AND3x1_ASAP7_75t_R _23926_ (.A(_15184_),
    .B(net900),
    .C(_15138_),
    .Y(_15512_));
 NOR2x1_ASAP7_75t_R _23927_ (.A(_15512_),
    .B(_15301_),
    .Y(_15513_));
 NAND2x1_ASAP7_75t_R _23928_ (.A(_15190_),
    .B(_15184_),
    .Y(_15514_));
 OAI21x1_ASAP7_75t_R _23929_ (.A1(_15333_),
    .A2(_15514_),
    .B(_15213_),
    .Y(_15515_));
 NOR2x1_ASAP7_75t_R _23930_ (.A(_15463_),
    .B(_15505_),
    .Y(_15516_));
 NOR2x1_ASAP7_75t_R _23931_ (.A(_15515_),
    .B(_15516_),
    .Y(_15517_));
 OAI21x1_ASAP7_75t_R _23932_ (.A1(_15513_),
    .A2(_15517_),
    .B(_15233_),
    .Y(_15518_));
 NAND2x1_ASAP7_75t_R _23933_ (.A(_15260_),
    .B(_15518_),
    .Y(_15519_));
 NAND2x1_ASAP7_75t_R _23934_ (.A(_15913_),
    .B(_15290_),
    .Y(_15520_));
 AOI21x1_ASAP7_75t_R _23935_ (.A1(_15112_),
    .A2(_15413_),
    .B(_15207_),
    .Y(_15521_));
 AOI21x1_ASAP7_75t_R _23936_ (.A1(_15520_),
    .A2(_15521_),
    .B(_15156_),
    .Y(_15522_));
 AO21x1_ASAP7_75t_R _23937_ (.A1(_15212_),
    .A2(_15425_),
    .B(_15351_),
    .Y(_15523_));
 NAND2x1_ASAP7_75t_R _23938_ (.A(_15523_),
    .B(_15396_),
    .Y(_15524_));
 NAND2x1_ASAP7_75t_R _23939_ (.A(_15522_),
    .B(_15524_),
    .Y(_15525_));
 OAI21x1_ASAP7_75t_R _23940_ (.A1(_15193_),
    .A2(_15368_),
    .B(_15185_),
    .Y(_15526_));
 AOI21x1_ASAP7_75t_R _23941_ (.A1(_15292_),
    .A2(_15526_),
    .B(_15233_),
    .Y(_15527_));
 AO21x1_ASAP7_75t_R _23942_ (.A1(_15270_),
    .A2(_15447_),
    .B(_15351_),
    .Y(_15528_));
 AOI21x1_ASAP7_75t_R _23943_ (.A1(_15318_),
    .A2(_15331_),
    .B(_15135_),
    .Y(_15529_));
 NAND2x1_ASAP7_75t_R _23944_ (.A(_15528_),
    .B(_15529_),
    .Y(_15530_));
 AOI21x1_ASAP7_75t_R _23945_ (.A1(_15527_),
    .A2(_15530_),
    .B(_15260_),
    .Y(_15531_));
 AOI21x1_ASAP7_75t_R _23946_ (.A1(_15525_),
    .A2(_15531_),
    .B(_15244_),
    .Y(_15532_));
 OAI21x1_ASAP7_75t_R _23947_ (.A1(_15519_),
    .A2(_15511_),
    .B(_15532_),
    .Y(_15533_));
 NAND2x1_ASAP7_75t_R _23948_ (.A(_15504_),
    .B(_15533_),
    .Y(_00083_));
 OAI21x1_ASAP7_75t_R _23949_ (.A1(net620),
    .A2(_15913_),
    .B(_15185_),
    .Y(_15534_));
 NAND2x1_ASAP7_75t_R _23950_ (.A(_15144_),
    .B(_15293_),
    .Y(_15535_));
 AOI21x1_ASAP7_75t_R _23951_ (.A1(_15534_),
    .A2(_15535_),
    .B(_15315_),
    .Y(_15536_));
 NOR2x1_ASAP7_75t_R _23952_ (.A(_15213_),
    .B(_15115_),
    .Y(_15537_));
 AOI21x1_ASAP7_75t_R _23953_ (.A1(_15111_),
    .A2(_15537_),
    .B(_15392_),
    .Y(_15538_));
 OAI21x1_ASAP7_75t_R _23954_ (.A1(_15252_),
    .A2(_15536_),
    .B(_15538_),
    .Y(_15539_));
 NAND2x1_ASAP7_75t_R _23955_ (.A(_15282_),
    .B(_15539_),
    .Y(_15540_));
 AOI21x1_ASAP7_75t_R _23956_ (.A1(_15112_),
    .A2(_15318_),
    .B(_15304_),
    .Y(_15541_));
 NOR2x1_ASAP7_75t_R _23957_ (.A(net9),
    .B(_15916_),
    .Y(_15542_));
 OA21x2_ASAP7_75t_R _23958_ (.A1(_15542_),
    .A2(_15183_),
    .B(_15145_),
    .Y(_15543_));
 OAI21x1_ASAP7_75t_R _23959_ (.A1(_15541_),
    .A2(_15543_),
    .B(_15187_),
    .Y(_15544_));
 OA21x2_ASAP7_75t_R _23960_ (.A1(_15368_),
    .A2(_15379_),
    .B(_15145_),
    .Y(_15545_));
 OA21x2_ASAP7_75t_R _23961_ (.A1(_15315_),
    .A2(_15278_),
    .B(_15121_),
    .Y(_15546_));
 OAI21x1_ASAP7_75t_R _23962_ (.A1(_15545_),
    .A2(_15546_),
    .B(_15196_),
    .Y(_15547_));
 AOI21x1_ASAP7_75t_R _23963_ (.A1(_15544_),
    .A2(_15547_),
    .B(_15173_),
    .Y(_15548_));
 OAI21x1_ASAP7_75t_R _23964_ (.A1(_15540_),
    .A2(_15548_),
    .B(_15245_),
    .Y(_15549_));
 OAI21x1_ASAP7_75t_R _23965_ (.A1(_15251_),
    .A2(_15408_),
    .B(_15258_),
    .Y(_15550_));
 NOR2x1_ASAP7_75t_R _23966_ (.A(_15113_),
    .B(_15463_),
    .Y(_15551_));
 OAI21x1_ASAP7_75t_R _23967_ (.A1(_15550_),
    .A2(_15551_),
    .B(_15392_),
    .Y(_15552_));
 NAND2x1_ASAP7_75t_R _23968_ (.A(_15225_),
    .B(_15293_),
    .Y(_15553_));
 AOI211x1_ASAP7_75t_R _23969_ (.A1(_15142_),
    .A2(_15553_),
    .B(_15252_),
    .C(_15221_),
    .Y(_15554_));
 NOR2x1_ASAP7_75t_R _23970_ (.A(_15552_),
    .B(_15554_),
    .Y(_15555_));
 OA21x2_ASAP7_75t_R _23971_ (.A1(_15222_),
    .A2(_15190_),
    .B(_15215_),
    .Y(_15556_));
 AO21x1_ASAP7_75t_R _23972_ (.A1(_15367_),
    .A2(_15556_),
    .B(_15392_),
    .Y(_15557_));
 OAI21x1_ASAP7_75t_R _23973_ (.A1(_15363_),
    .A2(_15326_),
    .B(_15418_),
    .Y(_15558_));
 NOR2x1_ASAP7_75t_R _23974_ (.A(_15114_),
    .B(_15558_),
    .Y(_15559_));
 OAI21x1_ASAP7_75t_R _23975_ (.A1(_15557_),
    .A2(_15559_),
    .B(_15198_),
    .Y(_15560_));
 NOR2x1_ASAP7_75t_R _23976_ (.A(_15555_),
    .B(_15560_),
    .Y(_15561_));
 NOR2x1_ASAP7_75t_R _23977_ (.A(_15227_),
    .B(_15300_),
    .Y(_15562_));
 OAI21x1_ASAP7_75t_R _23978_ (.A1(_15562_),
    .A2(_15186_),
    .B(_15322_),
    .Y(_15563_));
 NOR2x1_ASAP7_75t_R _23979_ (.A(_15193_),
    .B(_15111_),
    .Y(_15564_));
 AND3x1_ASAP7_75t_R _23980_ (.A(_15318_),
    .B(_15334_),
    .C(_15112_),
    .Y(_15565_));
 OAI21x1_ASAP7_75t_R _23981_ (.A1(_15564_),
    .A2(_15565_),
    .B(_15252_),
    .Y(_15566_));
 AOI21x1_ASAP7_75t_R _23982_ (.A1(_15563_),
    .A2(_15566_),
    .B(_15173_),
    .Y(_15567_));
 AO21x1_ASAP7_75t_R _23983_ (.A1(_15118_),
    .A2(_15117_),
    .B(_00557_),
    .Y(_15568_));
 OAI21x1_ASAP7_75t_R _23984_ (.A1(_15121_),
    .A2(net5),
    .B(_15568_),
    .Y(_15569_));
 AO21x1_ASAP7_75t_R _23985_ (.A1(_15569_),
    .A2(_15322_),
    .B(_15392_),
    .Y(_15570_));
 NOR2x1_ASAP7_75t_R _23986_ (.A(_15369_),
    .B(_15111_),
    .Y(_15571_));
 NOR2x1_ASAP7_75t_R _23987_ (.A(_15286_),
    .B(_15370_),
    .Y(_15572_));
 OAI21x1_ASAP7_75t_R _23988_ (.A1(_15145_),
    .A2(_15413_),
    .B(_15258_),
    .Y(_15573_));
 NOR3x1_ASAP7_75t_R _23989_ (.A(_15571_),
    .B(_15572_),
    .C(_15573_),
    .Y(_15574_));
 OAI21x1_ASAP7_75t_R _23990_ (.A1(_15570_),
    .A2(_15574_),
    .B(_15198_),
    .Y(_15575_));
 NOR2x1_ASAP7_75t_R _23991_ (.A(_15567_),
    .B(_15575_),
    .Y(_15576_));
 NAND2x1_ASAP7_75t_R _23992_ (.A(_15225_),
    .B(_15318_),
    .Y(_15577_));
 AOI22x1_ASAP7_75t_R _23993_ (.A1(_15577_),
    .A2(_15274_),
    .B1(_15179_),
    .B2(_15318_),
    .Y(_15578_));
 AOI21x1_ASAP7_75t_R _23994_ (.A1(_15428_),
    .A2(_15350_),
    .B(_15304_),
    .Y(_15579_));
 AO21x1_ASAP7_75t_R _23995_ (.A1(_15286_),
    .A2(_15916_),
    .B(_15135_),
    .Y(_15580_));
 OAI21x1_ASAP7_75t_R _23996_ (.A1(_15579_),
    .A2(_15580_),
    .B(_15432_),
    .Y(_15581_));
 AOI21x1_ASAP7_75t_R _23997_ (.A1(_15187_),
    .A2(_15578_),
    .B(_15581_),
    .Y(_15582_));
 OAI21x1_ASAP7_75t_R _23998_ (.A1(_15142_),
    .A2(_15324_),
    .B(_15345_),
    .Y(_15583_));
 OA21x2_ASAP7_75t_R _23999_ (.A1(_15200_),
    .A2(_15913_),
    .B(_15286_),
    .Y(_15584_));
 OAI21x1_ASAP7_75t_R _24000_ (.A1(_15583_),
    .A2(_15584_),
    .B(_15260_),
    .Y(_15585_));
 OAI21x1_ASAP7_75t_R _24001_ (.A1(_15231_),
    .A2(_15408_),
    .B(_15418_),
    .Y(_15586_));
 NOR2x1_ASAP7_75t_R _24002_ (.A(_15277_),
    .B(_15586_),
    .Y(_15587_));
 OAI21x1_ASAP7_75t_R _24003_ (.A1(_15585_),
    .A2(_15587_),
    .B(_15282_),
    .Y(_15588_));
 OAI21x1_ASAP7_75t_R _24004_ (.A1(_15582_),
    .A2(_15588_),
    .B(_15244_),
    .Y(_15589_));
 OAI22x1_ASAP7_75t_R _24005_ (.A1(_15549_),
    .A2(_15561_),
    .B1(_15576_),
    .B2(_15589_),
    .Y(_00084_));
 AO21x1_ASAP7_75t_R _24006_ (.A1(_15231_),
    .A2(_15210_),
    .B(_15149_),
    .Y(_15590_));
 OA21x2_ASAP7_75t_R _24007_ (.A1(_15369_),
    .A2(_15223_),
    .B(_15121_),
    .Y(_15591_));
 OAI21x1_ASAP7_75t_R _24008_ (.A1(_15590_),
    .A2(_15591_),
    .B(_15392_),
    .Y(_15592_));
 NOR2x1_ASAP7_75t_R _24009_ (.A(_15183_),
    .B(_15248_),
    .Y(_15593_));
 OA21x2_ASAP7_75t_R _24010_ (.A1(_15593_),
    .A2(_15485_),
    .B(_15418_),
    .Y(_15594_));
 OAI21x1_ASAP7_75t_R _24011_ (.A1(_15592_),
    .A2(_15594_),
    .B(_15198_),
    .Y(_15595_));
 NOR2x1_ASAP7_75t_R _24012_ (.A(net9),
    .B(_15256_),
    .Y(_15596_));
 OAI21x1_ASAP7_75t_R _24013_ (.A1(_15596_),
    .A2(_15541_),
    .B(_15196_),
    .Y(_15597_));
 AOI21x1_ASAP7_75t_R _24014_ (.A1(_15200_),
    .A2(_15202_),
    .B(_15142_),
    .Y(_15598_));
 OA21x2_ASAP7_75t_R _24015_ (.A1(_15333_),
    .A2(_15194_),
    .B(_15286_),
    .Y(_15599_));
 OAI21x1_ASAP7_75t_R _24016_ (.A1(_15598_),
    .A2(_15599_),
    .B(_15187_),
    .Y(_15600_));
 AOI21x1_ASAP7_75t_R _24017_ (.A1(_15597_),
    .A2(_15600_),
    .B(_15432_),
    .Y(_15601_));
 NOR2x1_ASAP7_75t_R _24018_ (.A(_15595_),
    .B(_15601_),
    .Y(_15602_));
 AO21x1_ASAP7_75t_R _24019_ (.A1(_15121_),
    .A2(net900),
    .B(_15258_),
    .Y(_15603_));
 OAI21x1_ASAP7_75t_R _24020_ (.A1(_15478_),
    .A2(_15603_),
    .B(_15432_),
    .Y(_15604_));
 AOI211x1_ASAP7_75t_R _24021_ (.A1(_15381_),
    .A2(_15112_),
    .B(_15376_),
    .C(_15322_),
    .Y(_15605_));
 OAI21x1_ASAP7_75t_R _24022_ (.A1(_15604_),
    .A2(_15605_),
    .B(_15282_),
    .Y(_15606_));
 AOI21x1_ASAP7_75t_R _24023_ (.A1(_15220_),
    .A2(_15469_),
    .B(_15256_),
    .Y(_15607_));
 OAI21x1_ASAP7_75t_R _24024_ (.A1(_15093_),
    .A2(_15913_),
    .B(_15204_),
    .Y(_15608_));
 NOR2x1_ASAP7_75t_R _24025_ (.A(_15608_),
    .B(_15113_),
    .Y(_15609_));
 OAI21x1_ASAP7_75t_R _24026_ (.A1(_15607_),
    .A2(_15609_),
    .B(_15187_),
    .Y(_15610_));
 AOI21x1_ASAP7_75t_R _24027_ (.A1(_15428_),
    .A2(_15254_),
    .B(_15274_),
    .Y(_15611_));
 OAI21x1_ASAP7_75t_R _24028_ (.A1(_15611_),
    .A2(_15279_),
    .B(_15196_),
    .Y(_15612_));
 AOI21x1_ASAP7_75t_R _24029_ (.A1(_15610_),
    .A2(_15612_),
    .B(_15432_),
    .Y(_15613_));
 OAI21x1_ASAP7_75t_R _24030_ (.A1(_15606_),
    .A2(_15613_),
    .B(_15245_),
    .Y(_15614_));
 NOR2x1_ASAP7_75t_R _24031_ (.A(_15142_),
    .B(_15201_),
    .Y(_15615_));
 AO21x1_ASAP7_75t_R _24032_ (.A1(_15304_),
    .A2(_00551_),
    .B(_15345_),
    .Y(_15616_));
 OA21x2_ASAP7_75t_R _24033_ (.A1(_15615_),
    .A2(_15616_),
    .B(_15432_),
    .Y(_15617_));
 INVx1_ASAP7_75t_R _24034_ (.A(_00551_),
    .Y(_15618_));
 NAND2x1_ASAP7_75t_R _24035_ (.A(_15618_),
    .B(_15916_),
    .Y(_15619_));
 INVx1_ASAP7_75t_R _24036_ (.A(_15251_),
    .Y(_15620_));
 AO221x1_ASAP7_75t_R _24037_ (.A1(_15619_),
    .A2(_15331_),
    .B1(_15295_),
    .B2(_15620_),
    .C(_15322_),
    .Y(_15621_));
 NAND2x1_ASAP7_75t_R _24038_ (.A(_15467_),
    .B(_15913_),
    .Y(_15622_));
 AOI21x1_ASAP7_75t_R _24039_ (.A1(_15145_),
    .A2(_15622_),
    .B(_15258_),
    .Y(_15623_));
 OA21x2_ASAP7_75t_R _24040_ (.A1(_15201_),
    .A2(_15419_),
    .B(_15623_),
    .Y(_15624_));
 INVx1_ASAP7_75t_R _24041_ (.A(_15395_),
    .Y(_15625_));
 AO21x1_ASAP7_75t_R _24042_ (.A1(_15367_),
    .A2(_15625_),
    .B(_15392_),
    .Y(_15626_));
 OAI21x1_ASAP7_75t_R _24043_ (.A1(_15624_),
    .A2(_15626_),
    .B(_15198_),
    .Y(_15627_));
 AOI21x1_ASAP7_75t_R _24044_ (.A1(_15621_),
    .A2(_15617_),
    .B(_15627_),
    .Y(_15628_));
 AO21x1_ASAP7_75t_R _24045_ (.A1(_15194_),
    .A2(_15210_),
    .B(_15149_),
    .Y(_15629_));
 AOI21x1_ASAP7_75t_R _24046_ (.A1(_15428_),
    .A2(_15342_),
    .B(_15304_),
    .Y(_15630_));
 OAI21x1_ASAP7_75t_R _24047_ (.A1(_15629_),
    .A2(_15630_),
    .B(_15392_),
    .Y(_15631_));
 NOR2x2_ASAP7_75t_R _24048_ (.A(_15144_),
    .B(_15340_),
    .Y(_15632_));
 NOR2x1_ASAP7_75t_R _24049_ (.A(_15632_),
    .B(_15209_),
    .Y(_15633_));
 NOR2x1_ASAP7_75t_R _24050_ (.A(_15631_),
    .B(_15633_),
    .Y(_15634_));
 AO21x1_ASAP7_75t_R _24051_ (.A1(_15908_),
    .A2(_15286_),
    .B(_15258_),
    .Y(_15635_));
 OAI21x1_ASAP7_75t_R _24052_ (.A1(_15299_),
    .A2(_15635_),
    .B(_15260_),
    .Y(_15636_));
 AOI21x1_ASAP7_75t_R _24053_ (.A1(net558),
    .A2(_15255_),
    .B(_15256_),
    .Y(_15637_));
 OAI21x1_ASAP7_75t_R _24054_ (.A1(_15369_),
    .A2(_15608_),
    .B(_15345_),
    .Y(_15638_));
 NOR2x1_ASAP7_75t_R _24055_ (.A(_15637_),
    .B(_15638_),
    .Y(_15639_));
 OAI21x1_ASAP7_75t_R _24056_ (.A1(_15636_),
    .A2(_15639_),
    .B(_15282_),
    .Y(_15640_));
 OAI21x1_ASAP7_75t_R _24057_ (.A1(_15634_),
    .A2(_15640_),
    .B(_15244_),
    .Y(_15641_));
 OAI22x1_ASAP7_75t_R _24058_ (.A1(_15602_),
    .A2(_15614_),
    .B1(_15641_),
    .B2(_15628_),
    .Y(_00085_));
 NAND2x1_ASAP7_75t_R _24059_ (.A(_01205_),
    .B(_01203_),
    .Y(_15642_));
 AO21x1_ASAP7_75t_R _24060_ (.A1(_15185_),
    .A2(_15642_),
    .B(_15135_),
    .Y(_15643_));
 NOR2x1_ASAP7_75t_R _24061_ (.A(_15452_),
    .B(_15463_),
    .Y(_15644_));
 OAI21x1_ASAP7_75t_R _24062_ (.A1(_15643_),
    .A2(_15644_),
    .B(_15260_),
    .Y(_15645_));
 OA21x2_ASAP7_75t_R _24063_ (.A1(_15223_),
    .A2(_15216_),
    .B(_15210_),
    .Y(_15646_));
 AOI211x1_ASAP7_75t_R _24064_ (.A1(_15274_),
    .A2(_15226_),
    .B(_15646_),
    .C(_15322_),
    .Y(_15647_));
 OAI21x1_ASAP7_75t_R _24065_ (.A1(_15645_),
    .A2(_15647_),
    .B(_15282_),
    .Y(_15648_));
 AND2x2_ASAP7_75t_R _24066_ (.A(_15220_),
    .B(_15215_),
    .Y(_15649_));
 OAI21x1_ASAP7_75t_R _24067_ (.A1(_15145_),
    .A2(_15413_),
    .B(_15232_),
    .Y(_15650_));
 AO21x1_ASAP7_75t_R _24068_ (.A1(_15649_),
    .A2(_15414_),
    .B(_15650_),
    .Y(_15651_));
 AO21x1_ASAP7_75t_R _24069_ (.A1(_15490_),
    .A2(_15303_),
    .B(_15334_),
    .Y(_15652_));
 INVx1_ASAP7_75t_R _24070_ (.A(_15425_),
    .Y(_15653_));
 OAI21x1_ASAP7_75t_R _24071_ (.A1(_15653_),
    .A2(_15271_),
    .B(_15334_),
    .Y(_15654_));
 AO21x1_ASAP7_75t_R _24072_ (.A1(_15652_),
    .A2(_15654_),
    .B(_15252_),
    .Y(_15655_));
 AOI21x1_ASAP7_75t_R _24073_ (.A1(_15651_),
    .A2(_15655_),
    .B(_15173_),
    .Y(_15656_));
 NOR2x1_ASAP7_75t_R _24074_ (.A(_15648_),
    .B(_15656_),
    .Y(_15657_));
 NOR2x1_ASAP7_75t_R _24075_ (.A(_15324_),
    .B(_15294_),
    .Y(_15658_));
 AOI21x1_ASAP7_75t_R _24076_ (.A1(_15268_),
    .A2(_15255_),
    .B(_15274_),
    .Y(_15659_));
 OAI21x1_ASAP7_75t_R _24077_ (.A1(_15658_),
    .A2(_15659_),
    .B(_15196_),
    .Y(_15660_));
 AND2x2_ASAP7_75t_R _24078_ (.A(_15489_),
    .B(_15258_),
    .Y(_15661_));
 OAI21x1_ASAP7_75t_R _24079_ (.A1(_15453_),
    .A2(_15451_),
    .B(_15661_),
    .Y(_15662_));
 AOI21x1_ASAP7_75t_R _24080_ (.A1(_15660_),
    .A2(_15662_),
    .B(_15432_),
    .Y(_15663_));
 AO21x1_ASAP7_75t_R _24081_ (.A1(_15413_),
    .A2(_15906_),
    .B(_15185_),
    .Y(_15664_));
 OA21x2_ASAP7_75t_R _24082_ (.A1(_15290_),
    .A2(_15138_),
    .B(_15135_),
    .Y(_15665_));
 AO21x1_ASAP7_75t_R _24083_ (.A1(_15664_),
    .A2(_15665_),
    .B(_15172_),
    .Y(_15666_));
 AOI21x1_ASAP7_75t_R _24084_ (.A1(net904),
    .A2(_15381_),
    .B(_15135_),
    .Y(_15667_));
 AO21x1_ASAP7_75t_R _24085_ (.A1(_15413_),
    .A2(_15447_),
    .B(_15334_),
    .Y(_15668_));
 AO21x1_ASAP7_75t_R _24086_ (.A1(_15291_),
    .A2(_15469_),
    .B(_15290_),
    .Y(_15669_));
 AND3x1_ASAP7_75t_R _24087_ (.A(_15667_),
    .B(_15668_),
    .C(_15669_),
    .Y(_15670_));
 OAI21x1_ASAP7_75t_R _24088_ (.A1(_15666_),
    .A2(_15670_),
    .B(_15198_),
    .Y(_15671_));
 OAI21x1_ASAP7_75t_R _24089_ (.A1(_15663_),
    .A2(_15671_),
    .B(_15245_),
    .Y(_15672_));
 NOR2x1_ASAP7_75t_R _24090_ (.A(_15369_),
    .B(_15608_),
    .Y(_15673_));
 AO21x1_ASAP7_75t_R _24091_ (.A1(_15286_),
    .A2(_00558_),
    .B(_15258_),
    .Y(_15674_));
 AO21x1_ASAP7_75t_R _24092_ (.A1(_15212_),
    .A2(_15428_),
    .B(_15222_),
    .Y(_15675_));
 OA21x2_ASAP7_75t_R _24093_ (.A1(_15270_),
    .A2(_15351_),
    .B(_15207_),
    .Y(_15676_));
 AOI21x1_ASAP7_75t_R _24094_ (.A1(_15675_),
    .A2(_15676_),
    .B(_15233_),
    .Y(_15677_));
 OAI21x1_ASAP7_75t_R _24095_ (.A1(_15673_),
    .A2(_15674_),
    .B(_15677_),
    .Y(_15678_));
 NAND2x1_ASAP7_75t_R _24096_ (.A(net9),
    .B(_15334_),
    .Y(_15679_));
 AOI21x1_ASAP7_75t_R _24097_ (.A1(_15679_),
    .A2(_15521_),
    .B(_15157_),
    .Y(_15680_));
 AOI21x1_ASAP7_75t_R _24098_ (.A1(net9),
    .A2(net904),
    .B(_15273_),
    .Y(_15681_));
 OAI21x1_ASAP7_75t_R _24099_ (.A1(_15681_),
    .A2(_15325_),
    .B(_15270_),
    .Y(_15682_));
 NAND2x1_ASAP7_75t_R _24100_ (.A(_15345_),
    .B(_15682_),
    .Y(_15683_));
 AOI21x1_ASAP7_75t_R _24101_ (.A1(_15680_),
    .A2(_15683_),
    .B(_15432_),
    .Y(_15684_));
 NAND2x1_ASAP7_75t_R _24102_ (.A(_15684_),
    .B(_15678_),
    .Y(_15685_));
 AOI21x1_ASAP7_75t_R _24103_ (.A1(_15210_),
    .A2(_15293_),
    .B(_15149_),
    .Y(_15686_));
 AOI21x1_ASAP7_75t_R _24104_ (.A1(_15686_),
    .A2(_15247_),
    .B(_15157_),
    .Y(_15687_));
 OAI21x1_ASAP7_75t_R _24105_ (.A1(_15185_),
    .A2(_15216_),
    .B(_15294_),
    .Y(_15688_));
 NAND2x1_ASAP7_75t_R _24106_ (.A(_15667_),
    .B(_15688_),
    .Y(_15689_));
 AOI21x1_ASAP7_75t_R _24107_ (.A1(_15687_),
    .A2(_15689_),
    .B(_15260_),
    .Y(_15690_));
 AOI21x1_ASAP7_75t_R _24108_ (.A1(_15142_),
    .A2(_15361_),
    .B(_15252_),
    .Y(_15691_));
 NAND2x1_ASAP7_75t_R _24109_ (.A(_15185_),
    .B(_15619_),
    .Y(_15692_));
 AO21x1_ASAP7_75t_R _24110_ (.A1(_15268_),
    .A2(_15425_),
    .B(_15273_),
    .Y(_15693_));
 AOI21x1_ASAP7_75t_R _24111_ (.A1(_15692_),
    .A2(_15693_),
    .B(_15418_),
    .Y(_15694_));
 OAI21x1_ASAP7_75t_R _24112_ (.A1(_15691_),
    .A2(_15694_),
    .B(_15157_),
    .Y(_15695_));
 AOI21x1_ASAP7_75t_R _24113_ (.A1(_15690_),
    .A2(_15695_),
    .B(_15245_),
    .Y(_15696_));
 NAND2x1_ASAP7_75t_R _24114_ (.A(_15696_),
    .B(_15685_),
    .Y(_15697_));
 OAI21x1_ASAP7_75t_R _24115_ (.A1(_15657_),
    .A2(_15672_),
    .B(_15697_),
    .Y(_00086_));
 AO21x1_ASAP7_75t_R _24116_ (.A1(_15303_),
    .A2(_15268_),
    .B(_15110_),
    .Y(_15698_));
 NAND2x1_ASAP7_75t_R _24117_ (.A(_15698_),
    .B(_15449_),
    .Y(_15699_));
 AO21x1_ASAP7_75t_R _24118_ (.A1(_15118_),
    .A2(_15117_),
    .B(_15908_),
    .Y(_15700_));
 OAI21x1_ASAP7_75t_R _24119_ (.A1(_15315_),
    .A2(_15535_),
    .B(_15700_),
    .Y(_15701_));
 AOI21x1_ASAP7_75t_R _24120_ (.A1(_15258_),
    .A2(_15701_),
    .B(_15170_),
    .Y(_15702_));
 NAND2x1_ASAP7_75t_R _24121_ (.A(_15699_),
    .B(_15702_),
    .Y(_15703_));
 OA21x2_ASAP7_75t_R _24122_ (.A1(_15342_),
    .A2(_15184_),
    .B(_15148_),
    .Y(_15704_));
 NAND2x1_ASAP7_75t_R _24123_ (.A(_15489_),
    .B(_15704_),
    .Y(_15705_));
 AO21x1_ASAP7_75t_R _24124_ (.A1(_15303_),
    .A2(net900),
    .B(_15351_),
    .Y(_15706_));
 NAND2x1_ASAP7_75t_R _24125_ (.A(_15094_),
    .B(_15452_),
    .Y(_15707_));
 AOI21x1_ASAP7_75t_R _24126_ (.A1(_15290_),
    .A2(_15707_),
    .B(_15213_),
    .Y(_15708_));
 AOI21x1_ASAP7_75t_R _24127_ (.A1(_15706_),
    .A2(_15708_),
    .B(_15172_),
    .Y(_15709_));
 AOI21x1_ASAP7_75t_R _24128_ (.A1(_15705_),
    .A2(_15709_),
    .B(_15233_),
    .Y(_15710_));
 NAND2x1_ASAP7_75t_R _24129_ (.A(_15703_),
    .B(_15710_),
    .Y(_15711_));
 AOI21x1_ASAP7_75t_R _24130_ (.A1(_15204_),
    .A2(_15362_),
    .B(_15135_),
    .Y(_15712_));
 AOI21x1_ASAP7_75t_R _24131_ (.A1(_15712_),
    .A2(_15693_),
    .B(_15170_),
    .Y(_15713_));
 AO21x1_ASAP7_75t_R _24132_ (.A1(_15303_),
    .A2(_15225_),
    .B(_15273_),
    .Y(_15714_));
 AO21x1_ASAP7_75t_R _24133_ (.A1(_15094_),
    .A2(net9),
    .B(_15908_),
    .Y(_15715_));
 AOI21x1_ASAP7_75t_R _24134_ (.A1(_15334_),
    .A2(_15715_),
    .B(_15213_),
    .Y(_15716_));
 NAND2x1_ASAP7_75t_R _24135_ (.A(_15714_),
    .B(_15716_),
    .Y(_15717_));
 AOI21x1_ASAP7_75t_R _24136_ (.A1(_15713_),
    .A2(_15717_),
    .B(_15157_),
    .Y(_15718_));
 NAND2x1_ASAP7_75t_R _24137_ (.A(_15374_),
    .B(_15204_),
    .Y(_15719_));
 NAND2x1_ASAP7_75t_R _24138_ (.A(_15364_),
    .B(_15362_),
    .Y(_15720_));
 AOI21x1_ASAP7_75t_R _24139_ (.A1(_15719_),
    .A2(_15720_),
    .B(_15418_),
    .Y(_15721_));
 AO21x1_ASAP7_75t_R _24140_ (.A1(_15293_),
    .A2(_15413_),
    .B(_15222_),
    .Y(_15722_));
 AOI21x1_ASAP7_75t_R _24141_ (.A1(_15654_),
    .A2(_15722_),
    .B(_15345_),
    .Y(_15723_));
 OAI21x1_ASAP7_75t_R _24142_ (.A1(_15721_),
    .A2(_15723_),
    .B(_15432_),
    .Y(_15724_));
 AOI21x1_ASAP7_75t_R _24143_ (.A1(_15718_),
    .A2(_15724_),
    .B(_15245_),
    .Y(_15725_));
 NAND2x1_ASAP7_75t_R _24144_ (.A(_15711_),
    .B(_15725_),
    .Y(_15726_));
 INVx1_ASAP7_75t_R _24145_ (.A(_00557_),
    .Y(_15727_));
 OAI21x1_ASAP7_75t_R _24146_ (.A1(_15727_),
    .A2(_15256_),
    .B(_15224_),
    .Y(_15728_));
 OAI21x1_ASAP7_75t_R _24147_ (.A1(_15906_),
    .A2(_15144_),
    .B(_15134_),
    .Y(_01427_));
 NOR2x1_ASAP7_75t_R _24148_ (.A(_01427_),
    .B(_15632_),
    .Y(_01428_));
 NAND2x1_ASAP7_75t_R _24149_ (.A(_15319_),
    .B(_01428_),
    .Y(_01429_));
 AOI21x1_ASAP7_75t_R _24150_ (.A1(_15728_),
    .A2(_01429_),
    .B(_15392_),
    .Y(_01430_));
 AND3x1_ASAP7_75t_R _24151_ (.A(_15118_),
    .B(_15117_),
    .C(_01205_),
    .Y(_01431_));
 NAND2x1_ASAP7_75t_R _24152_ (.A(_15215_),
    .B(_15291_),
    .Y(_01432_));
 OAI21x1_ASAP7_75t_R _24153_ (.A1(_15210_),
    .A2(_01432_),
    .B(_15149_),
    .Y(_01433_));
 OAI21x1_ASAP7_75t_R _24154_ (.A1(_01431_),
    .A2(_01433_),
    .B(_15170_),
    .Y(_01434_));
 AO21x1_ASAP7_75t_R _24155_ (.A1(_15190_),
    .A2(_15212_),
    .B(_15222_),
    .Y(_01435_));
 AO21x1_ASAP7_75t_R _24156_ (.A1(_15270_),
    .A2(_15268_),
    .B(_15351_),
    .Y(_01436_));
 AOI21x1_ASAP7_75t_R _24157_ (.A1(_01435_),
    .A2(_01436_),
    .B(_15418_),
    .Y(_01437_));
 OAI21x1_ASAP7_75t_R _24158_ (.A1(_01434_),
    .A2(_01437_),
    .B(_15157_),
    .Y(_01438_));
 NOR2x1_ASAP7_75t_R _24159_ (.A(_01430_),
    .B(_01438_),
    .Y(_01439_));
 OA21x2_ASAP7_75t_R _24160_ (.A1(_15351_),
    .A2(_01200_),
    .B(_15207_),
    .Y(_01440_));
 OAI21x1_ASAP7_75t_R _24161_ (.A1(_15452_),
    .A2(_15463_),
    .B(_01440_),
    .Y(_01441_));
 OA21x2_ASAP7_75t_R _24162_ (.A1(_15317_),
    .A2(_15273_),
    .B(_15225_),
    .Y(_01442_));
 AOI21x1_ASAP7_75t_R _24163_ (.A1(_15224_),
    .A2(_01442_),
    .B(_15172_),
    .Y(_01443_));
 NAND2x1_ASAP7_75t_R _24164_ (.A(_01441_),
    .B(_01443_),
    .Y(_01444_));
 NAND2x1_ASAP7_75t_R _24165_ (.A(_15225_),
    .B(_15184_),
    .Y(_01445_));
 NOR2x1_ASAP7_75t_R _24166_ (.A(_15328_),
    .B(_01445_),
    .Y(_01446_));
 AND3x1_ASAP7_75t_R _24167_ (.A(_15110_),
    .B(net900),
    .C(_15138_),
    .Y(_01447_));
 OAI21x1_ASAP7_75t_R _24168_ (.A1(_01446_),
    .A2(_01447_),
    .B(_15418_),
    .Y(_01448_));
 NOR2x1_ASAP7_75t_R _24169_ (.A(_15110_),
    .B(_15202_),
    .Y(_01449_));
 NOR2x1_ASAP7_75t_R _24170_ (.A(_01427_),
    .B(_01449_),
    .Y(_01450_));
 AOI21x1_ASAP7_75t_R _24171_ (.A1(_15483_),
    .A2(_01450_),
    .B(_15392_),
    .Y(_01451_));
 NAND2x1_ASAP7_75t_R _24172_ (.A(_01448_),
    .B(_01451_),
    .Y(_01452_));
 AOI21x1_ASAP7_75t_R _24173_ (.A1(_01444_),
    .A2(_01452_),
    .B(_15198_),
    .Y(_01453_));
 OAI21x1_ASAP7_75t_R _24174_ (.A1(_01439_),
    .A2(_01453_),
    .B(_15245_),
    .Y(_01454_));
 NAND2x2_ASAP7_75t_R _24175_ (.A(_15726_),
    .B(_01454_),
    .Y(_00087_));
 NOR2x2_ASAP7_75t_R _24176_ (.A(net641),
    .B(_00559_),
    .Y(_01455_));
 INVx1_ASAP7_75t_R _24177_ (.A(_12870_),
    .Y(_01456_));
 XOR2x1_ASAP7_75t_R _24178_ (.A(net645),
    .Y(_01457_),
    .B(_01456_));
 XNOR2x2_ASAP7_75t_R _24179_ (.A(net911),
    .B(_13011_),
    .Y(_01458_));
 XOR2x2_ASAP7_75t_R _24180_ (.A(_12831_),
    .B(_12836_),
    .Y(_01459_));
 XOR2x1_ASAP7_75t_R _24181_ (.A(_01458_),
    .Y(_01460_),
    .B(_01459_));
 NAND2x1_ASAP7_75t_R _24182_ (.A(_01457_),
    .B(_01460_),
    .Y(_01461_));
 XOR2x1_ASAP7_75t_R _24183_ (.A(net646),
    .Y(_01462_),
    .B(_12870_));
 XOR2x2_ASAP7_75t_R _24184_ (.A(_13011_),
    .B(_00820_),
    .Y(_01463_));
 XOR2x1_ASAP7_75t_R _24185_ (.A(_01463_),
    .Y(_01464_),
    .B(_01459_));
 NAND2x1_ASAP7_75t_R _24186_ (.A(_01462_),
    .B(_01464_),
    .Y(_01465_));
 AOI21x1_ASAP7_75t_R _24187_ (.A1(_01461_),
    .A2(_01465_),
    .B(_11370_),
    .Y(_01466_));
 OAI21x1_ASAP7_75t_R _24188_ (.A1(_01455_),
    .A2(_01466_),
    .B(_07973_),
    .Y(_01467_));
 AND2x2_ASAP7_75t_R _24189_ (.A(_10640_),
    .B(_00559_),
    .Y(_01468_));
 NAND2x1_ASAP7_75t_R _24190_ (.A(_01462_),
    .B(_01460_),
    .Y(_01469_));
 NAND2x1_ASAP7_75t_R _24191_ (.A(_01457_),
    .B(_01464_),
    .Y(_01470_));
 AOI21x1_ASAP7_75t_R _24192_ (.A1(_01469_),
    .A2(_01470_),
    .B(_11370_),
    .Y(_01471_));
 INVx1_ASAP7_75t_R _24193_ (.A(_07973_),
    .Y(_01472_));
 OAI21x1_ASAP7_75t_R _24194_ (.A1(_01468_),
    .A2(_01471_),
    .B(_01472_),
    .Y(_01473_));
 NAND2x2_ASAP7_75t_R _24195_ (.A(_01473_),
    .B(_01467_),
    .Y(_01474_));
 BUFx12f_ASAP7_75t_R _24196_ (.A(_01474_),
    .Y(_15923_));
 NOR2x1_ASAP7_75t_R _24197_ (.A(_10742_),
    .B(_00560_),
    .Y(_01475_));
 INVx1_ASAP7_75t_R _24198_ (.A(_01475_),
    .Y(_01476_));
 NOR2x1_ASAP7_75t_R _24199_ (.A(net35),
    .B(net72),
    .Y(_01477_));
 AND2x2_ASAP7_75t_R _24200_ (.A(_00756_),
    .B(net72),
    .Y(_01478_));
 OAI21x1_ASAP7_75t_R _24201_ (.A1(_01477_),
    .A2(_01478_),
    .B(_12848_),
    .Y(_01479_));
 XOR2x1_ASAP7_75t_R _24202_ (.A(net658),
    .Y(_01480_),
    .B(_12850_));
 NAND2x1_ASAP7_75t_R _24203_ (.A(_12849_),
    .B(_01480_),
    .Y(_01481_));
 AOI21x1_ASAP7_75t_R _24204_ (.A1(_01479_),
    .A2(_01481_),
    .B(_01458_),
    .Y(_01482_));
 XOR2x1_ASAP7_75t_R _24205_ (.A(_12850_),
    .Y(_01483_),
    .B(net664));
 NAND2x1_ASAP7_75t_R _24206_ (.A(net35),
    .B(_01483_),
    .Y(_01484_));
 INVx1_ASAP7_75t_R _24207_ (.A(net35),
    .Y(_01485_));
 XNOR2x1_ASAP7_75t_R _24208_ (.B(net664),
    .Y(_01486_),
    .A(_12850_));
 NAND2x1_ASAP7_75t_R _24209_ (.A(_01485_),
    .B(_01486_),
    .Y(_01487_));
 AOI21x1_ASAP7_75t_R _24210_ (.A1(_01484_),
    .A2(_01487_),
    .B(net907),
    .Y(_01488_));
 OAI21x1_ASAP7_75t_R _24211_ (.A1(_01482_),
    .A2(_01488_),
    .B(_10621_),
    .Y(_01489_));
 NAND2x2_ASAP7_75t_R _24212_ (.A(_01476_),
    .B(_01489_),
    .Y(_01490_));
 XNOR2x2_ASAP7_75t_R _24213_ (.A(_01098_),
    .B(_01490_),
    .Y(_01491_));
 BUFx12f_ASAP7_75t_R _24214_ (.A(_01491_),
    .Y(_15925_));
 NOR2x2_ASAP7_75t_R _24215_ (.A(net667),
    .B(_00562_),
    .Y(_01492_));
 INVx4_ASAP7_75t_R _24216_ (.A(_01492_),
    .Y(_01493_));
 NAND2x1_ASAP7_75t_R _24217_ (.A(_12879_),
    .B(_12880_),
    .Y(_01494_));
 INVx1_ASAP7_75t_R _24218_ (.A(_12879_),
    .Y(_01495_));
 INVx3_ASAP7_75t_R _24219_ (.A(_12880_),
    .Y(_01496_));
 NAND2x1_ASAP7_75t_R _24220_ (.A(_01495_),
    .B(_01496_),
    .Y(_01497_));
 INVx2_ASAP7_75t_R _24221_ (.A(_12910_),
    .Y(_01498_));
 AOI21x1_ASAP7_75t_R _24222_ (.A1(_01494_),
    .A2(_01497_),
    .B(_01498_),
    .Y(_01499_));
 NOR2x2_ASAP7_75t_R _24223_ (.A(_12910_),
    .B(_12875_),
    .Y(_01500_));
 OAI21x1_ASAP7_75t_R _24224_ (.A1(_01499_),
    .A2(_01500_),
    .B(net642),
    .Y(_01501_));
 INVx1_ASAP7_75t_R _24225_ (.A(_01501_),
    .Y(_01502_));
 NOR3x1_ASAP7_75t_R _24226_ (.A(_01500_),
    .B(net643),
    .C(_01499_),
    .Y(_01503_));
 OAI21x1_ASAP7_75t_R _24227_ (.A1(_01502_),
    .A2(_01503_),
    .B(_10668_),
    .Y(_01504_));
 INVx2_ASAP7_75t_R _24228_ (.A(_08008_),
    .Y(_01505_));
 AOI21x1_ASAP7_75t_R _24229_ (.A1(_01504_),
    .A2(_01493_),
    .B(_01505_),
    .Y(_01506_));
 NAND2x1_ASAP7_75t_R _24230_ (.A(_00562_),
    .B(_11373_),
    .Y(_01507_));
 NAND2x2_ASAP7_75t_R _24231_ (.A(_01498_),
    .B(_12881_),
    .Y(_01508_));
 INVx1_ASAP7_75t_R _24232_ (.A(net644),
    .Y(_01509_));
 NOR2x1_ASAP7_75t_R _24233_ (.A(_12879_),
    .B(_12880_),
    .Y(_01510_));
 AND2x2_ASAP7_75t_R _24234_ (.A(_12879_),
    .B(_12880_),
    .Y(_01511_));
 OAI21x1_ASAP7_75t_R _24235_ (.A1(_01510_),
    .A2(_01511_),
    .B(_12910_),
    .Y(_01512_));
 NAND3x2_ASAP7_75t_R _24236_ (.B(_01509_),
    .C(_01512_),
    .Y(_01513_),
    .A(_01508_));
 NAND3x2_ASAP7_75t_R _24237_ (.B(net650),
    .C(_01501_),
    .Y(_01514_),
    .A(_01513_));
 AOI21x1_ASAP7_75t_R _24238_ (.A1(_01507_),
    .A2(_01514_),
    .B(_08008_),
    .Y(_01515_));
 NOR2x2_ASAP7_75t_R _24239_ (.A(_01506_),
    .B(_01515_),
    .Y(_01516_));
 BUFx12f_ASAP7_75t_R _24240_ (.A(_01516_),
    .Y(_01517_));
 BUFx10_ASAP7_75t_R _24241_ (.A(_01517_),
    .Y(_15933_));
 XOR2x2_ASAP7_75t_R _24242_ (.A(_01490_),
    .B(_01098_),
    .Y(_01518_));
 BUFx6f_ASAP7_75t_R _24243_ (.A(_01518_),
    .Y(_15920_));
 AOI21x1_ASAP7_75t_R _24244_ (.A1(_01493_),
    .A2(_01504_),
    .B(_08008_),
    .Y(_01519_));
 AOI21x1_ASAP7_75t_R _24245_ (.A1(_01507_),
    .A2(_01514_),
    .B(_01505_),
    .Y(_01520_));
 NOR2x2_ASAP7_75t_R _24246_ (.A(_01520_),
    .B(_01519_),
    .Y(_01521_));
 BUFx10_ASAP7_75t_R _24247_ (.A(_01521_),
    .Y(_15930_));
 NAND3x2_ASAP7_75t_R _24248_ (.B(_01505_),
    .C(_01493_),
    .Y(_01522_),
    .A(_01504_));
 AOI21x1_ASAP7_75t_R _24249_ (.A1(_01501_),
    .A2(_01513_),
    .B(_12161_),
    .Y(_01523_));
 OAI21x1_ASAP7_75t_R _24250_ (.A1(_01492_),
    .A2(_01523_),
    .B(_08008_),
    .Y(_01524_));
 AO21x2_ASAP7_75t_R _24251_ (.A1(_01522_),
    .A2(_01524_),
    .B(_00564_),
    .Y(_01525_));
 OAI21x1_ASAP7_75t_R _24252_ (.A1(_01519_),
    .A2(_01520_),
    .B(_00563_),
    .Y(_01526_));
 NOR2x2_ASAP7_75t_R _24253_ (.A(net651),
    .B(_00700_),
    .Y(_01527_));
 XOR2x1_ASAP7_75t_R _24254_ (.A(_12915_),
    .Y(_01528_),
    .B(_00759_));
 XOR2x2_ASAP7_75t_R _24255_ (.A(_12879_),
    .B(net908),
    .Y(_01529_));
 XOR2x1_ASAP7_75t_R _24256_ (.A(_12919_),
    .Y(_01530_),
    .B(_01529_));
 NAND2x1_ASAP7_75t_R _24257_ (.A(_01528_),
    .B(_01530_),
    .Y(_01531_));
 NOR2x1_ASAP7_75t_R _24258_ (.A(_01528_),
    .B(_01530_),
    .Y(_01532_));
 INVx1_ASAP7_75t_R _24259_ (.A(_01532_),
    .Y(_01533_));
 AOI21x1_ASAP7_75t_R _24260_ (.A1(_01531_),
    .A2(_01533_),
    .B(_12092_),
    .Y(_01534_));
 INVx2_ASAP7_75t_R _24261_ (.A(_07945_),
    .Y(_01535_));
 OAI21x1_ASAP7_75t_R _24262_ (.A1(_01527_),
    .A2(_01534_),
    .B(_01535_),
    .Y(_01536_));
 INVx1_ASAP7_75t_R _24263_ (.A(_00759_),
    .Y(_01537_));
 XOR2x1_ASAP7_75t_R _24264_ (.A(_12915_),
    .Y(_01538_),
    .B(_01537_));
 XOR2x1_ASAP7_75t_R _24265_ (.A(_12914_),
    .Y(_01539_),
    .B(_01529_));
 NOR2x1_ASAP7_75t_R _24266_ (.A(_01538_),
    .B(_01539_),
    .Y(_01540_));
 OAI21x1_ASAP7_75t_R _24267_ (.A1(_01540_),
    .A2(_01532_),
    .B(_10761_),
    .Y(_01541_));
 INVx2_ASAP7_75t_R _24268_ (.A(_01527_),
    .Y(_01542_));
 NAND3x2_ASAP7_75t_R _24269_ (.B(_07945_),
    .C(_01542_),
    .Y(_01543_),
    .A(_01541_));
 NAND2x2_ASAP7_75t_R _24270_ (.A(_01536_),
    .B(_01543_),
    .Y(_01544_));
 BUFx6f_ASAP7_75t_R _24271_ (.A(_01544_),
    .Y(_01545_));
 AO21x1_ASAP7_75t_R _24272_ (.A1(_01525_),
    .A2(_01526_),
    .B(_01545_),
    .Y(_01546_));
 NAND3x2_ASAP7_75t_R _24273_ (.B(_08008_),
    .C(_01493_),
    .Y(_01547_),
    .A(_01504_));
 INVx2_ASAP7_75t_R _24274_ (.A(_01519_),
    .Y(_01548_));
 INVx1_ASAP7_75t_R _24275_ (.A(_00561_),
    .Y(_01549_));
 AO21x2_ASAP7_75t_R _24276_ (.A1(_01547_),
    .A2(_01548_),
    .B(_01549_),
    .Y(_01550_));
 OAI21x1_ASAP7_75t_R _24277_ (.A1(net887),
    .A2(_01515_),
    .B(_00563_),
    .Y(_01551_));
 OAI21x1_ASAP7_75t_R _24278_ (.A1(_01527_),
    .A2(_01534_),
    .B(_07945_),
    .Y(_01552_));
 NAND3x2_ASAP7_75t_R _24279_ (.B(_01535_),
    .C(_01542_),
    .Y(_01553_),
    .A(_01541_));
 NAND2x2_ASAP7_75t_R _24280_ (.A(_01552_),
    .B(_01553_),
    .Y(_01554_));
 BUFx6f_ASAP7_75t_R _24281_ (.A(_01554_),
    .Y(_01555_));
 AO21x1_ASAP7_75t_R _24282_ (.A1(_01550_),
    .A2(_01551_),
    .B(_01555_),
    .Y(_01556_));
 INVx1_ASAP7_75t_R _24283_ (.A(_00699_),
    .Y(_01557_));
 NOR2x1_ASAP7_75t_R _24284_ (.A(_10743_),
    .B(_01557_),
    .Y(_01558_));
 XOR2x2_ASAP7_75t_R _24285_ (.A(_12913_),
    .B(net908),
    .Y(_01559_));
 INVx1_ASAP7_75t_R _24286_ (.A(_00856_),
    .Y(_01560_));
 XOR2x2_ASAP7_75t_R _24287_ (.A(_01559_),
    .B(_01560_),
    .Y(_01561_));
 XOR2x2_ASAP7_75t_R _24288_ (.A(_12952_),
    .B(_00824_),
    .Y(_01562_));
 XOR2x1_ASAP7_75t_R _24289_ (.A(_12930_),
    .Y(_01563_),
    .B(_01562_));
 NAND2x1_ASAP7_75t_R _24290_ (.A(_01561_),
    .B(_01563_),
    .Y(_01564_));
 XOR2x2_ASAP7_75t_R _24291_ (.A(_01559_),
    .B(_00856_),
    .Y(_01565_));
 XNOR2x1_ASAP7_75t_R _24292_ (.B(_01562_),
    .Y(_01566_),
    .A(_12930_));
 NAND2x1_ASAP7_75t_R _24293_ (.A(_01565_),
    .B(_01566_),
    .Y(_01567_));
 AOI21x1_ASAP7_75t_R _24294_ (.A1(_01564_),
    .A2(_01567_),
    .B(_11370_),
    .Y(_01568_));
 OAI21x1_ASAP7_75t_R _24295_ (.A1(_01558_),
    .A2(_01568_),
    .B(_07996_),
    .Y(_01569_));
 NOR2x1_ASAP7_75t_R _24296_ (.A(_10743_),
    .B(_00699_),
    .Y(_01570_));
 XOR2x1_ASAP7_75t_R _24297_ (.A(_12930_),
    .Y(_01571_),
    .B(_12952_));
 XOR2x2_ASAP7_75t_R _24298_ (.A(_12931_),
    .B(_01559_),
    .Y(_01572_));
 NAND2x1_ASAP7_75t_R _24299_ (.A(_01571_),
    .B(_01572_),
    .Y(_01573_));
 XNOR2x1_ASAP7_75t_R _24300_ (.B(_12930_),
    .Y(_01574_),
    .A(_12952_));
 INVx1_ASAP7_75t_R _24301_ (.A(_01572_),
    .Y(_01575_));
 NAND2x1_ASAP7_75t_R _24302_ (.A(_01574_),
    .B(_01575_),
    .Y(_01576_));
 AOI21x1_ASAP7_75t_R _24303_ (.A1(_01573_),
    .A2(_01576_),
    .B(_11370_),
    .Y(_01577_));
 INVx1_ASAP7_75t_R _24304_ (.A(_07996_),
    .Y(_01578_));
 OAI21x1_ASAP7_75t_R _24305_ (.A1(_01570_),
    .A2(_01577_),
    .B(_01578_),
    .Y(_01579_));
 NAND2x2_ASAP7_75t_R _24306_ (.A(_01569_),
    .B(_01579_),
    .Y(_01580_));
 CKINVDCx6p67_ASAP7_75t_R _24307_ (.A(_01580_),
    .Y(_01581_));
 BUFx6f_ASAP7_75t_R _24308_ (.A(_01581_),
    .Y(_01582_));
 AO21x1_ASAP7_75t_R _24309_ (.A1(_01546_),
    .A2(_01556_),
    .B(_01582_),
    .Y(_01583_));
 NAND2x2_ASAP7_75t_R _24310_ (.A(_01517_),
    .B(net571),
    .Y(_01584_));
 AO21x1_ASAP7_75t_R _24311_ (.A1(_01584_),
    .A2(_01525_),
    .B(_01555_),
    .Y(_01585_));
 BUFx6f_ASAP7_75t_R _24312_ (.A(_01554_),
    .Y(_01586_));
 OAI21x1_ASAP7_75t_R _24313_ (.A1(_01519_),
    .A2(_01520_),
    .B(net504),
    .Y(_01587_));
 INVx4_ASAP7_75t_R _24314_ (.A(_01587_),
    .Y(_01588_));
 NAND2x2_ASAP7_75t_R _24315_ (.A(_01586_),
    .B(_01588_),
    .Y(_01589_));
 BUFx6f_ASAP7_75t_R _24316_ (.A(_01580_),
    .Y(_01590_));
 BUFx6f_ASAP7_75t_R _24317_ (.A(_01590_),
    .Y(_01591_));
 AO21x1_ASAP7_75t_R _24318_ (.A1(_01585_),
    .A2(_01589_),
    .B(_01591_),
    .Y(_01592_));
 NOR2x2_ASAP7_75t_R _24319_ (.A(net585),
    .B(_00698_),
    .Y(_01593_));
 INVx1_ASAP7_75t_R _24320_ (.A(_01593_),
    .Y(_01594_));
 XNOR2x1_ASAP7_75t_R _24321_ (.B(_00792_),
    .Y(_01595_),
    .A(_12902_));
 XOR2x2_ASAP7_75t_R _24322_ (.A(_00824_),
    .B(_00825_),
    .Y(_01596_));
 XOR2x1_ASAP7_75t_R _24323_ (.A(_01596_),
    .Y(_01597_),
    .B(_12956_));
 NAND2x1_ASAP7_75t_R _24324_ (.A(_01595_),
    .B(_01597_),
    .Y(_01598_));
 INVx1_ASAP7_75t_R _24325_ (.A(_01595_),
    .Y(_01599_));
 XOR2x1_ASAP7_75t_R _24326_ (.A(_01596_),
    .Y(_01600_),
    .B(_12955_));
 NAND2x1_ASAP7_75t_R _24327_ (.A(_01599_),
    .B(_01600_),
    .Y(_01601_));
 AOI21x1_ASAP7_75t_R _24328_ (.A1(_01598_),
    .A2(_01601_),
    .B(_11374_),
    .Y(_01602_));
 INVx1_ASAP7_75t_R _24329_ (.A(_01602_),
    .Y(_01603_));
 INVx1_ASAP7_75t_R _24330_ (.A(_01104_),
    .Y(_01604_));
 AOI21x1_ASAP7_75t_R _24331_ (.A1(_01594_),
    .A2(_01603_),
    .B(_01604_),
    .Y(_01605_));
 NOR3x2_ASAP7_75t_R _24332_ (.B(_01104_),
    .C(_01593_),
    .Y(_01606_),
    .A(_01602_));
 NOR2x2_ASAP7_75t_R _24333_ (.A(_01605_),
    .B(_01606_),
    .Y(_01607_));
 CKINVDCx5p33_ASAP7_75t_R _24334_ (.A(_01607_),
    .Y(_01608_));
 BUFx10_ASAP7_75t_R _24335_ (.A(_01608_),
    .Y(_01609_));
 AOI21x1_ASAP7_75t_R _24336_ (.A1(_01583_),
    .A2(_01592_),
    .B(_01609_),
    .Y(_01610_));
 BUFx6f_ASAP7_75t_R _24337_ (.A(_01580_),
    .Y(_01611_));
 OAI21x1_ASAP7_75t_R _24338_ (.A1(net887),
    .A2(_01515_),
    .B(_00561_),
    .Y(_01612_));
 BUFx6f_ASAP7_75t_R _24339_ (.A(_01544_),
    .Y(_01613_));
 AO21x1_ASAP7_75t_R _24340_ (.A1(_01526_),
    .A2(_01612_),
    .B(_01613_),
    .Y(_01614_));
 NAND2x1_ASAP7_75t_R _24341_ (.A(_01611_),
    .B(_01614_),
    .Y(_01615_));
 BUFx12_ASAP7_75t_R _24342_ (.A(_01521_),
    .Y(_01616_));
 AOI21x1_ASAP7_75t_R _24343_ (.A1(_15925_),
    .A2(_15923_),
    .B(_01616_),
    .Y(_01617_));
 INVx1_ASAP7_75t_R _24344_ (.A(_00564_),
    .Y(_01618_));
 OA21x2_ASAP7_75t_R _24345_ (.A1(_01515_),
    .A2(net887),
    .B(_01618_),
    .Y(_01619_));
 BUFx4f_ASAP7_75t_R _24346_ (.A(_01619_),
    .Y(_01620_));
 BUFx6f_ASAP7_75t_R _24347_ (.A(_01544_),
    .Y(_01621_));
 OA21x2_ASAP7_75t_R _24348_ (.A1(_01617_),
    .A2(_01620_),
    .B(_01621_),
    .Y(_01622_));
 OAI21x1_ASAP7_75t_R _24349_ (.A1(_01615_),
    .A2(_01622_),
    .B(_01609_),
    .Y(_01623_));
 NOR2x2_ASAP7_75t_R _24350_ (.A(_15925_),
    .B(_15923_),
    .Y(_01624_));
 BUFx10_ASAP7_75t_R _24351_ (.A(_01544_),
    .Y(_01625_));
 NAND2x2_ASAP7_75t_R _24352_ (.A(_01491_),
    .B(net885),
    .Y(_01626_));
 NAND2x2_ASAP7_75t_R _24353_ (.A(_01625_),
    .B(_01626_),
    .Y(_01627_));
 NOR2x2_ASAP7_75t_R _24354_ (.A(_01624_),
    .B(_01627_),
    .Y(_01628_));
 OAI21x1_ASAP7_75t_R _24355_ (.A1(_01455_),
    .A2(_01466_),
    .B(_01472_),
    .Y(_01629_));
 OAI21x1_ASAP7_75t_R _24356_ (.A1(_01468_),
    .A2(_01471_),
    .B(_07973_),
    .Y(_01630_));
 NAND2x2_ASAP7_75t_R _24357_ (.A(_01630_),
    .B(_01629_),
    .Y(_01631_));
 BUFx6f_ASAP7_75t_R _24358_ (.A(_01631_),
    .Y(_15921_));
 NAND2x1_ASAP7_75t_R _24359_ (.A(net536),
    .B(net70),
    .Y(_01632_));
 NAND2x1_ASAP7_75t_R _24360_ (.A(_01626_),
    .B(_01632_),
    .Y(_01633_));
 BUFx6f_ASAP7_75t_R _24361_ (.A(_01554_),
    .Y(_01634_));
 BUFx6f_ASAP7_75t_R _24362_ (.A(_01580_),
    .Y(_01635_));
 AO21x1_ASAP7_75t_R _24363_ (.A1(_01633_),
    .A2(_01634_),
    .B(_01635_),
    .Y(_01636_));
 NOR2x1_ASAP7_75t_R _24364_ (.A(_01628_),
    .B(_01636_),
    .Y(_01637_));
 XOR2x2_ASAP7_75t_R _24365_ (.A(_00826_),
    .B(_00858_),
    .Y(_01638_));
 XOR2x1_ASAP7_75t_R _24366_ (.A(_12954_),
    .Y(_01639_),
    .B(_00762_));
 XNOR2x1_ASAP7_75t_R _24367_ (.B(_01639_),
    .Y(_01640_),
    .A(_01638_));
 NOR2x1_ASAP7_75t_R _24368_ (.A(_10787_),
    .B(_00697_),
    .Y(_01641_));
 AO21x1_ASAP7_75t_R _24369_ (.A1(_01640_),
    .A2(_11451_),
    .B(_01641_),
    .Y(_01642_));
 XOR2x2_ASAP7_75t_R _24370_ (.A(_01642_),
    .B(_01105_),
    .Y(_01643_));
 BUFx10_ASAP7_75t_R _24371_ (.A(_01643_),
    .Y(_01644_));
 OAI21x1_ASAP7_75t_R _24372_ (.A1(_01623_),
    .A2(_01637_),
    .B(_01644_),
    .Y(_01645_));
 NOR2x1_ASAP7_75t_R _24373_ (.A(_01610_),
    .B(_01645_),
    .Y(_01646_));
 BUFx10_ASAP7_75t_R _24374_ (.A(_01554_),
    .Y(_01647_));
 NAND2x2_ASAP7_75t_R _24375_ (.A(net535),
    .B(_01516_),
    .Y(_01648_));
 NAND2x2_ASAP7_75t_R _24376_ (.A(_01647_),
    .B(_01648_),
    .Y(_01649_));
 NAND2x2_ASAP7_75t_R _24377_ (.A(_01491_),
    .B(net571),
    .Y(_01650_));
 NOR2x2_ASAP7_75t_R _24378_ (.A(_01517_),
    .B(_01650_),
    .Y(_01651_));
 NOR2x1_ASAP7_75t_R _24379_ (.A(_01649_),
    .B(_01651_),
    .Y(_01652_));
 BUFx10_ASAP7_75t_R _24380_ (.A(_01544_),
    .Y(_01653_));
 NAND2x2_ASAP7_75t_R _24381_ (.A(_01516_),
    .B(net876),
    .Y(_01654_));
 INVx1_ASAP7_75t_R _24382_ (.A(_01654_),
    .Y(_01655_));
 INVx2_ASAP7_75t_R _24383_ (.A(_01207_),
    .Y(_01656_));
 OAI21x1_ASAP7_75t_R _24384_ (.A1(net887),
    .A2(_01515_),
    .B(_01656_),
    .Y(_01657_));
 OAI21x1_ASAP7_75t_R _24385_ (.A1(_01657_),
    .A2(_01586_),
    .B(_01590_),
    .Y(_01658_));
 AO21x1_ASAP7_75t_R _24386_ (.A1(_01653_),
    .A2(_01655_),
    .B(_01658_),
    .Y(_01659_));
 NOR2x1_ASAP7_75t_R _24387_ (.A(_01652_),
    .B(_01659_),
    .Y(_01660_));
 INVx3_ASAP7_75t_R _24388_ (.A(_01210_),
    .Y(_01661_));
 AO21x2_ASAP7_75t_R _24389_ (.A1(_01522_),
    .A2(_01524_),
    .B(_01661_),
    .Y(_01662_));
 BUFx6f_ASAP7_75t_R _24390_ (.A(_01544_),
    .Y(_01663_));
 NOR2x2_ASAP7_75t_R _24391_ (.A(_01491_),
    .B(net886),
    .Y(_01664_));
 NOR2x1_ASAP7_75t_R _24392_ (.A(_01663_),
    .B(_01664_),
    .Y(_01665_));
 AOI21x1_ASAP7_75t_R _24393_ (.A1(_01662_),
    .A2(_01665_),
    .B(_01611_),
    .Y(_01666_));
 OAI21x1_ASAP7_75t_R _24394_ (.A1(_15925_),
    .A2(net70),
    .B(_15933_),
    .Y(_01667_));
 NAND2x2_ASAP7_75t_R _24395_ (.A(_01521_),
    .B(net573),
    .Y(_01668_));
 BUFx6f_ASAP7_75t_R _24396_ (.A(_01554_),
    .Y(_01669_));
 AO21x1_ASAP7_75t_R _24397_ (.A1(_01667_),
    .A2(_01668_),
    .B(_01669_),
    .Y(_01670_));
 BUFx6f_ASAP7_75t_R _24398_ (.A(_01608_),
    .Y(_01671_));
 AO21x1_ASAP7_75t_R _24399_ (.A1(_01666_),
    .A2(_01670_),
    .B(_01671_),
    .Y(_01672_));
 NOR2x1_ASAP7_75t_R _24400_ (.A(_01660_),
    .B(_01672_),
    .Y(_01673_));
 OAI21x1_ASAP7_75t_R _24401_ (.A1(_01606_),
    .A2(_01605_),
    .B(_01580_),
    .Y(_01674_));
 AOI21x1_ASAP7_75t_R _24402_ (.A1(_01208_),
    .A2(_01616_),
    .B(_01544_),
    .Y(_01675_));
 NAND3x2_ASAP7_75t_R _24403_ (.B(_01517_),
    .C(net71),
    .Y(_01676_),
    .A(_15923_));
 NOR2x2_ASAP7_75t_R _24404_ (.A(_01586_),
    .B(_01664_),
    .Y(_01677_));
 AOI21x1_ASAP7_75t_R _24405_ (.A1(_01675_),
    .A2(_01676_),
    .B(_01677_),
    .Y(_01678_));
 INVx1_ASAP7_75t_R _24406_ (.A(_01570_),
    .Y(_01679_));
 NOR2x1_ASAP7_75t_R _24407_ (.A(_01571_),
    .B(_01572_),
    .Y(_01680_));
 INVx1_ASAP7_75t_R _24408_ (.A(_01573_),
    .Y(_01681_));
 OAI21x1_ASAP7_75t_R _24409_ (.A1(_01680_),
    .A2(_01681_),
    .B(_13017_),
    .Y(_01682_));
 AOI21x1_ASAP7_75t_R _24410_ (.A1(_01679_),
    .A2(_01682_),
    .B(_01578_),
    .Y(_01683_));
 INVx1_ASAP7_75t_R _24411_ (.A(_01558_),
    .Y(_01684_));
 NOR2x1_ASAP7_75t_R _24412_ (.A(_01565_),
    .B(_01566_),
    .Y(_01685_));
 INVx1_ASAP7_75t_R _24413_ (.A(_01567_),
    .Y(_01686_));
 OAI21x1_ASAP7_75t_R _24414_ (.A1(_01685_),
    .A2(_01686_),
    .B(_13017_),
    .Y(_01687_));
 AOI21x1_ASAP7_75t_R _24415_ (.A1(_01684_),
    .A2(_01687_),
    .B(_07996_),
    .Y(_01688_));
 OAI22x1_ASAP7_75t_R _24416_ (.A1(_01606_),
    .A2(_01605_),
    .B1(_01683_),
    .B2(_01688_),
    .Y(_01689_));
 INVx4_ASAP7_75t_R _24417_ (.A(_01689_),
    .Y(_01690_));
 NOR2x2_ASAP7_75t_R _24418_ (.A(_01491_),
    .B(_01516_),
    .Y(_01691_));
 OAI21x1_ASAP7_75t_R _24419_ (.A1(net70),
    .A2(_01648_),
    .B(_01545_),
    .Y(_01692_));
 AO21x1_ASAP7_75t_R _24420_ (.A1(_01522_),
    .A2(_01524_),
    .B(_01618_),
    .Y(_01693_));
 BUFx4f_ASAP7_75t_R _24421_ (.A(_01693_),
    .Y(_01694_));
 AOI21x1_ASAP7_75t_R _24422_ (.A1(_01548_),
    .A2(_01547_),
    .B(_01661_),
    .Y(_01695_));
 NOR2x1_ASAP7_75t_R _24423_ (.A(_01625_),
    .B(_01695_),
    .Y(_01696_));
 NAND2x1_ASAP7_75t_R _24424_ (.A(_01694_),
    .B(_01696_),
    .Y(_01697_));
 OAI21x1_ASAP7_75t_R _24425_ (.A1(_01691_),
    .A2(_01692_),
    .B(_01697_),
    .Y(_01698_));
 AOI21x1_ASAP7_75t_R _24426_ (.A1(_01690_),
    .A2(_01698_),
    .B(_01644_),
    .Y(_01699_));
 OAI21x1_ASAP7_75t_R _24427_ (.A1(_01674_),
    .A2(_01678_),
    .B(_01699_),
    .Y(_01700_));
 XOR2x1_ASAP7_75t_R _24428_ (.A(_13013_),
    .Y(_01701_),
    .B(_00826_));
 INVx1_ASAP7_75t_R _24429_ (.A(_13011_),
    .Y(_01702_));
 XOR2x1_ASAP7_75t_R _24430_ (.A(_01701_),
    .Y(_01703_),
    .B(_01702_));
 XOR2x1_ASAP7_75t_R _24431_ (.A(net647),
    .Y(_01704_),
    .B(_00794_));
 XOR2x1_ASAP7_75t_R _24432_ (.A(_01703_),
    .Y(_01705_),
    .B(_01704_));
 NAND2x1_ASAP7_75t_R _24433_ (.A(_11451_),
    .B(_01705_),
    .Y(_01706_));
 OA21x2_ASAP7_75t_R _24434_ (.A1(_13017_),
    .A2(_00696_),
    .B(_01706_),
    .Y(_01707_));
 XOR2x2_ASAP7_75t_R _24435_ (.A(_01707_),
    .B(_01106_),
    .Y(_01708_));
 INVx4_ASAP7_75t_R _24436_ (.A(_01708_),
    .Y(_01709_));
 BUFx10_ASAP7_75t_R _24437_ (.A(_01709_),
    .Y(_01710_));
 OAI21x1_ASAP7_75t_R _24438_ (.A1(_01673_),
    .A2(_01700_),
    .B(_01710_),
    .Y(_01711_));
 OAI21x1_ASAP7_75t_R _24439_ (.A1(_15923_),
    .A2(_15933_),
    .B(_01587_),
    .Y(_01712_));
 NAND2x1_ASAP7_75t_R _24440_ (.A(_01545_),
    .B(_01712_),
    .Y(_01713_));
 AO21x1_ASAP7_75t_R _24441_ (.A1(_01626_),
    .A2(_01550_),
    .B(_01663_),
    .Y(_01714_));
 AOI21x1_ASAP7_75t_R _24442_ (.A1(_01713_),
    .A2(_01714_),
    .B(_01674_),
    .Y(_01715_));
 INVx6_ASAP7_75t_R _24443_ (.A(_01643_),
    .Y(_01716_));
 AOI21x1_ASAP7_75t_R _24444_ (.A1(_01657_),
    .A2(_01526_),
    .B(_01647_),
    .Y(_01717_));
 OAI21x1_ASAP7_75t_R _24445_ (.A1(_01675_),
    .A2(_01717_),
    .B(_01690_),
    .Y(_01718_));
 NAND2x1_ASAP7_75t_R _24446_ (.A(_01716_),
    .B(_01718_),
    .Y(_01719_));
 NOR2x1_ASAP7_75t_R _24447_ (.A(_01715_),
    .B(_01719_),
    .Y(_01720_));
 INVx2_ASAP7_75t_R _24448_ (.A(_01208_),
    .Y(_01721_));
 OA21x2_ASAP7_75t_R _24449_ (.A1(_01520_),
    .A2(_01519_),
    .B(_01721_),
    .Y(_01722_));
 BUFx6f_ASAP7_75t_R _24450_ (.A(_01722_),
    .Y(_01723_));
 AOI21x1_ASAP7_75t_R _24451_ (.A1(_01613_),
    .A2(_01723_),
    .B(_01581_),
    .Y(_01724_));
 OAI21x1_ASAP7_75t_R _24452_ (.A1(_01649_),
    .A2(_01651_),
    .B(_01724_),
    .Y(_01725_));
 AOI21x1_ASAP7_75t_R _24453_ (.A1(_01613_),
    .A2(_01722_),
    .B(_01590_),
    .Y(_01726_));
 INVx1_ASAP7_75t_R _24454_ (.A(_01209_),
    .Y(_01727_));
 OAI21x1_ASAP7_75t_R _24455_ (.A1(net887),
    .A2(_01515_),
    .B(_01727_),
    .Y(_01728_));
 NOR2x1_ASAP7_75t_R _24456_ (.A(_01728_),
    .B(_01647_),
    .Y(_01729_));
 OA21x2_ASAP7_75t_R _24457_ (.A1(_01515_),
    .A2(net887),
    .B(net503),
    .Y(_01730_));
 BUFx6f_ASAP7_75t_R _24458_ (.A(_01730_),
    .Y(_01731_));
 NOR2x2_ASAP7_75t_R _24459_ (.A(_01544_),
    .B(_01731_),
    .Y(_01732_));
 NOR2x1_ASAP7_75t_R _24460_ (.A(_01729_),
    .B(_01732_),
    .Y(_01733_));
 BUFx6f_ASAP7_75t_R _24461_ (.A(_01608_),
    .Y(_01734_));
 AOI21x1_ASAP7_75t_R _24462_ (.A1(_01726_),
    .A2(_01733_),
    .B(_01734_),
    .Y(_01735_));
 NAND2x1_ASAP7_75t_R _24463_ (.A(_01725_),
    .B(_01735_),
    .Y(_01736_));
 AOI21x1_ASAP7_75t_R _24464_ (.A1(_01720_),
    .A2(_01736_),
    .B(_01709_),
    .Y(_01737_));
 AOI21x1_ASAP7_75t_R _24465_ (.A1(net534),
    .A2(net573),
    .B(_01517_),
    .Y(_01738_));
 OAI21x1_ASAP7_75t_R _24466_ (.A1(_01723_),
    .A2(_01738_),
    .B(_01545_),
    .Y(_01739_));
 INVx2_ASAP7_75t_R _24467_ (.A(_01739_),
    .Y(_01740_));
 OAI21x1_ASAP7_75t_R _24468_ (.A1(_01519_),
    .A2(_01520_),
    .B(_01656_),
    .Y(_01741_));
 OA21x2_ASAP7_75t_R _24469_ (.A1(_01647_),
    .A2(_01741_),
    .B(_01590_),
    .Y(_01742_));
 OAI21x1_ASAP7_75t_R _24470_ (.A1(net71),
    .A2(_15930_),
    .B(_01551_),
    .Y(_01743_));
 NAND2x1_ASAP7_75t_R _24471_ (.A(_01555_),
    .B(_01743_),
    .Y(_01744_));
 NAND2x1_ASAP7_75t_R _24472_ (.A(_01742_),
    .B(_01744_),
    .Y(_01745_));
 OAI21x1_ASAP7_75t_R _24473_ (.A1(_01519_),
    .A2(_01520_),
    .B(_01618_),
    .Y(_01746_));
 INVx1_ASAP7_75t_R _24474_ (.A(_01746_),
    .Y(_01747_));
 AO21x1_ASAP7_75t_R _24475_ (.A1(_01747_),
    .A2(_01625_),
    .B(_01590_),
    .Y(_01748_));
 NOR2x1_ASAP7_75t_R _24476_ (.A(_01212_),
    .B(_01663_),
    .Y(_01749_));
 BUFx6f_ASAP7_75t_R _24477_ (.A(_01607_),
    .Y(_01750_));
 OA21x2_ASAP7_75t_R _24478_ (.A1(_01748_),
    .A2(_01749_),
    .B(_01750_),
    .Y(_01751_));
 OAI21x1_ASAP7_75t_R _24479_ (.A1(_01740_),
    .A2(_01745_),
    .B(_01751_),
    .Y(_01752_));
 NAND2x2_ASAP7_75t_R _24480_ (.A(net536),
    .B(net571),
    .Y(_01753_));
 NOR2x1_ASAP7_75t_R _24481_ (.A(_15933_),
    .B(_01753_),
    .Y(_01754_));
 AO21x1_ASAP7_75t_R _24482_ (.A1(_01547_),
    .A2(_01548_),
    .B(_00561_),
    .Y(_01755_));
 NAND2x2_ASAP7_75t_R _24483_ (.A(_01545_),
    .B(_01755_),
    .Y(_01756_));
 OA21x2_ASAP7_75t_R _24484_ (.A1(_01613_),
    .A2(_01657_),
    .B(_01581_),
    .Y(_01757_));
 OAI21x1_ASAP7_75t_R _24485_ (.A1(_01754_),
    .A2(_01756_),
    .B(_01757_),
    .Y(_01758_));
 INVx1_ASAP7_75t_R _24486_ (.A(_01658_),
    .Y(_01759_));
 AOI21x1_ASAP7_75t_R _24487_ (.A1(_01209_),
    .A2(_01517_),
    .B(_01625_),
    .Y(_01760_));
 AOI22x1_ASAP7_75t_R _24488_ (.A1(_01522_),
    .A2(_01524_),
    .B1(_01467_),
    .B2(_01473_),
    .Y(_01761_));
 NAND2x2_ASAP7_75t_R _24489_ (.A(_15920_),
    .B(_01761_),
    .Y(_01762_));
 NAND2x1_ASAP7_75t_R _24490_ (.A(_01760_),
    .B(_01762_),
    .Y(_01763_));
 BUFx10_ASAP7_75t_R _24491_ (.A(_01607_),
    .Y(_01764_));
 AOI21x1_ASAP7_75t_R _24492_ (.A1(_01759_),
    .A2(_01763_),
    .B(_01764_),
    .Y(_01765_));
 AOI21x1_ASAP7_75t_R _24493_ (.A1(_01758_),
    .A2(_01765_),
    .B(_01716_),
    .Y(_01766_));
 NAND2x1_ASAP7_75t_R _24494_ (.A(_01752_),
    .B(_01766_),
    .Y(_01767_));
 NAND2x1_ASAP7_75t_R _24495_ (.A(_01737_),
    .B(_01767_),
    .Y(_01768_));
 OAI21x1_ASAP7_75t_R _24496_ (.A1(_01646_),
    .A2(_01711_),
    .B(_01768_),
    .Y(_00088_));
 BUFx10_ASAP7_75t_R _24497_ (.A(_01716_),
    .Y(_01769_));
 BUFx10_ASAP7_75t_R _24498_ (.A(_01750_),
    .Y(_01770_));
 NOR2x2_ASAP7_75t_R _24499_ (.A(_01517_),
    .B(net574),
    .Y(_01771_));
 BUFx6f_ASAP7_75t_R _24500_ (.A(_01554_),
    .Y(_01772_));
 OAI21x1_ASAP7_75t_R _24501_ (.A1(_01661_),
    .A2(_15930_),
    .B(_01772_),
    .Y(_01773_));
 OAI21x1_ASAP7_75t_R _24502_ (.A1(_01771_),
    .A2(_01773_),
    .B(_01582_),
    .Y(_01774_));
 BUFx6f_ASAP7_75t_R _24503_ (.A(_01647_),
    .Y(_01775_));
 AOI21x1_ASAP7_75t_R _24504_ (.A1(_15925_),
    .A2(net573),
    .B(_01517_),
    .Y(_01776_));
 INVx1_ASAP7_75t_R _24505_ (.A(_01776_),
    .Y(_01777_));
 NOR2x1_ASAP7_75t_R _24506_ (.A(_01775_),
    .B(_01777_),
    .Y(_01778_));
 OAI21x1_ASAP7_75t_R _24507_ (.A1(net888),
    .A2(_01515_),
    .B(_01721_),
    .Y(_01779_));
 INVx2_ASAP7_75t_R _24508_ (.A(_01779_),
    .Y(_01780_));
 BUFx6f_ASAP7_75t_R _24509_ (.A(_01625_),
    .Y(_01781_));
 BUFx6f_ASAP7_75t_R _24510_ (.A(_01581_),
    .Y(_01782_));
 AO21x1_ASAP7_75t_R _24511_ (.A1(_01780_),
    .A2(_01781_),
    .B(_01782_),
    .Y(_01783_));
 OAI21x1_ASAP7_75t_R _24512_ (.A1(net71),
    .A2(net70),
    .B(_15933_),
    .Y(_01784_));
 AOI21x1_ASAP7_75t_R _24513_ (.A1(_01694_),
    .A2(_01784_),
    .B(_01781_),
    .Y(_01785_));
 OAI22x1_ASAP7_75t_R _24514_ (.A1(_01774_),
    .A2(_01778_),
    .B1(_01783_),
    .B2(_01785_),
    .Y(_01786_));
 OAI21x1_ASAP7_75t_R _24515_ (.A1(_01731_),
    .A2(_01723_),
    .B(_01634_),
    .Y(_01787_));
 INVx2_ASAP7_75t_R _24516_ (.A(_01551_),
    .Y(_01788_));
 NOR2x2_ASAP7_75t_R _24517_ (.A(net535),
    .B(net885),
    .Y(_01789_));
 OAI21x1_ASAP7_75t_R _24518_ (.A1(_01788_),
    .A2(_01789_),
    .B(_01621_),
    .Y(_01790_));
 BUFx10_ASAP7_75t_R _24519_ (.A(_01590_),
    .Y(_01791_));
 AOI21x1_ASAP7_75t_R _24520_ (.A1(_01787_),
    .A2(_01790_),
    .B(_01791_),
    .Y(_01792_));
 NOR2x2_ASAP7_75t_R _24521_ (.A(net534),
    .B(_01517_),
    .Y(_01793_));
 OAI21x1_ASAP7_75t_R _24522_ (.A1(_01588_),
    .A2(_01793_),
    .B(_01621_),
    .Y(_01794_));
 NOR2x2_ASAP7_75t_R _24523_ (.A(_15920_),
    .B(net70),
    .Y(_01795_));
 OAI21x1_ASAP7_75t_R _24524_ (.A1(_01691_),
    .A2(_01795_),
    .B(_01634_),
    .Y(_01796_));
 AOI21x1_ASAP7_75t_R _24525_ (.A1(_01794_),
    .A2(_01796_),
    .B(_01582_),
    .Y(_01797_));
 OAI21x1_ASAP7_75t_R _24526_ (.A1(_01792_),
    .A2(_01797_),
    .B(_01770_),
    .Y(_01798_));
 OAI21x1_ASAP7_75t_R _24527_ (.A1(_01770_),
    .A2(_01786_),
    .B(_01798_),
    .Y(_01799_));
 AO21x1_ASAP7_75t_R _24528_ (.A1(_01551_),
    .A2(_01746_),
    .B(_01663_),
    .Y(_01800_));
 INVx1_ASAP7_75t_R _24529_ (.A(_01657_),
    .Y(_01801_));
 BUFx6f_ASAP7_75t_R _24530_ (.A(_01625_),
    .Y(_01802_));
 OAI21x1_ASAP7_75t_R _24531_ (.A1(_01801_),
    .A2(_01789_),
    .B(_01802_),
    .Y(_01803_));
 AOI21x1_ASAP7_75t_R _24532_ (.A1(_01800_),
    .A2(_01803_),
    .B(_01791_),
    .Y(_01804_));
 INVx1_ASAP7_75t_R _24533_ (.A(_01526_),
    .Y(_01805_));
 OAI21x1_ASAP7_75t_R _24534_ (.A1(_01805_),
    .A2(_01691_),
    .B(_01802_),
    .Y(_01806_));
 NOR2x2_ASAP7_75t_R _24535_ (.A(_01616_),
    .B(net875),
    .Y(_01807_));
 OAI21x1_ASAP7_75t_R _24536_ (.A1(_01780_),
    .A2(_01807_),
    .B(_01669_),
    .Y(_01808_));
 AOI21x1_ASAP7_75t_R _24537_ (.A1(_01806_),
    .A2(_01808_),
    .B(_01582_),
    .Y(_01809_));
 OAI21x1_ASAP7_75t_R _24538_ (.A1(_01804_),
    .A2(_01809_),
    .B(_01609_),
    .Y(_01810_));
 BUFx6f_ASAP7_75t_R _24539_ (.A(_01554_),
    .Y(_01811_));
 OAI21x1_ASAP7_75t_R _24540_ (.A1(_01731_),
    .A2(_01617_),
    .B(_01811_),
    .Y(_01812_));
 OAI21x1_ASAP7_75t_R _24541_ (.A1(net889),
    .A2(_15933_),
    .B(_01741_),
    .Y(_01813_));
 AOI21x1_ASAP7_75t_R _24542_ (.A1(_01653_),
    .A2(_01813_),
    .B(_01635_),
    .Y(_01814_));
 NAND2x1_ASAP7_75t_R _24543_ (.A(_01812_),
    .B(_01814_),
    .Y(_01815_));
 BUFx6f_ASAP7_75t_R _24544_ (.A(_01581_),
    .Y(_01816_));
 AOI21x1_ASAP7_75t_R _24545_ (.A1(_01772_),
    .A2(_01694_),
    .B(_01816_),
    .Y(_01817_));
 OAI21x1_ASAP7_75t_R _24546_ (.A1(_01789_),
    .A2(_01776_),
    .B(_01621_),
    .Y(_01818_));
 AOI21x1_ASAP7_75t_R _24547_ (.A1(_01817_),
    .A2(_01818_),
    .B(_01734_),
    .Y(_01819_));
 AOI21x1_ASAP7_75t_R _24548_ (.A1(_01815_),
    .A2(_01819_),
    .B(_01708_),
    .Y(_01820_));
 NAND2x1_ASAP7_75t_R _24549_ (.A(_01810_),
    .B(_01820_),
    .Y(_01821_));
 OAI21x1_ASAP7_75t_R _24550_ (.A1(_01710_),
    .A2(_01799_),
    .B(_01821_),
    .Y(_01822_));
 OAI21x1_ASAP7_75t_R _24551_ (.A1(_01620_),
    .A2(_01789_),
    .B(_01555_),
    .Y(_01823_));
 OAI21x1_ASAP7_75t_R _24552_ (.A1(_01780_),
    .A2(_01664_),
    .B(_01545_),
    .Y(_01824_));
 AOI21x1_ASAP7_75t_R _24553_ (.A1(_01823_),
    .A2(_01824_),
    .B(_01689_),
    .Y(_01825_));
 NOR2x2_ASAP7_75t_R _24554_ (.A(_01616_),
    .B(_01544_),
    .Y(_01826_));
 NAND2x1_ASAP7_75t_R _24555_ (.A(_01753_),
    .B(_01826_),
    .Y(_01827_));
 NOR2x2_ASAP7_75t_R _24556_ (.A(_15920_),
    .B(net572),
    .Y(_01828_));
 OAI21x1_ASAP7_75t_R _24557_ (.A1(_01828_),
    .A2(_01807_),
    .B(_01545_),
    .Y(_01829_));
 AOI21x1_ASAP7_75t_R _24558_ (.A1(_01827_),
    .A2(_01829_),
    .B(_01674_),
    .Y(_01830_));
 NOR2x1_ASAP7_75t_R _24559_ (.A(_01825_),
    .B(_01830_),
    .Y(_01831_));
 OAI21x1_ASAP7_75t_R _24560_ (.A1(_01210_),
    .A2(_15933_),
    .B(_01746_),
    .Y(_01832_));
 AO21x1_ASAP7_75t_R _24561_ (.A1(_01832_),
    .A2(_01634_),
    .B(_01782_),
    .Y(_01833_));
 AOI21x1_ASAP7_75t_R _24562_ (.A1(_01669_),
    .A2(_01584_),
    .B(_01771_),
    .Y(_01834_));
 AOI21x1_ASAP7_75t_R _24563_ (.A1(_01726_),
    .A2(_01834_),
    .B(_01734_),
    .Y(_01835_));
 OAI21x1_ASAP7_75t_R _24564_ (.A1(_01740_),
    .A2(_01833_),
    .B(_01835_),
    .Y(_01836_));
 AOI21x1_ASAP7_75t_R _24565_ (.A1(_01831_),
    .A2(_01836_),
    .B(_01709_),
    .Y(_01837_));
 INVx1_ASAP7_75t_R _24566_ (.A(_01691_),
    .Y(_01838_));
 INVx1_ASAP7_75t_R _24567_ (.A(net606),
    .Y(_01839_));
 AOI21x1_ASAP7_75t_R _24568_ (.A1(_01839_),
    .A2(_15933_),
    .B(_01647_),
    .Y(_01840_));
 OAI21x1_ASAP7_75t_R _24569_ (.A1(_01781_),
    .A2(_01667_),
    .B(_01690_),
    .Y(_01841_));
 AOI22x1_ASAP7_75t_R _24570_ (.A1(_01553_),
    .A2(_01552_),
    .B1(_01522_),
    .B2(_01524_),
    .Y(_01842_));
 INVx2_ASAP7_75t_R _24571_ (.A(_01842_),
    .Y(_01843_));
 NOR2x2_ASAP7_75t_R _24572_ (.A(_01795_),
    .B(_01843_),
    .Y(_01844_));
 AOI211x1_ASAP7_75t_R _24573_ (.A1(_01838_),
    .A2(_01840_),
    .B(_01841_),
    .C(_01844_),
    .Y(_01845_));
 NOR2x2_ASAP7_75t_R _24574_ (.A(_01549_),
    .B(_01616_),
    .Y(_01846_));
 OAI21x1_ASAP7_75t_R _24575_ (.A1(_01846_),
    .A2(_01776_),
    .B(_01663_),
    .Y(_01847_));
 INVx1_ASAP7_75t_R _24576_ (.A(_00565_),
    .Y(_01848_));
 NOR2x1_ASAP7_75t_R _24577_ (.A(_01848_),
    .B(_01613_),
    .Y(_01849_));
 AOI21x1_ASAP7_75t_R _24578_ (.A1(_01750_),
    .A2(_01849_),
    .B(_01816_),
    .Y(_01850_));
 AOI21x1_ASAP7_75t_R _24579_ (.A1(_01847_),
    .A2(_01850_),
    .B(_01708_),
    .Y(_01851_));
 AOI21x1_ASAP7_75t_R _24580_ (.A1(_01654_),
    .A2(_01675_),
    .B(_01590_),
    .Y(_01852_));
 AOI21x1_ASAP7_75t_R _24581_ (.A1(_15925_),
    .A2(_01616_),
    .B(_01647_),
    .Y(_01853_));
 AOI21x1_ASAP7_75t_R _24582_ (.A1(_01584_),
    .A2(_01853_),
    .B(_01608_),
    .Y(_01854_));
 NAND2x1_ASAP7_75t_R _24583_ (.A(_01852_),
    .B(_01854_),
    .Y(_01855_));
 NAND2x1_ASAP7_75t_R _24584_ (.A(_01851_),
    .B(_01855_),
    .Y(_01856_));
 OAI21x1_ASAP7_75t_R _24585_ (.A1(_01845_),
    .A2(_01856_),
    .B(_01644_),
    .Y(_01857_));
 NOR2x1_ASAP7_75t_R _24586_ (.A(_01837_),
    .B(_01857_),
    .Y(_01858_));
 AOI21x1_ASAP7_75t_R _24587_ (.A1(_01769_),
    .A2(_01822_),
    .B(_01858_),
    .Y(_00089_));
 AND2x2_ASAP7_75t_R _24588_ (.A(_01208_),
    .B(_01207_),
    .Y(_01859_));
 NOR2x1_ASAP7_75t_R _24589_ (.A(_01859_),
    .B(_15933_),
    .Y(_01860_));
 OA21x2_ASAP7_75t_R _24590_ (.A1(_01617_),
    .A2(_01860_),
    .B(_01772_),
    .Y(_01861_));
 NAND2x1_ASAP7_75t_R _24591_ (.A(_01782_),
    .B(_01847_),
    .Y(_01862_));
 OAI21x1_ASAP7_75t_R _24592_ (.A1(_01723_),
    .A2(_01620_),
    .B(_01669_),
    .Y(_01863_));
 OA21x2_ASAP7_75t_R _24593_ (.A1(_01586_),
    .A2(_01551_),
    .B(_01590_),
    .Y(_01864_));
 AOI21x1_ASAP7_75t_R _24594_ (.A1(_01863_),
    .A2(_01864_),
    .B(_01750_),
    .Y(_01865_));
 OAI21x1_ASAP7_75t_R _24595_ (.A1(_01861_),
    .A2(_01862_),
    .B(_01865_),
    .Y(_01866_));
 BUFx10_ASAP7_75t_R _24596_ (.A(_01581_),
    .Y(_01867_));
 AND3x2_ASAP7_75t_R _24597_ (.A(_01543_),
    .B(_00566_),
    .C(_01536_),
    .Y(_01868_));
 AO21x1_ASAP7_75t_R _24598_ (.A1(_01676_),
    .A2(_01621_),
    .B(_01868_),
    .Y(_01869_));
 OA21x2_ASAP7_75t_R _24599_ (.A1(_01586_),
    .A2(_01214_),
    .B(_01581_),
    .Y(_01870_));
 OAI21x1_ASAP7_75t_R _24600_ (.A1(net71),
    .A2(_01616_),
    .B(_15923_),
    .Y(_01871_));
 NAND2x1_ASAP7_75t_R _24601_ (.A(_01555_),
    .B(_01871_),
    .Y(_01872_));
 AOI21x1_ASAP7_75t_R _24602_ (.A1(_01870_),
    .A2(_01872_),
    .B(_01734_),
    .Y(_01873_));
 OAI21x1_ASAP7_75t_R _24603_ (.A1(_01867_),
    .A2(_01869_),
    .B(_01873_),
    .Y(_01874_));
 AOI21x1_ASAP7_75t_R _24604_ (.A1(_01866_),
    .A2(_01874_),
    .B(_01716_),
    .Y(_01875_));
 AO21x1_ASAP7_75t_R _24605_ (.A1(_01746_),
    .A2(_01612_),
    .B(_01613_),
    .Y(_01876_));
 OAI21x1_ASAP7_75t_R _24606_ (.A1(_01805_),
    .A2(_01761_),
    .B(_01653_),
    .Y(_01877_));
 AOI21x1_ASAP7_75t_R _24607_ (.A1(_01876_),
    .A2(_01877_),
    .B(_01791_),
    .Y(_01878_));
 AO21x1_ASAP7_75t_R _24608_ (.A1(_01543_),
    .A2(_01536_),
    .B(_01848_),
    .Y(_01879_));
 BUFx6f_ASAP7_75t_R _24609_ (.A(_01554_),
    .Y(_01880_));
 OAI21x1_ASAP7_75t_R _24610_ (.A1(_01828_),
    .A2(_01807_),
    .B(_01880_),
    .Y(_01881_));
 AOI21x1_ASAP7_75t_R _24611_ (.A1(_01879_),
    .A2(_01881_),
    .B(_01582_),
    .Y(_01882_));
 OAI21x1_ASAP7_75t_R _24612_ (.A1(_01878_),
    .A2(_01882_),
    .B(_01764_),
    .Y(_01883_));
 OA21x2_ASAP7_75t_R _24613_ (.A1(_01586_),
    .A2(_01212_),
    .B(_01590_),
    .Y(_01884_));
 OAI21x1_ASAP7_75t_R _24614_ (.A1(_01747_),
    .A2(_01738_),
    .B(_01669_),
    .Y(_01885_));
 AOI21x1_ASAP7_75t_R _24615_ (.A1(_01884_),
    .A2(_01885_),
    .B(_01750_),
    .Y(_01886_));
 OAI21x1_ASAP7_75t_R _24616_ (.A1(net573),
    .A2(_01616_),
    .B(_01554_),
    .Y(_01887_));
 AOI21x1_ASAP7_75t_R _24617_ (.A1(_01653_),
    .A2(_01712_),
    .B(_01635_),
    .Y(_01888_));
 OAI21x1_ASAP7_75t_R _24618_ (.A1(_01691_),
    .A2(_01887_),
    .B(_01888_),
    .Y(_01889_));
 NAND2x1_ASAP7_75t_R _24619_ (.A(_01886_),
    .B(_01889_),
    .Y(_01890_));
 AOI21x1_ASAP7_75t_R _24620_ (.A1(_01883_),
    .A2(_01890_),
    .B(_01644_),
    .Y(_01891_));
 OAI21x1_ASAP7_75t_R _24621_ (.A1(_01875_),
    .A2(_01891_),
    .B(_01708_),
    .Y(_01892_));
 OAI21x1_ASAP7_75t_R _24622_ (.A1(_01588_),
    .A2(_01620_),
    .B(_01669_),
    .Y(_01893_));
 OA21x2_ASAP7_75t_R _24623_ (.A1(_01520_),
    .A2(_01519_),
    .B(_01727_),
    .Y(_01894_));
 OAI21x1_ASAP7_75t_R _24624_ (.A1(_01894_),
    .A2(_01793_),
    .B(_01653_),
    .Y(_01895_));
 AOI21x1_ASAP7_75t_R _24625_ (.A1(_01893_),
    .A2(_01895_),
    .B(_01782_),
    .Y(_01896_));
 INVx3_ASAP7_75t_R _24626_ (.A(_01728_),
    .Y(_01897_));
 NOR2x1_ASAP7_75t_R _24627_ (.A(_01897_),
    .B(_01887_),
    .Y(_01898_));
 OAI21x1_ASAP7_75t_R _24628_ (.A1(_01519_),
    .A2(_01520_),
    .B(_01661_),
    .Y(_01899_));
 NAND2x1_ASAP7_75t_R _24629_ (.A(_01899_),
    .B(_01625_),
    .Y(_01900_));
 OAI21x1_ASAP7_75t_R _24630_ (.A1(_01793_),
    .A2(_01900_),
    .B(_01816_),
    .Y(_01901_));
 NOR2x1_ASAP7_75t_R _24631_ (.A(_01898_),
    .B(_01901_),
    .Y(_01902_));
 OAI21x1_ASAP7_75t_R _24632_ (.A1(_01896_),
    .A2(_01902_),
    .B(_01671_),
    .Y(_01903_));
 AO21x1_ASAP7_75t_R _24633_ (.A1(_01728_),
    .A2(_01899_),
    .B(_01586_),
    .Y(_01904_));
 OAI21x1_ASAP7_75t_R _24634_ (.A1(_01723_),
    .A2(_01793_),
    .B(_01811_),
    .Y(_01905_));
 AOI21x1_ASAP7_75t_R _24635_ (.A1(_01904_),
    .A2(_01905_),
    .B(_01791_),
    .Y(_01906_));
 OAI21x1_ASAP7_75t_R _24636_ (.A1(_01897_),
    .A2(_01723_),
    .B(_01653_),
    .Y(_01907_));
 OAI21x1_ASAP7_75t_R _24637_ (.A1(_01723_),
    .A2(_01761_),
    .B(_01811_),
    .Y(_01908_));
 AOI21x1_ASAP7_75t_R _24638_ (.A1(_01907_),
    .A2(_01908_),
    .B(_01582_),
    .Y(_01909_));
 OAI21x1_ASAP7_75t_R _24639_ (.A1(_01906_),
    .A2(_01909_),
    .B(_01764_),
    .Y(_01910_));
 AOI21x1_ASAP7_75t_R _24640_ (.A1(_01903_),
    .A2(_01910_),
    .B(_01644_),
    .Y(_01911_));
 OAI21x1_ASAP7_75t_R _24641_ (.A1(_01723_),
    .A2(_01738_),
    .B(_01880_),
    .Y(_01912_));
 AO21x1_ASAP7_75t_R _24642_ (.A1(_01668_),
    .A2(_01746_),
    .B(_01586_),
    .Y(_01913_));
 AOI21x1_ASAP7_75t_R _24643_ (.A1(_01912_),
    .A2(_01913_),
    .B(_01782_),
    .Y(_01914_));
 AOI21x1_ASAP7_75t_R _24644_ (.A1(_01779_),
    .A2(_01899_),
    .B(_01647_),
    .Y(_01915_));
 AOI21x1_ASAP7_75t_R _24645_ (.A1(_01555_),
    .A2(_01871_),
    .B(_01915_),
    .Y(_01916_));
 OAI21x1_ASAP7_75t_R _24646_ (.A1(_01611_),
    .A2(_01916_),
    .B(_01750_),
    .Y(_01917_));
 NOR2x1_ASAP7_75t_R _24647_ (.A(_01914_),
    .B(_01917_),
    .Y(_01918_));
 NAND2x2_ASAP7_75t_R _24648_ (.A(_01544_),
    .B(_01525_),
    .Y(_01919_));
 NOR2x1_ASAP7_75t_R _24649_ (.A(_01655_),
    .B(_01919_),
    .Y(_01920_));
 AND3x1_ASAP7_75t_R _24650_ (.A(_01626_),
    .B(_01647_),
    .C(_01741_),
    .Y(_01921_));
 OAI21x1_ASAP7_75t_R _24651_ (.A1(_01920_),
    .A2(_01921_),
    .B(_01690_),
    .Y(_01922_));
 NOR2x2_ASAP7_75t_R _24652_ (.A(net890),
    .B(_01517_),
    .Y(_01923_));
 OAI21x1_ASAP7_75t_R _24653_ (.A1(_01923_),
    .A2(_01617_),
    .B(_01669_),
    .Y(_01924_));
 AOI21x1_ASAP7_75t_R _24654_ (.A1(_01653_),
    .A2(_01676_),
    .B(_01674_),
    .Y(_01925_));
 AOI21x1_ASAP7_75t_R _24655_ (.A1(_01924_),
    .A2(_01925_),
    .B(_01716_),
    .Y(_01926_));
 NAND2x1_ASAP7_75t_R _24656_ (.A(_01922_),
    .B(_01926_),
    .Y(_01927_));
 NOR2x1_ASAP7_75t_R _24657_ (.A(_01918_),
    .B(_01927_),
    .Y(_01928_));
 OAI21x1_ASAP7_75t_R _24658_ (.A1(_01911_),
    .A2(_01928_),
    .B(_01710_),
    .Y(_01929_));
 NAND2x1_ASAP7_75t_R _24659_ (.A(_01892_),
    .B(_01929_),
    .Y(_00090_));
 NOR2x2_ASAP7_75t_R _24660_ (.A(_01586_),
    .B(_01694_),
    .Y(_01930_));
 AOI22x1_ASAP7_75t_R _24661_ (.A1(_01930_),
    .A2(_01671_),
    .B1(_01775_),
    .B2(_01801_),
    .Y(_01931_));
 NAND2x2_ASAP7_75t_R _24662_ (.A(net885),
    .B(net877),
    .Y(_01932_));
 AO21x1_ASAP7_75t_R _24663_ (.A1(_01932_),
    .A2(_01550_),
    .B(_01555_),
    .Y(_01933_));
 AO21x1_ASAP7_75t_R _24664_ (.A1(_01933_),
    .A2(_01589_),
    .B(_01671_),
    .Y(_01934_));
 AOI21x1_ASAP7_75t_R _24665_ (.A1(_01931_),
    .A2(_01934_),
    .B(_01591_),
    .Y(_01935_));
 OA21x2_ASAP7_75t_R _24666_ (.A1(_01545_),
    .A2(_01728_),
    .B(_01608_),
    .Y(_01936_));
 AO21x1_ASAP7_75t_R _24667_ (.A1(_01936_),
    .A2(_01895_),
    .B(_01867_),
    .Y(_01937_));
 NAND2x2_ASAP7_75t_R _24668_ (.A(_01859_),
    .B(_01616_),
    .Y(_01938_));
 INVx1_ASAP7_75t_R _24669_ (.A(_01695_),
    .Y(_01939_));
 AND3x1_ASAP7_75t_R _24670_ (.A(_01938_),
    .B(_01939_),
    .C(_01555_),
    .Y(_01940_));
 NAND2x2_ASAP7_75t_R _24671_ (.A(_01625_),
    .B(_01648_),
    .Y(_01941_));
 NOR2x2_ASAP7_75t_R _24672_ (.A(_01731_),
    .B(_01941_),
    .Y(_01942_));
 NOR3x1_ASAP7_75t_R _24673_ (.A(_01940_),
    .B(_01942_),
    .C(_01671_),
    .Y(_01943_));
 OAI21x1_ASAP7_75t_R _24674_ (.A1(_01937_),
    .A2(_01943_),
    .B(_01644_),
    .Y(_01944_));
 NOR2x1_ASAP7_75t_R _24675_ (.A(_01935_),
    .B(_01944_),
    .Y(_01945_));
 AND3x1_ASAP7_75t_R _24676_ (.A(_01694_),
    .B(_01939_),
    .C(_01802_),
    .Y(_01946_));
 OAI21x1_ASAP7_75t_R _24677_ (.A1(_15925_),
    .A2(_15930_),
    .B(_01728_),
    .Y(_01947_));
 AO21x1_ASAP7_75t_R _24678_ (.A1(_01947_),
    .A2(_01634_),
    .B(_01689_),
    .Y(_01948_));
 AOI21x1_ASAP7_75t_R _24679_ (.A1(_01811_),
    .A2(_01743_),
    .B(_01674_),
    .Y(_01949_));
 NAND2x1_ASAP7_75t_R _24680_ (.A(_01829_),
    .B(_01949_),
    .Y(_01950_));
 OAI21x1_ASAP7_75t_R _24681_ (.A1(_01946_),
    .A2(_01948_),
    .B(_01950_),
    .Y(_01951_));
 NAND2x1_ASAP7_75t_R _24682_ (.A(_01938_),
    .B(_01760_),
    .Y(_01952_));
 NAND2x1_ASAP7_75t_R _24683_ (.A(_01847_),
    .B(_01952_),
    .Y(_01953_));
 NAND2x1_ASAP7_75t_R _24684_ (.A(_01750_),
    .B(_01901_),
    .Y(_01954_));
 AOI21x1_ASAP7_75t_R _24685_ (.A1(_01591_),
    .A2(_01953_),
    .B(_01954_),
    .Y(_01955_));
 OAI21x1_ASAP7_75t_R _24686_ (.A1(_01951_),
    .A2(_01955_),
    .B(_01769_),
    .Y(_01956_));
 NAND2x1_ASAP7_75t_R _24687_ (.A(_01710_),
    .B(_01956_),
    .Y(_01957_));
 OAI21x1_ASAP7_75t_R _24688_ (.A1(_01731_),
    .A2(_01846_),
    .B(_01802_),
    .Y(_01958_));
 NOR2x2_ASAP7_75t_R _24689_ (.A(_15925_),
    .B(_15921_),
    .Y(_01959_));
 OAI21x1_ASAP7_75t_R _24690_ (.A1(_01789_),
    .A2(_01959_),
    .B(_01772_),
    .Y(_01960_));
 AOI21x1_ASAP7_75t_R _24691_ (.A1(_01958_),
    .A2(_01960_),
    .B(_01791_),
    .Y(_01961_));
 OAI21x1_ASAP7_75t_R _24692_ (.A1(net71),
    .A2(_01616_),
    .B(_01612_),
    .Y(_01962_));
 NOR2x1_ASAP7_75t_R _24693_ (.A(_01962_),
    .B(_01887_),
    .Y(_01963_));
 NAND2x1_ASAP7_75t_R _24694_ (.A(_01746_),
    .B(_01613_),
    .Y(_01964_));
 OAI21x1_ASAP7_75t_R _24695_ (.A1(_01964_),
    .A2(_01776_),
    .B(_01635_),
    .Y(_01965_));
 NOR2x1_ASAP7_75t_R _24696_ (.A(_01963_),
    .B(_01965_),
    .Y(_01966_));
 OAI21x1_ASAP7_75t_R _24697_ (.A1(_01961_),
    .A2(_01966_),
    .B(_01609_),
    .Y(_01967_));
 OAI21x1_ASAP7_75t_R _24698_ (.A1(net71),
    .A2(_15930_),
    .B(_01580_),
    .Y(_01968_));
 NOR2x2_ASAP7_75t_R _24699_ (.A(_01624_),
    .B(_01968_),
    .Y(_01969_));
 AOI21x1_ASAP7_75t_R _24700_ (.A1(_01843_),
    .A2(_01969_),
    .B(_01734_),
    .Y(_01970_));
 AOI21x1_ASAP7_75t_R _24701_ (.A1(_01932_),
    .A2(_01696_),
    .B(_01635_),
    .Y(_01971_));
 AO21x2_ASAP7_75t_R _24702_ (.A1(_01547_),
    .A2(_01548_),
    .B(_01727_),
    .Y(_01972_));
 NOR2x1_ASAP7_75t_R _24703_ (.A(_01647_),
    .B(_01620_),
    .Y(_01973_));
 NAND2x1_ASAP7_75t_R _24704_ (.A(_01972_),
    .B(_01973_),
    .Y(_01974_));
 NAND2x1_ASAP7_75t_R _24705_ (.A(_01971_),
    .B(_01974_),
    .Y(_01975_));
 AOI21x1_ASAP7_75t_R _24706_ (.A1(_01970_),
    .A2(_01975_),
    .B(_01643_),
    .Y(_01976_));
 AOI21x1_ASAP7_75t_R _24707_ (.A1(_01967_),
    .A2(_01976_),
    .B(_01709_),
    .Y(_01977_));
 AOI21x1_ASAP7_75t_R _24708_ (.A1(_01654_),
    .A2(_01732_),
    .B(_01608_),
    .Y(_01978_));
 OAI21x1_ASAP7_75t_R _24709_ (.A1(_01959_),
    .A2(_01627_),
    .B(_01978_),
    .Y(_01979_));
 OAI21x1_ASAP7_75t_R _24710_ (.A1(_01723_),
    .A2(_01923_),
    .B(_01811_),
    .Y(_01980_));
 AOI21x1_ASAP7_75t_R _24711_ (.A1(_01654_),
    .A2(_01973_),
    .B(_01750_),
    .Y(_01981_));
 AOI21x1_ASAP7_75t_R _24712_ (.A1(_01980_),
    .A2(_01981_),
    .B(_01582_),
    .Y(_01982_));
 NAND2x1_ASAP7_75t_R _24713_ (.A(_01979_),
    .B(_01982_),
    .Y(_01983_));
 NOR2x2_ASAP7_75t_R _24714_ (.A(_01625_),
    .B(_01588_),
    .Y(_01984_));
 NOR2x1_ASAP7_75t_R _24715_ (.A(_01608_),
    .B(_01984_),
    .Y(_01985_));
 AO21x1_ASAP7_75t_R _24716_ (.A1(_01584_),
    .A2(_01626_),
    .B(_01880_),
    .Y(_01986_));
 AOI21x1_ASAP7_75t_R _24717_ (.A1(_01985_),
    .A2(_01986_),
    .B(_01791_),
    .Y(_01987_));
 AOI21x1_ASAP7_75t_R _24718_ (.A1(net607),
    .A2(_01842_),
    .B(_01750_),
    .Y(_01988_));
 NAND2x1_ASAP7_75t_R _24719_ (.A(_01545_),
    .B(_01962_),
    .Y(_01989_));
 NAND3x1_ASAP7_75t_R _24720_ (.A(_01988_),
    .B(_01989_),
    .C(_01589_),
    .Y(_01990_));
 AOI21x1_ASAP7_75t_R _24721_ (.A1(_01987_),
    .A2(_01990_),
    .B(_01716_),
    .Y(_01991_));
 NAND2x1_ASAP7_75t_R _24722_ (.A(_01983_),
    .B(_01991_),
    .Y(_01992_));
 NAND2x1_ASAP7_75t_R _24723_ (.A(_01977_),
    .B(_01992_),
    .Y(_01993_));
 OAI21x1_ASAP7_75t_R _24724_ (.A1(_01945_),
    .A2(_01957_),
    .B(_01993_),
    .Y(_00091_));
 OAI21x1_ASAP7_75t_R _24725_ (.A1(_01894_),
    .A2(_01761_),
    .B(_01555_),
    .Y(_01994_));
 NAND2x1_ASAP7_75t_R _24726_ (.A(_01613_),
    .B(_01793_),
    .Y(_01995_));
 INVx1_ASAP7_75t_R _24727_ (.A(_01995_),
    .Y(_01996_));
 AOI211x1_ASAP7_75t_R _24728_ (.A1(_01781_),
    .A2(_01771_),
    .B(_01996_),
    .C(_01689_),
    .Y(_01997_));
 NOR2x2_ASAP7_75t_R _24729_ (.A(_01746_),
    .B(_01625_),
    .Y(_01998_));
 NOR2x1_ASAP7_75t_R _24730_ (.A(_00567_),
    .B(_01669_),
    .Y(_01999_));
 OA211x2_ASAP7_75t_R _24731_ (.A1(_01998_),
    .A2(_01999_),
    .B(_01611_),
    .C(_01734_),
    .Y(_02000_));
 AOI21x1_ASAP7_75t_R _24732_ (.A1(_01994_),
    .A2(_01997_),
    .B(_02000_),
    .Y(_02001_));
 AOI211x1_ASAP7_75t_R _24733_ (.A1(_01633_),
    .A2(_01775_),
    .B(_01717_),
    .C(_01867_),
    .Y(_02002_));
 AND3x1_ASAP7_75t_R _24734_ (.A(_01626_),
    .B(_01972_),
    .C(_01811_),
    .Y(_02003_));
 AO21x1_ASAP7_75t_R _24735_ (.A1(_01932_),
    .A2(_01650_),
    .B(_01586_),
    .Y(_02004_));
 NAND2x1_ASAP7_75t_R _24736_ (.A(_01582_),
    .B(_02004_),
    .Y(_02005_));
 NOR2x1_ASAP7_75t_R _24737_ (.A(_02003_),
    .B(_02005_),
    .Y(_02006_));
 OAI21x1_ASAP7_75t_R _24738_ (.A1(_02002_),
    .A2(_02006_),
    .B(_01770_),
    .Y(_02007_));
 AOI21x1_ASAP7_75t_R _24739_ (.A1(_02001_),
    .A2(_02007_),
    .B(_01769_),
    .Y(_02008_));
 AO21x1_ASAP7_75t_R _24740_ (.A1(_01788_),
    .A2(_01653_),
    .B(_01635_),
    .Y(_02009_));
 OAI21x1_ASAP7_75t_R _24741_ (.A1(_01775_),
    .A2(_01654_),
    .B(_01808_),
    .Y(_02010_));
 NOR2x1_ASAP7_75t_R _24742_ (.A(_01816_),
    .B(_01826_),
    .Y(_02011_));
 OAI21x1_ASAP7_75t_R _24743_ (.A1(_01627_),
    .A2(_01695_),
    .B(_02011_),
    .Y(_02012_));
 OAI21x1_ASAP7_75t_R _24744_ (.A1(_02009_),
    .A2(_02010_),
    .B(_02012_),
    .Y(_02013_));
 OAI21x1_ASAP7_75t_R _24745_ (.A1(_01649_),
    .A2(_01651_),
    .B(_01791_),
    .Y(_02014_));
 AO21x1_ASAP7_75t_R _24746_ (.A1(_01587_),
    .A2(_01779_),
    .B(_01880_),
    .Y(_02015_));
 NAND2x1_ASAP7_75t_R _24747_ (.A(_01734_),
    .B(_02015_),
    .Y(_02016_));
 OAI21x1_ASAP7_75t_R _24748_ (.A1(_15930_),
    .A2(_01650_),
    .B(_01772_),
    .Y(_02017_));
 AO21x1_ASAP7_75t_R _24749_ (.A1(_01547_),
    .A2(_01548_),
    .B(_01656_),
    .Y(_02018_));
 AOI21x1_ASAP7_75t_R _24750_ (.A1(_01802_),
    .A2(_02018_),
    .B(_01689_),
    .Y(_02019_));
 NAND2x1_ASAP7_75t_R _24751_ (.A(_02017_),
    .B(_02019_),
    .Y(_02020_));
 OAI21x1_ASAP7_75t_R _24752_ (.A1(_02014_),
    .A2(_02016_),
    .B(_02020_),
    .Y(_02021_));
 AOI21x1_ASAP7_75t_R _24753_ (.A1(_01770_),
    .A2(_02013_),
    .B(_02021_),
    .Y(_02022_));
 OAI21x1_ASAP7_75t_R _24754_ (.A1(_01644_),
    .A2(_02022_),
    .B(_01710_),
    .Y(_02023_));
 NAND2x1_ASAP7_75t_R _24755_ (.A(_01657_),
    .B(_01581_),
    .Y(_02024_));
 OA21x2_ASAP7_75t_R _24756_ (.A1(_01760_),
    .A2(_02024_),
    .B(_01734_),
    .Y(_02025_));
 AO21x1_ASAP7_75t_R _24757_ (.A1(_01654_),
    .A2(_01626_),
    .B(_01613_),
    .Y(_02026_));
 AOI21x1_ASAP7_75t_R _24758_ (.A1(_01838_),
    .A2(_01840_),
    .B(_01816_),
    .Y(_02027_));
 NAND2x1_ASAP7_75t_R _24759_ (.A(_02026_),
    .B(_02027_),
    .Y(_02028_));
 AOI21x1_ASAP7_75t_R _24760_ (.A1(_02025_),
    .A2(_02028_),
    .B(_01643_),
    .Y(_02029_));
 NAND2x1_ASAP7_75t_R _24761_ (.A(_01584_),
    .B(_01853_),
    .Y(_02030_));
 AOI21x1_ASAP7_75t_R _24762_ (.A1(_01881_),
    .A2(_02030_),
    .B(_01582_),
    .Y(_02031_));
 AO21x1_ASAP7_75t_R _24763_ (.A1(_01654_),
    .A2(_01753_),
    .B(_01880_),
    .Y(_02032_));
 AO21x1_ASAP7_75t_R _24764_ (.A1(_01668_),
    .A2(_01526_),
    .B(_01663_),
    .Y(_02033_));
 AOI21x1_ASAP7_75t_R _24765_ (.A1(_02032_),
    .A2(_02033_),
    .B(_01791_),
    .Y(_02034_));
 OAI21x1_ASAP7_75t_R _24766_ (.A1(_02031_),
    .A2(_02034_),
    .B(_01770_),
    .Y(_02035_));
 NAND2x1_ASAP7_75t_R _24767_ (.A(_02029_),
    .B(_02035_),
    .Y(_02036_));
 OAI21x1_ASAP7_75t_R _24768_ (.A1(net70),
    .A2(_15930_),
    .B(_01551_),
    .Y(_02037_));
 AOI21x1_ASAP7_75t_R _24769_ (.A1(_01669_),
    .A2(_02037_),
    .B(_01816_),
    .Y(_02038_));
 NAND2x1_ASAP7_75t_R _24770_ (.A(_01739_),
    .B(_02038_),
    .Y(_02039_));
 OAI21x1_ASAP7_75t_R _24771_ (.A1(_01807_),
    .A2(_01738_),
    .B(_01772_),
    .Y(_02040_));
 NOR2x1_ASAP7_75t_R _24772_ (.A(_01635_),
    .B(_01915_),
    .Y(_02041_));
 AOI21x1_ASAP7_75t_R _24773_ (.A1(_02040_),
    .A2(_02041_),
    .B(_01734_),
    .Y(_02042_));
 NAND2x1_ASAP7_75t_R _24774_ (.A(_02039_),
    .B(_02042_),
    .Y(_02043_));
 NOR2x1_ASAP7_75t_R _24775_ (.A(_01897_),
    .B(_01998_),
    .Y(_02044_));
 AOI21x1_ASAP7_75t_R _24776_ (.A1(_01726_),
    .A2(_02044_),
    .B(_01764_),
    .Y(_02045_));
 AOI21x1_ASAP7_75t_R _24777_ (.A1(_01802_),
    .A2(_01832_),
    .B(_01816_),
    .Y(_02046_));
 NAND2x1_ASAP7_75t_R _24778_ (.A(_02046_),
    .B(_01763_),
    .Y(_02047_));
 AOI21x1_ASAP7_75t_R _24779_ (.A1(_02045_),
    .A2(_02047_),
    .B(_01716_),
    .Y(_02048_));
 AOI21x1_ASAP7_75t_R _24780_ (.A1(_02043_),
    .A2(_02048_),
    .B(_01710_),
    .Y(_02049_));
 NAND2x1_ASAP7_75t_R _24781_ (.A(_02036_),
    .B(_02049_),
    .Y(_02050_));
 OAI21x1_ASAP7_75t_R _24782_ (.A1(_02008_),
    .A2(_02023_),
    .B(_02050_),
    .Y(_00092_));
 OA21x2_ASAP7_75t_R _24783_ (.A1(_01721_),
    .A2(_15933_),
    .B(_01802_),
    .Y(_02051_));
 AOI211x1_ASAP7_75t_R _24784_ (.A1(_01753_),
    .A2(_01826_),
    .B(_02051_),
    .C(_01591_),
    .Y(_02052_));
 AO21x1_ASAP7_75t_R _24785_ (.A1(_01694_),
    .A2(_01621_),
    .B(_01782_),
    .Y(_02053_));
 NAND2x1_ASAP7_75t_R _24786_ (.A(_01555_),
    .B(_01947_),
    .Y(_02054_));
 INVx1_ASAP7_75t_R _24787_ (.A(_02054_),
    .Y(_02055_));
 OAI21x1_ASAP7_75t_R _24788_ (.A1(_02053_),
    .A2(_02055_),
    .B(_01770_),
    .Y(_02056_));
 OAI21x1_ASAP7_75t_R _24789_ (.A1(_02052_),
    .A2(_02056_),
    .B(_01769_),
    .Y(_02057_));
 INVx2_ASAP7_75t_R _24790_ (.A(_01899_),
    .Y(_02058_));
 OA21x2_ASAP7_75t_R _24791_ (.A1(_01780_),
    .A2(_02058_),
    .B(_01811_),
    .Y(_02059_));
 NOR2x1_ASAP7_75t_R _24792_ (.A(_02059_),
    .B(_01659_),
    .Y(_02060_));
 NAND2x1_ASAP7_75t_R _24793_ (.A(_01663_),
    .B(_01972_),
    .Y(_02061_));
 NOR2x1_ASAP7_75t_R _24794_ (.A(_02061_),
    .B(_01754_),
    .Y(_02062_));
 AO21x1_ASAP7_75t_R _24795_ (.A1(_01553_),
    .A2(_01552_),
    .B(_01208_),
    .Y(_02063_));
 NAND2x1_ASAP7_75t_R _24796_ (.A(_02063_),
    .B(_01757_),
    .Y(_02064_));
 OAI21x1_ASAP7_75t_R _24797_ (.A1(_02062_),
    .A2(_02064_),
    .B(_01609_),
    .Y(_02065_));
 NOR2x1_ASAP7_75t_R _24798_ (.A(_02060_),
    .B(_02065_),
    .Y(_02066_));
 OAI21x1_ASAP7_75t_R _24799_ (.A1(_02057_),
    .A2(_02066_),
    .B(_01708_),
    .Y(_02067_));
 AND2x2_ASAP7_75t_R _24800_ (.A(_01900_),
    .B(_01590_),
    .Y(_02068_));
 NAND2x1_ASAP7_75t_R _24801_ (.A(_01526_),
    .B(_01732_),
    .Y(_02069_));
 AOI21x1_ASAP7_75t_R _24802_ (.A1(_02068_),
    .A2(_02069_),
    .B(_01671_),
    .Y(_02070_));
 INVx1_ASAP7_75t_R _24803_ (.A(_01741_),
    .Y(_02071_));
 OA21x2_ASAP7_75t_R _24804_ (.A1(_01771_),
    .A2(_02071_),
    .B(_01621_),
    .Y(_02072_));
 OAI21x1_ASAP7_75t_R _24805_ (.A1(_01998_),
    .A2(_02072_),
    .B(_01867_),
    .Y(_02073_));
 NAND2x1_ASAP7_75t_R _24806_ (.A(_02070_),
    .B(_02073_),
    .Y(_02074_));
 AO21x1_ASAP7_75t_R _24807_ (.A1(_01677_),
    .A2(_01650_),
    .B(_01591_),
    .Y(_02075_));
 AND3x1_ASAP7_75t_R _24808_ (.A(_01777_),
    .B(_01775_),
    .C(_01550_),
    .Y(_02076_));
 OA21x2_ASAP7_75t_R _24809_ (.A1(_01802_),
    .A2(_15923_),
    .B(_01611_),
    .Y(_02077_));
 AOI21x1_ASAP7_75t_R _24810_ (.A1(_02077_),
    .A2(_02004_),
    .B(_01764_),
    .Y(_02078_));
 OAI21x1_ASAP7_75t_R _24811_ (.A1(_02075_),
    .A2(_02076_),
    .B(_02078_),
    .Y(_02079_));
 AOI21x1_ASAP7_75t_R _24812_ (.A1(_02074_),
    .A2(_02079_),
    .B(_01769_),
    .Y(_02080_));
 AND3x1_ASAP7_75t_R _24813_ (.A(_01755_),
    .B(_01694_),
    .C(_01880_),
    .Y(_02081_));
 OAI21x1_ASAP7_75t_R _24814_ (.A1(_01695_),
    .A2(_01919_),
    .B(_01782_),
    .Y(_02082_));
 NOR2x1_ASAP7_75t_R _24815_ (.A(_02081_),
    .B(_02082_),
    .Y(_02083_));
 AO21x1_ASAP7_75t_R _24816_ (.A1(_01772_),
    .A2(_00561_),
    .B(_01782_),
    .Y(_02084_));
 NOR2x1_ASAP7_75t_R _24817_ (.A(_01775_),
    .B(_01651_),
    .Y(_02085_));
 OAI21x1_ASAP7_75t_R _24818_ (.A1(_02084_),
    .A2(_02085_),
    .B(_01764_),
    .Y(_02086_));
 NOR2x1_ASAP7_75t_R _24819_ (.A(_02083_),
    .B(_02086_),
    .Y(_02087_));
 AO21x1_ASAP7_75t_R _24820_ (.A1(_01726_),
    .A2(_01773_),
    .B(_01764_),
    .Y(_02088_));
 AOI21x1_ASAP7_75t_R _24821_ (.A1(_01775_),
    .A2(_01938_),
    .B(_01782_),
    .Y(_02089_));
 OA21x2_ASAP7_75t_R _24822_ (.A1(_01692_),
    .A2(_01651_),
    .B(_02089_),
    .Y(_02090_));
 OAI21x1_ASAP7_75t_R _24823_ (.A1(_02088_),
    .A2(_02090_),
    .B(_01644_),
    .Y(_02091_));
 OAI21x1_ASAP7_75t_R _24824_ (.A1(_02087_),
    .A2(_02091_),
    .B(_01710_),
    .Y(_02092_));
 NOR2x1_ASAP7_75t_R _24825_ (.A(_01996_),
    .B(_01725_),
    .Y(_02093_));
 AO21x1_ASAP7_75t_R _24826_ (.A1(_01846_),
    .A2(_01669_),
    .B(_01635_),
    .Y(_02094_));
 OA21x2_ASAP7_75t_R _24827_ (.A1(_01776_),
    .A2(_02058_),
    .B(_01802_),
    .Y(_02095_));
 OAI21x1_ASAP7_75t_R _24828_ (.A1(_02094_),
    .A2(_02095_),
    .B(_01764_),
    .Y(_02096_));
 NOR2x1_ASAP7_75t_R _24829_ (.A(_02093_),
    .B(_02096_),
    .Y(_02097_));
 AO21x1_ASAP7_75t_R _24830_ (.A1(_01772_),
    .A2(_15925_),
    .B(_01816_),
    .Y(_02098_));
 OAI21x1_ASAP7_75t_R _24831_ (.A1(_02098_),
    .A2(_01628_),
    .B(_01671_),
    .Y(_02099_));
 AND2x2_ASAP7_75t_R _24832_ (.A(_01732_),
    .B(_01676_),
    .Y(_02100_));
 OAI21x1_ASAP7_75t_R _24833_ (.A1(_01894_),
    .A2(_01761_),
    .B(_01545_),
    .Y(_02101_));
 NAND2x1_ASAP7_75t_R _24834_ (.A(_01782_),
    .B(_02101_),
    .Y(_02102_));
 NOR2x1_ASAP7_75t_R _24835_ (.A(_02100_),
    .B(_02102_),
    .Y(_02103_));
 OAI21x1_ASAP7_75t_R _24836_ (.A1(_02099_),
    .A2(_02103_),
    .B(_01769_),
    .Y(_02104_));
 NOR2x1_ASAP7_75t_R _24837_ (.A(_02097_),
    .B(_02104_),
    .Y(_02105_));
 OAI22x1_ASAP7_75t_R _24838_ (.A1(_02067_),
    .A2(_02080_),
    .B1(_02092_),
    .B2(_02105_),
    .Y(_00093_));
 AOI21x1_ASAP7_75t_R _24839_ (.A1(_01657_),
    .A2(_01784_),
    .B(_01781_),
    .Y(_02106_));
 OA21x2_ASAP7_75t_R _24840_ (.A1(_01923_),
    .A2(_01894_),
    .B(_01621_),
    .Y(_02107_));
 OAI21x1_ASAP7_75t_R _24841_ (.A1(_02106_),
    .A2(_02107_),
    .B(_01591_),
    .Y(_02108_));
 NOR2x1_ASAP7_75t_R _24842_ (.A(_01859_),
    .B(_15930_),
    .Y(_02109_));
 OA21x2_ASAP7_75t_R _24843_ (.A1(_02109_),
    .A2(_01897_),
    .B(_01775_),
    .Y(_02110_));
 OA21x2_ASAP7_75t_R _24844_ (.A1(_01691_),
    .A2(_01588_),
    .B(_01781_),
    .Y(_02111_));
 OAI21x1_ASAP7_75t_R _24845_ (.A1(_02110_),
    .A2(_02111_),
    .B(_01867_),
    .Y(_02112_));
 AOI21x1_ASAP7_75t_R _24846_ (.A1(_02108_),
    .A2(_02112_),
    .B(_01609_),
    .Y(_02113_));
 OA21x2_ASAP7_75t_R _24847_ (.A1(_02071_),
    .A2(_01897_),
    .B(_01634_),
    .Y(_02114_));
 OAI21x1_ASAP7_75t_R _24848_ (.A1(_02009_),
    .A2(_02114_),
    .B(_01609_),
    .Y(_02115_));
 AND2x2_ASAP7_75t_R _24849_ (.A(_01213_),
    .B(_01211_),
    .Y(_02116_));
 OA21x2_ASAP7_75t_R _24850_ (.A1(_01880_),
    .A2(_02116_),
    .B(_01635_),
    .Y(_02117_));
 OA21x2_ASAP7_75t_R _24851_ (.A1(_01887_),
    .A2(_01959_),
    .B(_02117_),
    .Y(_02118_));
 OAI21x1_ASAP7_75t_R _24852_ (.A1(_02115_),
    .A2(_02118_),
    .B(_01769_),
    .Y(_02119_));
 AOI21x1_ASAP7_75t_R _24853_ (.A1(_01663_),
    .A2(_01588_),
    .B(_01581_),
    .Y(_02120_));
 NAND2x1_ASAP7_75t_R _24854_ (.A(_01663_),
    .B(_01860_),
    .Y(_02121_));
 NAND2x1_ASAP7_75t_R _24855_ (.A(_02121_),
    .B(_02120_),
    .Y(_02122_));
 INVx1_ASAP7_75t_R _24856_ (.A(_01738_),
    .Y(_02123_));
 AOI21x1_ASAP7_75t_R _24857_ (.A1(_01648_),
    .A2(_02123_),
    .B(_01781_),
    .Y(_02124_));
 NOR2x1_ASAP7_75t_R _24858_ (.A(_02124_),
    .B(_02122_),
    .Y(_02125_));
 AOI21x1_ASAP7_75t_R _24859_ (.A1(_15923_),
    .A2(_01626_),
    .B(_01781_),
    .Y(_02126_));
 AO21x1_ASAP7_75t_R _24860_ (.A1(_01846_),
    .A2(_01781_),
    .B(_01611_),
    .Y(_02127_));
 OAI21x1_ASAP7_75t_R _24861_ (.A1(_02126_),
    .A2(_02127_),
    .B(_01770_),
    .Y(_02128_));
 OAI21x1_ASAP7_75t_R _24862_ (.A1(_02125_),
    .A2(_02128_),
    .B(_01644_),
    .Y(_02129_));
 AOI21x1_ASAP7_75t_R _24863_ (.A1(_01668_),
    .A2(_01667_),
    .B(_01781_),
    .Y(_02130_));
 OA21x2_ASAP7_75t_R _24864_ (.A1(_01731_),
    .A2(_02071_),
    .B(_01621_),
    .Y(_02131_));
 OAI21x1_ASAP7_75t_R _24865_ (.A1(_02130_),
    .A2(_02131_),
    .B(_01591_),
    .Y(_02132_));
 INVx1_ASAP7_75t_R _24866_ (.A(_01692_),
    .Y(_02133_));
 NOR2x1_ASAP7_75t_R _24867_ (.A(_01611_),
    .B(_01930_),
    .Y(_02134_));
 OAI21x1_ASAP7_75t_R _24868_ (.A1(_01868_),
    .A2(_02133_),
    .B(_02134_),
    .Y(_02135_));
 AOI21x1_ASAP7_75t_R _24869_ (.A1(_02132_),
    .A2(_02135_),
    .B(_01770_),
    .Y(_02136_));
 OAI22x1_ASAP7_75t_R _24870_ (.A1(_02113_),
    .A2(_02119_),
    .B1(_02129_),
    .B2(_02136_),
    .Y(_02137_));
 AOI21x1_ASAP7_75t_R _24871_ (.A1(_01811_),
    .A2(_01584_),
    .B(_01635_),
    .Y(_02138_));
 OAI21x1_ASAP7_75t_R _24872_ (.A1(_01691_),
    .A2(_01692_),
    .B(_02138_),
    .Y(_02139_));
 AOI21x1_ASAP7_75t_R _24873_ (.A1(_01802_),
    .A2(_01620_),
    .B(_01816_),
    .Y(_02140_));
 AOI21x1_ASAP7_75t_R _24874_ (.A1(_02140_),
    .A2(_02054_),
    .B(_01734_),
    .Y(_02141_));
 NAND2x1_ASAP7_75t_R _24875_ (.A(_02139_),
    .B(_02141_),
    .Y(_02142_));
 NAND2x2_ASAP7_75t_R _24876_ (.A(_01663_),
    .B(_01662_),
    .Y(_02143_));
 NAND2x1_ASAP7_75t_R _24877_ (.A(_01772_),
    .B(_01632_),
    .Y(_02144_));
 AOI21x1_ASAP7_75t_R _24878_ (.A1(_02143_),
    .A2(_02144_),
    .B(_01789_),
    .Y(_02145_));
 NAND2x1_ASAP7_75t_R _24879_ (.A(net70),
    .B(_01621_),
    .Y(_02146_));
 AOI21x1_ASAP7_75t_R _24880_ (.A1(_02146_),
    .A2(_01969_),
    .B(_01764_),
    .Y(_02147_));
 OAI21x1_ASAP7_75t_R _24881_ (.A1(_01591_),
    .A2(_02145_),
    .B(_02147_),
    .Y(_02148_));
 AOI21x1_ASAP7_75t_R _24882_ (.A1(_02142_),
    .A2(_02148_),
    .B(_01644_),
    .Y(_02149_));
 NAND2x1_ASAP7_75t_R _24883_ (.A(_01653_),
    .B(_01789_),
    .Y(_02150_));
 OAI21x1_ASAP7_75t_R _24884_ (.A1(_02058_),
    .A2(_01731_),
    .B(_01634_),
    .Y(_02151_));
 AOI21x1_ASAP7_75t_R _24885_ (.A1(_02150_),
    .A2(_02151_),
    .B(_01791_),
    .Y(_02152_));
 NAND2x1_ASAP7_75t_R _24886_ (.A(_00568_),
    .B(_01772_),
    .Y(_02153_));
 AOI21x1_ASAP7_75t_R _24887_ (.A1(_02153_),
    .A2(_02101_),
    .B(_01867_),
    .Y(_02154_));
 OAI21x1_ASAP7_75t_R _24888_ (.A1(_02152_),
    .A2(_02154_),
    .B(_01609_),
    .Y(_02155_));
 AOI21x1_ASAP7_75t_R _24889_ (.A1(_15930_),
    .A2(_01753_),
    .B(_01723_),
    .Y(_02156_));
 AOI21x1_ASAP7_75t_R _24890_ (.A1(_01775_),
    .A2(_02156_),
    .B(_01867_),
    .Y(_02157_));
 AOI21x1_ASAP7_75t_R _24891_ (.A1(_01756_),
    .A2(_01994_),
    .B(_01591_),
    .Y(_02158_));
 OAI21x1_ASAP7_75t_R _24892_ (.A1(_02157_),
    .A2(_02158_),
    .B(_01770_),
    .Y(_02159_));
 AOI21x1_ASAP7_75t_R _24893_ (.A1(_02155_),
    .A2(_02159_),
    .B(_01769_),
    .Y(_02160_));
 OAI21x1_ASAP7_75t_R _24894_ (.A1(_02149_),
    .A2(_02160_),
    .B(_01710_),
    .Y(_02161_));
 OAI21x1_ASAP7_75t_R _24895_ (.A1(_01710_),
    .A2(_02137_),
    .B(_02161_),
    .Y(_00094_));
 OAI21x1_ASAP7_75t_R _24896_ (.A1(_15925_),
    .A2(_01775_),
    .B(_02026_),
    .Y(_02162_));
 AND2x2_ASAP7_75t_R _24897_ (.A(_01881_),
    .B(_01791_),
    .Y(_02163_));
 NAND2x1_ASAP7_75t_R _24898_ (.A(_01653_),
    .B(_01932_),
    .Y(_02164_));
 NOR2x1_ASAP7_75t_R _24899_ (.A(_15930_),
    .B(_01650_),
    .Y(_02165_));
 OA21x2_ASAP7_75t_R _24900_ (.A1(_02164_),
    .A2(_02165_),
    .B(_01671_),
    .Y(_02166_));
 AOI22x1_ASAP7_75t_R _24901_ (.A1(_02162_),
    .A2(_01690_),
    .B1(_02163_),
    .B2(_02166_),
    .Y(_02167_));
 NOR3x1_ASAP7_75t_R _24902_ (.A(_01844_),
    .B(_01867_),
    .C(_01930_),
    .Y(_02168_));
 NOR2x1_ASAP7_75t_R _24903_ (.A(_01919_),
    .B(_02165_),
    .Y(_02169_));
 AO21x1_ASAP7_75t_R _24904_ (.A1(_01762_),
    .A2(_01634_),
    .B(_01611_),
    .Y(_02170_));
 NOR2x1_ASAP7_75t_R _24905_ (.A(_02169_),
    .B(_02170_),
    .Y(_02171_));
 OAI21x1_ASAP7_75t_R _24906_ (.A1(_02168_),
    .A2(_02171_),
    .B(_01770_),
    .Y(_02172_));
 AOI21x1_ASAP7_75t_R _24907_ (.A1(_02167_),
    .A2(_02172_),
    .B(_01769_),
    .Y(_02173_));
 NOR2x1_ASAP7_75t_R _24908_ (.A(_01691_),
    .B(_01887_),
    .Y(_02174_));
 OAI21x1_ASAP7_75t_R _24909_ (.A1(_02174_),
    .A2(_02107_),
    .B(_01591_),
    .Y(_02175_));
 AND2x2_ASAP7_75t_R _24910_ (.A(_01832_),
    .B(_01634_),
    .Y(_02176_));
 OAI21x1_ASAP7_75t_R _24911_ (.A1(_02176_),
    .A2(_01942_),
    .B(_01867_),
    .Y(_02177_));
 AOI21x1_ASAP7_75t_R _24912_ (.A1(_02175_),
    .A2(_02177_),
    .B(_01609_),
    .Y(_02178_));
 NAND2x1_ASAP7_75t_R _24913_ (.A(_02143_),
    .B(_01994_),
    .Y(_02179_));
 OAI21x1_ASAP7_75t_R _24914_ (.A1(_01867_),
    .A2(_02179_),
    .B(_01609_),
    .Y(_02180_));
 OA21x2_ASAP7_75t_R _24915_ (.A1(_01617_),
    .A2(_01788_),
    .B(_01634_),
    .Y(_02181_));
 AO21x1_ASAP7_75t_R _24916_ (.A1(_01677_),
    .A2(_01762_),
    .B(_01611_),
    .Y(_02182_));
 NOR2x1_ASAP7_75t_R _24917_ (.A(_02181_),
    .B(_02182_),
    .Y(_02183_));
 OAI21x1_ASAP7_75t_R _24918_ (.A1(_02180_),
    .A2(_02183_),
    .B(_01769_),
    .Y(_02184_));
 OAI21x1_ASAP7_75t_R _24919_ (.A1(_02178_),
    .A2(_02184_),
    .B(_01710_),
    .Y(_02185_));
 AO21x1_ASAP7_75t_R _24920_ (.A1(_01648_),
    .A2(_15923_),
    .B(_01880_),
    .Y(_02186_));
 AND3x1_ASAP7_75t_R _24921_ (.A(_02186_),
    .B(_01952_),
    .C(_01582_),
    .Y(_02187_));
 AOI21x1_ASAP7_75t_R _24922_ (.A1(_01550_),
    .A2(_01732_),
    .B(_01750_),
    .Y(_02188_));
 OR3x1_ASAP7_75t_R _24923_ (.A(_01617_),
    .B(_01811_),
    .C(_01788_),
    .Y(_02189_));
 AOI21x1_ASAP7_75t_R _24924_ (.A1(_02188_),
    .A2(_02189_),
    .B(_01690_),
    .Y(_02190_));
 OA21x2_ASAP7_75t_R _24925_ (.A1(_01880_),
    .A2(_01208_),
    .B(_01816_),
    .Y(_02191_));
 OAI21x1_ASAP7_75t_R _24926_ (.A1(_01959_),
    .A2(_01887_),
    .B(_02191_),
    .Y(_02192_));
 AOI21x1_ASAP7_75t_R _24927_ (.A1(net70),
    .A2(_01826_),
    .B(_01788_),
    .Y(_02193_));
 AOI21x1_ASAP7_75t_R _24928_ (.A1(_01742_),
    .A2(_02193_),
    .B(_01671_),
    .Y(_02194_));
 AOI21x1_ASAP7_75t_R _24929_ (.A1(_02192_),
    .A2(_02194_),
    .B(_01643_),
    .Y(_02195_));
 OAI21x1_ASAP7_75t_R _24930_ (.A1(_02187_),
    .A2(_02190_),
    .B(_02195_),
    .Y(_02196_));
 NOR2x1_ASAP7_75t_R _24931_ (.A(_01771_),
    .B(_01941_),
    .Y(_02197_));
 AO21x1_ASAP7_75t_R _24932_ (.A1(_01984_),
    .A2(_01525_),
    .B(_01611_),
    .Y(_02198_));
 NOR2x1_ASAP7_75t_R _24933_ (.A(_01213_),
    .B(_01613_),
    .Y(_02199_));
 NOR2x1_ASAP7_75t_R _24934_ (.A(_02199_),
    .B(_01729_),
    .Y(_02200_));
 AOI21x1_ASAP7_75t_R _24935_ (.A1(_02120_),
    .A2(_02200_),
    .B(_01671_),
    .Y(_02201_));
 OAI21x1_ASAP7_75t_R _24936_ (.A1(_02197_),
    .A2(_02198_),
    .B(_02201_),
    .Y(_02202_));
 NAND2x1_ASAP7_75t_R _24937_ (.A(_00567_),
    .B(_01811_),
    .Y(_02203_));
 AOI21x1_ASAP7_75t_R _24938_ (.A1(_02203_),
    .A2(_01742_),
    .B(_01764_),
    .Y(_02204_));
 AO21x1_ASAP7_75t_R _24939_ (.A1(_01626_),
    .A2(_15923_),
    .B(_01880_),
    .Y(_02205_));
 NAND2x1_ASAP7_75t_R _24940_ (.A(_02205_),
    .B(_01852_),
    .Y(_02206_));
 AOI21x1_ASAP7_75t_R _24941_ (.A1(_02204_),
    .A2(_02206_),
    .B(_01716_),
    .Y(_02207_));
 AOI21x1_ASAP7_75t_R _24942_ (.A1(_02202_),
    .A2(_02207_),
    .B(_01709_),
    .Y(_02208_));
 NAND2x1_ASAP7_75t_R _24943_ (.A(_02196_),
    .B(_02208_),
    .Y(_02209_));
 OAI21x1_ASAP7_75t_R _24944_ (.A1(_02173_),
    .A2(_02185_),
    .B(_02209_),
    .Y(_00095_));
 NOR2x1_ASAP7_75t_R _24945_ (.A(_10621_),
    .B(_00569_),
    .Y(_02210_));
 XOR2x2_ASAP7_75t_R _24946_ (.A(_10651_),
    .B(_10822_),
    .Y(_02211_));
 XOR2x1_ASAP7_75t_R _24947_ (.A(_10632_),
    .Y(_02212_),
    .B(_02211_));
 XOR2x1_ASAP7_75t_R _24948_ (.A(_10679_),
    .Y(_02213_),
    .B(_13584_));
 NAND2x1_ASAP7_75t_R _24949_ (.A(_02213_),
    .B(_02212_),
    .Y(_02214_));
 XOR2x1_ASAP7_75t_R _24950_ (.A(_10624_),
    .Y(_02215_),
    .B(_02211_));
 XOR2x1_ASAP7_75t_R _24951_ (.A(_10677_),
    .Y(_02216_),
    .B(_13584_));
 NAND2x1_ASAP7_75t_R _24952_ (.A(_02216_),
    .B(_02215_),
    .Y(_02217_));
 AOI21x1_ASAP7_75t_R _24953_ (.A1(_02214_),
    .A2(_02217_),
    .B(_12160_),
    .Y(_02218_));
 INVx1_ASAP7_75t_R _24954_ (.A(_08101_),
    .Y(_02219_));
 OAI21x1_ASAP7_75t_R _24955_ (.A1(_02210_),
    .A2(_02218_),
    .B(_02219_),
    .Y(_02220_));
 AND2x2_ASAP7_75t_R _24956_ (.A(_10643_),
    .B(_00569_),
    .Y(_02221_));
 NAND2x1_ASAP7_75t_R _24957_ (.A(_02215_),
    .B(_02213_),
    .Y(_02222_));
 NAND2x1_ASAP7_75t_R _24958_ (.A(_02212_),
    .B(_02216_),
    .Y(_02223_));
 AOI21x1_ASAP7_75t_R _24959_ (.A1(_02222_),
    .A2(_02223_),
    .B(_12160_),
    .Y(_02224_));
 OAI21x1_ASAP7_75t_R _24960_ (.A1(_02221_),
    .A2(_02224_),
    .B(_08101_),
    .Y(_02225_));
 NAND2x2_ASAP7_75t_R _24961_ (.A(_02220_),
    .B(_02225_),
    .Y(_02226_));
 CKINVDCx9p33_ASAP7_75t_R _24962_ (.A(net547),
    .Y(_15940_));
 NOR2x1_ASAP7_75t_R _24963_ (.A(_10723_),
    .B(_00570_),
    .Y(_02227_));
 INVx1_ASAP7_75t_R _24964_ (.A(_02227_),
    .Y(_02228_));
 INVx1_ASAP7_75t_R _24965_ (.A(_10826_),
    .Y(_02229_));
 XOR2x1_ASAP7_75t_R _24966_ (.A(_10634_),
    .Y(_02230_),
    .B(_10658_));
 NAND2x1_ASAP7_75t_R _24967_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 XNOR2x1_ASAP7_75t_R _24968_ (.B(_10658_),
    .Y(_02232_),
    .A(_10634_));
 NAND2x1_ASAP7_75t_R _24969_ (.A(_10826_),
    .B(_02232_),
    .Y(_02233_));
 INVx1_ASAP7_75t_R _24970_ (.A(_02211_),
    .Y(_02234_));
 AOI21x1_ASAP7_75t_R _24971_ (.A1(_02231_),
    .A2(_02233_),
    .B(_02234_),
    .Y(_02235_));
 XOR2x1_ASAP7_75t_R _24972_ (.A(net49),
    .Y(_02236_),
    .B(net761));
 NAND2x1_ASAP7_75t_R _24973_ (.A(net25),
    .B(_02236_),
    .Y(_02237_));
 XNOR2x1_ASAP7_75t_R _24974_ (.B(net761),
    .Y(_02238_),
    .A(_10658_));
 NAND2x1_ASAP7_75t_R _24975_ (.A(_13604_),
    .B(_02238_),
    .Y(_02239_));
 AOI21x1_ASAP7_75t_R _24976_ (.A1(_02237_),
    .A2(_02239_),
    .B(_02211_),
    .Y(_02240_));
 OAI21x1_ASAP7_75t_R _24977_ (.A1(_02235_),
    .A2(_02240_),
    .B(_10763_),
    .Y(_02241_));
 NAND2x1_ASAP7_75t_R _24978_ (.A(_02241_),
    .B(_02228_),
    .Y(_02242_));
 XNOR2x2_ASAP7_75t_R _24979_ (.A(_01025_),
    .B(_02242_),
    .Y(_02243_));
 BUFx12_ASAP7_75t_R _24980_ (.A(_02243_),
    .Y(_15943_));
 NOR2x2_ASAP7_75t_R _24981_ (.A(net668),
    .B(_00572_),
    .Y(_02244_));
 INVx2_ASAP7_75t_R _24982_ (.A(_02244_),
    .Y(_02245_));
 XOR2x2_ASAP7_75t_R _24983_ (.A(_10711_),
    .B(_00766_),
    .Y(_02246_));
 XOR2x1_ASAP7_75t_R _24984_ (.A(_02246_),
    .Y(_02247_),
    .B(_10682_));
 NOR2x1_ASAP7_75t_R _24985_ (.A(net613),
    .B(_02247_),
    .Y(_02248_));
 XNOR2x1_ASAP7_75t_R _24986_ (.B(_10624_),
    .Y(_02249_),
    .A(_10628_));
 INVx2_ASAP7_75t_R _24987_ (.A(_10682_),
    .Y(_02250_));
 XOR2x1_ASAP7_75t_R _24988_ (.A(_02246_),
    .Y(_02251_),
    .B(_02250_));
 NOR2x1_ASAP7_75t_R _24989_ (.A(_02249_),
    .B(_02251_),
    .Y(_02252_));
 OAI21x1_ASAP7_75t_R _24990_ (.A1(_02248_),
    .A2(_02252_),
    .B(net650),
    .Y(_02253_));
 INVx2_ASAP7_75t_R _24991_ (.A(_08106_),
    .Y(_02254_));
 AOI21x1_ASAP7_75t_R _24992_ (.A1(_02245_),
    .A2(_02253_),
    .B(_02254_),
    .Y(_02255_));
 NAND2x2_ASAP7_75t_R _24993_ (.A(_00572_),
    .B(_11373_),
    .Y(_02256_));
 NAND2x2_ASAP7_75t_R _24994_ (.A(_02250_),
    .B(net612),
    .Y(_02257_));
 INVx3_ASAP7_75t_R _24995_ (.A(_02246_),
    .Y(_02258_));
 NOR2x1_ASAP7_75t_R _24996_ (.A(_10628_),
    .B(_10624_),
    .Y(_02259_));
 AND2x2_ASAP7_75t_R _24997_ (.A(_10628_),
    .B(_10624_),
    .Y(_02260_));
 OAI21x1_ASAP7_75t_R _24998_ (.A1(_02259_),
    .A2(_02260_),
    .B(_10682_),
    .Y(_02261_));
 NAND3x2_ASAP7_75t_R _24999_ (.B(_02258_),
    .C(_02261_),
    .Y(_02262_),
    .A(_02257_));
 NOR2x1_ASAP7_75t_R _25000_ (.A(_02250_),
    .B(net612),
    .Y(_02263_));
 NOR2x1_ASAP7_75t_R _25001_ (.A(_10682_),
    .B(_02249_),
    .Y(_02264_));
 OAI21x1_ASAP7_75t_R _25002_ (.A1(_02263_),
    .A2(_02264_),
    .B(_02246_),
    .Y(_02265_));
 NAND3x2_ASAP7_75t_R _25003_ (.B(net650),
    .C(_02265_),
    .Y(_02266_),
    .A(_02262_));
 AOI21x1_ASAP7_75t_R _25004_ (.A1(_02256_),
    .A2(_02266_),
    .B(_08106_),
    .Y(_02267_));
 NOR2x2_ASAP7_75t_R _25005_ (.A(_02255_),
    .B(_02267_),
    .Y(_02268_));
 BUFx10_ASAP7_75t_R _25006_ (.A(_02268_),
    .Y(_15951_));
 BUFx6f_ASAP7_75t_R _25007_ (.A(_02226_),
    .Y(_15938_));
 AOI21x1_ASAP7_75t_R _25008_ (.A1(_02245_),
    .A2(_02253_),
    .B(_08106_),
    .Y(_02269_));
 AOI21x1_ASAP7_75t_R _25009_ (.A1(_02256_),
    .A2(_02266_),
    .B(_02254_),
    .Y(_02270_));
 NOR2x2_ASAP7_75t_R _25010_ (.A(_02269_),
    .B(_02270_),
    .Y(_02271_));
 BUFx12f_ASAP7_75t_R _25011_ (.A(_02271_),
    .Y(_02272_));
 BUFx6f_ASAP7_75t_R _25012_ (.A(_02272_),
    .Y(_15948_));
 XOR2x2_ASAP7_75t_R _25013_ (.A(_01025_),
    .B(_02242_),
    .Y(_02273_));
 XNOR2x1_ASAP7_75t_R _25014_ (.B(_13656_),
    .Y(_02274_),
    .A(_10715_));
 XNOR2x2_ASAP7_75t_R _25015_ (.A(_10682_),
    .B(_10822_),
    .Y(_02275_));
 XOR2x2_ASAP7_75t_R _25016_ (.A(_00735_),
    .B(_10710_),
    .Y(_02276_));
 XOR2x1_ASAP7_75t_R _25017_ (.A(_02275_),
    .Y(_02277_),
    .B(_02276_));
 NOR2x1_ASAP7_75t_R _25018_ (.A(_02274_),
    .B(_02277_),
    .Y(_02278_));
 XOR2x1_ASAP7_75t_R _25019_ (.A(_13656_),
    .Y(_02279_),
    .B(_10715_));
 XNOR2x1_ASAP7_75t_R _25020_ (.B(_02275_),
    .Y(_02280_),
    .A(_02276_));
 OAI21x1_ASAP7_75t_R _25021_ (.A1(_02279_),
    .A2(_02280_),
    .B(_12921_),
    .Y(_02281_));
 NAND2x1_ASAP7_75t_R _25022_ (.A(_00720_),
    .B(_10689_),
    .Y(_02282_));
 OAI21x1_ASAP7_75t_R _25023_ (.A1(_02278_),
    .A2(_02281_),
    .B(_02282_),
    .Y(_02283_));
 XNOR2x2_ASAP7_75t_R _25024_ (.A(_00997_),
    .B(_02283_),
    .Y(_02284_));
 BUFx6f_ASAP7_75t_R _25025_ (.A(_02284_),
    .Y(_02285_));
 OAI21x1_ASAP7_75t_R _25026_ (.A1(net530),
    .A2(_02268_),
    .B(_02285_),
    .Y(_02286_));
 AOI21x1_ASAP7_75t_R _25027_ (.A1(_02220_),
    .A2(_02225_),
    .B(_02243_),
    .Y(_02287_));
 NOR2x1_ASAP7_75t_R _25028_ (.A(_02286_),
    .B(_02287_),
    .Y(_02288_));
 NAND2x2_ASAP7_75t_R _25029_ (.A(net531),
    .B(_15938_),
    .Y(_02289_));
 BUFx10_ASAP7_75t_R _25030_ (.A(_02272_),
    .Y(_02290_));
 NAND2x1_ASAP7_75t_R _25031_ (.A(_15943_),
    .B(_02290_),
    .Y(_02291_));
 BUFx6f_ASAP7_75t_R _25032_ (.A(_02284_),
    .Y(_02292_));
 AOI21x1_ASAP7_75t_R _25033_ (.A1(_02289_),
    .A2(_02291_),
    .B(_02292_),
    .Y(_02293_));
 XOR2x2_ASAP7_75t_R _25034_ (.A(_10715_),
    .B(_10822_),
    .Y(_02294_));
 XOR2x1_ASAP7_75t_R _25035_ (.A(_10757_),
    .Y(_02295_),
    .B(_02294_));
 NAND2x1_ASAP7_75t_R _25036_ (.A(_13677_),
    .B(_02295_),
    .Y(_02296_));
 OA21x2_ASAP7_75t_R _25037_ (.A1(_02295_),
    .A2(_13677_),
    .B(net585),
    .Y(_02297_));
 AND2x2_ASAP7_75t_R _25038_ (.A(_10640_),
    .B(_00719_),
    .Y(_02298_));
 AOI21x1_ASAP7_75t_R _25039_ (.A1(_02296_),
    .A2(_02297_),
    .B(_02298_),
    .Y(_02299_));
 XNOR2x2_ASAP7_75t_R _25040_ (.A(_00998_),
    .B(_02299_),
    .Y(_02300_));
 BUFx6f_ASAP7_75t_R _25041_ (.A(_02300_),
    .Y(_02301_));
 OA21x2_ASAP7_75t_R _25042_ (.A1(_02288_),
    .A2(_02293_),
    .B(_02301_),
    .Y(_02302_));
 BUFx10_ASAP7_75t_R _25043_ (.A(_02268_),
    .Y(_02303_));
 NAND2x2_ASAP7_75t_R _25044_ (.A(net738),
    .B(_02303_),
    .Y(_02304_));
 INVx1_ASAP7_75t_R _25045_ (.A(_00574_),
    .Y(_02305_));
 OAI21x1_ASAP7_75t_R _25046_ (.A1(_02255_),
    .A2(_02267_),
    .B(_02305_),
    .Y(_02306_));
 BUFx3_ASAP7_75t_R _25047_ (.A(_02306_),
    .Y(_02307_));
 XOR2x2_ASAP7_75t_R _25048_ (.A(_02283_),
    .B(_00997_),
    .Y(_02308_));
 BUFx10_ASAP7_75t_R _25049_ (.A(_02308_),
    .Y(_02309_));
 BUFx6f_ASAP7_75t_R _25050_ (.A(_02309_),
    .Y(_02310_));
 AO21x1_ASAP7_75t_R _25051_ (.A1(_02304_),
    .A2(net73),
    .B(_02310_),
    .Y(_02311_));
 BUFx10_ASAP7_75t_R _25052_ (.A(_02268_),
    .Y(_02312_));
 NAND2x2_ASAP7_75t_R _25053_ (.A(net489),
    .B(_02312_),
    .Y(_02313_));
 NAND2x2_ASAP7_75t_R _25054_ (.A(_00571_),
    .B(_02272_),
    .Y(_02314_));
 BUFx4f_ASAP7_75t_R _25055_ (.A(_02285_),
    .Y(_02315_));
 AO21x1_ASAP7_75t_R _25056_ (.A1(_02313_),
    .A2(_02314_),
    .B(_02315_),
    .Y(_02316_));
 BUFx6f_ASAP7_75t_R _25057_ (.A(_02300_),
    .Y(_02317_));
 BUFx6f_ASAP7_75t_R _25058_ (.A(_02317_),
    .Y(_02318_));
 AOI21x1_ASAP7_75t_R _25059_ (.A1(_02311_),
    .A2(_02316_),
    .B(_02318_),
    .Y(_02319_));
 NOR2x1_ASAP7_75t_R _25060_ (.A(net650),
    .B(_00718_),
    .Y(_02320_));
 INVx1_ASAP7_75t_R _25061_ (.A(_02320_),
    .Y(_02321_));
 XOR2x1_ASAP7_75t_R _25062_ (.A(_10783_),
    .Y(_02322_),
    .B(_00769_));
 NAND2x1_ASAP7_75t_R _25063_ (.A(_13714_),
    .B(_02322_),
    .Y(_02323_));
 NAND2x1_ASAP7_75t_R _25064_ (.A(_10758_),
    .B(_10784_),
    .Y(_02324_));
 INVx1_ASAP7_75t_R _25065_ (.A(_10736_),
    .Y(_02325_));
 AOI21x1_ASAP7_75t_R _25066_ (.A1(_02323_),
    .A2(_02324_),
    .B(_02325_),
    .Y(_02326_));
 NAND2x1_ASAP7_75t_R _25067_ (.A(_10758_),
    .B(_02322_),
    .Y(_02327_));
 NAND2x1_ASAP7_75t_R _25068_ (.A(_13714_),
    .B(_10784_),
    .Y(_02328_));
 AOI21x1_ASAP7_75t_R _25069_ (.A1(_02327_),
    .A2(_02328_),
    .B(_10736_),
    .Y(_02329_));
 OAI21x1_ASAP7_75t_R _25070_ (.A1(_02326_),
    .A2(_02329_),
    .B(_12921_),
    .Y(_02330_));
 NAND2x1_ASAP7_75t_R _25071_ (.A(_02321_),
    .B(_02330_),
    .Y(_02331_));
 XNOR2x2_ASAP7_75t_R _25072_ (.A(_00999_),
    .B(_02331_),
    .Y(_02332_));
 BUFx6f_ASAP7_75t_R _25073_ (.A(_02332_),
    .Y(_02333_));
 OA21x2_ASAP7_75t_R _25074_ (.A1(_02302_),
    .A2(_02319_),
    .B(_02333_),
    .Y(_02334_));
 INVx1_ASAP7_75t_R _25075_ (.A(net489),
    .Y(_02335_));
 NAND2x2_ASAP7_75t_R _25076_ (.A(_02335_),
    .B(_02303_),
    .Y(_02336_));
 OAI21x1_ASAP7_75t_R _25077_ (.A1(_02255_),
    .A2(_02267_),
    .B(net457),
    .Y(_02337_));
 NAND2x2_ASAP7_75t_R _25078_ (.A(_02337_),
    .B(_02308_),
    .Y(_02338_));
 INVx2_ASAP7_75t_R _25079_ (.A(_02338_),
    .Y(_02339_));
 NAND2x1_ASAP7_75t_R _25080_ (.A(_02336_),
    .B(_02339_),
    .Y(_02340_));
 INVx2_ASAP7_75t_R _25081_ (.A(_00571_),
    .Y(_02341_));
 NOR2x2_ASAP7_75t_R _25082_ (.A(_02341_),
    .B(_02272_),
    .Y(_02342_));
 NAND2x1_ASAP7_75t_R _25083_ (.A(_02315_),
    .B(_02342_),
    .Y(_02343_));
 OAI21x1_ASAP7_75t_R _25084_ (.A1(_02255_),
    .A2(_02267_),
    .B(_00573_),
    .Y(_02344_));
 BUFx4f_ASAP7_75t_R _25085_ (.A(_02308_),
    .Y(_02345_));
 XOR2x2_ASAP7_75t_R _25086_ (.A(_02299_),
    .B(_00998_),
    .Y(_02346_));
 OA21x2_ASAP7_75t_R _25087_ (.A1(_02344_),
    .A2(_02345_),
    .B(_02346_),
    .Y(_02347_));
 NAND3x1_ASAP7_75t_R _25088_ (.A(_02340_),
    .B(_02343_),
    .C(_02347_),
    .Y(_02348_));
 BUFx6f_ASAP7_75t_R _25089_ (.A(_02317_),
    .Y(_02349_));
 BUFx6f_ASAP7_75t_R _25090_ (.A(_02284_),
    .Y(_02350_));
 BUFx6f_ASAP7_75t_R _25091_ (.A(_02350_),
    .Y(_02351_));
 OAI21x1_ASAP7_75t_R _25092_ (.A1(net57),
    .A2(_15948_),
    .B(_02307_),
    .Y(_02352_));
 OAI21x1_ASAP7_75t_R _25093_ (.A1(_02269_),
    .A2(_02270_),
    .B(net456),
    .Y(_02353_));
 NOR2x1_ASAP7_75t_R _25094_ (.A(_02292_),
    .B(_02353_),
    .Y(_02354_));
 AOI21x1_ASAP7_75t_R _25095_ (.A1(_02351_),
    .A2(_02352_),
    .B(_02354_),
    .Y(_02355_));
 BUFx6f_ASAP7_75t_R _25096_ (.A(_02332_),
    .Y(_02356_));
 AOI21x1_ASAP7_75t_R _25097_ (.A1(_02349_),
    .A2(_02355_),
    .B(_02356_),
    .Y(_02357_));
 XOR2x1_ASAP7_75t_R _25098_ (.A(_10758_),
    .Y(_02358_),
    .B(_00834_));
 XOR2x1_ASAP7_75t_R _25099_ (.A(_02358_),
    .Y(_02359_),
    .B(_00801_));
 XOR2x1_ASAP7_75t_R _25100_ (.A(_02359_),
    .Y(_02360_),
    .B(_10821_));
 NOR2x1_ASAP7_75t_R _25101_ (.A(_10829_),
    .B(_00717_),
    .Y(_02361_));
 AO21x1_ASAP7_75t_R _25102_ (.A1(_02360_),
    .A2(_11451_),
    .B(_02361_),
    .Y(_02362_));
 XOR2x2_ASAP7_75t_R _25103_ (.A(_02362_),
    .B(_01000_),
    .Y(_02363_));
 CKINVDCx8_ASAP7_75t_R _25104_ (.A(_02363_),
    .Y(_02364_));
 AO21x1_ASAP7_75t_R _25105_ (.A1(_02348_),
    .A2(_02357_),
    .B(_02364_),
    .Y(_02365_));
 BUFx16f_ASAP7_75t_R _25106_ (.A(_02273_),
    .Y(_15937_));
 AOI21x1_ASAP7_75t_R _25107_ (.A1(_15937_),
    .A2(_02312_),
    .B(_02285_),
    .Y(_02366_));
 INVx2_ASAP7_75t_R _25108_ (.A(_01218_),
    .Y(_02367_));
 NOR2x2_ASAP7_75t_R _25109_ (.A(_02367_),
    .B(_02268_),
    .Y(_02368_));
 INVx2_ASAP7_75t_R _25110_ (.A(_02368_),
    .Y(_02369_));
 NAND2x1_ASAP7_75t_R _25111_ (.A(_02366_),
    .B(_02369_),
    .Y(_02370_));
 NAND2x2_ASAP7_75t_R _25112_ (.A(_02271_),
    .B(net546),
    .Y(_02371_));
 BUFx6f_ASAP7_75t_R _25113_ (.A(_02371_),
    .Y(_02372_));
 INVx5_ASAP7_75t_R _25114_ (.A(_00576_),
    .Y(_02373_));
 AOI21x1_ASAP7_75t_R _25115_ (.A1(_02373_),
    .A2(_02312_),
    .B(_02309_),
    .Y(_02374_));
 BUFx6f_ASAP7_75t_R _25116_ (.A(_02346_),
    .Y(_02375_));
 AOI21x1_ASAP7_75t_R _25117_ (.A1(_02372_),
    .A2(_02374_),
    .B(_02375_),
    .Y(_02376_));
 AOI21x1_ASAP7_75t_R _25118_ (.A1(_02370_),
    .A2(_02376_),
    .B(_02332_),
    .Y(_02377_));
 INVx3_ASAP7_75t_R _25119_ (.A(_00575_),
    .Y(_02378_));
 OAI21x1_ASAP7_75t_R _25120_ (.A1(_02255_),
    .A2(_02267_),
    .B(_02378_),
    .Y(_02379_));
 NAND2x1_ASAP7_75t_R _25121_ (.A(_02379_),
    .B(_02366_),
    .Y(_02380_));
 BUFx10_ASAP7_75t_R _25122_ (.A(_02308_),
    .Y(_02381_));
 INVx1_ASAP7_75t_R _25123_ (.A(_01215_),
    .Y(_02382_));
 OAI21x1_ASAP7_75t_R _25124_ (.A1(_02255_),
    .A2(_02267_),
    .B(_02382_),
    .Y(_02383_));
 OAI21x1_ASAP7_75t_R _25125_ (.A1(_02381_),
    .A2(_02383_),
    .B(_02346_),
    .Y(_02384_));
 NAND2x2_ASAP7_75t_R _25126_ (.A(_02268_),
    .B(net548),
    .Y(_02385_));
 NOR2x2_ASAP7_75t_R _25127_ (.A(_02309_),
    .B(_02385_),
    .Y(_02386_));
 NOR2x1_ASAP7_75t_R _25128_ (.A(_02384_),
    .B(_02386_),
    .Y(_02387_));
 NAND2x1_ASAP7_75t_R _25129_ (.A(_02380_),
    .B(_02387_),
    .Y(_02388_));
 NAND2x1_ASAP7_75t_R _25130_ (.A(_02377_),
    .B(_02388_),
    .Y(_02389_));
 NAND2x1_ASAP7_75t_R _25131_ (.A(_02373_),
    .B(_02303_),
    .Y(_02390_));
 BUFx3_ASAP7_75t_R _25132_ (.A(_01216_),
    .Y(_02391_));
 AOI21x1_ASAP7_75t_R _25133_ (.A1(_02391_),
    .A2(_02290_),
    .B(_02350_),
    .Y(_02392_));
 NAND2x1_ASAP7_75t_R _25134_ (.A(_02390_),
    .B(_02392_),
    .Y(_02393_));
 BUFx6f_ASAP7_75t_R _25135_ (.A(_02300_),
    .Y(_02394_));
 AOI21x1_ASAP7_75t_R _25136_ (.A1(_15937_),
    .A2(_02303_),
    .B(_02309_),
    .Y(_02395_));
 NOR2x1_ASAP7_75t_R _25137_ (.A(_02394_),
    .B(_02395_),
    .Y(_02396_));
 INVx1_ASAP7_75t_R _25138_ (.A(_02332_),
    .Y(_02397_));
 BUFx6f_ASAP7_75t_R _25139_ (.A(_02397_),
    .Y(_02398_));
 BUFx6f_ASAP7_75t_R _25140_ (.A(_02398_),
    .Y(_02399_));
 AOI21x1_ASAP7_75t_R _25141_ (.A1(_02393_),
    .A2(_02396_),
    .B(_02399_),
    .Y(_02400_));
 INVx2_ASAP7_75t_R _25142_ (.A(_02337_),
    .Y(_02401_));
 AO21x1_ASAP7_75t_R _25143_ (.A1(_02312_),
    .A2(_01218_),
    .B(_02285_),
    .Y(_02402_));
 BUFx4f_ASAP7_75t_R _25144_ (.A(_02402_),
    .Y(_02403_));
 NAND2x2_ASAP7_75t_R _25145_ (.A(net530),
    .B(_02272_),
    .Y(_02404_));
 BUFx6f_ASAP7_75t_R _25146_ (.A(_02346_),
    .Y(_02405_));
 AOI21x1_ASAP7_75t_R _25147_ (.A1(_02404_),
    .A2(_02374_),
    .B(_02405_),
    .Y(_02406_));
 OAI21x1_ASAP7_75t_R _25148_ (.A1(_02401_),
    .A2(_02403_),
    .B(_02406_),
    .Y(_02407_));
 AOI21x1_ASAP7_75t_R _25149_ (.A1(_02400_),
    .A2(_02407_),
    .B(_02363_),
    .Y(_02408_));
 XOR2x1_ASAP7_75t_R _25150_ (.A(_13758_),
    .Y(_02409_),
    .B(_10823_));
 XOR2x1_ASAP7_75t_R _25151_ (.A(_02409_),
    .Y(_02410_),
    .B(_10654_));
 NOR2x1_ASAP7_75t_R _25152_ (.A(_10831_),
    .B(_00716_),
    .Y(_02411_));
 AO21x1_ASAP7_75t_R _25153_ (.A1(_02410_),
    .A2(_10830_),
    .B(_02411_),
    .Y(_02412_));
 XOR2x2_ASAP7_75t_R _25154_ (.A(_02412_),
    .B(_01001_),
    .Y(_02413_));
 CKINVDCx5p33_ASAP7_75t_R _25155_ (.A(_02413_),
    .Y(_02414_));
 AOI21x1_ASAP7_75t_R _25156_ (.A1(_02389_),
    .A2(_02408_),
    .B(_02414_),
    .Y(_02415_));
 OAI21x1_ASAP7_75t_R _25157_ (.A1(_02334_),
    .A2(_02365_),
    .B(_02415_),
    .Y(_02416_));
 AOI21x1_ASAP7_75t_R _25158_ (.A1(_02292_),
    .A2(_02342_),
    .B(_02375_),
    .Y(_02417_));
 INVx1_ASAP7_75t_R _25159_ (.A(_02417_),
    .Y(_02418_));
 BUFx6f_ASAP7_75t_R _25160_ (.A(_02309_),
    .Y(_02419_));
 INVx2_ASAP7_75t_R _25161_ (.A(_02383_),
    .Y(_02420_));
 NOR2x2_ASAP7_75t_R _25162_ (.A(_02373_),
    .B(_02268_),
    .Y(_02421_));
 NAND2x1_ASAP7_75t_R _25163_ (.A(_02285_),
    .B(_02421_),
    .Y(_02422_));
 INVx1_ASAP7_75t_R _25164_ (.A(_02422_),
    .Y(_02423_));
 AO21x1_ASAP7_75t_R _25165_ (.A1(_02419_),
    .A2(_02420_),
    .B(_02423_),
    .Y(_02424_));
 INVx1_ASAP7_75t_R _25166_ (.A(_02384_),
    .Y(_02425_));
 NAND2x2_ASAP7_75t_R _25167_ (.A(_02373_),
    .B(_02272_),
    .Y(_02426_));
 AOI21x1_ASAP7_75t_R _25168_ (.A1(_01217_),
    .A2(_02312_),
    .B(_02285_),
    .Y(_02427_));
 NAND2x1_ASAP7_75t_R _25169_ (.A(_02426_),
    .B(_02427_),
    .Y(_02428_));
 AOI21x1_ASAP7_75t_R _25170_ (.A1(_02425_),
    .A2(_02428_),
    .B(_02398_),
    .Y(_02429_));
 OAI21x1_ASAP7_75t_R _25171_ (.A1(_02418_),
    .A2(_02424_),
    .B(_02429_),
    .Y(_02430_));
 OAI21x1_ASAP7_75t_R _25172_ (.A1(net623),
    .A2(_02290_),
    .B(_02344_),
    .Y(_02431_));
 OAI21x1_ASAP7_75t_R _25173_ (.A1(_02269_),
    .A2(_02270_),
    .B(_02382_),
    .Y(_02432_));
 NOR2x1_ASAP7_75t_R _25174_ (.A(_02381_),
    .B(_02432_),
    .Y(_02433_));
 AOI21x1_ASAP7_75t_R _25175_ (.A1(_02310_),
    .A2(_02431_),
    .B(_02433_),
    .Y(_02434_));
 INVx1_ASAP7_75t_R _25176_ (.A(_02391_),
    .Y(_02435_));
 OAI21x1_ASAP7_75t_R _25177_ (.A1(_02269_),
    .A2(_02270_),
    .B(_02435_),
    .Y(_02436_));
 OAI21x1_ASAP7_75t_R _25178_ (.A1(_02308_),
    .A2(_02436_),
    .B(_02346_),
    .Y(_02437_));
 INVx1_ASAP7_75t_R _25179_ (.A(_02437_),
    .Y(_02438_));
 NAND2x1_ASAP7_75t_R _25180_ (.A(_02438_),
    .B(_02422_),
    .Y(_02439_));
 INVx1_ASAP7_75t_R _25181_ (.A(_02439_),
    .Y(_02440_));
 NAND2x1_ASAP7_75t_R _25182_ (.A(_02434_),
    .B(_02440_),
    .Y(_02441_));
 AOI21x1_ASAP7_75t_R _25183_ (.A1(_02265_),
    .A2(_02262_),
    .B(_12161_),
    .Y(_02442_));
 OAI21x1_ASAP7_75t_R _25184_ (.A1(_02244_),
    .A2(_02442_),
    .B(_02254_),
    .Y(_02443_));
 NAND3x1_ASAP7_75t_R _25185_ (.A(_02253_),
    .B(_08106_),
    .C(_02245_),
    .Y(_02444_));
 AOI21x1_ASAP7_75t_R _25186_ (.A1(_02443_),
    .A2(_02444_),
    .B(net457),
    .Y(_02445_));
 NOR2x1_ASAP7_75t_R _25187_ (.A(_01220_),
    .B(_02285_),
    .Y(_02446_));
 AO21x1_ASAP7_75t_R _25188_ (.A1(net463),
    .A2(_02350_),
    .B(_02446_),
    .Y(_02447_));
 OA21x2_ASAP7_75t_R _25189_ (.A1(_02447_),
    .A2(_02375_),
    .B(_02398_),
    .Y(_02448_));
 AOI21x1_ASAP7_75t_R _25190_ (.A1(_02441_),
    .A2(_02448_),
    .B(_02364_),
    .Y(_02449_));
 NAND2x1_ASAP7_75t_R _25191_ (.A(_02430_),
    .B(_02449_),
    .Y(_02450_));
 NOR2x2_ASAP7_75t_R _25192_ (.A(_02381_),
    .B(_02436_),
    .Y(_02451_));
 AO21x1_ASAP7_75t_R _25193_ (.A1(_02366_),
    .A2(_02379_),
    .B(_02394_),
    .Y(_02452_));
 INVx1_ASAP7_75t_R _25194_ (.A(_01217_),
    .Y(_02453_));
 OAI21x1_ASAP7_75t_R _25195_ (.A1(_02255_),
    .A2(_02267_),
    .B(_02453_),
    .Y(_02454_));
 AOI21x1_ASAP7_75t_R _25196_ (.A1(_02436_),
    .A2(_02454_),
    .B(_02381_),
    .Y(_02455_));
 NOR2x1_ASAP7_75t_R _25197_ (.A(_02339_),
    .B(_02455_),
    .Y(_02456_));
 AOI21x1_ASAP7_75t_R _25198_ (.A1(_02301_),
    .A2(_02456_),
    .B(_02332_),
    .Y(_02457_));
 OAI21x1_ASAP7_75t_R _25199_ (.A1(_02451_),
    .A2(_02452_),
    .B(_02457_),
    .Y(_02458_));
 NOR2x1_ASAP7_75t_R _25200_ (.A(_02375_),
    .B(_02392_),
    .Y(_02459_));
 BUFx6f_ASAP7_75t_R _25201_ (.A(_02308_),
    .Y(_02460_));
 AOI21x1_ASAP7_75t_R _25202_ (.A1(_02383_),
    .A2(_02313_),
    .B(_02460_),
    .Y(_02461_));
 INVx1_ASAP7_75t_R _25203_ (.A(_02461_),
    .Y(_02462_));
 AOI21x1_ASAP7_75t_R _25204_ (.A1(_02459_),
    .A2(_02462_),
    .B(_02398_),
    .Y(_02463_));
 AOI21x1_ASAP7_75t_R _25205_ (.A1(_02353_),
    .A2(_02372_),
    .B(_02460_),
    .Y(_02464_));
 INVx1_ASAP7_75t_R _25206_ (.A(_02464_),
    .Y(_02465_));
 NAND2x2_ASAP7_75t_R _25207_ (.A(_02341_),
    .B(_02312_),
    .Y(_02466_));
 OA21x2_ASAP7_75t_R _25208_ (.A1(_02303_),
    .A2(_15943_),
    .B(_02381_),
    .Y(_02467_));
 AOI21x1_ASAP7_75t_R _25209_ (.A1(_02466_),
    .A2(_02467_),
    .B(_02394_),
    .Y(_02468_));
 NAND2x1_ASAP7_75t_R _25210_ (.A(_02465_),
    .B(_02468_),
    .Y(_02469_));
 AOI21x1_ASAP7_75t_R _25211_ (.A1(_02463_),
    .A2(_02469_),
    .B(_02363_),
    .Y(_02470_));
 BUFx10_ASAP7_75t_R _25212_ (.A(_02413_),
    .Y(_02471_));
 AOI21x1_ASAP7_75t_R _25213_ (.A1(_02458_),
    .A2(_02470_),
    .B(_02471_),
    .Y(_02472_));
 NAND2x1_ASAP7_75t_R _25214_ (.A(_02450_),
    .B(_02472_),
    .Y(_02473_));
 NAND2x1_ASAP7_75t_R _25215_ (.A(_02416_),
    .B(_02473_),
    .Y(_00096_));
 INVx3_ASAP7_75t_R _25216_ (.A(_02371_),
    .Y(_02474_));
 OR3x1_ASAP7_75t_R _25217_ (.A(_15951_),
    .B(_02378_),
    .C(_02310_),
    .Y(_02475_));
 OAI21x1_ASAP7_75t_R _25218_ (.A1(_02474_),
    .A2(_02403_),
    .B(_02475_),
    .Y(_02476_));
 BUFx6f_ASAP7_75t_R _25219_ (.A(_02375_),
    .Y(_02477_));
 NOR2x1_ASAP7_75t_R _25220_ (.A(_02391_),
    .B(_02345_),
    .Y(_02478_));
 AOI21x1_ASAP7_75t_R _25221_ (.A1(_15948_),
    .A2(_02478_),
    .B(_02301_),
    .Y(_02479_));
 AOI21x1_ASAP7_75t_R _25222_ (.A1(_02378_),
    .A2(_15951_),
    .B(_02350_),
    .Y(_02480_));
 NAND2x1_ASAP7_75t_R _25223_ (.A(net73),
    .B(_02480_),
    .Y(_02481_));
 BUFx6f_ASAP7_75t_R _25224_ (.A(_02398_),
    .Y(_02482_));
 AOI21x1_ASAP7_75t_R _25225_ (.A1(_02479_),
    .A2(_02481_),
    .B(_02482_),
    .Y(_02483_));
 OA21x2_ASAP7_75t_R _25226_ (.A1(_02476_),
    .A2(_02477_),
    .B(_02483_),
    .Y(_02484_));
 INVx3_ASAP7_75t_R _25227_ (.A(net463),
    .Y(_02485_));
 AOI21x1_ASAP7_75t_R _25228_ (.A1(net623),
    .A2(_15948_),
    .B(_02345_),
    .Y(_02486_));
 NAND2x1_ASAP7_75t_R _25229_ (.A(_02486_),
    .B(_02485_),
    .Y(_02487_));
 OAI21x1_ASAP7_75t_R _25230_ (.A1(_15940_),
    .A2(net623),
    .B(_02366_),
    .Y(_02488_));
 AOI21x1_ASAP7_75t_R _25231_ (.A1(_02487_),
    .A2(_02488_),
    .B(_02349_),
    .Y(_02489_));
 INVx4_ASAP7_75t_R _25232_ (.A(_02344_),
    .Y(_02490_));
 OAI21x1_ASAP7_75t_R _25233_ (.A1(_15937_),
    .A2(_02290_),
    .B(_02350_),
    .Y(_02491_));
 NOR2x1_ASAP7_75t_R _25234_ (.A(_02490_),
    .B(_02491_),
    .Y(_02492_));
 INVx2_ASAP7_75t_R _25235_ (.A(net739),
    .Y(_02493_));
 OAI21x1_ASAP7_75t_R _25236_ (.A1(_02493_),
    .A2(_02338_),
    .B(_02301_),
    .Y(_02494_));
 NOR2x1_ASAP7_75t_R _25237_ (.A(_02492_),
    .B(_02494_),
    .Y(_02495_));
 BUFx10_ASAP7_75t_R _25238_ (.A(_02398_),
    .Y(_02496_));
 OA21x2_ASAP7_75t_R _25239_ (.A1(_02489_),
    .A2(_02495_),
    .B(_02496_),
    .Y(_02497_));
 BUFx10_ASAP7_75t_R _25240_ (.A(_02364_),
    .Y(_02498_));
 OAI21x1_ASAP7_75t_R _25241_ (.A1(_02484_),
    .A2(_02497_),
    .B(_02498_),
    .Y(_02499_));
 NOR2x2_ASAP7_75t_R _25242_ (.A(_01218_),
    .B(_15951_),
    .Y(_02500_));
 OAI21x1_ASAP7_75t_R _25243_ (.A1(_02445_),
    .A2(_02500_),
    .B(_02419_),
    .Y(_02501_));
 BUFx4f_ASAP7_75t_R _25244_ (.A(_02350_),
    .Y(_02502_));
 OAI21x1_ASAP7_75t_R _25245_ (.A1(_02493_),
    .A2(_02421_),
    .B(_02502_),
    .Y(_02503_));
 AOI21x1_ASAP7_75t_R _25246_ (.A1(_02501_),
    .A2(_02503_),
    .B(_02318_),
    .Y(_02504_));
 INVx1_ASAP7_75t_R _25247_ (.A(_00578_),
    .Y(_02505_));
 NOR2x1_ASAP7_75t_R _25248_ (.A(_02505_),
    .B(_02350_),
    .Y(_02506_));
 NOR2x1_ASAP7_75t_R _25249_ (.A(_02506_),
    .B(_02451_),
    .Y(_02507_));
 NAND2x1_ASAP7_75t_R _25250_ (.A(_02502_),
    .B(_02474_),
    .Y(_02508_));
 BUFx6f_ASAP7_75t_R _25251_ (.A(_02346_),
    .Y(_02509_));
 AOI21x1_ASAP7_75t_R _25252_ (.A1(_02507_),
    .A2(_02508_),
    .B(_02509_),
    .Y(_02510_));
 OAI21x1_ASAP7_75t_R _25253_ (.A1(_02504_),
    .A2(_02510_),
    .B(_02496_),
    .Y(_02511_));
 INVx1_ASAP7_75t_R _25254_ (.A(_02366_),
    .Y(_02512_));
 NAND2x2_ASAP7_75t_R _25255_ (.A(_15943_),
    .B(_02312_),
    .Y(_02513_));
 AOI21x1_ASAP7_75t_R _25256_ (.A1(_02391_),
    .A2(_02290_),
    .B(_02309_),
    .Y(_02514_));
 AOI21x1_ASAP7_75t_R _25257_ (.A1(_02513_),
    .A2(_02514_),
    .B(_02405_),
    .Y(_02515_));
 OAI21x1_ASAP7_75t_R _25258_ (.A1(_02401_),
    .A2(_02512_),
    .B(_02515_),
    .Y(_02516_));
 NAND2x2_ASAP7_75t_R _25259_ (.A(net685),
    .B(_02312_),
    .Y(_02517_));
 OA21x2_ASAP7_75t_R _25260_ (.A1(_02517_),
    .A2(_02292_),
    .B(_02375_),
    .Y(_02518_));
 OA21x2_ASAP7_75t_R _25261_ (.A1(net57),
    .A2(_02303_),
    .B(_02350_),
    .Y(_02519_));
 NAND2x1_ASAP7_75t_R _25262_ (.A(_02289_),
    .B(_02519_),
    .Y(_02520_));
 AOI21x1_ASAP7_75t_R _25263_ (.A1(_02518_),
    .A2(_02520_),
    .B(_02399_),
    .Y(_02521_));
 NAND2x1_ASAP7_75t_R _25264_ (.A(_02516_),
    .B(_02521_),
    .Y(_02522_));
 AOI21x1_ASAP7_75t_R _25265_ (.A1(_02511_),
    .A2(_02522_),
    .B(_02498_),
    .Y(_02523_));
 NOR2x1_ASAP7_75t_R _25266_ (.A(_02471_),
    .B(_02523_),
    .Y(_02524_));
 AOI21x1_ASAP7_75t_R _25267_ (.A1(_15943_),
    .A2(_02290_),
    .B(_02381_),
    .Y(_02525_));
 AND2x2_ASAP7_75t_R _25268_ (.A(_02392_),
    .B(_02385_),
    .Y(_02526_));
 BUFx6f_ASAP7_75t_R _25269_ (.A(_02300_),
    .Y(_02527_));
 BUFx10_ASAP7_75t_R _25270_ (.A(_02527_),
    .Y(_02528_));
 AOI211x1_ASAP7_75t_R _25271_ (.A1(_02336_),
    .A2(_02525_),
    .B(_02526_),
    .C(_02528_),
    .Y(_02529_));
 NOR2x2_ASAP7_75t_R _25272_ (.A(net623),
    .B(_02290_),
    .Y(_02530_));
 AO21x1_ASAP7_75t_R _25273_ (.A1(_02530_),
    .A2(_02502_),
    .B(_02405_),
    .Y(_02531_));
 NAND2x1_ASAP7_75t_R _25274_ (.A(_02315_),
    .B(_02420_),
    .Y(_02532_));
 NAND2x1_ASAP7_75t_R _25275_ (.A(_02310_),
    .B(_02490_),
    .Y(_02533_));
 NAND2x2_ASAP7_75t_R _25276_ (.A(net463),
    .B(_02309_),
    .Y(_02534_));
 NAND3x1_ASAP7_75t_R _25277_ (.A(_02534_),
    .B(_02533_),
    .C(_02532_),
    .Y(_02535_));
 OAI21x1_ASAP7_75t_R _25278_ (.A1(_02531_),
    .A2(_02535_),
    .B(_02333_),
    .Y(_02536_));
 AO21x1_ASAP7_75t_R _25279_ (.A1(_15951_),
    .A2(_01215_),
    .B(_02460_),
    .Y(_02537_));
 NOR2x1_ASAP7_75t_R _25280_ (.A(_02368_),
    .B(_02537_),
    .Y(_02538_));
 AO21x1_ASAP7_75t_R _25281_ (.A1(_02480_),
    .A2(net73),
    .B(_02405_),
    .Y(_02539_));
 BUFx6f_ASAP7_75t_R _25282_ (.A(_02381_),
    .Y(_02540_));
 BUFx6f_ASAP7_75t_R _25283_ (.A(_02337_),
    .Y(_02541_));
 AOI21x1_ASAP7_75t_R _25284_ (.A1(net679),
    .A2(_02540_),
    .B(_02527_),
    .Y(_02542_));
 NAND2x1_ASAP7_75t_R _25285_ (.A(_02379_),
    .B(_02395_),
    .Y(_02543_));
 AOI21x1_ASAP7_75t_R _25286_ (.A1(_02543_),
    .A2(_02542_),
    .B(_02356_),
    .Y(_02544_));
 OAI21x1_ASAP7_75t_R _25287_ (.A1(_02538_),
    .A2(_02539_),
    .B(_02544_),
    .Y(_02545_));
 OAI21x1_ASAP7_75t_R _25288_ (.A1(_02529_),
    .A2(_02536_),
    .B(_02545_),
    .Y(_02546_));
 AOI21x1_ASAP7_75t_R _25289_ (.A1(_02373_),
    .A2(_02312_),
    .B(_02285_),
    .Y(_02547_));
 NAND2x1_ASAP7_75t_R _25290_ (.A(_02332_),
    .B(_02301_),
    .Y(_02548_));
 AOI221x1_ASAP7_75t_R _25291_ (.A1(_02379_),
    .A2(_02547_),
    .B1(_02336_),
    .B2(_02486_),
    .C(_02548_),
    .Y(_02549_));
 NOR2x1_ASAP7_75t_R _25292_ (.A(_02350_),
    .B(_02332_),
    .Y(_02550_));
 AOI21x1_ASAP7_75t_R _25293_ (.A1(_00577_),
    .A2(_02550_),
    .B(_02394_),
    .Y(_02551_));
 AOI21x1_ASAP7_75t_R _25294_ (.A1(_02378_),
    .A2(_02272_),
    .B(_02308_),
    .Y(_02552_));
 NAND2x1_ASAP7_75t_R _25295_ (.A(_02466_),
    .B(_02552_),
    .Y(_02553_));
 AOI21x1_ASAP7_75t_R _25296_ (.A1(_02551_),
    .A2(_02553_),
    .B(_02364_),
    .Y(_02554_));
 NOR2x2_ASAP7_75t_R _25297_ (.A(_02272_),
    .B(_15938_),
    .Y(_02555_));
 NOR2x1_ASAP7_75t_R _25298_ (.A(_02555_),
    .B(_02286_),
    .Y(_02556_));
 INVx1_ASAP7_75t_R _25299_ (.A(_02556_),
    .Y(_02557_));
 NAND2x1_ASAP7_75t_R _25300_ (.A(_02397_),
    .B(_02317_),
    .Y(_02558_));
 AOI21x1_ASAP7_75t_R _25301_ (.A1(_02385_),
    .A2(_02392_),
    .B(_02558_),
    .Y(_02559_));
 NAND2x1_ASAP7_75t_R _25302_ (.A(_02557_),
    .B(_02559_),
    .Y(_02560_));
 NAND2x1_ASAP7_75t_R _25303_ (.A(_02554_),
    .B(_02560_),
    .Y(_02561_));
 OAI21x1_ASAP7_75t_R _25304_ (.A1(_02549_),
    .A2(_02561_),
    .B(_02471_),
    .Y(_02562_));
 AOI21x1_ASAP7_75t_R _25305_ (.A1(_02498_),
    .A2(_02546_),
    .B(_02562_),
    .Y(_02563_));
 AOI21x1_ASAP7_75t_R _25306_ (.A1(_02499_),
    .A2(_02524_),
    .B(_02563_),
    .Y(_00097_));
 OA21x2_ASAP7_75t_R _25307_ (.A1(_15948_),
    .A2(_02435_),
    .B(_02310_),
    .Y(_02564_));
 AOI211x1_ASAP7_75t_R _25308_ (.A1(_02564_),
    .A2(_02372_),
    .B(_02455_),
    .C(_02349_),
    .Y(_02565_));
 INVx2_ASAP7_75t_R _25309_ (.A(_02454_),
    .Y(_02566_));
 AO21x1_ASAP7_75t_R _25310_ (.A1(_02566_),
    .A2(_02502_),
    .B(_02405_),
    .Y(_02567_));
 NAND2x2_ASAP7_75t_R _25311_ (.A(_02367_),
    .B(_02268_),
    .Y(_02568_));
 NOR2x2_ASAP7_75t_R _25312_ (.A(_02309_),
    .B(_02568_),
    .Y(_02569_));
 AOI211x1_ASAP7_75t_R _25313_ (.A1(_02564_),
    .A2(_02404_),
    .B(_02567_),
    .C(_02569_),
    .Y(_02570_));
 OAI21x1_ASAP7_75t_R _25314_ (.A1(_02565_),
    .A2(_02570_),
    .B(_02496_),
    .Y(_02571_));
 AOI21x1_ASAP7_75t_R _25315_ (.A1(_01217_),
    .A2(_02303_),
    .B(_02309_),
    .Y(_02572_));
 NAND2x1_ASAP7_75t_R _25316_ (.A(_02404_),
    .B(_02572_),
    .Y(_02573_));
 AO21x1_ASAP7_75t_R _25317_ (.A1(_02307_),
    .A2(_02353_),
    .B(_02315_),
    .Y(_02574_));
 AO21x1_ASAP7_75t_R _25318_ (.A1(_02573_),
    .A2(_02574_),
    .B(_02349_),
    .Y(_02575_));
 AND3x1_ASAP7_75t_R _25319_ (.A(_02385_),
    .B(_02310_),
    .C(_02454_),
    .Y(_02576_));
 INVx1_ASAP7_75t_R _25320_ (.A(_02568_),
    .Y(_02577_));
 OAI21x1_ASAP7_75t_R _25321_ (.A1(_02286_),
    .A2(_02577_),
    .B(_02527_),
    .Y(_02578_));
 OA21x2_ASAP7_75t_R _25322_ (.A1(_02576_),
    .A2(_02578_),
    .B(_02356_),
    .Y(_02579_));
 NAND2x1_ASAP7_75t_R _25323_ (.A(_02575_),
    .B(_02579_),
    .Y(_02580_));
 BUFx10_ASAP7_75t_R _25324_ (.A(_02363_),
    .Y(_02581_));
 AOI21x1_ASAP7_75t_R _25325_ (.A1(_02571_),
    .A2(_02580_),
    .B(_02581_),
    .Y(_02582_));
 AOI21x1_ASAP7_75t_R _25326_ (.A1(_02303_),
    .A2(net57),
    .B(_02381_),
    .Y(_02583_));
 AND2x2_ASAP7_75t_R _25327_ (.A(_02583_),
    .B(_02307_),
    .Y(_02584_));
 NOR2x2_ASAP7_75t_R _25328_ (.A(net623),
    .B(_02303_),
    .Y(_02585_));
 NAND2x2_ASAP7_75t_R _25329_ (.A(_02460_),
    .B(_02432_),
    .Y(_02586_));
 NOR2x1_ASAP7_75t_R _25330_ (.A(_02585_),
    .B(_02586_),
    .Y(_02587_));
 OA21x2_ASAP7_75t_R _25331_ (.A1(_02584_),
    .A2(_02587_),
    .B(_02349_),
    .Y(_02588_));
 AOI21x1_ASAP7_75t_R _25332_ (.A1(_02369_),
    .A2(_02480_),
    .B(_02374_),
    .Y(_02589_));
 AO21x1_ASAP7_75t_R _25333_ (.A1(_02589_),
    .A2(_02477_),
    .B(_02482_),
    .Y(_02590_));
 NAND2x1_ASAP7_75t_R _25334_ (.A(_02460_),
    .B(net739),
    .Y(_02591_));
 OAI21x1_ASAP7_75t_R _25335_ (.A1(_02421_),
    .A2(_02591_),
    .B(_02405_),
    .Y(_02592_));
 NOR2x1_ASAP7_75t_R _25336_ (.A(_02464_),
    .B(_02592_),
    .Y(_02593_));
 NAND2x2_ASAP7_75t_R _25337_ (.A(_01218_),
    .B(_02268_),
    .Y(_02594_));
 NAND2x2_ASAP7_75t_R _25338_ (.A(_02594_),
    .B(_02514_),
    .Y(_02595_));
 NAND2x2_ASAP7_75t_R _25339_ (.A(_02290_),
    .B(_15940_),
    .Y(_02596_));
 NAND2x2_ASAP7_75t_R _25340_ (.A(_02547_),
    .B(_02596_),
    .Y(_02597_));
 AOI21x1_ASAP7_75t_R _25341_ (.A1(_02595_),
    .A2(_02597_),
    .B(_02509_),
    .Y(_02598_));
 OAI21x1_ASAP7_75t_R _25342_ (.A1(_02593_),
    .A2(_02598_),
    .B(_02496_),
    .Y(_02599_));
 OAI21x1_ASAP7_75t_R _25343_ (.A1(_02588_),
    .A2(_02590_),
    .B(_02599_),
    .Y(_02600_));
 OAI21x1_ASAP7_75t_R _25344_ (.A1(_02498_),
    .A2(_02600_),
    .B(_02471_),
    .Y(_02601_));
 OA21x2_ASAP7_75t_R _25345_ (.A1(_01222_),
    .A2(_02345_),
    .B(_02317_),
    .Y(_02602_));
 NAND2x1_ASAP7_75t_R _25346_ (.A(_02602_),
    .B(_02597_),
    .Y(_02603_));
 AOI21x1_ASAP7_75t_R _25347_ (.A1(_00579_),
    .A2(_02310_),
    .B(_02374_),
    .Y(_02604_));
 AOI21x1_ASAP7_75t_R _25348_ (.A1(_02509_),
    .A2(_02604_),
    .B(_02356_),
    .Y(_02605_));
 NAND2x1_ASAP7_75t_R _25349_ (.A(_02603_),
    .B(_02605_),
    .Y(_02606_));
 AO21x1_ASAP7_75t_R _25350_ (.A1(_02307_),
    .A2(net739),
    .B(_02315_),
    .Y(_02607_));
 AOI21x1_ASAP7_75t_R _25351_ (.A1(_02607_),
    .A2(_02347_),
    .B(_02399_),
    .Y(_02608_));
 INVx1_ASAP7_75t_R _25352_ (.A(_02480_),
    .Y(_02609_));
 AND2x2_ASAP7_75t_R _25353_ (.A(_02391_),
    .B(_01215_),
    .Y(_02610_));
 NAND2x2_ASAP7_75t_R _25354_ (.A(_02610_),
    .B(_02272_),
    .Y(_02611_));
 INVx1_ASAP7_75t_R _25355_ (.A(_02611_),
    .Y(_02612_));
 AOI21x1_ASAP7_75t_R _25356_ (.A1(_02466_),
    .A2(_02552_),
    .B(_02405_),
    .Y(_02613_));
 OAI21x1_ASAP7_75t_R _25357_ (.A1(_02609_),
    .A2(_02612_),
    .B(_02613_),
    .Y(_02614_));
 AOI21x1_ASAP7_75t_R _25358_ (.A1(_02608_),
    .A2(_02614_),
    .B(_02364_),
    .Y(_02615_));
 AOI21x1_ASAP7_75t_R _25359_ (.A1(_02606_),
    .A2(_02615_),
    .B(_02471_),
    .Y(_02616_));
 NOR2x1_ASAP7_75t_R _25360_ (.A(_02285_),
    .B(_02445_),
    .Y(_02617_));
 AND2x2_ASAP7_75t_R _25361_ (.A(_02617_),
    .B(_02314_),
    .Y(_02618_));
 NOR2x2_ASAP7_75t_R _25362_ (.A(_02303_),
    .B(net57),
    .Y(_02619_));
 AOI211x1_ASAP7_75t_R _25363_ (.A1(_00573_),
    .A2(_15951_),
    .B(_02619_),
    .C(_02419_),
    .Y(_02620_));
 OAI21x1_ASAP7_75t_R _25364_ (.A1(_02618_),
    .A2(_02620_),
    .B(_02318_),
    .Y(_02621_));
 OAI21x1_ASAP7_75t_R _25365_ (.A1(_02312_),
    .A2(net57),
    .B(_02309_),
    .Y(_02622_));
 OAI21x1_ASAP7_75t_R _25366_ (.A1(_02287_),
    .A2(_02622_),
    .B(_02346_),
    .Y(_02623_));
 AND2x2_ASAP7_75t_R _25367_ (.A(_02350_),
    .B(_00577_),
    .Y(_02624_));
 OA21x2_ASAP7_75t_R _25368_ (.A1(_02623_),
    .A2(_02624_),
    .B(_02398_),
    .Y(_02625_));
 NAND2x1_ASAP7_75t_R _25369_ (.A(_02621_),
    .B(_02625_),
    .Y(_02626_));
 OA21x2_ASAP7_75t_R _25370_ (.A1(_01220_),
    .A2(_02345_),
    .B(_02375_),
    .Y(_02627_));
 NAND2x2_ASAP7_75t_R _25371_ (.A(net685),
    .B(_02290_),
    .Y(_02628_));
 AO21x1_ASAP7_75t_R _25372_ (.A1(_02485_),
    .A2(_02628_),
    .B(_02315_),
    .Y(_02629_));
 AOI21x1_ASAP7_75t_R _25373_ (.A1(_02627_),
    .A2(_02629_),
    .B(_02399_),
    .Y(_02630_));
 OAI21x1_ASAP7_75t_R _25374_ (.A1(_02585_),
    .A2(_02555_),
    .B(_02419_),
    .Y(_02631_));
 NOR2x1_ASAP7_75t_R _25375_ (.A(_02375_),
    .B(_02464_),
    .Y(_02632_));
 NAND2x1_ASAP7_75t_R _25376_ (.A(_02631_),
    .B(_02632_),
    .Y(_02633_));
 AOI21x1_ASAP7_75t_R _25377_ (.A1(_02630_),
    .A2(_02633_),
    .B(_02581_),
    .Y(_02634_));
 NAND2x1_ASAP7_75t_R _25378_ (.A(_02626_),
    .B(_02634_),
    .Y(_02635_));
 NAND2x1_ASAP7_75t_R _25379_ (.A(_02616_),
    .B(_02635_),
    .Y(_02636_));
 OAI21x1_ASAP7_75t_R _25380_ (.A1(_02582_),
    .A2(_02601_),
    .B(_02636_),
    .Y(_00098_));
 AOI21x1_ASAP7_75t_R _25381_ (.A1(_02314_),
    .A2(_02517_),
    .B(_02351_),
    .Y(_02637_));
 AND3x1_ASAP7_75t_R _25382_ (.A(_02353_),
    .B(_02379_),
    .C(_02315_),
    .Y(_02638_));
 OAI21x1_ASAP7_75t_R _25383_ (.A1(_02637_),
    .A2(_02638_),
    .B(_02477_),
    .Y(_02639_));
 NAND2x1_ASAP7_75t_R _25384_ (.A(net623),
    .B(_15940_),
    .Y(_02640_));
 AOI21x1_ASAP7_75t_R _25385_ (.A1(_02513_),
    .A2(_02640_),
    .B(_02351_),
    .Y(_02641_));
 INVx1_ASAP7_75t_R _25386_ (.A(_02342_),
    .Y(_02642_));
 BUFx6f_ASAP7_75t_R _25387_ (.A(_02460_),
    .Y(_02643_));
 AOI21x1_ASAP7_75t_R _25388_ (.A1(_02541_),
    .A2(_02642_),
    .B(_02643_),
    .Y(_02644_));
 OAI21x1_ASAP7_75t_R _25389_ (.A1(_02641_),
    .A2(_02644_),
    .B(_02349_),
    .Y(_02645_));
 NAND2x1_ASAP7_75t_R _25390_ (.A(_02639_),
    .B(_02645_),
    .Y(_02646_));
 AOI21x1_ASAP7_75t_R _25391_ (.A1(_02289_),
    .A2(_02513_),
    .B(_02643_),
    .Y(_02647_));
 OAI21x1_ASAP7_75t_R _25392_ (.A1(_02547_),
    .A2(_02647_),
    .B(_02477_),
    .Y(_02648_));
 AND2x2_ASAP7_75t_R _25393_ (.A(_02572_),
    .B(net73),
    .Y(_02649_));
 NOR2x1_ASAP7_75t_R _25394_ (.A(_02474_),
    .B(_02403_),
    .Y(_02650_));
 OAI21x1_ASAP7_75t_R _25395_ (.A1(_02649_),
    .A2(_02650_),
    .B(_02528_),
    .Y(_02651_));
 AOI21x1_ASAP7_75t_R _25396_ (.A1(_02648_),
    .A2(_02651_),
    .B(_02333_),
    .Y(_02652_));
 AOI211x1_ASAP7_75t_R _25397_ (.A1(_02646_),
    .A2(_02333_),
    .B(_02652_),
    .C(_02581_),
    .Y(_02653_));
 INVx1_ASAP7_75t_R _25398_ (.A(_02314_),
    .Y(_02654_));
 NOR2x1_ASAP7_75t_R _25399_ (.A(_02491_),
    .B(_02654_),
    .Y(_02655_));
 NAND2x1_ASAP7_75t_R _25400_ (.A(_02460_),
    .B(_02353_),
    .Y(_02656_));
 OAI21x1_ASAP7_75t_R _25401_ (.A1(_02490_),
    .A2(_02656_),
    .B(_02527_),
    .Y(_02657_));
 NOR2x1_ASAP7_75t_R _25402_ (.A(_02655_),
    .B(_02657_),
    .Y(_02658_));
 OAI21x1_ASAP7_75t_R _25403_ (.A1(_02493_),
    .A2(_02500_),
    .B(_02540_),
    .Y(_02659_));
 NAND2x1_ASAP7_75t_R _25404_ (.A(net73),
    .B(_02583_),
    .Y(_02660_));
 AOI21x1_ASAP7_75t_R _25405_ (.A1(_02659_),
    .A2(_02660_),
    .B(_02318_),
    .Y(_02661_));
 OAI21x1_ASAP7_75t_R _25406_ (.A1(_02658_),
    .A2(_02661_),
    .B(_02333_),
    .Y(_02662_));
 NAND2x1_ASAP7_75t_R _25407_ (.A(_02404_),
    .B(_02583_),
    .Y(_02663_));
 AOI21x1_ASAP7_75t_R _25408_ (.A1(_02656_),
    .A2(_02663_),
    .B(_02509_),
    .Y(_02664_));
 NAND2x1_ASAP7_75t_R _25409_ (.A(_02419_),
    .B(_02352_),
    .Y(_02665_));
 OAI21x1_ASAP7_75t_R _25410_ (.A1(_02530_),
    .A2(_02287_),
    .B(_02502_),
    .Y(_02666_));
 AOI21x1_ASAP7_75t_R _25411_ (.A1(_02665_),
    .A2(_02666_),
    .B(_02318_),
    .Y(_02667_));
 OAI21x1_ASAP7_75t_R _25412_ (.A1(_02664_),
    .A2(_02667_),
    .B(_02496_),
    .Y(_02668_));
 NAND2x1_ASAP7_75t_R _25413_ (.A(_02662_),
    .B(_02668_),
    .Y(_02669_));
 OAI21x1_ASAP7_75t_R _25414_ (.A1(_02498_),
    .A2(_02669_),
    .B(_02414_),
    .Y(_02670_));
 INVx1_ASAP7_75t_R _25415_ (.A(_02353_),
    .Y(_02671_));
 NAND2x1_ASAP7_75t_R _25416_ (.A(_02671_),
    .B(_02550_),
    .Y(_02672_));
 OA21x2_ASAP7_75t_R _25417_ (.A1(_02383_),
    .A2(_02292_),
    .B(_02394_),
    .Y(_02673_));
 NAND2x1_ASAP7_75t_R _25418_ (.A(_02672_),
    .B(_02673_),
    .Y(_02674_));
 AO21x1_ASAP7_75t_R _25419_ (.A1(_15951_),
    .A2(_02341_),
    .B(_02345_),
    .Y(_02675_));
 OAI21x1_ASAP7_75t_R _25420_ (.A1(_15951_),
    .A2(net57),
    .B(_02398_),
    .Y(_02676_));
 NAND2x1_ASAP7_75t_R _25421_ (.A(_02315_),
    .B(_02401_),
    .Y(_02677_));
 OAI22x1_ASAP7_75t_R _25422_ (.A1(_02675_),
    .A2(_02676_),
    .B1(_02399_),
    .B2(_02677_),
    .Y(_02678_));
 OAI21x1_ASAP7_75t_R _25423_ (.A1(_02674_),
    .A2(_02678_),
    .B(_02581_),
    .Y(_02679_));
 OA21x2_ASAP7_75t_R _25424_ (.A1(_02454_),
    .A2(_02292_),
    .B(_02332_),
    .Y(_02680_));
 NAND2x1_ASAP7_75t_R _25425_ (.A(_02680_),
    .B(_02573_),
    .Y(_02681_));
 AOI21x1_ASAP7_75t_R _25426_ (.A1(_02541_),
    .A2(_02395_),
    .B(_02332_),
    .Y(_02682_));
 OAI21x1_ASAP7_75t_R _25427_ (.A1(_02403_),
    .A2(_02612_),
    .B(_02682_),
    .Y(_02683_));
 AOI21x1_ASAP7_75t_R _25428_ (.A1(_02683_),
    .A2(_02681_),
    .B(_02528_),
    .Y(_02684_));
 NOR2x1_ASAP7_75t_R _25429_ (.A(_02679_),
    .B(_02684_),
    .Y(_02685_));
 NAND2x1_ASAP7_75t_R _25430_ (.A(_02611_),
    .B(_02427_),
    .Y(_02686_));
 AOI21x1_ASAP7_75t_R _25431_ (.A1(_02553_),
    .A2(_02686_),
    .B(_02318_),
    .Y(_02687_));
 NAND2x1_ASAP7_75t_R _25432_ (.A(_02399_),
    .B(_02578_),
    .Y(_02688_));
 OAI21x1_ASAP7_75t_R _25433_ (.A1(_02687_),
    .A2(_02688_),
    .B(_02364_),
    .Y(_02689_));
 AO21x1_ASAP7_75t_R _25434_ (.A1(_02568_),
    .A2(_02307_),
    .B(_02310_),
    .Y(_02690_));
 OAI21x1_ASAP7_75t_R _25435_ (.A1(_15943_),
    .A2(_15948_),
    .B(_02454_),
    .Y(_02691_));
 AOI21x1_ASAP7_75t_R _25436_ (.A1(_02540_),
    .A2(_02691_),
    .B(_02405_),
    .Y(_02692_));
 NAND2x1_ASAP7_75t_R _25437_ (.A(_02690_),
    .B(_02692_),
    .Y(_02693_));
 AOI21x1_ASAP7_75t_R _25438_ (.A1(_02540_),
    .A2(_02431_),
    .B(_02527_),
    .Y(_02694_));
 NAND2x1_ASAP7_75t_R _25439_ (.A(_02694_),
    .B(_02520_),
    .Y(_02695_));
 AOI21x1_ASAP7_75t_R _25440_ (.A1(_02693_),
    .A2(_02695_),
    .B(_02496_),
    .Y(_02696_));
 NOR2x1_ASAP7_75t_R _25441_ (.A(_02689_),
    .B(_02696_),
    .Y(_02697_));
 OAI21x1_ASAP7_75t_R _25442_ (.A1(_02697_),
    .A2(_02685_),
    .B(_02471_),
    .Y(_02698_));
 OAI21x1_ASAP7_75t_R _25443_ (.A1(_02653_),
    .A2(_02670_),
    .B(_02698_),
    .Y(_00099_));
 AO21x1_ASAP7_75t_R _25444_ (.A1(_02372_),
    .A2(_02336_),
    .B(_02502_),
    .Y(_02699_));
 NAND2x1_ASAP7_75t_R _25445_ (.A(_15943_),
    .B(_15940_),
    .Y(_02700_));
 AOI21x1_ASAP7_75t_R _25446_ (.A1(_02372_),
    .A2(_02700_),
    .B(_02310_),
    .Y(_02701_));
 INVx1_ASAP7_75t_R _25447_ (.A(_02701_),
    .Y(_02702_));
 NAND2x1_ASAP7_75t_R _25448_ (.A(_02699_),
    .B(_02702_),
    .Y(_02703_));
 OAI21x1_ASAP7_75t_R _25449_ (.A1(_02556_),
    .A2(_02623_),
    .B(_02482_),
    .Y(_02704_));
 AOI21x1_ASAP7_75t_R _25450_ (.A1(_02528_),
    .A2(_02703_),
    .B(_02704_),
    .Y(_02705_));
 NOR2x1_ASAP7_75t_R _25451_ (.A(_02420_),
    .B(_02427_),
    .Y(_02706_));
 AO21x1_ASAP7_75t_R _25452_ (.A1(_02706_),
    .A2(_02349_),
    .B(_02482_),
    .Y(_02707_));
 AO21x1_ASAP7_75t_R _25453_ (.A1(_02486_),
    .A2(_02336_),
    .B(_02527_),
    .Y(_02708_));
 INVx1_ASAP7_75t_R _25454_ (.A(_02555_),
    .Y(_02709_));
 AND2x2_ASAP7_75t_R _25455_ (.A(_02467_),
    .B(_02709_),
    .Y(_02710_));
 NOR2x1_ASAP7_75t_R _25456_ (.A(_02708_),
    .B(_02710_),
    .Y(_02711_));
 OAI21x1_ASAP7_75t_R _25457_ (.A1(_02707_),
    .A2(_02711_),
    .B(_02414_),
    .Y(_02712_));
 OAI21x1_ASAP7_75t_R _25458_ (.A1(_02705_),
    .A2(_02712_),
    .B(_02498_),
    .Y(_02713_));
 NAND2x1_ASAP7_75t_R _25459_ (.A(_02301_),
    .B(_02537_),
    .Y(_02714_));
 OAI21x1_ASAP7_75t_R _25460_ (.A1(_02480_),
    .A2(_02714_),
    .B(_02356_),
    .Y(_02715_));
 INVx1_ASAP7_75t_R _25461_ (.A(_02514_),
    .Y(_02716_));
 NOR2x1_ASAP7_75t_R _25462_ (.A(net463),
    .B(_02716_),
    .Y(_02717_));
 NOR2x1_ASAP7_75t_R _25463_ (.A(_02717_),
    .B(_02452_),
    .Y(_02718_));
 OAI21x1_ASAP7_75t_R _25464_ (.A1(_02715_),
    .A2(_02718_),
    .B(_02413_),
    .Y(_02719_));
 NOR2x1_ASAP7_75t_R _25465_ (.A(_02386_),
    .B(_02526_),
    .Y(_02720_));
 OA21x2_ASAP7_75t_R _25466_ (.A1(_02344_),
    .A2(_02643_),
    .B(_02349_),
    .Y(_02721_));
 NAND2x1_ASAP7_75t_R _25467_ (.A(_02594_),
    .B(_02525_),
    .Y(_02722_));
 OA21x2_ASAP7_75t_R _25468_ (.A1(_15948_),
    .A2(_02315_),
    .B(_02375_),
    .Y(_02723_));
 AO21x1_ASAP7_75t_R _25469_ (.A1(_02722_),
    .A2(_02723_),
    .B(_02356_),
    .Y(_02724_));
 AOI21x1_ASAP7_75t_R _25470_ (.A1(_02720_),
    .A2(_02721_),
    .B(_02724_),
    .Y(_02725_));
 NOR2x1_ASAP7_75t_R _25471_ (.A(_02719_),
    .B(_02725_),
    .Y(_02726_));
 OA21x2_ASAP7_75t_R _25472_ (.A1(_02566_),
    .A2(net463),
    .B(_02540_),
    .Y(_02727_));
 OAI21x1_ASAP7_75t_R _25473_ (.A1(_02455_),
    .A2(_02727_),
    .B(_02528_),
    .Y(_02728_));
 AOI21x1_ASAP7_75t_R _25474_ (.A1(_01218_),
    .A2(_02290_),
    .B(_02381_),
    .Y(_02729_));
 NAND2x1_ASAP7_75t_R _25475_ (.A(_02353_),
    .B(_02729_),
    .Y(_02730_));
 AO21x1_ASAP7_75t_R _25476_ (.A1(_02428_),
    .A2(_02730_),
    .B(_02349_),
    .Y(_02731_));
 AOI21x1_ASAP7_75t_R _25477_ (.A1(_02728_),
    .A2(_02731_),
    .B(_02496_),
    .Y(_02732_));
 OA21x2_ASAP7_75t_R _25478_ (.A1(_02555_),
    .A2(_02490_),
    .B(_02643_),
    .Y(_02733_));
 OAI21x1_ASAP7_75t_R _25479_ (.A1(_02733_),
    .A2(_02439_),
    .B(_02482_),
    .Y(_02734_));
 AOI21x1_ASAP7_75t_R _25480_ (.A1(_02373_),
    .A2(_02272_),
    .B(_02285_),
    .Y(_02735_));
 NAND2x1_ASAP7_75t_R _25481_ (.A(_02385_),
    .B(_02735_),
    .Y(_02736_));
 AND3x1_ASAP7_75t_R _25482_ (.A(_02595_),
    .B(_02736_),
    .C(_02318_),
    .Y(_02737_));
 OAI21x1_ASAP7_75t_R _25483_ (.A1(_02734_),
    .A2(_02737_),
    .B(_02414_),
    .Y(_02738_));
 NOR2x1_ASAP7_75t_R _25484_ (.A(_02738_),
    .B(_02732_),
    .Y(_02739_));
 AO21x1_ASAP7_75t_R _25485_ (.A1(_00575_),
    .A2(_02502_),
    .B(_02527_),
    .Y(_02740_));
 OAI21x1_ASAP7_75t_R _25486_ (.A1(_02617_),
    .A2(_02740_),
    .B(_02356_),
    .Y(_02741_));
 OAI21x1_ASAP7_75t_R _25487_ (.A1(_02643_),
    .A2(_02628_),
    .B(_02301_),
    .Y(_02742_));
 AOI21x1_ASAP7_75t_R _25488_ (.A1(_02372_),
    .A2(_02427_),
    .B(_02742_),
    .Y(_02743_));
 OAI21x1_ASAP7_75t_R _25489_ (.A1(_02741_),
    .A2(_02743_),
    .B(_02471_),
    .Y(_02744_));
 OAI21x1_ASAP7_75t_R _25490_ (.A1(_02461_),
    .A2(_02293_),
    .B(_02477_),
    .Y(_02745_));
 AND2x2_ASAP7_75t_R _25491_ (.A(_02427_),
    .B(_02291_),
    .Y(_02746_));
 OAI21x1_ASAP7_75t_R _25492_ (.A1(_02701_),
    .A2(_02746_),
    .B(_02528_),
    .Y(_02747_));
 AOI21x1_ASAP7_75t_R _25493_ (.A1(_02745_),
    .A2(_02747_),
    .B(_02333_),
    .Y(_02748_));
 OAI21x1_ASAP7_75t_R _25494_ (.A1(_02744_),
    .A2(_02748_),
    .B(_02581_),
    .Y(_02749_));
 OAI22x1_ASAP7_75t_R _25495_ (.A1(_02713_),
    .A2(_02726_),
    .B1(_02739_),
    .B2(_02749_),
    .Y(_00100_));
 NAND2x1_ASAP7_75t_R _25496_ (.A(_02426_),
    .B(_02572_),
    .Y(_02750_));
 INVx1_ASAP7_75t_R _25497_ (.A(_02610_),
    .Y(_02751_));
 AOI21x1_ASAP7_75t_R _25498_ (.A1(_02751_),
    .A2(_02564_),
    .B(_02477_),
    .Y(_02752_));
 AO21x1_ASAP7_75t_R _25499_ (.A1(_02391_),
    .A2(_15948_),
    .B(_02403_),
    .Y(_02753_));
 AOI221x1_ASAP7_75t_R _25500_ (.A1(_02750_),
    .A2(_02752_),
    .B1(_02387_),
    .B2(_02753_),
    .C(_02581_),
    .Y(_02754_));
 OA21x2_ASAP7_75t_R _25501_ (.A1(_15940_),
    .A2(_02502_),
    .B(_02405_),
    .Y(_02755_));
 OAI21x1_ASAP7_75t_R _25502_ (.A1(_00571_),
    .A2(_15948_),
    .B(_02379_),
    .Y(_02756_));
 AOI21x1_ASAP7_75t_R _25503_ (.A1(_02643_),
    .A2(_02756_),
    .B(_02509_),
    .Y(_02757_));
 NAND2x1_ASAP7_75t_R _25504_ (.A(_02395_),
    .B(_02700_),
    .Y(_02758_));
 AOI22x1_ASAP7_75t_R _25505_ (.A1(_02702_),
    .A2(_02755_),
    .B1(_02757_),
    .B2(_02758_),
    .Y(_02759_));
 OAI21x1_ASAP7_75t_R _25506_ (.A1(_02498_),
    .A2(_02759_),
    .B(_02333_),
    .Y(_02760_));
 AND2x2_ASAP7_75t_R _25507_ (.A(_02517_),
    .B(_02317_),
    .Y(_02761_));
 AOI21x1_ASAP7_75t_R _25508_ (.A1(_02716_),
    .A2(_02761_),
    .B(_02363_),
    .Y(_02762_));
 AO21x1_ASAP7_75t_R _25509_ (.A1(_02337_),
    .A2(_02292_),
    .B(_02317_),
    .Y(_02763_));
 AO21x1_ASAP7_75t_R _25510_ (.A1(_02540_),
    .A2(_02691_),
    .B(_02763_),
    .Y(_02764_));
 AOI21x1_ASAP7_75t_R _25511_ (.A1(_02762_),
    .A2(_02764_),
    .B(_02356_),
    .Y(_02765_));
 AO21x1_ASAP7_75t_R _25512_ (.A1(_02313_),
    .A2(_02541_),
    .B(_02292_),
    .Y(_02766_));
 NOR2x1_ASAP7_75t_R _25513_ (.A(_02394_),
    .B(_02569_),
    .Y(_02767_));
 NAND2x1_ASAP7_75t_R _25514_ (.A(_02766_),
    .B(_02767_),
    .Y(_02768_));
 AO21x1_ASAP7_75t_R _25515_ (.A1(_02372_),
    .A2(_02432_),
    .B(_02345_),
    .Y(_02769_));
 AND2x2_ASAP7_75t_R _25516_ (.A(_02534_),
    .B(_02317_),
    .Y(_02770_));
 AOI21x1_ASAP7_75t_R _25517_ (.A1(_02770_),
    .A2(_02769_),
    .B(_02364_),
    .Y(_02771_));
 NAND2x1_ASAP7_75t_R _25518_ (.A(_02771_),
    .B(_02768_),
    .Y(_02772_));
 AOI21x1_ASAP7_75t_R _25519_ (.A1(_02765_),
    .A2(_02772_),
    .B(_02471_),
    .Y(_02773_));
 OAI21x1_ASAP7_75t_R _25520_ (.A1(_02754_),
    .A2(_02760_),
    .B(_02773_),
    .Y(_02774_));
 OA21x2_ASAP7_75t_R _25521_ (.A1(_02585_),
    .A2(_02493_),
    .B(_02351_),
    .Y(_02775_));
 AO21x1_ASAP7_75t_R _25522_ (.A1(_02342_),
    .A2(_02345_),
    .B(_02346_),
    .Y(_02776_));
 AND2x2_ASAP7_75t_R _25523_ (.A(_02552_),
    .B(_02594_),
    .Y(_02777_));
 OA21x2_ASAP7_75t_R _25524_ (.A1(_02776_),
    .A2(_02777_),
    .B(_02398_),
    .Y(_02778_));
 OA21x2_ASAP7_75t_R _25525_ (.A1(_02452_),
    .A2(_02775_),
    .B(_02778_),
    .Y(_02779_));
 AO21x1_ASAP7_75t_R _25526_ (.A1(_15943_),
    .A2(_02540_),
    .B(_02527_),
    .Y(_02780_));
 OAI21x1_ASAP7_75t_R _25527_ (.A1(_02780_),
    .A2(_02288_),
    .B(_02356_),
    .Y(_02781_));
 NAND2x1_ASAP7_75t_R _25528_ (.A(_02541_),
    .B(_02547_),
    .Y(_02782_));
 NAND2x1_ASAP7_75t_R _25529_ (.A(_02372_),
    .B(_02572_),
    .Y(_02783_));
 AND3x1_ASAP7_75t_R _25530_ (.A(_02782_),
    .B(_02783_),
    .C(_02318_),
    .Y(_02784_));
 OAI21x1_ASAP7_75t_R _25531_ (.A1(_02781_),
    .A2(_02784_),
    .B(_02498_),
    .Y(_02785_));
 AO21x1_ASAP7_75t_R _25532_ (.A1(_02643_),
    .A2(_02594_),
    .B(_02451_),
    .Y(_02786_));
 AOI21x1_ASAP7_75t_R _25533_ (.A1(_02419_),
    .A2(_02611_),
    .B(_02394_),
    .Y(_02787_));
 NAND2x1_ASAP7_75t_R _25534_ (.A(_02390_),
    .B(_02552_),
    .Y(_02788_));
 AOI21x1_ASAP7_75t_R _25535_ (.A1(_02787_),
    .A2(_02788_),
    .B(_02399_),
    .Y(_02789_));
 OAI21x1_ASAP7_75t_R _25536_ (.A1(_02477_),
    .A2(_02786_),
    .B(_02789_),
    .Y(_02790_));
 AO21x1_ASAP7_75t_R _25537_ (.A1(_00571_),
    .A2(_02460_),
    .B(_02317_),
    .Y(_02791_));
 OA21x2_ASAP7_75t_R _25538_ (.A1(_02791_),
    .A2(_02552_),
    .B(_02398_),
    .Y(_02792_));
 NAND2x1_ASAP7_75t_R _25539_ (.A(_02466_),
    .B(_02339_),
    .Y(_02793_));
 OAI21x1_ASAP7_75t_R _25540_ (.A1(_02460_),
    .A2(_02337_),
    .B(_02317_),
    .Y(_02794_));
 NOR2x1_ASAP7_75t_R _25541_ (.A(_02794_),
    .B(_02569_),
    .Y(_02795_));
 NAND2x1_ASAP7_75t_R _25542_ (.A(_02793_),
    .B(_02795_),
    .Y(_02796_));
 AOI21x1_ASAP7_75t_R _25543_ (.A1(_02792_),
    .A2(_02796_),
    .B(_02364_),
    .Y(_02797_));
 AOI21x1_ASAP7_75t_R _25544_ (.A1(_02790_),
    .A2(_02797_),
    .B(_02414_),
    .Y(_02798_));
 OAI21x1_ASAP7_75t_R _25545_ (.A1(_02779_),
    .A2(_02785_),
    .B(_02798_),
    .Y(_02799_));
 NAND2x1_ASAP7_75t_R _25546_ (.A(_02799_),
    .B(_02774_),
    .Y(_00101_));
 NAND2x1_ASAP7_75t_R _25547_ (.A(_02735_),
    .B(_02709_),
    .Y(_02800_));
 NAND2x1_ASAP7_75t_R _25548_ (.A(_02417_),
    .B(_02800_),
    .Y(_02801_));
 AOI21x1_ASAP7_75t_R _25549_ (.A1(_02513_),
    .A2(_02735_),
    .B(_02394_),
    .Y(_02802_));
 NOR2x1_ASAP7_75t_R _25550_ (.A(_02460_),
    .B(net463),
    .Y(_02803_));
 NAND2x1_ASAP7_75t_R _25551_ (.A(_02611_),
    .B(_02803_),
    .Y(_02804_));
 AOI21x1_ASAP7_75t_R _25552_ (.A1(_02802_),
    .A2(_02804_),
    .B(_02332_),
    .Y(_02805_));
 NAND2x1_ASAP7_75t_R _25553_ (.A(_02801_),
    .B(_02805_),
    .Y(_02806_));
 AO21x1_ASAP7_75t_R _25554_ (.A1(_02541_),
    .A2(_02432_),
    .B(_02345_),
    .Y(_02807_));
 NAND2x1_ASAP7_75t_R _25555_ (.A(_02372_),
    .B(_02547_),
    .Y(_02808_));
 AOI21x1_ASAP7_75t_R _25556_ (.A1(_02808_),
    .A2(_02807_),
    .B(_02301_),
    .Y(_02809_));
 NOR2x1_ASAP7_75t_R _25557_ (.A(_02794_),
    .B(_02604_),
    .Y(_02810_));
 OAI21x1_ASAP7_75t_R _25558_ (.A1(_02810_),
    .A2(_02809_),
    .B(_02356_),
    .Y(_02811_));
 AOI21x1_ASAP7_75t_R _25559_ (.A1(_02811_),
    .A2(_02806_),
    .B(_02364_),
    .Y(_02812_));
 NAND2x1_ASAP7_75t_R _25560_ (.A(_02385_),
    .B(_02640_),
    .Y(_02813_));
 AO21x1_ASAP7_75t_R _25561_ (.A1(_01221_),
    .A2(_01219_),
    .B(_02310_),
    .Y(_02814_));
 OAI21x1_ASAP7_75t_R _25562_ (.A1(_02351_),
    .A2(_02813_),
    .B(_02814_),
    .Y(_02815_));
 OA21x2_ASAP7_75t_R _25563_ (.A1(_02454_),
    .A2(_02292_),
    .B(_02317_),
    .Y(_02816_));
 OAI21x1_ASAP7_75t_R _25564_ (.A1(_02419_),
    .A2(_02490_),
    .B(_02586_),
    .Y(_02817_));
 AOI21x1_ASAP7_75t_R _25565_ (.A1(_02816_),
    .A2(_02817_),
    .B(_02399_),
    .Y(_02818_));
 OAI21x1_ASAP7_75t_R _25566_ (.A1(_02349_),
    .A2(_02815_),
    .B(_02818_),
    .Y(_02819_));
 OA21x2_ASAP7_75t_R _25567_ (.A1(_02270_),
    .A2(_02269_),
    .B(_00575_),
    .Y(_02820_));
 OAI21x1_ASAP7_75t_R _25568_ (.A1(_02420_),
    .A2(_02820_),
    .B(_02419_),
    .Y(_02821_));
 NAND2x1_ASAP7_75t_R _25569_ (.A(_02572_),
    .B(_02369_),
    .Y(_02822_));
 AOI21x1_ASAP7_75t_R _25570_ (.A1(_02821_),
    .A2(_02822_),
    .B(_02301_),
    .Y(_02823_));
 NAND2x1_ASAP7_75t_R _25571_ (.A(_02485_),
    .B(_02525_),
    .Y(_02824_));
 NOR2x1_ASAP7_75t_R _25572_ (.A(_02610_),
    .B(_15948_),
    .Y(_02825_));
 OAI21x1_ASAP7_75t_R _25573_ (.A1(_02566_),
    .A2(_02825_),
    .B(_02540_),
    .Y(_02826_));
 AOI21x1_ASAP7_75t_R _25574_ (.A1(_02824_),
    .A2(_02826_),
    .B(_02509_),
    .Y(_02827_));
 OAI21x1_ASAP7_75t_R _25575_ (.A1(_02823_),
    .A2(_02827_),
    .B(_02482_),
    .Y(_02828_));
 AOI21x1_ASAP7_75t_R _25576_ (.A1(_02819_),
    .A2(_02828_),
    .B(_02581_),
    .Y(_02829_));
 OAI21x1_ASAP7_75t_R _25577_ (.A1(_02812_),
    .A2(_02829_),
    .B(_02414_),
    .Y(_02830_));
 INVx1_ASAP7_75t_R _25578_ (.A(_02306_),
    .Y(_02831_));
 NOR2x1_ASAP7_75t_R _25579_ (.A(_02831_),
    .B(_02403_),
    .Y(_02832_));
 AOI21x1_ASAP7_75t_R _25580_ (.A1(_00580_),
    .A2(_02419_),
    .B(_02394_),
    .Y(_02833_));
 AOI21x1_ASAP7_75t_R _25581_ (.A1(_02833_),
    .A2(_02783_),
    .B(_02399_),
    .Y(_02834_));
 OAI21x1_ASAP7_75t_R _25582_ (.A1(_02531_),
    .A2(_02832_),
    .B(_02834_),
    .Y(_02835_));
 INVx1_ASAP7_75t_R _25583_ (.A(_02592_),
    .Y(_02836_));
 NAND2x1_ASAP7_75t_R _25584_ (.A(_02372_),
    .B(_02427_),
    .Y(_02837_));
 AOI21x1_ASAP7_75t_R _25585_ (.A1(_02675_),
    .A2(_02837_),
    .B(_02509_),
    .Y(_02838_));
 OAI21x1_ASAP7_75t_R _25586_ (.A1(_02836_),
    .A2(_02838_),
    .B(_02482_),
    .Y(_02839_));
 AOI21x1_ASAP7_75t_R _25587_ (.A1(_02835_),
    .A2(_02839_),
    .B(_02364_),
    .Y(_02840_));
 INVx1_ASAP7_75t_R _25588_ (.A(_02506_),
    .Y(_02841_));
 NAND2x1_ASAP7_75t_R _25589_ (.A(_02404_),
    .B(_02374_),
    .Y(_02842_));
 AOI21x1_ASAP7_75t_R _25590_ (.A1(_02841_),
    .A2(_02842_),
    .B(_02509_),
    .Y(_02843_));
 NAND2x1_ASAP7_75t_R _25591_ (.A(_02315_),
    .B(_02831_),
    .Y(_02844_));
 NAND2x1_ASAP7_75t_R _25592_ (.A(_02419_),
    .B(_02691_),
    .Y(_02845_));
 AOI21x1_ASAP7_75t_R _25593_ (.A1(_02844_),
    .A2(_02845_),
    .B(_02301_),
    .Y(_02846_));
 OAI21x1_ASAP7_75t_R _25594_ (.A1(_02843_),
    .A2(_02846_),
    .B(_02482_),
    .Y(_02847_));
 NAND2x1_ASAP7_75t_R _25595_ (.A(_02513_),
    .B(_02729_),
    .Y(_02848_));
 NOR2x1_ASAP7_75t_R _25596_ (.A(_15943_),
    .B(net57),
    .Y(_02849_));
 OAI21x1_ASAP7_75t_R _25597_ (.A1(_02585_),
    .A2(_02849_),
    .B(_02540_),
    .Y(_02850_));
 AOI21x1_ASAP7_75t_R _25598_ (.A1(_02848_),
    .A2(_02850_),
    .B(_02509_),
    .Y(_02851_));
 NAND2x1_ASAP7_75t_R _25599_ (.A(_02374_),
    .B(_02596_),
    .Y(_02852_));
 OAI21x1_ASAP7_75t_R _25600_ (.A1(_02530_),
    .A2(_02287_),
    .B(_02540_),
    .Y(_02853_));
 AOI21x1_ASAP7_75t_R _25601_ (.A1(_02852_),
    .A2(_02853_),
    .B(_02318_),
    .Y(_02854_));
 OAI21x1_ASAP7_75t_R _25602_ (.A1(_02851_),
    .A2(_02854_),
    .B(_02333_),
    .Y(_02855_));
 AOI21x1_ASAP7_75t_R _25603_ (.A1(_02847_),
    .A2(_02855_),
    .B(_02581_),
    .Y(_02856_));
 OAI21x1_ASAP7_75t_R _25604_ (.A1(_02840_),
    .A2(_02856_),
    .B(_02471_),
    .Y(_02857_));
 NAND2x1_ASAP7_75t_R _25605_ (.A(_02857_),
    .B(_02830_),
    .Y(_00102_));
 AOI21x1_ASAP7_75t_R _25606_ (.A1(net679),
    .A2(_02642_),
    .B(_02351_),
    .Y(_02858_));
 OA21x2_ASAP7_75t_R _25607_ (.A1(_02820_),
    .A2(_02490_),
    .B(_02351_),
    .Y(_02859_));
 OAI21x1_ASAP7_75t_R _25608_ (.A1(_02858_),
    .A2(_02859_),
    .B(_02477_),
    .Y(_02860_));
 INVx1_ASAP7_75t_R _25609_ (.A(_02686_),
    .Y(_02861_));
 AO21x1_ASAP7_75t_R _25610_ (.A1(_15951_),
    .A2(_02378_),
    .B(_02345_),
    .Y(_02862_));
 NOR2x1_ASAP7_75t_R _25611_ (.A(_02619_),
    .B(_02862_),
    .Y(_02863_));
 OAI21x1_ASAP7_75t_R _25612_ (.A1(_02861_),
    .A2(_02863_),
    .B(_02528_),
    .Y(_02864_));
 AOI21x1_ASAP7_75t_R _25613_ (.A1(_02860_),
    .A2(_02864_),
    .B(_02496_),
    .Y(_02865_));
 NOR2x1_ASAP7_75t_R _25614_ (.A(_02351_),
    .B(_02385_),
    .Y(_02866_));
 NOR2x1_ASAP7_75t_R _25615_ (.A(_02394_),
    .B(_02490_),
    .Y(_02867_));
 INVx1_ASAP7_75t_R _25616_ (.A(_02433_),
    .Y(_02868_));
 NAND2x1_ASAP7_75t_R _25617_ (.A(_02867_),
    .B(_02868_),
    .Y(_02869_));
 OAI21x1_ASAP7_75t_R _25618_ (.A1(_02866_),
    .A2(_02869_),
    .B(_02496_),
    .Y(_02870_));
 NOR2x1_ASAP7_75t_R _25619_ (.A(_02405_),
    .B(_02478_),
    .Y(_02871_));
 OA21x2_ASAP7_75t_R _25620_ (.A1(_02813_),
    .A2(_02351_),
    .B(_02871_),
    .Y(_02872_));
 OAI21x1_ASAP7_75t_R _25621_ (.A1(_02870_),
    .A2(_02872_),
    .B(_02498_),
    .Y(_02873_));
 OAI21x1_ASAP7_75t_R _25622_ (.A1(_02865_),
    .A2(_02873_),
    .B(_02414_),
    .Y(_02874_));
 NAND2x1_ASAP7_75t_R _25623_ (.A(net738),
    .B(_02381_),
    .Y(_02875_));
 AND2x2_ASAP7_75t_R _25624_ (.A(_02875_),
    .B(_02375_),
    .Y(_02876_));
 AO21x1_ASAP7_75t_R _25625_ (.A1(_02876_),
    .A2(_02868_),
    .B(_02399_),
    .Y(_02877_));
 AOI211x1_ASAP7_75t_R _25626_ (.A1(_02385_),
    .A2(_02392_),
    .B(_02742_),
    .C(_02386_),
    .Y(_02878_));
 OAI21x1_ASAP7_75t_R _25627_ (.A1(_02877_),
    .A2(_02878_),
    .B(_02581_),
    .Y(_02879_));
 AO22x2_ASAP7_75t_R _25628_ (.A1(_02485_),
    .A2(_02339_),
    .B1(_02519_),
    .B2(_02513_),
    .Y(_02880_));
 AO21x1_ASAP7_75t_R _25629_ (.A1(_02566_),
    .A2(_02502_),
    .B(_02527_),
    .Y(_02881_));
 NOR2x1_ASAP7_75t_R _25630_ (.A(_01221_),
    .B(_02292_),
    .Y(_02882_));
 AO21x1_ASAP7_75t_R _25631_ (.A1(_02671_),
    .A2(_02502_),
    .B(_02882_),
    .Y(_02883_));
 OAI21x1_ASAP7_75t_R _25632_ (.A1(_02881_),
    .A2(_02883_),
    .B(_02482_),
    .Y(_02884_));
 AOI21x1_ASAP7_75t_R _25633_ (.A1(_02528_),
    .A2(_02880_),
    .B(_02884_),
    .Y(_02885_));
 NOR2x1_ASAP7_75t_R _25634_ (.A(_02879_),
    .B(_02885_),
    .Y(_02886_));
 OAI22x1_ASAP7_75t_R _25635_ (.A1(_02875_),
    .A2(_15951_),
    .B1(_02643_),
    .B2(net679),
    .Y(_02887_));
 OAI21x1_ASAP7_75t_R _25636_ (.A1(_02528_),
    .A2(_02887_),
    .B(_02496_),
    .Y(_02888_));
 AOI21x1_ASAP7_75t_R _25637_ (.A1(net679),
    .A2(_02304_),
    .B(_02643_),
    .Y(_02889_));
 NOR3x1_ASAP7_75t_R _25638_ (.A(_02889_),
    .B(_02477_),
    .C(_02735_),
    .Y(_02890_));
 OAI21x1_ASAP7_75t_R _25639_ (.A1(_02888_),
    .A2(_02890_),
    .B(_02581_),
    .Y(_02891_));
 NOR2x1_ASAP7_75t_R _25640_ (.A(_02643_),
    .B(_15943_),
    .Y(_02892_));
 AO21x1_ASAP7_75t_R _25641_ (.A1(_02467_),
    .A2(_02709_),
    .B(_02892_),
    .Y(_02893_));
 NOR2x1_ASAP7_75t_R _25642_ (.A(_02474_),
    .B(_02862_),
    .Y(_02894_));
 OAI21x1_ASAP7_75t_R _25643_ (.A1(_02623_),
    .A2(_02894_),
    .B(_02333_),
    .Y(_02895_));
 AOI21x1_ASAP7_75t_R _25644_ (.A1(_02528_),
    .A2(_02893_),
    .B(_02895_),
    .Y(_02896_));
 OAI21x1_ASAP7_75t_R _25645_ (.A1(_02891_),
    .A2(_02896_),
    .B(_02471_),
    .Y(_02897_));
 NAND2x1_ASAP7_75t_R _25646_ (.A(net679),
    .B(_02395_),
    .Y(_02898_));
 AO21x1_ASAP7_75t_R _25647_ (.A1(_02501_),
    .A2(_02898_),
    .B(_02509_),
    .Y(_02899_));
 AO21x1_ASAP7_75t_R _25648_ (.A1(_02631_),
    .A2(_02822_),
    .B(_02318_),
    .Y(_02900_));
 AOI21x1_ASAP7_75t_R _25649_ (.A1(_02899_),
    .A2(_02900_),
    .B(_02333_),
    .Y(_02901_));
 NOR2x1_ASAP7_75t_R _25650_ (.A(_02527_),
    .B(_02729_),
    .Y(_02902_));
 AO21x1_ASAP7_75t_R _25651_ (.A1(_02902_),
    .A2(_02837_),
    .B(_02482_),
    .Y(_02903_));
 AOI21x1_ASAP7_75t_R _25652_ (.A1(_02344_),
    .A2(_02304_),
    .B(_02351_),
    .Y(_02904_));
 AOI211x1_ASAP7_75t_R _25653_ (.A1(_02395_),
    .A2(_02426_),
    .B(_02904_),
    .C(_02477_),
    .Y(_02905_));
 OAI21x1_ASAP7_75t_R _25654_ (.A1(_02903_),
    .A2(_02905_),
    .B(_02498_),
    .Y(_02906_));
 NOR2x1_ASAP7_75t_R _25655_ (.A(_02901_),
    .B(_02906_),
    .Y(_02907_));
 OAI22x1_ASAP7_75t_R _25656_ (.A1(_02886_),
    .A2(_02874_),
    .B1(_02897_),
    .B2(_02907_),
    .Y(_00103_));
 NOR2x1_ASAP7_75t_R _25657_ (.A(_11450_),
    .B(_00581_),
    .Y(_02908_));
 XOR2x2_ASAP7_75t_R _25658_ (.A(_11381_),
    .B(_11536_),
    .Y(_02909_));
 INVx1_ASAP7_75t_R _25659_ (.A(net700),
    .Y(_02910_));
 XOR2x1_ASAP7_75t_R _25660_ (.A(_02910_),
    .Y(_02911_),
    .B(net774));
 XOR2x1_ASAP7_75t_R _25661_ (.A(_14322_),
    .Y(_02912_),
    .B(net787));
 NAND2x1_ASAP7_75t_R _25662_ (.A(_02911_),
    .B(_02912_),
    .Y(_02913_));
 XOR2x1_ASAP7_75t_R _25663_ (.A(net701),
    .Y(_02914_),
    .B(net774));
 XOR2x1_ASAP7_75t_R _25664_ (.A(net788),
    .Y(_02915_),
    .B(_14322_));
 NAND2x1_ASAP7_75t_R _25665_ (.A(_02914_),
    .B(_02915_),
    .Y(_02916_));
 AOI21x1_ASAP7_75t_R _25666_ (.A1(_02916_),
    .A2(_02913_),
    .B(_12092_),
    .Y(_02917_));
 OAI21x1_ASAP7_75t_R _25667_ (.A1(_02908_),
    .A2(_02917_),
    .B(net929),
    .Y(_02918_));
 AND2x2_ASAP7_75t_R _25668_ (.A(_11370_),
    .B(_00581_),
    .Y(_02919_));
 NAND2x1_ASAP7_75t_R _25669_ (.A(_02914_),
    .B(_02912_),
    .Y(_02920_));
 NAND2x1_ASAP7_75t_R _25670_ (.A(_02911_),
    .B(_02915_),
    .Y(_02921_));
 AOI21x1_ASAP7_75t_R _25671_ (.A1(_02921_),
    .A2(_02920_),
    .B(_12092_),
    .Y(_02922_));
 INVx1_ASAP7_75t_R _25672_ (.A(net928),
    .Y(_02923_));
 OAI21x1_ASAP7_75t_R _25673_ (.A1(_02919_),
    .A2(_02922_),
    .B(_02923_),
    .Y(_02924_));
 NAND2x2_ASAP7_75t_R _25674_ (.A(_02924_),
    .B(_02918_),
    .Y(_15959_));
 INVx1_ASAP7_75t_R _25675_ (.A(net704),
    .Y(_02925_));
 XOR2x1_ASAP7_75t_R _25676_ (.A(_11362_),
    .Y(_02926_),
    .B(net688));
 NAND2x1_ASAP7_75t_R _25677_ (.A(_02925_),
    .B(_02926_),
    .Y(_02927_));
 XNOR2x1_ASAP7_75t_R _25678_ (.B(net688),
    .Y(_02928_),
    .A(_11362_));
 NAND2x1_ASAP7_75t_R _25679_ (.A(net28),
    .B(_02928_),
    .Y(_02929_));
 INVx2_ASAP7_75t_R _25680_ (.A(net774),
    .Y(_02930_));
 AOI21x1_ASAP7_75t_R _25681_ (.A1(_02927_),
    .A2(_02929_),
    .B(_02930_),
    .Y(_02931_));
 XOR2x1_ASAP7_75t_R _25682_ (.A(net688),
    .Y(_02932_),
    .B(net704));
 NAND2x1_ASAP7_75t_R _25683_ (.A(net19),
    .B(_02932_),
    .Y(_02933_));
 XNOR2x1_ASAP7_75t_R _25684_ (.B(net704),
    .Y(_02934_),
    .A(net688));
 NAND2x1_ASAP7_75t_R _25685_ (.A(_14335_),
    .B(_02934_),
    .Y(_02935_));
 AOI21x1_ASAP7_75t_R _25686_ (.A1(_02933_),
    .A2(_02935_),
    .B(net576),
    .Y(_02936_));
 OAI21x1_ASAP7_75t_R _25687_ (.A1(_02931_),
    .A2(_02936_),
    .B(_12921_),
    .Y(_02937_));
 NOR2x1_ASAP7_75t_R _25688_ (.A(_10762_),
    .B(_00582_),
    .Y(_02938_));
 INVx2_ASAP7_75t_R _25689_ (.A(_02938_),
    .Y(_02939_));
 NAND3x2_ASAP7_75t_R _25690_ (.B(_01057_),
    .C(_02939_),
    .Y(_02940_),
    .A(_02937_));
 AO21x2_ASAP7_75t_R _25691_ (.A1(_02939_),
    .A2(_02937_),
    .B(_01057_),
    .Y(_02941_));
 NAND2x2_ASAP7_75t_R _25692_ (.A(_02941_),
    .B(_02940_),
    .Y(_02942_));
 INVx2_ASAP7_75t_R _25693_ (.A(_02942_),
    .Y(_02943_));
 BUFx12f_ASAP7_75t_R _25694_ (.A(_02943_),
    .Y(_15962_));
 NOR2x1_ASAP7_75t_R _25695_ (.A(net668),
    .B(_00584_),
    .Y(_02944_));
 INVx2_ASAP7_75t_R _25696_ (.A(_02944_),
    .Y(_02945_));
 INVx2_ASAP7_75t_R _25697_ (.A(_11410_),
    .Y(_02946_));
 NOR2x2_ASAP7_75t_R _25698_ (.A(_02946_),
    .B(net694),
    .Y(_02947_));
 XNOR2x2_ASAP7_75t_R _25699_ (.A(_11365_),
    .B(net700),
    .Y(_02948_));
 NOR2x2_ASAP7_75t_R _25700_ (.A(_11410_),
    .B(_02948_),
    .Y(_02949_));
 XOR2x2_ASAP7_75t_R _25701_ (.A(_11433_),
    .B(_11402_),
    .Y(_02950_));
 OAI21x1_ASAP7_75t_R _25702_ (.A1(_02947_),
    .A2(_02949_),
    .B(_02950_),
    .Y(_02951_));
 INVx1_ASAP7_75t_R _25703_ (.A(_02951_),
    .Y(_02952_));
 NOR3x1_ASAP7_75t_R _25704_ (.A(_02949_),
    .B(_02947_),
    .C(_02950_),
    .Y(_02953_));
 OAI21x1_ASAP7_75t_R _25705_ (.A1(_02952_),
    .A2(_02953_),
    .B(net780),
    .Y(_02954_));
 INVx2_ASAP7_75t_R _25706_ (.A(_08108_),
    .Y(_02955_));
 AOI21x1_ASAP7_75t_R _25707_ (.A1(_02945_),
    .A2(_02954_),
    .B(_02955_),
    .Y(_02956_));
 NAND2x1_ASAP7_75t_R _25708_ (.A(_00584_),
    .B(net866),
    .Y(_02957_));
 NAND2x2_ASAP7_75t_R _25709_ (.A(_11410_),
    .B(_02948_),
    .Y(_02958_));
 NAND2x2_ASAP7_75t_R _25710_ (.A(_02946_),
    .B(net694),
    .Y(_02959_));
 INVx2_ASAP7_75t_R _25711_ (.A(_02950_),
    .Y(_02960_));
 NAND3x2_ASAP7_75t_R _25712_ (.B(_02959_),
    .C(_02960_),
    .Y(_02961_),
    .A(_02958_));
 NAND3x2_ASAP7_75t_R _25713_ (.B(net767),
    .C(_02951_),
    .Y(_02962_),
    .A(_02961_));
 AOI21x1_ASAP7_75t_R _25714_ (.A1(_02957_),
    .A2(_02962_),
    .B(_08108_),
    .Y(_02963_));
 NOR2x2_ASAP7_75t_R _25715_ (.A(_02956_),
    .B(_02963_),
    .Y(_02964_));
 BUFx10_ASAP7_75t_R _25716_ (.A(_02964_),
    .Y(_02965_));
 BUFx10_ASAP7_75t_R _25717_ (.A(_02965_),
    .Y(_15970_));
 OAI21x1_ASAP7_75t_R _25718_ (.A1(_02908_),
    .A2(_02917_),
    .B(_02923_),
    .Y(_02966_));
 OAI21x1_ASAP7_75t_R _25719_ (.A1(_02919_),
    .A2(_02922_),
    .B(net929),
    .Y(_02967_));
 NAND2x2_ASAP7_75t_R _25720_ (.A(_02966_),
    .B(_02967_),
    .Y(_15957_));
 AOI21x1_ASAP7_75t_R _25721_ (.A1(_02945_),
    .A2(_02954_),
    .B(_08108_),
    .Y(_02968_));
 AOI21x1_ASAP7_75t_R _25722_ (.A1(_02957_),
    .A2(_02962_),
    .B(_02955_),
    .Y(_02969_));
 NOR2x2_ASAP7_75t_R _25723_ (.A(_02968_),
    .B(_02969_),
    .Y(_02970_));
 BUFx12f_ASAP7_75t_R _25724_ (.A(_02970_),
    .Y(_15967_));
 NAND2x2_ASAP7_75t_R _25725_ (.A(_15957_),
    .B(_02964_),
    .Y(_02971_));
 BUFx10_ASAP7_75t_R _25726_ (.A(_02956_),
    .Y(_02972_));
 OAI21x1_ASAP7_75t_R _25727_ (.A1(_02972_),
    .A2(_02963_),
    .B(net474),
    .Y(_02973_));
 XOR2x1_ASAP7_75t_R _25728_ (.A(_14375_),
    .Y(_02974_),
    .B(_00839_));
 XOR2x2_ASAP7_75t_R _25729_ (.A(_00743_),
    .B(_00775_),
    .Y(_02975_));
 XNOR2x2_ASAP7_75t_R _25730_ (.A(_11410_),
    .B(net615),
    .Y(_02976_));
 XNOR2x2_ASAP7_75t_R _25731_ (.A(_02975_),
    .B(_02976_),
    .Y(_02977_));
 OAI21x1_ASAP7_75t_R _25732_ (.A1(_02974_),
    .A2(_02977_),
    .B(_12921_),
    .Y(_02978_));
 AND2x2_ASAP7_75t_R _25733_ (.A(_02977_),
    .B(_02974_),
    .Y(_02979_));
 NAND2x1_ASAP7_75t_R _25734_ (.A(_00661_),
    .B(net849),
    .Y(_02980_));
 OAI21x1_ASAP7_75t_R _25735_ (.A1(_02978_),
    .A2(_02979_),
    .B(_02980_),
    .Y(_02981_));
 XOR2x2_ASAP7_75t_R _25736_ (.A(_02981_),
    .B(_01029_),
    .Y(_02982_));
 BUFx10_ASAP7_75t_R _25737_ (.A(_02982_),
    .Y(_02983_));
 BUFx6f_ASAP7_75t_R _25738_ (.A(_02983_),
    .Y(_02984_));
 AO21x1_ASAP7_75t_R _25739_ (.A1(_02971_),
    .A2(_02973_),
    .B(_02984_),
    .Y(_02985_));
 XOR2x1_ASAP7_75t_R _25740_ (.A(_00839_),
    .Y(_02986_),
    .B(net615));
 XOR2x2_ASAP7_75t_R _25741_ (.A(_11484_),
    .B(_02986_),
    .Y(_02987_));
 NAND2x1_ASAP7_75t_R _25742_ (.A(_14403_),
    .B(_02987_),
    .Y(_02988_));
 OA21x2_ASAP7_75t_R _25743_ (.A1(_02987_),
    .A2(_14403_),
    .B(net651),
    .Y(_02989_));
 AND2x2_ASAP7_75t_R _25744_ (.A(_11373_),
    .B(_00660_),
    .Y(_02990_));
 AOI21x1_ASAP7_75t_R _25745_ (.A1(_02988_),
    .A2(_02989_),
    .B(_02990_),
    .Y(_02991_));
 XOR2x2_ASAP7_75t_R _25746_ (.A(_02991_),
    .B(_01030_),
    .Y(_02992_));
 INVx6_ASAP7_75t_R _25747_ (.A(_02992_),
    .Y(_02993_));
 BUFx6f_ASAP7_75t_R _25748_ (.A(_02993_),
    .Y(_02994_));
 BUFx6f_ASAP7_75t_R _25749_ (.A(_02994_),
    .Y(_02995_));
 OAI21x1_ASAP7_75t_R _25750_ (.A1(_02968_),
    .A2(_02969_),
    .B(net476),
    .Y(_02996_));
 NAND2x2_ASAP7_75t_R _25751_ (.A(_02983_),
    .B(_02996_),
    .Y(_02997_));
 NAND3x1_ASAP7_75t_R _25752_ (.A(_02985_),
    .B(_02995_),
    .C(_02997_),
    .Y(_02998_));
 OA21x2_ASAP7_75t_R _25753_ (.A1(_02969_),
    .A2(_02968_),
    .B(_00583_),
    .Y(_02999_));
 INVx1_ASAP7_75t_R _25754_ (.A(_02999_),
    .Y(_03000_));
 OAI21x1_ASAP7_75t_R _25755_ (.A1(_02972_),
    .A2(_02963_),
    .B(_00585_),
    .Y(_03001_));
 BUFx4f_ASAP7_75t_R _25756_ (.A(_02983_),
    .Y(_03002_));
 AO21x1_ASAP7_75t_R _25757_ (.A1(_03000_),
    .A2(_03001_),
    .B(_03002_),
    .Y(_03003_));
 NAND2x2_ASAP7_75t_R _25758_ (.A(net543),
    .B(_02965_),
    .Y(_03004_));
 INVx4_ASAP7_75t_R _25759_ (.A(net476),
    .Y(_03005_));
 OAI21x1_ASAP7_75t_R _25760_ (.A1(_02972_),
    .A2(_02963_),
    .B(_03005_),
    .Y(_03006_));
 XOR2x2_ASAP7_75t_R _25761_ (.A(_02981_),
    .B(_08121_),
    .Y(_03007_));
 BUFx6f_ASAP7_75t_R _25762_ (.A(_03007_),
    .Y(_03008_));
 AO21x1_ASAP7_75t_R _25763_ (.A1(_03004_),
    .A2(net33),
    .B(_03008_),
    .Y(_03009_));
 AO21x1_ASAP7_75t_R _25764_ (.A1(_03003_),
    .A2(_03009_),
    .B(_02995_),
    .Y(_03010_));
 INVx1_ASAP7_75t_R _25765_ (.A(_11466_),
    .Y(_03011_));
 XOR2x1_ASAP7_75t_R _25766_ (.A(_11496_),
    .Y(_03012_),
    .B(_11485_));
 NOR2x1_ASAP7_75t_R _25767_ (.A(_03011_),
    .B(_03012_),
    .Y(_03013_));
 XOR2x1_ASAP7_75t_R _25768_ (.A(_11496_),
    .Y(_03014_),
    .B(_00841_));
 NOR2x1_ASAP7_75t_R _25769_ (.A(_11466_),
    .B(_03014_),
    .Y(_03015_));
 OAI21x1_ASAP7_75t_R _25770_ (.A1(_03013_),
    .A2(_03015_),
    .B(net641),
    .Y(_03016_));
 NOR2x1_ASAP7_75t_R _25771_ (.A(net621),
    .B(_00659_),
    .Y(_03017_));
 INVx2_ASAP7_75t_R _25772_ (.A(_03017_),
    .Y(_03018_));
 NAND3x2_ASAP7_75t_R _25773_ (.B(_08139_),
    .C(_03018_),
    .Y(_03019_),
    .A(_03016_));
 AO21x1_ASAP7_75t_R _25774_ (.A1(_03016_),
    .A2(_03018_),
    .B(_08139_),
    .Y(_03020_));
 NAND2x2_ASAP7_75t_R _25775_ (.A(_03019_),
    .B(_03020_),
    .Y(_03021_));
 BUFx6f_ASAP7_75t_R _25776_ (.A(_03021_),
    .Y(_03022_));
 BUFx10_ASAP7_75t_R _25777_ (.A(_03022_),
    .Y(_03023_));
 AOI21x1_ASAP7_75t_R _25778_ (.A1(_02998_),
    .A2(_03010_),
    .B(_03023_),
    .Y(_03024_));
 BUFx6f_ASAP7_75t_R _25779_ (.A(_02942_),
    .Y(_15956_));
 NAND2x2_ASAP7_75t_R _25780_ (.A(_15956_),
    .B(net7),
    .Y(_03025_));
 BUFx10_ASAP7_75t_R _25781_ (.A(_02970_),
    .Y(_03026_));
 AOI21x1_ASAP7_75t_R _25782_ (.A1(_15962_),
    .A2(_03026_),
    .B(_02983_),
    .Y(_03027_));
 NAND2x1_ASAP7_75t_R _25783_ (.A(_03025_),
    .B(_03027_),
    .Y(_03028_));
 INVx1_ASAP7_75t_R _25784_ (.A(_03028_),
    .Y(_03029_));
 BUFx6f_ASAP7_75t_R _25785_ (.A(_03007_),
    .Y(_03030_));
 BUFx6f_ASAP7_75t_R _25786_ (.A(_03030_),
    .Y(_03031_));
 NOR2x2_ASAP7_75t_R _25787_ (.A(_15959_),
    .B(_15962_),
    .Y(_03032_));
 BUFx12_ASAP7_75t_R _25788_ (.A(_02964_),
    .Y(_03033_));
 NOR2x2_ASAP7_75t_R _25789_ (.A(net27),
    .B(_03033_),
    .Y(_03034_));
 NOR2x1_ASAP7_75t_R _25790_ (.A(_03032_),
    .B(_03034_),
    .Y(_03035_));
 BUFx6f_ASAP7_75t_R _25791_ (.A(_02993_),
    .Y(_03036_));
 OAI21x1_ASAP7_75t_R _25792_ (.A1(_03031_),
    .A2(_03035_),
    .B(_03036_),
    .Y(_03037_));
 BUFx10_ASAP7_75t_R _25793_ (.A(_03021_),
    .Y(_03038_));
 OAI21x1_ASAP7_75t_R _25794_ (.A1(_03029_),
    .A2(_03037_),
    .B(_03038_),
    .Y(_03039_));
 INVx3_ASAP7_75t_R _25795_ (.A(_00587_),
    .Y(_03040_));
 OAI21x1_ASAP7_75t_R _25796_ (.A1(_02968_),
    .A2(_02969_),
    .B(_03040_),
    .Y(_03041_));
 AND2x2_ASAP7_75t_R _25797_ (.A(_03041_),
    .B(_03007_),
    .Y(_03042_));
 INVx2_ASAP7_75t_R _25798_ (.A(_00585_),
    .Y(_03043_));
 NOR2x2_ASAP7_75t_R _25799_ (.A(_03043_),
    .B(_15967_),
    .Y(_03044_));
 INVx4_ASAP7_75t_R _25800_ (.A(_02972_),
    .Y(_03045_));
 NAND3x2_ASAP7_75t_R _25801_ (.B(_02955_),
    .C(_02945_),
    .Y(_03046_),
    .A(_02954_));
 INVx1_ASAP7_75t_R _25802_ (.A(_00583_),
    .Y(_03047_));
 AOI21x1_ASAP7_75t_R _25803_ (.A1(_03045_),
    .A2(_03046_),
    .B(_03047_),
    .Y(_03048_));
 BUFx6f_ASAP7_75t_R _25804_ (.A(_02982_),
    .Y(_03049_));
 BUFx10_ASAP7_75t_R _25805_ (.A(_03049_),
    .Y(_03050_));
 OA21x2_ASAP7_75t_R _25806_ (.A1(_03044_),
    .A2(_03048_),
    .B(_03050_),
    .Y(_03051_));
 AOI211x1_ASAP7_75t_R _25807_ (.A1(_02973_),
    .A2(_03042_),
    .B(_03051_),
    .C(_02995_),
    .Y(_03052_));
 XOR2x1_ASAP7_75t_R _25808_ (.A(_00841_),
    .Y(_03053_),
    .B(_00842_));
 XOR2x1_ASAP7_75t_R _25809_ (.A(_03053_),
    .Y(_03054_),
    .B(_00809_));
 XOR2x1_ASAP7_75t_R _25810_ (.A(_03054_),
    .Y(_03055_),
    .B(_11535_));
 NOR2x1_ASAP7_75t_R _25811_ (.A(_10787_),
    .B(_00658_),
    .Y(_03056_));
 AO21x1_ASAP7_75t_R _25812_ (.A1(_03055_),
    .A2(_10786_),
    .B(_03056_),
    .Y(_03057_));
 XOR2x2_ASAP7_75t_R _25813_ (.A(_03057_),
    .B(_08147_),
    .Y(_03058_));
 INVx8_ASAP7_75t_R _25814_ (.A(_03058_),
    .Y(_03059_));
 BUFx10_ASAP7_75t_R _25815_ (.A(_03059_),
    .Y(_03060_));
 OAI21x1_ASAP7_75t_R _25816_ (.A1(_03039_),
    .A2(_03052_),
    .B(_03060_),
    .Y(_03061_));
 NOR2x1_ASAP7_75t_R _25817_ (.A(_03024_),
    .B(_03061_),
    .Y(_03062_));
 NAND2x2_ASAP7_75t_R _25818_ (.A(net27),
    .B(_03026_),
    .Y(_03063_));
 BUFx4f_ASAP7_75t_R _25819_ (.A(_00588_),
    .Y(_03064_));
 INVx2_ASAP7_75t_R _25820_ (.A(_03064_),
    .Y(_03065_));
 AOI21x1_ASAP7_75t_R _25821_ (.A1(_03065_),
    .A2(_02965_),
    .B(_02983_),
    .Y(_03066_));
 NAND2x1_ASAP7_75t_R _25822_ (.A(_03063_),
    .B(_03066_),
    .Y(_03067_));
 BUFx4f_ASAP7_75t_R _25823_ (.A(_01226_),
    .Y(_03068_));
 AOI21x1_ASAP7_75t_R _25824_ (.A1(_03068_),
    .A2(_03033_),
    .B(_03030_),
    .Y(_03069_));
 NAND2x1_ASAP7_75t_R _25825_ (.A(_02973_),
    .B(_03069_),
    .Y(_03070_));
 BUFx6f_ASAP7_75t_R _25826_ (.A(_02992_),
    .Y(_03071_));
 AO21x1_ASAP7_75t_R _25827_ (.A1(_03067_),
    .A2(_03070_),
    .B(_03071_),
    .Y(_03072_));
 AOI21x1_ASAP7_75t_R _25828_ (.A1(net27),
    .A2(_02965_),
    .B(_02983_),
    .Y(_03073_));
 BUFx3_ASAP7_75t_R _25829_ (.A(_01224_),
    .Y(_03074_));
 BUFx10_ASAP7_75t_R _25830_ (.A(_03007_),
    .Y(_03075_));
 AOI21x1_ASAP7_75t_R _25831_ (.A1(_03074_),
    .A2(_03026_),
    .B(_03075_),
    .Y(_03076_));
 OA21x2_ASAP7_75t_R _25832_ (.A1(_03064_),
    .A2(_15967_),
    .B(_03076_),
    .Y(_03077_));
 BUFx6f_ASAP7_75t_R _25833_ (.A(_02992_),
    .Y(_03078_));
 BUFx6f_ASAP7_75t_R _25834_ (.A(_03078_),
    .Y(_03079_));
 OAI21x1_ASAP7_75t_R _25835_ (.A1(_03073_),
    .A2(_03077_),
    .B(_03079_),
    .Y(_03080_));
 INVx1_ASAP7_75t_R _25836_ (.A(_03021_),
    .Y(_03081_));
 BUFx6f_ASAP7_75t_R _25837_ (.A(_03081_),
    .Y(_03082_));
 BUFx10_ASAP7_75t_R _25838_ (.A(_03082_),
    .Y(_03083_));
 AOI21x1_ASAP7_75t_R _25839_ (.A1(_03072_),
    .A2(_03080_),
    .B(_03083_),
    .Y(_03084_));
 AOI21x1_ASAP7_75t_R _25840_ (.A1(_15956_),
    .A2(_02965_),
    .B(_03007_),
    .Y(_03085_));
 INVx1_ASAP7_75t_R _25841_ (.A(_03068_),
    .Y(_03086_));
 AO21x1_ASAP7_75t_R _25842_ (.A1(_03046_),
    .A2(_03045_),
    .B(_03086_),
    .Y(_03087_));
 BUFx4f_ASAP7_75t_R _25843_ (.A(_03087_),
    .Y(_03088_));
 NAND2x1_ASAP7_75t_R _25844_ (.A(_03064_),
    .B(_15970_),
    .Y(_03089_));
 NAND2x2_ASAP7_75t_R _25845_ (.A(net636),
    .B(_03026_),
    .Y(_03090_));
 AOI21x1_ASAP7_75t_R _25846_ (.A1(_03089_),
    .A2(_03090_),
    .B(_03050_),
    .Y(_03091_));
 AOI211x1_ASAP7_75t_R _25847_ (.A1(_03085_),
    .A2(_03088_),
    .B(_03091_),
    .C(_03079_),
    .Y(_03092_));
 AO21x2_ASAP7_75t_R _25848_ (.A1(_03046_),
    .A2(_03045_),
    .B(_00587_),
    .Y(_03093_));
 AO21x2_ASAP7_75t_R _25849_ (.A1(_03085_),
    .A2(_03093_),
    .B(_02994_),
    .Y(_03094_));
 INVx3_ASAP7_75t_R _25850_ (.A(_01223_),
    .Y(_03095_));
 OAI21x1_ASAP7_75t_R _25851_ (.A1(_02972_),
    .A2(_02963_),
    .B(_03095_),
    .Y(_03096_));
 AO21x1_ASAP7_75t_R _25852_ (.A1(_02971_),
    .A2(_03096_),
    .B(_03002_),
    .Y(_03097_));
 INVx1_ASAP7_75t_R _25853_ (.A(_03097_),
    .Y(_03098_));
 OAI21x1_ASAP7_75t_R _25854_ (.A1(_03094_),
    .A2(_03098_),
    .B(_03083_),
    .Y(_03099_));
 BUFx6f_ASAP7_75t_R _25855_ (.A(_03058_),
    .Y(_03100_));
 BUFx10_ASAP7_75t_R _25856_ (.A(_03100_),
    .Y(_03101_));
 OAI21x1_ASAP7_75t_R _25857_ (.A1(_03092_),
    .A2(_03099_),
    .B(_03101_),
    .Y(_03102_));
 XOR2x1_ASAP7_75t_R _25858_ (.A(_14461_),
    .Y(_03103_),
    .B(_11537_));
 XOR2x1_ASAP7_75t_R _25859_ (.A(_03103_),
    .Y(_03104_),
    .B(_11384_));
 NOR2x1_ASAP7_75t_R _25860_ (.A(_11451_),
    .B(_00657_),
    .Y(_03105_));
 AO21x1_ASAP7_75t_R _25861_ (.A1(_03104_),
    .A2(_10831_),
    .B(_03105_),
    .Y(_03106_));
 XOR2x2_ASAP7_75t_R _25862_ (.A(_03106_),
    .B(_01033_),
    .Y(_03107_));
 OAI21x1_ASAP7_75t_R _25863_ (.A1(_03084_),
    .A2(_03102_),
    .B(_03107_),
    .Y(_03108_));
 NOR2x1_ASAP7_75t_R _25864_ (.A(_03078_),
    .B(_03076_),
    .Y(_03109_));
 INVx3_ASAP7_75t_R _25865_ (.A(_03096_),
    .Y(_03110_));
 OAI21x1_ASAP7_75t_R _25866_ (.A1(_03110_),
    .A2(_03044_),
    .B(_03008_),
    .Y(_03111_));
 NAND2x1_ASAP7_75t_R _25867_ (.A(_03109_),
    .B(_03111_),
    .Y(_03112_));
 OAI21x1_ASAP7_75t_R _25868_ (.A1(_02968_),
    .A2(_02969_),
    .B(_03005_),
    .Y(_03113_));
 AOI21x1_ASAP7_75t_R _25869_ (.A1(_15959_),
    .A2(_02970_),
    .B(_02982_),
    .Y(_03114_));
 NAND2x2_ASAP7_75t_R _25870_ (.A(_03113_),
    .B(_03114_),
    .Y(_03115_));
 OAI21x1_ASAP7_75t_R _25871_ (.A1(_02968_),
    .A2(_02969_),
    .B(_03047_),
    .Y(_03116_));
 AOI21x1_ASAP7_75t_R _25872_ (.A1(net27),
    .A2(_03026_),
    .B(_03075_),
    .Y(_03117_));
 BUFx6f_ASAP7_75t_R _25873_ (.A(_02993_),
    .Y(_03118_));
 AOI21x1_ASAP7_75t_R _25874_ (.A1(_03116_),
    .A2(_03117_),
    .B(_03118_),
    .Y(_03119_));
 NAND2x1_ASAP7_75t_R _25875_ (.A(_03115_),
    .B(_03119_),
    .Y(_03120_));
 BUFx10_ASAP7_75t_R _25876_ (.A(_03082_),
    .Y(_03121_));
 AOI21x1_ASAP7_75t_R _25877_ (.A1(_03112_),
    .A2(_03120_),
    .B(_03121_),
    .Y(_03122_));
 INVx1_ASAP7_75t_R _25878_ (.A(_01225_),
    .Y(_03123_));
 OAI21x1_ASAP7_75t_R _25879_ (.A1(_02972_),
    .A2(_02963_),
    .B(_03123_),
    .Y(_03124_));
 BUFx6f_ASAP7_75t_R _25880_ (.A(_02992_),
    .Y(_03125_));
 AOI21x1_ASAP7_75t_R _25881_ (.A1(_03045_),
    .A2(_03046_),
    .B(_03005_),
    .Y(_03126_));
 NOR2x2_ASAP7_75t_R _25882_ (.A(_03075_),
    .B(_03126_),
    .Y(_03127_));
 NOR2x1_ASAP7_75t_R _25883_ (.A(_03127_),
    .B(_03125_),
    .Y(_03128_));
 OAI21x1_ASAP7_75t_R _25884_ (.A1(_03050_),
    .A2(_03124_),
    .B(_03128_),
    .Y(_03129_));
 INVx1_ASAP7_75t_R _25885_ (.A(_03074_),
    .Y(_03130_));
 OAI21x1_ASAP7_75t_R _25886_ (.A1(_02968_),
    .A2(_02969_),
    .B(_03130_),
    .Y(_03131_));
 INVx1_ASAP7_75t_R _25887_ (.A(_03131_),
    .Y(_03132_));
 AO21x1_ASAP7_75t_R _25888_ (.A1(_03132_),
    .A2(_03031_),
    .B(_03022_),
    .Y(_03133_));
 AOI21x1_ASAP7_75t_R _25889_ (.A1(_03094_),
    .A2(_03129_),
    .B(_03133_),
    .Y(_03134_));
 OAI21x1_ASAP7_75t_R _25890_ (.A1(_03134_),
    .A2(_03122_),
    .B(_03101_),
    .Y(_03135_));
 OAI21x1_ASAP7_75t_R _25891_ (.A1(_02972_),
    .A2(_02963_),
    .B(_03064_),
    .Y(_03136_));
 NOR2x2_ASAP7_75t_R _25892_ (.A(_02983_),
    .B(_03136_),
    .Y(_03137_));
 INVx1_ASAP7_75t_R _25893_ (.A(_03137_),
    .Y(_03138_));
 OA21x2_ASAP7_75t_R _25894_ (.A1(_03131_),
    .A2(_03049_),
    .B(_02992_),
    .Y(_03139_));
 NAND2x1_ASAP7_75t_R _25895_ (.A(_03138_),
    .B(_03139_),
    .Y(_03140_));
 BUFx4f_ASAP7_75t_R _25896_ (.A(_03007_),
    .Y(_03141_));
 OA21x2_ASAP7_75t_R _25897_ (.A1(_02969_),
    .A2(_02968_),
    .B(_03095_),
    .Y(_03142_));
 NAND2x1_ASAP7_75t_R _25898_ (.A(_03141_),
    .B(_03142_),
    .Y(_03143_));
 OAI21x1_ASAP7_75t_R _25899_ (.A1(_02972_),
    .A2(_02963_),
    .B(_03043_),
    .Y(_03144_));
 NAND2x1_ASAP7_75t_R _25900_ (.A(_03144_),
    .B(_03085_),
    .Y(_03145_));
 NAND2x1_ASAP7_75t_R _25901_ (.A(_03143_),
    .B(_03145_),
    .Y(_03146_));
 INVx1_ASAP7_75t_R _25902_ (.A(_01228_),
    .Y(_03147_));
 NOR2x1_ASAP7_75t_R _25903_ (.A(_03147_),
    .B(_03030_),
    .Y(_03148_));
 AO21x1_ASAP7_75t_R _25904_ (.A1(_03141_),
    .A2(_03113_),
    .B(_03148_),
    .Y(_03149_));
 AOI21x1_ASAP7_75t_R _25905_ (.A1(_03036_),
    .A2(_03149_),
    .B(_03038_),
    .Y(_03150_));
 OAI21x1_ASAP7_75t_R _25906_ (.A1(_03140_),
    .A2(_03146_),
    .B(_03150_),
    .Y(_03151_));
 AOI21x1_ASAP7_75t_R _25907_ (.A1(_03141_),
    .A2(_02999_),
    .B(_03078_),
    .Y(_03152_));
 NOR2x1_ASAP7_75t_R _25908_ (.A(_03030_),
    .B(_03096_),
    .Y(_03153_));
 NOR2x1_ASAP7_75t_R _25909_ (.A(_03137_),
    .B(_03153_),
    .Y(_03154_));
 AOI21x1_ASAP7_75t_R _25910_ (.A1(_03152_),
    .A2(_03154_),
    .B(_03121_),
    .Y(_03155_));
 OAI21x1_ASAP7_75t_R _25911_ (.A1(_02968_),
    .A2(_02969_),
    .B(_03123_),
    .Y(_03156_));
 BUFx6f_ASAP7_75t_R _25912_ (.A(_03007_),
    .Y(_03157_));
 AO21x1_ASAP7_75t_R _25913_ (.A1(_03136_),
    .A2(_03156_),
    .B(_03157_),
    .Y(_03158_));
 BUFx10_ASAP7_75t_R _25914_ (.A(_02992_),
    .Y(_03159_));
 NAND2x2_ASAP7_75t_R _25915_ (.A(_03157_),
    .B(_03110_),
    .Y(_03160_));
 NAND3x1_ASAP7_75t_R _25916_ (.A(_03158_),
    .B(_03159_),
    .C(_03160_),
    .Y(_03161_));
 AOI21x1_ASAP7_75t_R _25917_ (.A1(_03155_),
    .A2(_03161_),
    .B(_03100_),
    .Y(_03162_));
 AOI21x1_ASAP7_75t_R _25918_ (.A1(_03151_),
    .A2(_03162_),
    .B(_03107_),
    .Y(_03163_));
 NAND2x1_ASAP7_75t_R _25919_ (.A(_03135_),
    .B(_03163_),
    .Y(_03164_));
 OAI21x1_ASAP7_75t_R _25920_ (.A1(_03062_),
    .A2(_03108_),
    .B(_03164_),
    .Y(_00104_));
 AOI21x1_ASAP7_75t_R _25921_ (.A1(_03040_),
    .A2(_02965_),
    .B(_03075_),
    .Y(_03165_));
 NAND2x1_ASAP7_75t_R _25922_ (.A(_03006_),
    .B(_03165_),
    .Y(_03166_));
 AOI21x1_ASAP7_75t_R _25923_ (.A1(_01223_),
    .A2(_02965_),
    .B(_02983_),
    .Y(_03167_));
 NAND2x1_ASAP7_75t_R _25924_ (.A(_03088_),
    .B(_03167_),
    .Y(_03168_));
 AO21x1_ASAP7_75t_R _25925_ (.A1(_03166_),
    .A2(_03168_),
    .B(_03071_),
    .Y(_03169_));
 AO21x1_ASAP7_75t_R _25926_ (.A1(_03073_),
    .A2(_03093_),
    .B(_03127_),
    .Y(_03170_));
 NAND2x1_ASAP7_75t_R _25927_ (.A(_03170_),
    .B(_03079_),
    .Y(_03171_));
 AOI21x1_ASAP7_75t_R _25928_ (.A1(_03169_),
    .A2(_03171_),
    .B(_03023_),
    .Y(_03172_));
 NOR2x2_ASAP7_75t_R _25929_ (.A(_15956_),
    .B(_03026_),
    .Y(_03173_));
 AO21x1_ASAP7_75t_R _25930_ (.A1(_03173_),
    .A2(_03008_),
    .B(_03125_),
    .Y(_03174_));
 INVx1_ASAP7_75t_R _25931_ (.A(_03144_),
    .Y(_03175_));
 OAI21x1_ASAP7_75t_R _25932_ (.A1(_02997_),
    .A2(_03175_),
    .B(_03160_),
    .Y(_03176_));
 OAI21x1_ASAP7_75t_R _25933_ (.A1(_03174_),
    .A2(_03176_),
    .B(_03038_),
    .Y(_03177_));
 AO21x1_ASAP7_75t_R _25934_ (.A1(_03004_),
    .A2(_03063_),
    .B(_03002_),
    .Y(_03178_));
 NAND2x1_ASAP7_75t_R _25935_ (.A(_02971_),
    .B(_03076_),
    .Y(_03179_));
 AND3x1_ASAP7_75t_R _25936_ (.A(_03178_),
    .B(_03071_),
    .C(_03179_),
    .Y(_03180_));
 OAI21x1_ASAP7_75t_R _25937_ (.A1(_03177_),
    .A2(_03180_),
    .B(_03101_),
    .Y(_03181_));
 NOR2x1_ASAP7_75t_R _25938_ (.A(_03181_),
    .B(_03172_),
    .Y(_03182_));
 AOI21x1_ASAP7_75t_R _25939_ (.A1(_03040_),
    .A2(_02970_),
    .B(_02982_),
    .Y(_03183_));
 AOI21x1_ASAP7_75t_R _25940_ (.A1(_03116_),
    .A2(_03183_),
    .B(_02994_),
    .Y(_03184_));
 NOR2x1_ASAP7_75t_R _25941_ (.A(_03030_),
    .B(_03021_),
    .Y(_03185_));
 NAND2x1_ASAP7_75t_R _25942_ (.A(_00589_),
    .B(_03185_),
    .Y(_03186_));
 AND2x2_ASAP7_75t_R _25943_ (.A(_03184_),
    .B(_03186_),
    .Y(_03187_));
 NAND2x2_ASAP7_75t_R _25944_ (.A(net636),
    .B(_03033_),
    .Y(_03188_));
 AO21x1_ASAP7_75t_R _25945_ (.A1(_03027_),
    .A2(_03188_),
    .B(_03022_),
    .Y(_03189_));
 NOR2x2_ASAP7_75t_R _25946_ (.A(net636),
    .B(_15967_),
    .Y(_03190_));
 INVx1_ASAP7_75t_R _25947_ (.A(_03076_),
    .Y(_03191_));
 BUFx10_ASAP7_75t_R _25948_ (.A(_02993_),
    .Y(_03192_));
 OAI21x1_ASAP7_75t_R _25949_ (.A1(_03190_),
    .A2(_03191_),
    .B(_03192_),
    .Y(_03193_));
 NOR2x1_ASAP7_75t_R _25950_ (.A(_15962_),
    .B(_15970_),
    .Y(_03194_));
 AO21x1_ASAP7_75t_R _25951_ (.A1(_15970_),
    .A2(_03043_),
    .B(_03002_),
    .Y(_03195_));
 NOR2x1_ASAP7_75t_R _25952_ (.A(_03078_),
    .B(_03082_),
    .Y(_03196_));
 OAI21x1_ASAP7_75t_R _25953_ (.A1(_03194_),
    .A2(_03195_),
    .B(_03196_),
    .Y(_03197_));
 AOI21x1_ASAP7_75t_R _25954_ (.A1(_03065_),
    .A2(_03033_),
    .B(_03075_),
    .Y(_03198_));
 AND2x2_ASAP7_75t_R _25955_ (.A(_03198_),
    .B(_03093_),
    .Y(_03199_));
 OAI22x1_ASAP7_75t_R _25956_ (.A1(_03189_),
    .A2(_03193_),
    .B1(_03197_),
    .B2(_03199_),
    .Y(_03200_));
 OAI21x1_ASAP7_75t_R _25957_ (.A1(_03187_),
    .A2(_03200_),
    .B(_03060_),
    .Y(_03201_));
 NAND2x1_ASAP7_75t_R _25958_ (.A(_03107_),
    .B(_03201_),
    .Y(_03202_));
 OA21x2_ASAP7_75t_R _25959_ (.A1(_02969_),
    .A2(_02968_),
    .B(_03064_),
    .Y(_03203_));
 NAND2x1_ASAP7_75t_R _25960_ (.A(_03002_),
    .B(_03203_),
    .Y(_03204_));
 NAND2x2_ASAP7_75t_R _25961_ (.A(_03025_),
    .B(_03114_),
    .Y(_03205_));
 AOI21x1_ASAP7_75t_R _25962_ (.A1(_03204_),
    .A2(_03205_),
    .B(_03192_),
    .Y(_03206_));
 NAND2x2_ASAP7_75t_R _25963_ (.A(_15962_),
    .B(_03033_),
    .Y(_03207_));
 AOI21x1_ASAP7_75t_R _25964_ (.A1(_03074_),
    .A2(_15967_),
    .B(_03049_),
    .Y(_03208_));
 NAND2x1_ASAP7_75t_R _25965_ (.A(_03207_),
    .B(_03208_),
    .Y(_03209_));
 NAND2x1_ASAP7_75t_R _25966_ (.A(_02973_),
    .B(_03085_),
    .Y(_03210_));
 AOI21x1_ASAP7_75t_R _25967_ (.A1(_03209_),
    .A2(_03210_),
    .B(_03159_),
    .Y(_03211_));
 OAI21x1_ASAP7_75t_R _25968_ (.A1(_03206_),
    .A2(_03211_),
    .B(_03038_),
    .Y(_03212_));
 BUFx6f_ASAP7_75t_R _25969_ (.A(_02982_),
    .Y(_03213_));
 OA21x2_ASAP7_75t_R _25970_ (.A1(_03131_),
    .A2(_03213_),
    .B(_02993_),
    .Y(_03214_));
 BUFx6f_ASAP7_75t_R _25971_ (.A(_03075_),
    .Y(_03215_));
 NOR2x2_ASAP7_75t_R _25972_ (.A(_15959_),
    .B(_02965_),
    .Y(_03216_));
 AND2x2_ASAP7_75t_R _25973_ (.A(_03049_),
    .B(_00590_),
    .Y(_03217_));
 AOI21x1_ASAP7_75t_R _25974_ (.A1(_03215_),
    .A2(_03216_),
    .B(_03217_),
    .Y(_03218_));
 AOI21x1_ASAP7_75t_R _25975_ (.A1(_03214_),
    .A2(_03218_),
    .B(_03022_),
    .Y(_03219_));
 AOI21x1_ASAP7_75t_R _25976_ (.A1(net475),
    .A2(_03033_),
    .B(_03075_),
    .Y(_03220_));
 NAND2x1_ASAP7_75t_R _25977_ (.A(_03088_),
    .B(_03220_),
    .Y(_03221_));
 NAND3x1_ASAP7_75t_R _25978_ (.A(_03221_),
    .B(_03139_),
    .C(_03138_),
    .Y(_03222_));
 AOI21x1_ASAP7_75t_R _25979_ (.A1(_03219_),
    .A2(_03222_),
    .B(_03100_),
    .Y(_03223_));
 NAND2x1_ASAP7_75t_R _25980_ (.A(_03212_),
    .B(_03223_),
    .Y(_03224_));
 OR3x1_ASAP7_75t_R _25981_ (.A(_15970_),
    .B(_03040_),
    .C(_03049_),
    .Y(_03225_));
 NAND2x2_ASAP7_75t_R _25982_ (.A(net7),
    .B(_02970_),
    .Y(_03226_));
 AOI21x1_ASAP7_75t_R _25983_ (.A1(_03226_),
    .A2(_03069_),
    .B(_03125_),
    .Y(_03227_));
 NAND2x1_ASAP7_75t_R _25984_ (.A(_03225_),
    .B(_03227_),
    .Y(_03228_));
 NOR2x1_ASAP7_75t_R _25985_ (.A(_03074_),
    .B(_03049_),
    .Y(_03229_));
 AOI21x1_ASAP7_75t_R _25986_ (.A1(_15967_),
    .A2(_03229_),
    .B(_03118_),
    .Y(_03230_));
 AOI21x1_ASAP7_75t_R _25987_ (.A1(_03230_),
    .A2(_03166_),
    .B(_03121_),
    .Y(_03231_));
 AOI21x1_ASAP7_75t_R _25988_ (.A1(_03228_),
    .A2(_03231_),
    .B(_03059_),
    .Y(_03232_));
 AO21x1_ASAP7_75t_R _25989_ (.A1(_02973_),
    .A2(_03131_),
    .B(_03141_),
    .Y(_03233_));
 INVx1_ASAP7_75t_R _25990_ (.A(_03001_),
    .Y(_03234_));
 OAI21x1_ASAP7_75t_R _25991_ (.A1(_03234_),
    .A2(_03173_),
    .B(_03031_),
    .Y(_03235_));
 AOI21x1_ASAP7_75t_R _25992_ (.A1(_03233_),
    .A2(_03235_),
    .B(_03071_),
    .Y(_03236_));
 INVx1_ASAP7_75t_R _25993_ (.A(_02996_),
    .Y(_03237_));
 OAI21x1_ASAP7_75t_R _25994_ (.A1(_03237_),
    .A2(_03034_),
    .B(_03031_),
    .Y(_03238_));
 NOR2x2_ASAP7_75t_R _25995_ (.A(net27),
    .B(net7),
    .Y(_03239_));
 OAI21x1_ASAP7_75t_R _25996_ (.A1(_03239_),
    .A2(_03194_),
    .B(_03050_),
    .Y(_03240_));
 AOI21x1_ASAP7_75t_R _25997_ (.A1(_03238_),
    .A2(_03240_),
    .B(_02995_),
    .Y(_03241_));
 OAI21x1_ASAP7_75t_R _25998_ (.A1(_03236_),
    .A2(_03241_),
    .B(_03083_),
    .Y(_03242_));
 AOI21x1_ASAP7_75t_R _25999_ (.A1(_03232_),
    .A2(_03242_),
    .B(_03107_),
    .Y(_03243_));
 NAND2x1_ASAP7_75t_R _26000_ (.A(_03224_),
    .B(_03243_),
    .Y(_03244_));
 OAI21x1_ASAP7_75t_R _26001_ (.A1(_03202_),
    .A2(_03182_),
    .B(_03244_),
    .Y(_00105_));
 INVx1_ASAP7_75t_R _26002_ (.A(_03136_),
    .Y(_03245_));
 NOR2x1_ASAP7_75t_R _26003_ (.A(_03157_),
    .B(_03245_),
    .Y(_03246_));
 AOI21x1_ASAP7_75t_R _26004_ (.A1(_03131_),
    .A2(_03246_),
    .B(_03118_),
    .Y(_03247_));
 NAND2x1_ASAP7_75t_R _26005_ (.A(_03115_),
    .B(_03247_),
    .Y(_03248_));
 NAND2x1_ASAP7_75t_R _26006_ (.A(_03090_),
    .B(_03198_),
    .Y(_03249_));
 NAND2x2_ASAP7_75t_R _26007_ (.A(_03068_),
    .B(_02964_),
    .Y(_03250_));
 NAND2x1_ASAP7_75t_R _26008_ (.A(_03250_),
    .B(_03208_),
    .Y(_03251_));
 AO21x1_ASAP7_75t_R _26009_ (.A1(_03249_),
    .A2(_03251_),
    .B(_03071_),
    .Y(_03252_));
 AOI21x1_ASAP7_75t_R _26010_ (.A1(_03248_),
    .A2(_03252_),
    .B(_03023_),
    .Y(_03253_));
 INVx1_ASAP7_75t_R _26011_ (.A(_03088_),
    .Y(_03254_));
 NAND2x1_ASAP7_75t_R _26012_ (.A(_03213_),
    .B(_03041_),
    .Y(_03255_));
 INVx1_ASAP7_75t_R _26013_ (.A(_03066_),
    .Y(_03256_));
 OAI21x1_ASAP7_75t_R _26014_ (.A1(_03254_),
    .A2(_03255_),
    .B(_03256_),
    .Y(_03257_));
 OAI21x1_ASAP7_75t_R _26015_ (.A1(_02995_),
    .A2(_03257_),
    .B(_03038_),
    .Y(_03258_));
 AOI21x1_ASAP7_75t_R _26016_ (.A1(net7),
    .A2(_03033_),
    .B(_03049_),
    .Y(_03259_));
 NAND2x1_ASAP7_75t_R _26017_ (.A(_03006_),
    .B(_03259_),
    .Y(_03260_));
 INVx1_ASAP7_75t_R _26018_ (.A(_03142_),
    .Y(_03261_));
 NAND2x2_ASAP7_75t_R _26019_ (.A(_02943_),
    .B(_02970_),
    .Y(_03262_));
 NAND3x1_ASAP7_75t_R _26020_ (.A(_03261_),
    .B(_03262_),
    .C(_03050_),
    .Y(_03263_));
 AOI21x1_ASAP7_75t_R _26021_ (.A1(_03260_),
    .A2(_03263_),
    .B(_03071_),
    .Y(_03264_));
 NOR2x1_ASAP7_75t_R _26022_ (.A(_03258_),
    .B(_03264_),
    .Y(_03265_));
 NOR3x1_ASAP7_75t_R _26023_ (.A(_03253_),
    .B(_03265_),
    .C(_03101_),
    .Y(_03266_));
 AO21x1_ASAP7_75t_R _26024_ (.A1(_03006_),
    .A2(_02996_),
    .B(_03141_),
    .Y(_03267_));
 AOI21x1_ASAP7_75t_R _26025_ (.A1(_01225_),
    .A2(_02965_),
    .B(_02983_),
    .Y(_03268_));
 NAND2x1_ASAP7_75t_R _26026_ (.A(_03063_),
    .B(_03268_),
    .Y(_03269_));
 AOI21x1_ASAP7_75t_R _26027_ (.A1(_03267_),
    .A2(_03269_),
    .B(_03192_),
    .Y(_03270_));
 AOI21x1_ASAP7_75t_R _26028_ (.A1(_03045_),
    .A2(_03046_),
    .B(_01225_),
    .Y(_03271_));
 AOI211x1_ASAP7_75t_R _26029_ (.A1(_15970_),
    .A2(net7),
    .B(_03271_),
    .C(_03008_),
    .Y(_03272_));
 NOR2x2_ASAP7_75t_R _26030_ (.A(_03068_),
    .B(_03026_),
    .Y(_03273_));
 OAI21x1_ASAP7_75t_R _26031_ (.A1(net27),
    .A2(_03033_),
    .B(_03157_),
    .Y(_03274_));
 OAI21x1_ASAP7_75t_R _26032_ (.A1(_03273_),
    .A2(_03274_),
    .B(_03118_),
    .Y(_03275_));
 NOR2x1_ASAP7_75t_R _26033_ (.A(_03272_),
    .B(_03275_),
    .Y(_03276_));
 OAI21x1_ASAP7_75t_R _26034_ (.A1(_03270_),
    .A2(_03276_),
    .B(_03023_),
    .Y(_03277_));
 OAI21x1_ASAP7_75t_R _26035_ (.A1(_03271_),
    .A2(_03132_),
    .B(_03215_),
    .Y(_03278_));
 AOI21x1_ASAP7_75t_R _26036_ (.A1(_03074_),
    .A2(_03033_),
    .B(_03075_),
    .Y(_03279_));
 NAND2x1_ASAP7_75t_R _26037_ (.A(_03226_),
    .B(_03279_),
    .Y(_03280_));
 AOI21x1_ASAP7_75t_R _26038_ (.A1(_03278_),
    .A2(_03280_),
    .B(_03036_),
    .Y(_03281_));
 NAND2x1_ASAP7_75t_R _26039_ (.A(_03063_),
    .B(_03279_),
    .Y(_03282_));
 OAI21x1_ASAP7_75t_R _26040_ (.A1(_03271_),
    .A2(_03273_),
    .B(_03215_),
    .Y(_03283_));
 AOI21x1_ASAP7_75t_R _26041_ (.A1(_03282_),
    .A2(_03283_),
    .B(_03071_),
    .Y(_03284_));
 OAI21x1_ASAP7_75t_R _26042_ (.A1(_03281_),
    .A2(_03284_),
    .B(_03121_),
    .Y(_03285_));
 NAND2x1_ASAP7_75t_R _26043_ (.A(_03277_),
    .B(_03285_),
    .Y(_03286_));
 OAI21x1_ASAP7_75t_R _26044_ (.A1(_03060_),
    .A2(_03286_),
    .B(_03107_),
    .Y(_03287_));
 NAND2x1_ASAP7_75t_R _26045_ (.A(_00589_),
    .B(_03008_),
    .Y(_03288_));
 AOI21x1_ASAP7_75t_R _26046_ (.A1(net636),
    .A2(_03026_),
    .B(_03007_),
    .Y(_03289_));
 AOI21x1_ASAP7_75t_R _26047_ (.A1(_03025_),
    .A2(_03289_),
    .B(_02993_),
    .Y(_03290_));
 AOI21x1_ASAP7_75t_R _26048_ (.A1(_03288_),
    .A2(_03290_),
    .B(_03022_),
    .Y(_03291_));
 NAND2x2_ASAP7_75t_R _26049_ (.A(_03049_),
    .B(_03113_),
    .Y(_03292_));
 NOR2x1_ASAP7_75t_R _26050_ (.A(_03048_),
    .B(_03292_),
    .Y(_03293_));
 INVx2_ASAP7_75t_R _26051_ (.A(_03114_),
    .Y(_03294_));
 NOR2x1_ASAP7_75t_R _26052_ (.A(_03044_),
    .B(_03294_),
    .Y(_03295_));
 OAI21x1_ASAP7_75t_R _26053_ (.A1(_03295_),
    .A2(_03293_),
    .B(_03036_),
    .Y(_03296_));
 NAND2x1_ASAP7_75t_R _26054_ (.A(_03291_),
    .B(_03296_),
    .Y(_03297_));
 NAND2x1_ASAP7_75t_R _26055_ (.A(_03147_),
    .B(_03215_),
    .Y(_03298_));
 AO21x1_ASAP7_75t_R _26056_ (.A1(net32),
    .A2(_03136_),
    .B(_03008_),
    .Y(_03299_));
 AOI21x1_ASAP7_75t_R _26057_ (.A1(_03298_),
    .A2(_03299_),
    .B(_03036_),
    .Y(_03300_));
 NAND2x2_ASAP7_75t_R _26058_ (.A(_02971_),
    .B(_03117_),
    .Y(_03301_));
 AOI21x1_ASAP7_75t_R _26059_ (.A1(_03115_),
    .A2(_03301_),
    .B(_03071_),
    .Y(_03302_));
 OAI21x1_ASAP7_75t_R _26060_ (.A1(_03300_),
    .A2(_03302_),
    .B(_03023_),
    .Y(_03303_));
 NAND2x1_ASAP7_75t_R _26061_ (.A(_03303_),
    .B(_03297_),
    .Y(_03304_));
 AND2x2_ASAP7_75t_R _26062_ (.A(_03074_),
    .B(_01223_),
    .Y(_03305_));
 INVx1_ASAP7_75t_R _26063_ (.A(_03305_),
    .Y(_03306_));
 AO21x2_ASAP7_75t_R _26064_ (.A1(_03046_),
    .A2(_03045_),
    .B(_03306_),
    .Y(_03307_));
 INVx1_ASAP7_75t_R _26065_ (.A(_03307_),
    .Y(_03308_));
 NOR2x1_ASAP7_75t_R _26066_ (.A(_03308_),
    .B(_03255_),
    .Y(_03309_));
 AO21x1_ASAP7_75t_R _26067_ (.A1(_03183_),
    .A2(_03116_),
    .B(_03125_),
    .Y(_03310_));
 AO21x1_ASAP7_75t_R _26068_ (.A1(_03006_),
    .A2(_03131_),
    .B(_03008_),
    .Y(_03311_));
 NOR2x2_ASAP7_75t_R _26069_ (.A(_03049_),
    .B(_03001_),
    .Y(_03312_));
 NOR2x1_ASAP7_75t_R _26070_ (.A(_03118_),
    .B(_03312_),
    .Y(_03313_));
 AOI21x1_ASAP7_75t_R _26071_ (.A1(_03311_),
    .A2(_03313_),
    .B(_03121_),
    .Y(_03314_));
 OAI21x1_ASAP7_75t_R _26072_ (.A1(_03309_),
    .A2(_03310_),
    .B(_03314_),
    .Y(_03315_));
 AND2x2_ASAP7_75t_R _26073_ (.A(_02983_),
    .B(_00591_),
    .Y(_03316_));
 NOR2x2_ASAP7_75t_R _26074_ (.A(_03316_),
    .B(_03066_),
    .Y(_03317_));
 NAND2x1_ASAP7_75t_R _26075_ (.A(_03071_),
    .B(_03317_),
    .Y(_03318_));
 OA21x2_ASAP7_75t_R _26076_ (.A1(_01230_),
    .A2(_03002_),
    .B(_02994_),
    .Y(_03319_));
 AOI21x1_ASAP7_75t_R _26077_ (.A1(_03319_),
    .A2(_03249_),
    .B(_03038_),
    .Y(_03320_));
 AOI21x1_ASAP7_75t_R _26078_ (.A1(_03318_),
    .A2(_03320_),
    .B(_03100_),
    .Y(_03321_));
 AOI21x1_ASAP7_75t_R _26079_ (.A1(_03315_),
    .A2(_03321_),
    .B(_03107_),
    .Y(_03322_));
 OAI21x1_ASAP7_75t_R _26080_ (.A1(_03060_),
    .A2(_03304_),
    .B(_03322_),
    .Y(_03323_));
 OAI21x1_ASAP7_75t_R _26081_ (.A1(_03266_),
    .A2(_03287_),
    .B(_03323_),
    .Y(_00106_));
 INVx1_ASAP7_75t_R _26082_ (.A(_03069_),
    .Y(_03324_));
 NAND2x1_ASAP7_75t_R _26083_ (.A(_02973_),
    .B(_03073_),
    .Y(_03325_));
 OA21x2_ASAP7_75t_R _26084_ (.A1(_03324_),
    .A2(_03308_),
    .B(_03325_),
    .Y(_03326_));
 OA21x2_ASAP7_75t_R _26085_ (.A1(_03124_),
    .A2(_03141_),
    .B(_03022_),
    .Y(_03327_));
 AO21x1_ASAP7_75t_R _26086_ (.A1(_03269_),
    .A2(_03327_),
    .B(_03036_),
    .Y(_03328_));
 AOI21x1_ASAP7_75t_R _26087_ (.A1(_03083_),
    .A2(_03326_),
    .B(_03328_),
    .Y(_03329_));
 AO21x1_ASAP7_75t_R _26088_ (.A1(_03185_),
    .A2(_03237_),
    .B(_03153_),
    .Y(_03330_));
 NAND2x1_ASAP7_75t_R _26089_ (.A(_03116_),
    .B(_03081_),
    .Y(_03331_));
 NOR2x2_ASAP7_75t_R _26090_ (.A(_03331_),
    .B(_03294_),
    .Y(_03332_));
 AND3x4_ASAP7_75t_R _26091_ (.A(_03141_),
    .B(_03126_),
    .C(_03021_),
    .Y(_03333_));
 NOR3x2_ASAP7_75t_R _26092_ (.B(_03332_),
    .C(_03330_),
    .Y(_03334_),
    .A(_03333_));
 OAI21x1_ASAP7_75t_R _26093_ (.A1(_03334_),
    .A2(_03079_),
    .B(_03060_),
    .Y(_03335_));
 NOR2x1_ASAP7_75t_R _26094_ (.A(_15962_),
    .B(_03026_),
    .Y(_03336_));
 OAI21x1_ASAP7_75t_R _26095_ (.A1(_03271_),
    .A2(_03336_),
    .B(_03213_),
    .Y(_03337_));
 NOR2x2_ASAP7_75t_R _26096_ (.A(_02982_),
    .B(_03126_),
    .Y(_03338_));
 AOI21x1_ASAP7_75t_R _26097_ (.A1(_03250_),
    .A2(_03338_),
    .B(_03078_),
    .Y(_03339_));
 NAND2x1_ASAP7_75t_R _26098_ (.A(_03339_),
    .B(_03337_),
    .Y(_03340_));
 AOI21x1_ASAP7_75t_R _26099_ (.A1(_03144_),
    .A2(_03085_),
    .B(_02994_),
    .Y(_03341_));
 AOI21x1_ASAP7_75t_R _26100_ (.A1(_03205_),
    .A2(_03341_),
    .B(_03082_),
    .Y(_03342_));
 NAND2x1_ASAP7_75t_R _26101_ (.A(_03342_),
    .B(_03340_),
    .Y(_03343_));
 OAI21x1_ASAP7_75t_R _26102_ (.A1(_02972_),
    .A2(_02963_),
    .B(_03306_),
    .Y(_03344_));
 AO21x1_ASAP7_75t_R _26103_ (.A1(_03156_),
    .A2(_03344_),
    .B(_03157_),
    .Y(_03345_));
 NAND2x1_ASAP7_75t_R _26104_ (.A(_03345_),
    .B(_03184_),
    .Y(_03346_));
 NOR2x1_ASAP7_75t_R _26105_ (.A(_03273_),
    .B(_03274_),
    .Y(_03347_));
 AOI21x1_ASAP7_75t_R _26106_ (.A1(_03036_),
    .A2(_03347_),
    .B(_03022_),
    .Y(_03348_));
 AOI21x1_ASAP7_75t_R _26107_ (.A1(_03346_),
    .A2(_03348_),
    .B(_03059_),
    .Y(_03349_));
 INVx5_ASAP7_75t_R _26108_ (.A(_03107_),
    .Y(_03350_));
 AOI21x1_ASAP7_75t_R _26109_ (.A1(_03343_),
    .A2(_03349_),
    .B(_03350_),
    .Y(_03351_));
 OAI21x1_ASAP7_75t_R _26110_ (.A1(_03335_),
    .A2(_03329_),
    .B(_03351_),
    .Y(_03352_));
 OAI21x1_ASAP7_75t_R _26111_ (.A1(_03032_),
    .A2(_03173_),
    .B(_03141_),
    .Y(_03353_));
 NAND2x1_ASAP7_75t_R _26112_ (.A(_03125_),
    .B(_03353_),
    .Y(_03354_));
 AND3x1_ASAP7_75t_R _26113_ (.A(_02971_),
    .B(_02973_),
    .C(_02984_),
    .Y(_03355_));
 NAND2x1_ASAP7_75t_R _26114_ (.A(_03063_),
    .B(_03259_),
    .Y(_03356_));
 NOR2x1_ASAP7_75t_R _26115_ (.A(_03078_),
    .B(_03220_),
    .Y(_03357_));
 AOI21x1_ASAP7_75t_R _26116_ (.A1(_03356_),
    .A2(_03357_),
    .B(_03022_),
    .Y(_03358_));
 OAI21x1_ASAP7_75t_R _26117_ (.A1(_03354_),
    .A2(_03355_),
    .B(_03358_),
    .Y(_03359_));
 NOR2x1_ASAP7_75t_R _26118_ (.A(_03234_),
    .B(_02997_),
    .Y(_03360_));
 AOI211x1_ASAP7_75t_R _26119_ (.A1(_15970_),
    .A2(_15962_),
    .B(_03048_),
    .C(_03002_),
    .Y(_03361_));
 OAI21x1_ASAP7_75t_R _26120_ (.A1(_03360_),
    .A2(_03361_),
    .B(_03192_),
    .Y(_03362_));
 NAND2x1_ASAP7_75t_R _26121_ (.A(_03088_),
    .B(_03279_),
    .Y(_03363_));
 AOI21x1_ASAP7_75t_R _26122_ (.A1(net33),
    .A2(_03259_),
    .B(_03118_),
    .Y(_03364_));
 AOI21x1_ASAP7_75t_R _26123_ (.A1(_03363_),
    .A2(_03364_),
    .B(_03082_),
    .Y(_03365_));
 NAND2x1_ASAP7_75t_R _26124_ (.A(_03362_),
    .B(_03365_),
    .Y(_03366_));
 AOI21x1_ASAP7_75t_R _26125_ (.A1(_03359_),
    .A2(_03366_),
    .B(_03101_),
    .Y(_03367_));
 OAI21x1_ASAP7_75t_R _26126_ (.A1(_03048_),
    .A2(_03203_),
    .B(_02984_),
    .Y(_03368_));
 NAND2x1_ASAP7_75t_R _26127_ (.A(_02996_),
    .B(_03183_),
    .Y(_03369_));
 AOI21x1_ASAP7_75t_R _26128_ (.A1(_03368_),
    .A2(_03369_),
    .B(_03192_),
    .Y(_03370_));
 OAI21x1_ASAP7_75t_R _26129_ (.A1(net863),
    .A2(_02999_),
    .B(_03215_),
    .Y(_03371_));
 AOI22x1_ASAP7_75t_R _26130_ (.A1(_02918_),
    .A2(_02924_),
    .B1(_02940_),
    .B2(_02941_),
    .Y(_03372_));
 OAI21x1_ASAP7_75t_R _26131_ (.A1(_03372_),
    .A2(_03173_),
    .B(_02984_),
    .Y(_03373_));
 AOI21x1_ASAP7_75t_R _26132_ (.A1(_03371_),
    .A2(_03373_),
    .B(_03159_),
    .Y(_03374_));
 OAI21x1_ASAP7_75t_R _26133_ (.A1(_03370_),
    .A2(_03374_),
    .B(_03038_),
    .Y(_03375_));
 AO21x1_ASAP7_75t_R _26134_ (.A1(_02973_),
    .A2(_03156_),
    .B(_03213_),
    .Y(_03376_));
 NAND2x1_ASAP7_75t_R _26135_ (.A(_03226_),
    .B(_03069_),
    .Y(_03377_));
 AOI21x1_ASAP7_75t_R _26136_ (.A1(_03376_),
    .A2(_03377_),
    .B(_03159_),
    .Y(_03378_));
 INVx1_ASAP7_75t_R _26137_ (.A(_03198_),
    .Y(_03379_));
 AOI21x1_ASAP7_75t_R _26138_ (.A1(_03379_),
    .A2(_03353_),
    .B(_03036_),
    .Y(_03380_));
 OAI21x1_ASAP7_75t_R _26139_ (.A1(_03378_),
    .A2(_03380_),
    .B(_03121_),
    .Y(_03381_));
 AOI21x1_ASAP7_75t_R _26140_ (.A1(_03375_),
    .A2(_03381_),
    .B(_03060_),
    .Y(_03382_));
 OAI21x1_ASAP7_75t_R _26141_ (.A1(_03367_),
    .A2(_03382_),
    .B(_03350_),
    .Y(_03383_));
 NAND2x1_ASAP7_75t_R _26142_ (.A(_03352_),
    .B(_03383_),
    .Y(_00107_));
 NAND2x1_ASAP7_75t_R _26143_ (.A(net636),
    .B(_15962_),
    .Y(_03384_));
 AOI21x1_ASAP7_75t_R _26144_ (.A1(_03384_),
    .A2(_03226_),
    .B(_03002_),
    .Y(_03385_));
 INVx1_ASAP7_75t_R _26145_ (.A(_03385_),
    .Y(_03386_));
 NAND2x1_ASAP7_75t_R _26146_ (.A(_03004_),
    .B(_03289_),
    .Y(_03387_));
 AO21x1_ASAP7_75t_R _26147_ (.A1(_03386_),
    .A2(_03387_),
    .B(_03079_),
    .Y(_03388_));
 NAND2x1_ASAP7_75t_R _26148_ (.A(_03188_),
    .B(_03027_),
    .Y(_03389_));
 AOI21x1_ASAP7_75t_R _26149_ (.A1(_03389_),
    .A2(_03290_),
    .B(_03023_),
    .Y(_03390_));
 AOI21x1_ASAP7_75t_R _26150_ (.A1(_01225_),
    .A2(_02965_),
    .B(_03007_),
    .Y(_03391_));
 OAI21x1_ASAP7_75t_R _26151_ (.A1(_03110_),
    .A2(_03391_),
    .B(_02995_),
    .Y(_03392_));
 AOI21x1_ASAP7_75t_R _26152_ (.A1(_03004_),
    .A2(_03262_),
    .B(_03050_),
    .Y(_03393_));
 AOI21x1_ASAP7_75t_R _26153_ (.A1(_02971_),
    .A2(_03262_),
    .B(_03157_),
    .Y(_03394_));
 OAI21x1_ASAP7_75t_R _26154_ (.A1(_03393_),
    .A2(_03394_),
    .B(_03079_),
    .Y(_03395_));
 AOI21x1_ASAP7_75t_R _26155_ (.A1(_03392_),
    .A2(_03395_),
    .B(_03083_),
    .Y(_03396_));
 AOI211x1_ASAP7_75t_R _26156_ (.A1(_03388_),
    .A2(_03390_),
    .B(_03396_),
    .C(_03060_),
    .Y(_03397_));
 AND3x1_ASAP7_75t_R _26157_ (.A(_02971_),
    .B(_02984_),
    .C(_03144_),
    .Y(_03398_));
 NOR2x1_ASAP7_75t_R _26158_ (.A(_03398_),
    .B(_03140_),
    .Y(_03399_));
 AOI21x1_ASAP7_75t_R _26159_ (.A1(_03065_),
    .A2(_15967_),
    .B(_03030_),
    .Y(_03400_));
 AND2x2_ASAP7_75t_R _26160_ (.A(_03400_),
    .B(_02971_),
    .Y(_03401_));
 AO21x1_ASAP7_75t_R _26161_ (.A1(_03208_),
    .A2(_03250_),
    .B(_03125_),
    .Y(_03402_));
 OAI21x1_ASAP7_75t_R _26162_ (.A1(_03401_),
    .A2(_03402_),
    .B(_03083_),
    .Y(_03403_));
 AO21x1_ASAP7_75t_R _26163_ (.A1(net32),
    .A2(_03124_),
    .B(_03141_),
    .Y(_03404_));
 AOI21x1_ASAP7_75t_R _26164_ (.A1(_03278_),
    .A2(_03404_),
    .B(_03071_),
    .Y(_03405_));
 INVx2_ASAP7_75t_R _26165_ (.A(_03113_),
    .Y(_03406_));
 OA21x2_ASAP7_75t_R _26166_ (.A1(_02963_),
    .A2(_02972_),
    .B(_03086_),
    .Y(_03407_));
 OAI21x1_ASAP7_75t_R _26167_ (.A1(_03406_),
    .A2(_03407_),
    .B(_03031_),
    .Y(_03408_));
 AOI21x1_ASAP7_75t_R _26168_ (.A1(_03158_),
    .A2(_03408_),
    .B(_02995_),
    .Y(_03409_));
 OAI21x1_ASAP7_75t_R _26169_ (.A1(_03405_),
    .A2(_03409_),
    .B(_03023_),
    .Y(_03410_));
 OAI21x1_ASAP7_75t_R _26170_ (.A1(_03399_),
    .A2(_03403_),
    .B(_03410_),
    .Y(_03411_));
 OAI21x1_ASAP7_75t_R _26171_ (.A1(_03101_),
    .A2(_03411_),
    .B(_03350_),
    .Y(_03412_));
 AND3x1_ASAP7_75t_R _26172_ (.A(_03188_),
    .B(_03215_),
    .C(_03144_),
    .Y(_03413_));
 NOR2x1_ASAP7_75t_R _26173_ (.A(_03193_),
    .B(_03413_),
    .Y(_03414_));
 NOR2x2_ASAP7_75t_R _26174_ (.A(_03030_),
    .B(_15967_),
    .Y(_03415_));
 AOI21x1_ASAP7_75t_R _26175_ (.A1(_03250_),
    .A2(_03027_),
    .B(_03415_),
    .Y(_03416_));
 AO21x1_ASAP7_75t_R _26176_ (.A1(_03416_),
    .A2(_03079_),
    .B(_03059_),
    .Y(_03417_));
 OAI21x1_ASAP7_75t_R _26177_ (.A1(_03414_),
    .A2(_03417_),
    .B(_03083_),
    .Y(_03418_));
 NAND2x1_ASAP7_75t_R _26178_ (.A(_03262_),
    .B(_03391_),
    .Y(_03419_));
 AO21x1_ASAP7_75t_R _26179_ (.A1(_03386_),
    .A2(_03419_),
    .B(_03079_),
    .Y(_03420_));
 AO21x1_ASAP7_75t_R _26180_ (.A1(_03262_),
    .A2(_03025_),
    .B(_03215_),
    .Y(_03421_));
 AO21x1_ASAP7_75t_R _26181_ (.A1(_03421_),
    .A2(_03111_),
    .B(_02995_),
    .Y(_03422_));
 AOI21x1_ASAP7_75t_R _26182_ (.A1(_03420_),
    .A2(_03422_),
    .B(_03101_),
    .Y(_03423_));
 OA21x2_ASAP7_75t_R _26183_ (.A1(_03040_),
    .A2(_03002_),
    .B(_03078_),
    .Y(_03424_));
 AOI21x1_ASAP7_75t_R _26184_ (.A1(_03292_),
    .A2(_03424_),
    .B(_03100_),
    .Y(_03425_));
 NAND2x2_ASAP7_75t_R _26185_ (.A(_03226_),
    .B(_03391_),
    .Y(_03426_));
 NOR2x1_ASAP7_75t_R _26186_ (.A(_03125_),
    .B(_03137_),
    .Y(_03427_));
 NAND2x1_ASAP7_75t_R _26187_ (.A(_03426_),
    .B(_03427_),
    .Y(_03428_));
 AOI21x1_ASAP7_75t_R _26188_ (.A1(_03425_),
    .A2(_03428_),
    .B(_03083_),
    .Y(_03429_));
 AND2x2_ASAP7_75t_R _26189_ (.A(_03208_),
    .B(net32),
    .Y(_03430_));
 NOR2x1_ASAP7_75t_R _26190_ (.A(_03165_),
    .B(_03167_),
    .Y(_03431_));
 AOI21x1_ASAP7_75t_R _26191_ (.A1(_02995_),
    .A2(_03431_),
    .B(_03059_),
    .Y(_03432_));
 OAI21x1_ASAP7_75t_R _26192_ (.A1(_03094_),
    .A2(_03430_),
    .B(_03432_),
    .Y(_03433_));
 AOI21x1_ASAP7_75t_R _26193_ (.A1(_03429_),
    .A2(_03433_),
    .B(_03350_),
    .Y(_03434_));
 OAI21x1_ASAP7_75t_R _26194_ (.A1(_03418_),
    .A2(_03423_),
    .B(_03434_),
    .Y(_03435_));
 OAI21x1_ASAP7_75t_R _26195_ (.A1(_03397_),
    .A2(_03412_),
    .B(_03435_),
    .Y(_00108_));
 NAND2x1_ASAP7_75t_R _26196_ (.A(_03050_),
    .B(_15962_),
    .Y(_03436_));
 AOI21x1_ASAP7_75t_R _26197_ (.A1(_03436_),
    .A2(_03028_),
    .B(_02995_),
    .Y(_03437_));
 NAND2x2_ASAP7_75t_R _26198_ (.A(_03226_),
    .B(_03268_),
    .Y(_03438_));
 NAND2x1_ASAP7_75t_R _26199_ (.A(_02973_),
    .B(_03198_),
    .Y(_03439_));
 AOI21x1_ASAP7_75t_R _26200_ (.A1(_03438_),
    .A2(_03439_),
    .B(_03079_),
    .Y(_03440_));
 OAI21x1_ASAP7_75t_R _26201_ (.A1(_03437_),
    .A2(_03440_),
    .B(_03100_),
    .Y(_03441_));
 AOI21x1_ASAP7_75t_R _26202_ (.A1(_03050_),
    .A2(_03307_),
    .B(_03118_),
    .Y(_03442_));
 NAND2x1_ASAP7_75t_R _26203_ (.A(_03093_),
    .B(_03066_),
    .Y(_03443_));
 NAND2x1_ASAP7_75t_R _26204_ (.A(_03442_),
    .B(_03443_),
    .Y(_03444_));
 AOI21x1_ASAP7_75t_R _26205_ (.A1(_03324_),
    .A2(_03214_),
    .B(_03100_),
    .Y(_03445_));
 AOI21x1_ASAP7_75t_R _26206_ (.A1(_03444_),
    .A2(_03445_),
    .B(_03083_),
    .Y(_03446_));
 AO21x1_ASAP7_75t_R _26207_ (.A1(_03441_),
    .A2(_03446_),
    .B(_03350_),
    .Y(_03447_));
 OA21x2_ASAP7_75t_R _26208_ (.A1(_03034_),
    .A2(_03132_),
    .B(_03031_),
    .Y(_03448_));
 AND2x2_ASAP7_75t_R _26209_ (.A(_03183_),
    .B(_03250_),
    .Y(_03449_));
 AO21x1_ASAP7_75t_R _26210_ (.A1(_02999_),
    .A2(_03213_),
    .B(_02992_),
    .Y(_03450_));
 OA21x2_ASAP7_75t_R _26211_ (.A1(_03449_),
    .A2(_03450_),
    .B(_03100_),
    .Y(_03451_));
 OA21x2_ASAP7_75t_R _26212_ (.A1(_03094_),
    .A2(_03448_),
    .B(_03451_),
    .Y(_03452_));
 NAND2x1_ASAP7_75t_R _26213_ (.A(_03116_),
    .B(_03127_),
    .Y(_03453_));
 AO21x1_ASAP7_75t_R _26214_ (.A1(_03086_),
    .A2(_15970_),
    .B(_03126_),
    .Y(_03454_));
 AOI21x1_ASAP7_75t_R _26215_ (.A1(_03031_),
    .A2(_03454_),
    .B(_03125_),
    .Y(_03455_));
 NAND2x1_ASAP7_75t_R _26216_ (.A(_03453_),
    .B(_03455_),
    .Y(_03456_));
 AO21x1_ASAP7_75t_R _26217_ (.A1(_00583_),
    .A2(_03213_),
    .B(_02994_),
    .Y(_03457_));
 OA21x2_ASAP7_75t_R _26218_ (.A1(_03457_),
    .A2(_03183_),
    .B(_03059_),
    .Y(_03458_));
 AO21x1_ASAP7_75t_R _26219_ (.A1(_03456_),
    .A2(_03458_),
    .B(_03023_),
    .Y(_03459_));
 NOR2x1_ASAP7_75t_R _26220_ (.A(_03452_),
    .B(_03459_),
    .Y(_03460_));
 NAND2x1_ASAP7_75t_R _26221_ (.A(_02984_),
    .B(_03406_),
    .Y(_03461_));
 NAND2x1_ASAP7_75t_R _26222_ (.A(_03090_),
    .B(_03167_),
    .Y(_03462_));
 AOI21x1_ASAP7_75t_R _26223_ (.A1(_03461_),
    .A2(_03462_),
    .B(_03159_),
    .Y(_03463_));
 OAI21x1_ASAP7_75t_R _26224_ (.A1(_02984_),
    .A2(_03273_),
    .B(_03125_),
    .Y(_03464_));
 AOI21x1_ASAP7_75t_R _26225_ (.A1(_03127_),
    .A2(_03004_),
    .B(_03464_),
    .Y(_03465_));
 OAI21x1_ASAP7_75t_R _26226_ (.A1(_03463_),
    .A2(_03465_),
    .B(_03060_),
    .Y(_03466_));
 NOR2x1_ASAP7_75t_R _26227_ (.A(_02993_),
    .B(_03338_),
    .Y(_03467_));
 NAND2x1_ASAP7_75t_R _26228_ (.A(_03337_),
    .B(_03467_),
    .Y(_03468_));
 AO21x1_ASAP7_75t_R _26229_ (.A1(_03064_),
    .A2(_15970_),
    .B(_02992_),
    .Y(_03469_));
 OA21x2_ASAP7_75t_R _26230_ (.A1(_03469_),
    .A2(_03208_),
    .B(_03058_),
    .Y(_03470_));
 AOI21x1_ASAP7_75t_R _26231_ (.A1(_03468_),
    .A2(_03470_),
    .B(_03023_),
    .Y(_03471_));
 AOI21x1_ASAP7_75t_R _26232_ (.A1(_03466_),
    .A2(_03471_),
    .B(_03107_),
    .Y(_03472_));
 NAND2x1_ASAP7_75t_R _26233_ (.A(_03384_),
    .B(_03073_),
    .Y(_03473_));
 AO21x1_ASAP7_75t_R _26234_ (.A1(_03026_),
    .A2(_00587_),
    .B(_03075_),
    .Y(_03474_));
 OA21x2_ASAP7_75t_R _26235_ (.A1(_03474_),
    .A2(_02999_),
    .B(_03118_),
    .Y(_03475_));
 AO21x1_ASAP7_75t_R _26236_ (.A1(net7),
    .A2(_03002_),
    .B(_02994_),
    .Y(_03476_));
 OAI21x1_ASAP7_75t_R _26237_ (.A1(_03476_),
    .A2(_03385_),
    .B(_03059_),
    .Y(_03477_));
 AOI21x1_ASAP7_75t_R _26238_ (.A1(_03473_),
    .A2(_03475_),
    .B(_03477_),
    .Y(_03478_));
 AOI21x1_ASAP7_75t_R _26239_ (.A1(_03131_),
    .A2(_03344_),
    .B(_03157_),
    .Y(_03479_));
 AOI21x1_ASAP7_75t_R _26240_ (.A1(_03136_),
    .A2(_03156_),
    .B(_03213_),
    .Y(_03480_));
 OAI21x1_ASAP7_75t_R _26241_ (.A1(_03479_),
    .A2(_03480_),
    .B(_03118_),
    .Y(_03481_));
 NAND2x1_ASAP7_75t_R _26242_ (.A(_03100_),
    .B(_03481_),
    .Y(_03482_));
 NAND2x1_ASAP7_75t_R _26243_ (.A(_03250_),
    .B(_03076_),
    .Y(_03483_));
 AOI21x1_ASAP7_75t_R _26244_ (.A1(_03483_),
    .A2(_03097_),
    .B(_03036_),
    .Y(_03484_));
 NOR2x1_ASAP7_75t_R _26245_ (.A(_03482_),
    .B(_03484_),
    .Y(_03485_));
 OAI21x1_ASAP7_75t_R _26246_ (.A1(_03478_),
    .A2(_03485_),
    .B(_03023_),
    .Y(_03486_));
 NAND2x1_ASAP7_75t_R _26247_ (.A(_03486_),
    .B(_03472_),
    .Y(_03487_));
 OAI21x1_ASAP7_75t_R _26248_ (.A1(_03447_),
    .A2(_03460_),
    .B(_03487_),
    .Y(_00109_));
 AND3x1_ASAP7_75t_R _26249_ (.A(_03307_),
    .B(_03008_),
    .C(net32),
    .Y(_03488_));
 AO21x1_ASAP7_75t_R _26250_ (.A1(_03400_),
    .A2(_03207_),
    .B(_03118_),
    .Y(_03489_));
 AO21x1_ASAP7_75t_R _26251_ (.A1(_03046_),
    .A2(_03045_),
    .B(_03064_),
    .Y(_03490_));
 AOI21x1_ASAP7_75t_R _26252_ (.A1(_15959_),
    .A2(_03033_),
    .B(_03030_),
    .Y(_03491_));
 NAND2x1_ASAP7_75t_R _26253_ (.A(_03490_),
    .B(_03491_),
    .Y(_03492_));
 AOI21x1_ASAP7_75t_R _26254_ (.A1(_03152_),
    .A2(_03492_),
    .B(_03022_),
    .Y(_03493_));
 OAI21x1_ASAP7_75t_R _26255_ (.A1(_03488_),
    .A2(_03489_),
    .B(_03493_),
    .Y(_03494_));
 AO21x1_ASAP7_75t_R _26256_ (.A1(_03157_),
    .A2(net594),
    .B(_02992_),
    .Y(_03495_));
 NOR2x1_ASAP7_75t_R _26257_ (.A(_03495_),
    .B(_03317_),
    .Y(_03496_));
 OAI21x1_ASAP7_75t_R _26258_ (.A1(net594),
    .A2(_03142_),
    .B(_03215_),
    .Y(_03497_));
 NAND2x1_ASAP7_75t_R _26259_ (.A(_03226_),
    .B(_03198_),
    .Y(_03498_));
 AOI21x1_ASAP7_75t_R _26260_ (.A1(_03497_),
    .A2(_03498_),
    .B(_03192_),
    .Y(_03499_));
 OAI21x1_ASAP7_75t_R _26261_ (.A1(_03499_),
    .A2(_03496_),
    .B(_03038_),
    .Y(_03500_));
 AOI21x1_ASAP7_75t_R _26262_ (.A1(_03500_),
    .A2(_03494_),
    .B(_03101_),
    .Y(_03501_));
 NAND2x1_ASAP7_75t_R _26263_ (.A(net32),
    .B(_03027_),
    .Y(_03502_));
 OAI21x1_ASAP7_75t_R _26264_ (.A1(_03030_),
    .A2(_03124_),
    .B(_02993_),
    .Y(_03503_));
 NOR3x1_ASAP7_75t_R _26265_ (.A(_15967_),
    .B(_03075_),
    .C(_03305_),
    .Y(_03504_));
 NOR2x1_ASAP7_75t_R _26266_ (.A(_03503_),
    .B(_03504_),
    .Y(_03505_));
 NAND2x1_ASAP7_75t_R _26267_ (.A(_03502_),
    .B(_03505_),
    .Y(_03506_));
 OAI21x1_ASAP7_75t_R _26268_ (.A1(_03095_),
    .A2(_15970_),
    .B(_03165_),
    .Y(_03507_));
 AOI21x1_ASAP7_75t_R _26269_ (.A1(_03088_),
    .A2(_03268_),
    .B(_02994_),
    .Y(_03508_));
 AOI21x1_ASAP7_75t_R _26270_ (.A1(_03507_),
    .A2(_03508_),
    .B(_03022_),
    .Y(_03509_));
 NAND2x1_ASAP7_75t_R _26271_ (.A(_03506_),
    .B(_03509_),
    .Y(_03510_));
 NOR2x1_ASAP7_75t_R _26272_ (.A(_03239_),
    .B(_03216_),
    .Y(_03511_));
 AND2x2_ASAP7_75t_R _26273_ (.A(_01229_),
    .B(_01227_),
    .Y(_03512_));
 OA21x2_ASAP7_75t_R _26274_ (.A1(_03213_),
    .A2(_03512_),
    .B(_03078_),
    .Y(_03513_));
 OAI21x1_ASAP7_75t_R _26275_ (.A1(_03031_),
    .A2(_03511_),
    .B(_03513_),
    .Y(_03514_));
 INVx1_ASAP7_75t_R _26276_ (.A(_03503_),
    .Y(_03515_));
 AOI21x1_ASAP7_75t_R _26277_ (.A1(_03095_),
    .A2(_03415_),
    .B(_03312_),
    .Y(_03516_));
 AOI21x1_ASAP7_75t_R _26278_ (.A1(_03515_),
    .A2(_03516_),
    .B(_03082_),
    .Y(_03517_));
 NAND2x1_ASAP7_75t_R _26279_ (.A(_03514_),
    .B(_03517_),
    .Y(_03518_));
 AOI21x1_ASAP7_75t_R _26280_ (.A1(_03510_),
    .A2(_03518_),
    .B(_03060_),
    .Y(_03519_));
 OAI21x1_ASAP7_75t_R _26281_ (.A1(_03501_),
    .A2(_03519_),
    .B(_03350_),
    .Y(_03520_));
 AND3x1_ASAP7_75t_R _26282_ (.A(_03250_),
    .B(_02984_),
    .C(net33),
    .Y(_03521_));
 AOI21x1_ASAP7_75t_R _26283_ (.A1(_00592_),
    .A2(_02984_),
    .B(_02994_),
    .Y(_03522_));
 AOI21x1_ASAP7_75t_R _26284_ (.A1(_03522_),
    .A2(_03438_),
    .B(_03082_),
    .Y(_03523_));
 OAI21x1_ASAP7_75t_R _26285_ (.A1(_03174_),
    .A2(_03521_),
    .B(_03523_),
    .Y(_03524_));
 NAND2x1_ASAP7_75t_R _26286_ (.A(_03008_),
    .B(_03116_),
    .Y(_03525_));
 AOI21x1_ASAP7_75t_R _26287_ (.A1(_03525_),
    .A2(_03426_),
    .B(_03159_),
    .Y(_03526_));
 OAI21x1_ASAP7_75t_R _26288_ (.A1(_03247_),
    .A2(_03526_),
    .B(_03121_),
    .Y(_03527_));
 AOI21x1_ASAP7_75t_R _26289_ (.A1(_03524_),
    .A2(_03527_),
    .B(_03101_),
    .Y(_03528_));
 INVx1_ASAP7_75t_R _26290_ (.A(_03217_),
    .Y(_03529_));
 AOI21x1_ASAP7_75t_R _26291_ (.A1(_03529_),
    .A2(_03067_),
    .B(_03125_),
    .Y(_03530_));
 INVx1_ASAP7_75t_R _26292_ (.A(_03006_),
    .Y(_03531_));
 NAND2x1_ASAP7_75t_R _26293_ (.A(_03008_),
    .B(_03531_),
    .Y(_03532_));
 AOI21x1_ASAP7_75t_R _26294_ (.A1(_03532_),
    .A2(_03337_),
    .B(_03192_),
    .Y(_03533_));
 OAI21x1_ASAP7_75t_R _26295_ (.A1(_03530_),
    .A2(_03533_),
    .B(_03121_),
    .Y(_03534_));
 AOI21x1_ASAP7_75t_R _26296_ (.A1(_03068_),
    .A2(_15967_),
    .B(_03049_),
    .Y(_03535_));
 NAND2x1_ASAP7_75t_R _26297_ (.A(_03207_),
    .B(_03535_),
    .Y(_03536_));
 OAI21x1_ASAP7_75t_R _26298_ (.A1(_03372_),
    .A2(_03034_),
    .B(_03050_),
    .Y(_03537_));
 AOI21x1_ASAP7_75t_R _26299_ (.A1(_03536_),
    .A2(_03537_),
    .B(_03159_),
    .Y(_03538_));
 OAI21x1_ASAP7_75t_R _26300_ (.A1(_03203_),
    .A2(_03216_),
    .B(_03215_),
    .Y(_03539_));
 OAI21x1_ASAP7_75t_R _26301_ (.A1(_03032_),
    .A2(_03173_),
    .B(_03050_),
    .Y(_03540_));
 AOI21x1_ASAP7_75t_R _26302_ (.A1(_03539_),
    .A2(_03540_),
    .B(_03036_),
    .Y(_03541_));
 OAI21x1_ASAP7_75t_R _26303_ (.A1(_03538_),
    .A2(_03541_),
    .B(_03038_),
    .Y(_03542_));
 AOI21x1_ASAP7_75t_R _26304_ (.A1(_03534_),
    .A2(_03542_),
    .B(_03060_),
    .Y(_03543_));
 OAI21x1_ASAP7_75t_R _26305_ (.A1(_03528_),
    .A2(_03543_),
    .B(_03107_),
    .Y(_03544_));
 NAND2x1_ASAP7_75t_R _26306_ (.A(_03544_),
    .B(_03520_),
    .Y(_00110_));
 NOR2x1_ASAP7_75t_R _26307_ (.A(_03213_),
    .B(_15962_),
    .Y(_03545_));
 OAI21x1_ASAP7_75t_R _26308_ (.A1(_03545_),
    .A2(_03394_),
    .B(_03192_),
    .Y(_03546_));
 NAND2x1_ASAP7_75t_R _26309_ (.A(_03226_),
    .B(_03042_),
    .Y(_03547_));
 AOI21x1_ASAP7_75t_R _26310_ (.A1(_03290_),
    .A2(_03547_),
    .B(_03058_),
    .Y(_03548_));
 NAND2x1_ASAP7_75t_R _26311_ (.A(_03546_),
    .B(_03548_),
    .Y(_03549_));
 NAND2x1_ASAP7_75t_R _26312_ (.A(_03490_),
    .B(_03073_),
    .Y(_03550_));
 AOI21x1_ASAP7_75t_R _26313_ (.A1(_03144_),
    .A2(_03165_),
    .B(_03078_),
    .Y(_03551_));
 NAND2x1_ASAP7_75t_R _26314_ (.A(_03550_),
    .B(_03551_),
    .Y(_03552_));
 NOR2x1_ASAP7_75t_R _26315_ (.A(_02994_),
    .B(_03535_),
    .Y(_03553_));
 AOI21x1_ASAP7_75t_R _26316_ (.A1(_03426_),
    .A2(_03553_),
    .B(_03059_),
    .Y(_03554_));
 AOI21x1_ASAP7_75t_R _26317_ (.A1(_03552_),
    .A2(_03554_),
    .B(_03121_),
    .Y(_03555_));
 AOI21x1_ASAP7_75t_R _26318_ (.A1(_03549_),
    .A2(_03555_),
    .B(_03350_),
    .Y(_03556_));
 NAND2x1_ASAP7_75t_R _26319_ (.A(_03301_),
    .B(_03508_),
    .Y(_03557_));
 AOI21x1_ASAP7_75t_R _26320_ (.A1(_03088_),
    .A2(_03220_),
    .B(_03078_),
    .Y(_03558_));
 NAND2x1_ASAP7_75t_R _26321_ (.A(_03325_),
    .B(_03558_),
    .Y(_03559_));
 AOI21x1_ASAP7_75t_R _26322_ (.A1(_03557_),
    .A2(_03559_),
    .B(_03059_),
    .Y(_03560_));
 AND2x2_ASAP7_75t_R _26323_ (.A(_03467_),
    .B(_03474_),
    .Y(_03561_));
 AO21x1_ASAP7_75t_R _26324_ (.A1(_03531_),
    .A2(_03157_),
    .B(_02992_),
    .Y(_03562_));
 NOR2x1_ASAP7_75t_R _26325_ (.A(_03400_),
    .B(_03042_),
    .Y(_03563_));
 OAI21x1_ASAP7_75t_R _26326_ (.A1(_03562_),
    .A2(_03563_),
    .B(_03059_),
    .Y(_03564_));
 NOR2x1_ASAP7_75t_R _26327_ (.A(_03561_),
    .B(_03564_),
    .Y(_03565_));
 OAI21x1_ASAP7_75t_R _26328_ (.A1(_03560_),
    .A2(_03565_),
    .B(_03083_),
    .Y(_03566_));
 NAND2x1_ASAP7_75t_R _26329_ (.A(_03566_),
    .B(_03556_),
    .Y(_03567_));
 NOR2x1_ASAP7_75t_R _26330_ (.A(_03021_),
    .B(_03229_),
    .Y(_03568_));
 OAI21x1_ASAP7_75t_R _26331_ (.A1(_03031_),
    .A2(_03511_),
    .B(_03568_),
    .Y(_03569_));
 NAND2x1_ASAP7_75t_R _26332_ (.A(_03041_),
    .B(_03114_),
    .Y(_03570_));
 AOI21x1_ASAP7_75t_R _26333_ (.A1(_03307_),
    .A2(_03391_),
    .B(_03082_),
    .Y(_03571_));
 NAND2x1_ASAP7_75t_R _26334_ (.A(_03570_),
    .B(_03571_),
    .Y(_03572_));
 AOI21x1_ASAP7_75t_R _26335_ (.A1(_03569_),
    .A2(_03572_),
    .B(_03079_),
    .Y(_03573_));
 NAND2x1_ASAP7_75t_R _26336_ (.A(_03041_),
    .B(_03144_),
    .Y(_03574_));
 AOI21x1_ASAP7_75t_R _26337_ (.A1(net33),
    .A2(_03116_),
    .B(_03141_),
    .Y(_03575_));
 AOI211x1_ASAP7_75t_R _26338_ (.A1(_03574_),
    .A2(_03031_),
    .B(_03575_),
    .C(_03082_),
    .Y(_03576_));
 NAND2x1_ASAP7_75t_R _26339_ (.A(_03144_),
    .B(_03082_),
    .Y(_03577_));
 NOR2x1_ASAP7_75t_R _26340_ (.A(_03167_),
    .B(_03491_),
    .Y(_03578_));
 OAI21x1_ASAP7_75t_R _26341_ (.A1(_03577_),
    .A2(_03578_),
    .B(_03159_),
    .Y(_03579_));
 OAI21x1_ASAP7_75t_R _26342_ (.A1(_03576_),
    .A2(_03579_),
    .B(_03100_),
    .Y(_03580_));
 NOR2x1_ASAP7_75t_R _26343_ (.A(_03573_),
    .B(_03580_),
    .Y(_03581_));
 OR2x2_ASAP7_75t_R _26344_ (.A(_01229_),
    .B(_03030_),
    .Y(_03582_));
 AO21x1_ASAP7_75t_R _26345_ (.A1(_02996_),
    .A2(_03124_),
    .B(_03213_),
    .Y(_03583_));
 AOI21x1_ASAP7_75t_R _26346_ (.A1(_03582_),
    .A2(_03583_),
    .B(_03192_),
    .Y(_03584_));
 AO21x1_ASAP7_75t_R _26347_ (.A1(_02973_),
    .A2(_03113_),
    .B(_03157_),
    .Y(_03585_));
 NAND2x1_ASAP7_75t_R _26348_ (.A(_03226_),
    .B(_03073_),
    .Y(_03586_));
 AOI21x1_ASAP7_75t_R _26349_ (.A1(_03585_),
    .A2(_03586_),
    .B(_03159_),
    .Y(_03587_));
 OAI21x1_ASAP7_75t_R _26350_ (.A1(_03584_),
    .A2(_03587_),
    .B(_03121_),
    .Y(_03588_));
 NAND2x1_ASAP7_75t_R _26351_ (.A(_00587_),
    .B(_02984_),
    .Y(_03589_));
 AOI21x1_ASAP7_75t_R _26352_ (.A1(_03589_),
    .A2(_03143_),
    .B(_03192_),
    .Y(_03590_));
 OAI21x1_ASAP7_75t_R _26353_ (.A1(_03245_),
    .A2(_03190_),
    .B(_03215_),
    .Y(_03591_));
 AOI21x1_ASAP7_75t_R _26354_ (.A1(_03179_),
    .A2(_03591_),
    .B(_03159_),
    .Y(_03592_));
 OAI21x1_ASAP7_75t_R _26355_ (.A1(_03590_),
    .A2(_03592_),
    .B(_03038_),
    .Y(_03593_));
 AOI21x1_ASAP7_75t_R _26356_ (.A1(_03588_),
    .A2(_03593_),
    .B(_03101_),
    .Y(_03594_));
 OAI21x1_ASAP7_75t_R _26357_ (.A1(_03581_),
    .A2(_03594_),
    .B(_03350_),
    .Y(_03595_));
 NAND2x1_ASAP7_75t_R _26358_ (.A(_03567_),
    .B(_03595_),
    .Y(_00111_));
 NOR2x2_ASAP7_75t_R _26359_ (.A(net867),
    .B(_00593_),
    .Y(_03596_));
 XOR2x2_ASAP7_75t_R _26360_ (.A(_12104_),
    .B(_12275_),
    .Y(_03597_));
 XOR2x1_ASAP7_75t_R _26361_ (.A(_12097_),
    .Y(_03598_),
    .B(net835));
 XOR2x1_ASAP7_75t_R _26362_ (.A(_12130_),
    .Y(_03599_),
    .B(net903));
 NAND2x1_ASAP7_75t_R _26363_ (.A(_03599_),
    .B(_03598_),
    .Y(_03600_));
 XOR2x1_ASAP7_75t_R _26364_ (.A(net835),
    .Y(_03601_),
    .B(net905));
 XOR2x1_ASAP7_75t_R _26365_ (.A(net903),
    .Y(_03602_),
    .B(_12128_));
 NAND2x1_ASAP7_75t_R _26366_ (.A(_03601_),
    .B(_03602_),
    .Y(_03603_));
 AOI21x1_ASAP7_75t_R _26367_ (.A1(_03600_),
    .A2(_03603_),
    .B(_11374_),
    .Y(_03604_));
 OAI21x1_ASAP7_75t_R _26368_ (.A1(_03596_),
    .A2(_03604_),
    .B(_08099_),
    .Y(_03605_));
 AND2x2_ASAP7_75t_R _26369_ (.A(_10689_),
    .B(_00593_),
    .Y(_03606_));
 NAND2x1_ASAP7_75t_R _26370_ (.A(_03599_),
    .B(_03601_),
    .Y(_03607_));
 NAND2x1_ASAP7_75t_R _26371_ (.A(_03598_),
    .B(_03602_),
    .Y(_03608_));
 AOI21x1_ASAP7_75t_R _26372_ (.A1(_03607_),
    .A2(_03608_),
    .B(_12160_),
    .Y(_03609_));
 INVx1_ASAP7_75t_R _26373_ (.A(_08099_),
    .Y(_03610_));
 OAI21x1_ASAP7_75t_R _26374_ (.A1(_03606_),
    .A2(_03609_),
    .B(_03610_),
    .Y(_03611_));
 NAND2x2_ASAP7_75t_R _26375_ (.A(_03611_),
    .B(_03605_),
    .Y(_15978_));
 INVx1_ASAP7_75t_R _26376_ (.A(net830),
    .Y(_03612_));
 XOR2x1_ASAP7_75t_R _26377_ (.A(net921),
    .Y(_03613_),
    .B(_12115_));
 NAND2x1_ASAP7_75t_R _26378_ (.A(_03612_),
    .B(_03613_),
    .Y(_03614_));
 XNOR2x1_ASAP7_75t_R _26379_ (.B(_12115_),
    .Y(_03615_),
    .A(net921));
 NAND2x1_ASAP7_75t_R _26380_ (.A(net40),
    .B(_03615_),
    .Y(_03616_));
 INVx2_ASAP7_75t_R _26381_ (.A(net835),
    .Y(_03617_));
 AOI21x1_ASAP7_75t_R _26382_ (.A1(_03614_),
    .A2(_03616_),
    .B(_03617_),
    .Y(_03618_));
 XOR2x1_ASAP7_75t_R _26383_ (.A(_12115_),
    .Y(_03619_),
    .B(net830));
 NAND2x1_ASAP7_75t_R _26384_ (.A(net38),
    .B(_03619_),
    .Y(_03620_));
 XNOR2x1_ASAP7_75t_R _26385_ (.B(net830),
    .Y(_03621_),
    .A(_12115_));
 NAND2x1_ASAP7_75t_R _26386_ (.A(_15055_),
    .B(_03621_),
    .Y(_03622_));
 AOI21x1_ASAP7_75t_R _26387_ (.A1(_03620_),
    .A2(_03622_),
    .B(net835),
    .Y(_03623_));
 NOR2x1_ASAP7_75t_R _26388_ (.A(_03623_),
    .B(_03618_),
    .Y(_03624_));
 AND2x2_ASAP7_75t_R _26389_ (.A(_10643_),
    .B(_00594_),
    .Y(_03625_));
 AOI21x1_ASAP7_75t_R _26390_ (.A1(_03624_),
    .A2(_10743_),
    .B(_03625_),
    .Y(_03626_));
 XNOR2x2_ASAP7_75t_R _26391_ (.A(_03626_),
    .B(_01089_),
    .Y(_03627_));
 BUFx12f_ASAP7_75t_R _26392_ (.A(_03627_),
    .Y(_15981_));
 NOR2x2_ASAP7_75t_R _26393_ (.A(net668),
    .B(_00596_),
    .Y(_03628_));
 INVx4_ASAP7_75t_R _26394_ (.A(_03628_),
    .Y(_03629_));
 INVx2_ASAP7_75t_R _26395_ (.A(_12133_),
    .Y(_03630_));
 NOR2x2_ASAP7_75t_R _26396_ (.A(_03630_),
    .B(net899),
    .Y(_03631_));
 XNOR2x2_ASAP7_75t_R _26397_ (.A(_12087_),
    .B(net905),
    .Y(_03632_));
 NOR2x2_ASAP7_75t_R _26398_ (.A(_12133_),
    .B(_03632_),
    .Y(_03633_));
 XOR2x2_ASAP7_75t_R _26399_ (.A(_12169_),
    .B(_12125_),
    .Y(_03634_));
 OAI21x1_ASAP7_75t_R _26400_ (.A1(_03631_),
    .A2(_03633_),
    .B(_03634_),
    .Y(_03635_));
 INVx1_ASAP7_75t_R _26401_ (.A(_03635_),
    .Y(_03636_));
 NOR3x1_ASAP7_75t_R _26402_ (.A(_03633_),
    .B(_03631_),
    .C(_03634_),
    .Y(_03637_));
 OAI21x1_ASAP7_75t_R _26403_ (.A1(_03636_),
    .A2(_03637_),
    .B(_10668_),
    .Y(_03638_));
 AOI21x1_ASAP7_75t_R _26404_ (.A1(_03629_),
    .A2(_03638_),
    .B(_08279_),
    .Y(_03639_));
 BUFx6f_ASAP7_75t_R _26405_ (.A(_03639_),
    .Y(_03640_));
 NAND2x1_ASAP7_75t_R _26406_ (.A(_00596_),
    .B(_11373_),
    .Y(_03641_));
 NAND2x2_ASAP7_75t_R _26407_ (.A(_12133_),
    .B(_03632_),
    .Y(_03642_));
 NAND2x2_ASAP7_75t_R _26408_ (.A(_03630_),
    .B(net779),
    .Y(_03643_));
 INVx3_ASAP7_75t_R _26409_ (.A(_03634_),
    .Y(_03644_));
 NAND3x2_ASAP7_75t_R _26410_ (.B(_03643_),
    .C(_03644_),
    .Y(_03645_),
    .A(_03642_));
 NAND3x2_ASAP7_75t_R _26411_ (.B(_10762_),
    .C(_03635_),
    .Y(_03646_),
    .A(_03645_));
 AOI21x1_ASAP7_75t_R _26412_ (.A1(_03641_),
    .A2(_03646_),
    .B(_08110_),
    .Y(_03647_));
 NOR2x2_ASAP7_75t_R _26413_ (.A(_03647_),
    .B(_03640_),
    .Y(_03648_));
 BUFx12_ASAP7_75t_R _26414_ (.A(_03648_),
    .Y(_15989_));
 OAI21x1_ASAP7_75t_R _26415_ (.A1(_03596_),
    .A2(_03604_),
    .B(_03610_),
    .Y(_03649_));
 OAI21x1_ASAP7_75t_R _26416_ (.A1(_03606_),
    .A2(_03609_),
    .B(_08099_),
    .Y(_03650_));
 NAND2x2_ASAP7_75t_R _26417_ (.A(_03650_),
    .B(_03649_),
    .Y(_03651_));
 BUFx6f_ASAP7_75t_R _26418_ (.A(_03651_),
    .Y(_15976_));
 AOI21x1_ASAP7_75t_R _26419_ (.A1(_03638_),
    .A2(_03629_),
    .B(_08110_),
    .Y(_03652_));
 AOI21x1_ASAP7_75t_R _26420_ (.A1(_03641_),
    .A2(_03646_),
    .B(_08279_),
    .Y(_03653_));
 NOR2x2_ASAP7_75t_R _26421_ (.A(_03652_),
    .B(_03653_),
    .Y(_03654_));
 BUFx10_ASAP7_75t_R _26422_ (.A(_03654_),
    .Y(_03655_));
 BUFx10_ASAP7_75t_R _26423_ (.A(_03655_),
    .Y(_15986_));
 XOR2x2_ASAP7_75t_R _26424_ (.A(_15097_),
    .B(_00847_),
    .Y(_03656_));
 XOR2x2_ASAP7_75t_R _26425_ (.A(_00751_),
    .B(_00783_),
    .Y(_03657_));
 XNOR2x2_ASAP7_75t_R _26426_ (.A(_12133_),
    .B(_12275_),
    .Y(_03658_));
 XNOR2x2_ASAP7_75t_R _26427_ (.A(_03657_),
    .B(_03658_),
    .Y(_03659_));
 OAI21x1_ASAP7_75t_R _26428_ (.A1(_03656_),
    .A2(_03659_),
    .B(_12921_),
    .Y(_03660_));
 AND2x2_ASAP7_75t_R _26429_ (.A(_03659_),
    .B(_03656_),
    .Y(_03661_));
 NAND2x1_ASAP7_75t_R _26430_ (.A(_00684_),
    .B(net849),
    .Y(_03662_));
 OAI21x1_ASAP7_75t_R _26431_ (.A1(_03660_),
    .A2(_03661_),
    .B(_03662_),
    .Y(_03663_));
 XOR2x2_ASAP7_75t_R _26432_ (.A(_03663_),
    .B(_08955_),
    .Y(_03664_));
 BUFx10_ASAP7_75t_R _26433_ (.A(_03664_),
    .Y(_03665_));
 NOR2x2_ASAP7_75t_R _26434_ (.A(net586),
    .B(_03654_),
    .Y(_03666_));
 NAND2x2_ASAP7_75t_R _26435_ (.A(_03665_),
    .B(_03666_),
    .Y(_03667_));
 INVx1_ASAP7_75t_R _26436_ (.A(_03667_),
    .Y(_03668_));
 XOR2x2_ASAP7_75t_R _26437_ (.A(_03663_),
    .B(_01061_),
    .Y(_03669_));
 BUFx10_ASAP7_75t_R _26438_ (.A(_03669_),
    .Y(_03670_));
 OAI21x1_ASAP7_75t_R _26439_ (.A1(net872),
    .A2(_03653_),
    .B(net495),
    .Y(_03671_));
 NAND2x2_ASAP7_75t_R _26440_ (.A(_03670_),
    .B(_03671_),
    .Y(_03672_));
 BUFx6f_ASAP7_75t_R _26441_ (.A(_03664_),
    .Y(_03673_));
 INVx3_ASAP7_75t_R _26442_ (.A(_03640_),
    .Y(_03674_));
 NAND3x2_ASAP7_75t_R _26443_ (.B(_08279_),
    .C(_03629_),
    .Y(_03675_),
    .A(_03638_));
 INVx3_ASAP7_75t_R _26444_ (.A(net495),
    .Y(_03676_));
 AOI21x1_ASAP7_75t_R _26445_ (.A1(_03674_),
    .A2(_03675_),
    .B(_03676_),
    .Y(_03677_));
 NAND2x1_ASAP7_75t_R _26446_ (.A(_03677_),
    .B(_03673_),
    .Y(_03678_));
 NAND2x1_ASAP7_75t_R _26447_ (.A(_03672_),
    .B(_03678_),
    .Y(_03679_));
 XOR2x1_ASAP7_75t_R _26448_ (.A(_15124_),
    .Y(_03680_),
    .B(_00848_));
 XOR2x1_ASAP7_75t_R _26449_ (.A(_00847_),
    .Y(_03681_),
    .B(_12275_));
 XOR2x2_ASAP7_75t_R _26450_ (.A(_12256_),
    .B(_03681_),
    .Y(_03682_));
 NAND2x1_ASAP7_75t_R _26451_ (.A(_03680_),
    .B(_03682_),
    .Y(_03683_));
 OA21x2_ASAP7_75t_R _26452_ (.A1(_03682_),
    .A2(_03680_),
    .B(_10733_),
    .Y(_03684_));
 AND2x2_ASAP7_75t_R _26453_ (.A(_10640_),
    .B(_00683_),
    .Y(_03685_));
 AOI21x1_ASAP7_75t_R _26454_ (.A1(_03683_),
    .A2(_03684_),
    .B(_03685_),
    .Y(_03686_));
 XNOR2x2_ASAP7_75t_R _26455_ (.A(_01062_),
    .B(_03686_),
    .Y(_03687_));
 BUFx10_ASAP7_75t_R _26456_ (.A(_03687_),
    .Y(_03688_));
 OAI21x1_ASAP7_75t_R _26457_ (.A1(_03668_),
    .A2(_03679_),
    .B(_03688_),
    .Y(_03689_));
 OA21x2_ASAP7_75t_R _26458_ (.A1(_03647_),
    .A2(_03640_),
    .B(_03676_),
    .Y(_03690_));
 INVx2_ASAP7_75t_R _26459_ (.A(net512),
    .Y(_03691_));
 NOR2x2_ASAP7_75t_R _26460_ (.A(_03691_),
    .B(_03655_),
    .Y(_03692_));
 BUFx10_ASAP7_75t_R _26461_ (.A(_03669_),
    .Y(_03693_));
 BUFx6f_ASAP7_75t_R _26462_ (.A(_03693_),
    .Y(_03694_));
 OAI21x1_ASAP7_75t_R _26463_ (.A1(_03690_),
    .A2(_03692_),
    .B(_03694_),
    .Y(_03695_));
 OAI21x1_ASAP7_75t_R _26464_ (.A1(net874),
    .A2(_03653_),
    .B(_00595_),
    .Y(_03696_));
 NOR2x2_ASAP7_75t_R _26465_ (.A(_03670_),
    .B(_03696_),
    .Y(_03697_));
 OAI21x1_ASAP7_75t_R _26466_ (.A1(_03640_),
    .A2(_03647_),
    .B(_00597_),
    .Y(_03698_));
 XOR2x2_ASAP7_75t_R _26467_ (.A(_03686_),
    .B(_01062_),
    .Y(_03699_));
 OAI21x1_ASAP7_75t_R _26468_ (.A1(_03670_),
    .A2(_03698_),
    .B(_03699_),
    .Y(_03700_));
 NOR2x1_ASAP7_75t_R _26469_ (.A(_03697_),
    .B(_03700_),
    .Y(_03701_));
 NOR2x1_ASAP7_75t_R _26470_ (.A(net641),
    .B(_00682_),
    .Y(_03702_));
 INVx1_ASAP7_75t_R _26471_ (.A(_03702_),
    .Y(_03703_));
 INVx1_ASAP7_75t_R _26472_ (.A(_12188_),
    .Y(_03704_));
 XOR2x1_ASAP7_75t_R _26473_ (.A(_12219_),
    .Y(_03705_),
    .B(_12260_));
 NOR2x1_ASAP7_75t_R _26474_ (.A(_03704_),
    .B(_03705_),
    .Y(_03706_));
 XOR2x1_ASAP7_75t_R _26475_ (.A(_12219_),
    .Y(_03707_),
    .B(_12259_));
 NOR2x1_ASAP7_75t_R _26476_ (.A(_12188_),
    .B(_03707_),
    .Y(_03708_));
 OAI21x1_ASAP7_75t_R _26477_ (.A1(_03706_),
    .A2(_03708_),
    .B(_11450_),
    .Y(_03709_));
 NAND2x1_ASAP7_75t_R _26478_ (.A(_03703_),
    .B(_03709_),
    .Y(_03710_));
 XOR2x2_ASAP7_75t_R _26479_ (.A(_03710_),
    .B(_01063_),
    .Y(_03711_));
 INVx3_ASAP7_75t_R _26480_ (.A(_03711_),
    .Y(_03712_));
 BUFx6f_ASAP7_75t_R _26481_ (.A(_03712_),
    .Y(_03713_));
 AOI21x1_ASAP7_75t_R _26482_ (.A1(_03695_),
    .A2(_03701_),
    .B(_03713_),
    .Y(_03714_));
 XOR2x1_ASAP7_75t_R _26483_ (.A(_12259_),
    .Y(_03715_),
    .B(_00850_));
 XOR2x1_ASAP7_75t_R _26484_ (.A(_03715_),
    .Y(_03716_),
    .B(_00817_));
 XOR2x1_ASAP7_75t_R _26485_ (.A(_03716_),
    .Y(_03717_),
    .B(_12274_));
 NOR2x1_ASAP7_75t_R _26486_ (.A(_10734_),
    .B(_00681_),
    .Y(_03718_));
 AO21x1_ASAP7_75t_R _26487_ (.A1(_03717_),
    .A2(_10829_),
    .B(_03718_),
    .Y(_03719_));
 XOR2x2_ASAP7_75t_R _26488_ (.A(_03719_),
    .B(_01064_),
    .Y(_03720_));
 CKINVDCx6p67_ASAP7_75t_R _26489_ (.A(_03720_),
    .Y(_03721_));
 AOI21x1_ASAP7_75t_R _26490_ (.A1(_03689_),
    .A2(_03714_),
    .B(_03721_),
    .Y(_03722_));
 INVx1_ASAP7_75t_R _26491_ (.A(_00595_),
    .Y(_03723_));
 AOI21x1_ASAP7_75t_R _26492_ (.A1(_03674_),
    .A2(_03675_),
    .B(_03723_),
    .Y(_03724_));
 OAI21x1_ASAP7_75t_R _26493_ (.A1(_03724_),
    .A2(_03692_),
    .B(_03694_),
    .Y(_03725_));
 NAND3x2_ASAP7_75t_R _26494_ (.B(_08110_),
    .C(_03629_),
    .Y(_03726_),
    .A(_03638_));
 INVx2_ASAP7_75t_R _26495_ (.A(net872),
    .Y(_03727_));
 AO21x2_ASAP7_75t_R _26496_ (.A1(_03726_),
    .A2(_03727_),
    .B(_00599_),
    .Y(_03728_));
 NOR2x2_ASAP7_75t_R _26497_ (.A(_03670_),
    .B(_03677_),
    .Y(_03729_));
 NAND2x1_ASAP7_75t_R _26498_ (.A(_03728_),
    .B(_03729_),
    .Y(_03730_));
 AOI21x1_ASAP7_75t_R _26499_ (.A1(_03725_),
    .A2(_03730_),
    .B(_03688_),
    .Y(_03731_));
 XOR2x2_ASAP7_75t_R _26500_ (.A(_01089_),
    .B(_03626_),
    .Y(_03732_));
 NAND2x2_ASAP7_75t_R _26501_ (.A(net831),
    .B(_15976_),
    .Y(_03733_));
 AOI21x1_ASAP7_75t_R _26502_ (.A1(_03627_),
    .A2(_03655_),
    .B(_03693_),
    .Y(_03734_));
 NAND2x1_ASAP7_75t_R _26503_ (.A(_03733_),
    .B(_03734_),
    .Y(_03735_));
 NAND2x2_ASAP7_75t_R _26504_ (.A(_03627_),
    .B(_03655_),
    .Y(_03736_));
 BUFx6f_ASAP7_75t_R _26505_ (.A(_03664_),
    .Y(_03737_));
 AO21x1_ASAP7_75t_R _26506_ (.A1(_03736_),
    .A2(_03733_),
    .B(_03737_),
    .Y(_03738_));
 BUFx10_ASAP7_75t_R _26507_ (.A(_03699_),
    .Y(_03739_));
 AOI21x1_ASAP7_75t_R _26508_ (.A1(_03735_),
    .A2(_03738_),
    .B(_03739_),
    .Y(_03740_));
 BUFx10_ASAP7_75t_R _26509_ (.A(_03712_),
    .Y(_03741_));
 OAI21x1_ASAP7_75t_R _26510_ (.A1(_03740_),
    .A2(_03731_),
    .B(_03741_),
    .Y(_03742_));
 NAND2x1_ASAP7_75t_R _26511_ (.A(_03742_),
    .B(_03722_),
    .Y(_03743_));
 BUFx3_ASAP7_75t_R _26512_ (.A(_01232_),
    .Y(_03744_));
 AOI21x1_ASAP7_75t_R _26513_ (.A1(_03674_),
    .A2(_03675_),
    .B(_03744_),
    .Y(_03745_));
 OA21x2_ASAP7_75t_R _26514_ (.A1(_03653_),
    .A2(net873),
    .B(_00600_),
    .Y(_03746_));
 BUFx10_ASAP7_75t_R _26515_ (.A(_03670_),
    .Y(_03747_));
 OAI21x1_ASAP7_75t_R _26516_ (.A1(_03745_),
    .A2(_03746_),
    .B(_03747_),
    .Y(_03748_));
 BUFx6f_ASAP7_75t_R _26517_ (.A(_03687_),
    .Y(_03749_));
 BUFx12f_ASAP7_75t_R _26518_ (.A(_03732_),
    .Y(_15975_));
 AOI21x1_ASAP7_75t_R _26519_ (.A1(_15975_),
    .A2(net924),
    .B(_03693_),
    .Y(_03750_));
 NOR2x1_ASAP7_75t_R _26520_ (.A(_03749_),
    .B(_03750_),
    .Y(_03751_));
 BUFx6f_ASAP7_75t_R _26521_ (.A(_03711_),
    .Y(_03752_));
 BUFx6f_ASAP7_75t_R _26522_ (.A(_03752_),
    .Y(_03753_));
 AOI21x1_ASAP7_75t_R _26523_ (.A1(_03748_),
    .A2(_03751_),
    .B(_03753_),
    .Y(_03754_));
 BUFx6f_ASAP7_75t_R _26524_ (.A(_03648_),
    .Y(_03755_));
 AOI21x1_ASAP7_75t_R _26525_ (.A1(_01234_),
    .A2(_03755_),
    .B(_03665_),
    .Y(_03756_));
 INVx1_ASAP7_75t_R _26526_ (.A(_03756_),
    .Y(_03757_));
 BUFx12_ASAP7_75t_R _26527_ (.A(_03654_),
    .Y(_03758_));
 NAND2x2_ASAP7_75t_R _26528_ (.A(net833),
    .B(_03758_),
    .Y(_03759_));
 INVx2_ASAP7_75t_R _26529_ (.A(_00600_),
    .Y(_03760_));
 AOI21x1_ASAP7_75t_R _26530_ (.A1(_03760_),
    .A2(_03755_),
    .B(_03693_),
    .Y(_03761_));
 BUFx6f_ASAP7_75t_R _26531_ (.A(_03699_),
    .Y(_03762_));
 AOI21x1_ASAP7_75t_R _26532_ (.A1(_03759_),
    .A2(_03761_),
    .B(_03762_),
    .Y(_03763_));
 OAI21x1_ASAP7_75t_R _26533_ (.A1(_03677_),
    .A2(_03757_),
    .B(_03763_),
    .Y(_03764_));
 BUFx10_ASAP7_75t_R _26534_ (.A(_03720_),
    .Y(_03765_));
 AOI21x1_ASAP7_75t_R _26535_ (.A1(_03754_),
    .A2(_03764_),
    .B(_03765_),
    .Y(_03766_));
 AOI21x1_ASAP7_75t_R _26536_ (.A1(_15975_),
    .A2(_03755_),
    .B(_03665_),
    .Y(_03767_));
 INVx3_ASAP7_75t_R _26537_ (.A(_00599_),
    .Y(_03768_));
 OAI21x1_ASAP7_75t_R _26538_ (.A1(_03640_),
    .A2(_03647_),
    .B(_03768_),
    .Y(_03769_));
 AND2x2_ASAP7_75t_R _26539_ (.A(_03767_),
    .B(net915),
    .Y(_03770_));
 BUFx10_ASAP7_75t_R _26540_ (.A(_03664_),
    .Y(_03771_));
 INVx1_ASAP7_75t_R _26541_ (.A(_01231_),
    .Y(_03772_));
 OAI21x1_ASAP7_75t_R _26542_ (.A1(_03640_),
    .A2(_03647_),
    .B(_03772_),
    .Y(_03773_));
 INVx2_ASAP7_75t_R _26543_ (.A(_03773_),
    .Y(_03774_));
 BUFx6f_ASAP7_75t_R _26544_ (.A(_03687_),
    .Y(_03775_));
 AOI21x1_ASAP7_75t_R _26545_ (.A1(_03771_),
    .A2(_03774_),
    .B(_03775_),
    .Y(_03776_));
 NAND2x1_ASAP7_75t_R _26546_ (.A(_03776_),
    .B(_03667_),
    .Y(_03777_));
 INVx1_ASAP7_75t_R _26547_ (.A(_01234_),
    .Y(_03778_));
 AO21x2_ASAP7_75t_R _26548_ (.A1(_03675_),
    .A2(_03674_),
    .B(_03778_),
    .Y(_03779_));
 NAND2x1_ASAP7_75t_R _26549_ (.A(_03779_),
    .B(_03767_),
    .Y(_03780_));
 NAND2x2_ASAP7_75t_R _26550_ (.A(net832),
    .B(_03655_),
    .Y(_03781_));
 AOI21x1_ASAP7_75t_R _26551_ (.A1(_03781_),
    .A2(_03761_),
    .B(_03762_),
    .Y(_03782_));
 AOI21x1_ASAP7_75t_R _26552_ (.A1(_03780_),
    .A2(_03782_),
    .B(_03713_),
    .Y(_03783_));
 OAI21x1_ASAP7_75t_R _26553_ (.A1(_03770_),
    .A2(_03777_),
    .B(_03783_),
    .Y(_03784_));
 XOR2x1_ASAP7_75t_R _26554_ (.A(_15151_),
    .Y(_03785_),
    .B(_12276_));
 XOR2x1_ASAP7_75t_R _26555_ (.A(_03785_),
    .Y(_03786_),
    .B(_12106_));
 NOR2x1_ASAP7_75t_R _26556_ (.A(_11451_),
    .B(_00680_),
    .Y(_03787_));
 AO21x1_ASAP7_75t_R _26557_ (.A1(_03786_),
    .A2(_10831_),
    .B(_03787_),
    .Y(_03788_));
 XOR2x2_ASAP7_75t_R _26558_ (.A(_03788_),
    .B(_01065_),
    .Y(_03789_));
 CKINVDCx5p33_ASAP7_75t_R _26559_ (.A(_03789_),
    .Y(_03790_));
 AOI21x1_ASAP7_75t_R _26560_ (.A1(_03766_),
    .A2(_03784_),
    .B(_03790_),
    .Y(_03791_));
 NAND2x1_ASAP7_75t_R _26561_ (.A(_03791_),
    .B(_03743_),
    .Y(_03792_));
 AOI21x1_ASAP7_75t_R _26562_ (.A1(net916),
    .A2(_03767_),
    .B(_03749_),
    .Y(_03793_));
 INVx2_ASAP7_75t_R _26563_ (.A(_03793_),
    .Y(_03794_));
 OAI21x1_ASAP7_75t_R _26564_ (.A1(_03640_),
    .A2(_03647_),
    .B(net622),
    .Y(_03795_));
 NAND2x2_ASAP7_75t_R _26565_ (.A(_03795_),
    .B(_03693_),
    .Y(_03796_));
 INVx2_ASAP7_75t_R _26566_ (.A(_01233_),
    .Y(_03797_));
 OAI21x1_ASAP7_75t_R _26567_ (.A1(_03640_),
    .A2(_03647_),
    .B(_03797_),
    .Y(_03798_));
 BUFx6f_ASAP7_75t_R _26568_ (.A(_03669_),
    .Y(_03799_));
 OA21x2_ASAP7_75t_R _26569_ (.A1(_03798_),
    .A2(_03799_),
    .B(_03775_),
    .Y(_03800_));
 NAND2x1_ASAP7_75t_R _26570_ (.A(_03796_),
    .B(_03800_),
    .Y(_03801_));
 INVx2_ASAP7_75t_R _26571_ (.A(_03744_),
    .Y(_03802_));
 OAI21x1_ASAP7_75t_R _26572_ (.A1(net872),
    .A2(_03653_),
    .B(_03802_),
    .Y(_03803_));
 INVx1_ASAP7_75t_R _26573_ (.A(_03803_),
    .Y(_03804_));
 BUFx10_ASAP7_75t_R _26574_ (.A(_03665_),
    .Y(_03805_));
 AO21x1_ASAP7_75t_R _26575_ (.A1(_03804_),
    .A2(_03805_),
    .B(_03712_),
    .Y(_03806_));
 AOI21x1_ASAP7_75t_R _26576_ (.A1(_03794_),
    .A2(_03801_),
    .B(_03806_),
    .Y(_03807_));
 OAI21x1_ASAP7_75t_R _26577_ (.A1(net872),
    .A2(_03653_),
    .B(_03676_),
    .Y(_03808_));
 AOI21x1_ASAP7_75t_R _26578_ (.A1(net587),
    .A2(_03655_),
    .B(_03693_),
    .Y(_03809_));
 NAND2x2_ASAP7_75t_R _26579_ (.A(_03809_),
    .B(net836),
    .Y(_03810_));
 OAI21x1_ASAP7_75t_R _26580_ (.A1(net872),
    .A2(_03653_),
    .B(_03723_),
    .Y(_03811_));
 AOI21x1_ASAP7_75t_R _26581_ (.A1(_15975_),
    .A2(_03655_),
    .B(_03665_),
    .Y(_03812_));
 BUFx6f_ASAP7_75t_R _26582_ (.A(_03687_),
    .Y(_03813_));
 AOI21x1_ASAP7_75t_R _26583_ (.A1(_03811_),
    .A2(_03812_),
    .B(_03813_),
    .Y(_03814_));
 NAND2x1_ASAP7_75t_R _26584_ (.A(_03810_),
    .B(_03814_),
    .Y(_03815_));
 BUFx6f_ASAP7_75t_R _26585_ (.A(_03665_),
    .Y(_03816_));
 OAI21x1_ASAP7_75t_R _26586_ (.A1(_03774_),
    .A2(_03692_),
    .B(_03816_),
    .Y(_03817_));
 NOR2x1_ASAP7_75t_R _26587_ (.A(_03802_),
    .B(_03755_),
    .Y(_03818_));
 OA21x2_ASAP7_75t_R _26588_ (.A1(_03818_),
    .A2(_03737_),
    .B(_03749_),
    .Y(_03819_));
 NAND2x1_ASAP7_75t_R _26589_ (.A(_03817_),
    .B(_03819_),
    .Y(_03820_));
 BUFx10_ASAP7_75t_R _26590_ (.A(_03752_),
    .Y(_03821_));
 AOI21x1_ASAP7_75t_R _26591_ (.A1(_03815_),
    .A2(_03820_),
    .B(_03821_),
    .Y(_03822_));
 BUFx10_ASAP7_75t_R _26592_ (.A(_03721_),
    .Y(_03823_));
 OAI21x1_ASAP7_75t_R _26593_ (.A1(_03807_),
    .A2(_03822_),
    .B(_03823_),
    .Y(_03824_));
 BUFx6f_ASAP7_75t_R _26594_ (.A(_03699_),
    .Y(_03825_));
 NOR2x1_ASAP7_75t_R _26595_ (.A(_03825_),
    .B(_03697_),
    .Y(_03826_));
 INVx1_ASAP7_75t_R _26596_ (.A(_03826_),
    .Y(_03827_));
 BUFx6f_ASAP7_75t_R _26597_ (.A(_03673_),
    .Y(_03828_));
 OAI21x1_ASAP7_75t_R _26598_ (.A1(_03640_),
    .A2(_03647_),
    .B(_00600_),
    .Y(_03829_));
 INVx2_ASAP7_75t_R _26599_ (.A(_03829_),
    .Y(_03830_));
 NOR2x1_ASAP7_75t_R _26600_ (.A(_03673_),
    .B(_03773_),
    .Y(_03831_));
 AO21x1_ASAP7_75t_R _26601_ (.A1(_03828_),
    .A2(_03830_),
    .B(_03831_),
    .Y(_03832_));
 AO21x2_ASAP7_75t_R _26602_ (.A1(_03675_),
    .A2(_03674_),
    .B(_00600_),
    .Y(_03833_));
 OAI21x1_ASAP7_75t_R _26603_ (.A1(_03797_),
    .A2(_03655_),
    .B(_03669_),
    .Y(_03834_));
 INVx2_ASAP7_75t_R _26604_ (.A(_03834_),
    .Y(_03835_));
 NAND2x1_ASAP7_75t_R _26605_ (.A(_03833_),
    .B(_03835_),
    .Y(_03836_));
 AOI21x1_ASAP7_75t_R _26606_ (.A1(_03776_),
    .A2(_03836_),
    .B(_03753_),
    .Y(_03837_));
 OAI21x1_ASAP7_75t_R _26607_ (.A1(_03827_),
    .A2(_03832_),
    .B(_03837_),
    .Y(_03838_));
 BUFx10_ASAP7_75t_R _26608_ (.A(_03775_),
    .Y(_03839_));
 INVx1_ASAP7_75t_R _26609_ (.A(_01236_),
    .Y(_03840_));
 NOR2x1_ASAP7_75t_R _26610_ (.A(_03840_),
    .B(_03771_),
    .Y(_03841_));
 AO21x1_ASAP7_75t_R _26611_ (.A1(_03737_),
    .A2(net600),
    .B(_03841_),
    .Y(_03842_));
 AOI21x1_ASAP7_75t_R _26612_ (.A1(_03839_),
    .A2(_03842_),
    .B(_03713_),
    .Y(_03843_));
 AND2x4_ASAP7_75t_R _26613_ (.A(_01231_),
    .B(_03744_),
    .Y(_03844_));
 NOR2x2_ASAP7_75t_R _26614_ (.A(_03844_),
    .B(_03758_),
    .Y(_03845_));
 OAI21x1_ASAP7_75t_R _26615_ (.A1(_03830_),
    .A2(_03845_),
    .B(_03805_),
    .Y(_03846_));
 NOR2x2_ASAP7_75t_R _26616_ (.A(_03665_),
    .B(_03758_),
    .Y(_03847_));
 OAI21x1_ASAP7_75t_R _26617_ (.A1(_03771_),
    .A2(_03698_),
    .B(_03699_),
    .Y(_03848_));
 AOI21x1_ASAP7_75t_R _26618_ (.A1(_15981_),
    .A2(_03847_),
    .B(_03848_),
    .Y(_03849_));
 NAND2x1_ASAP7_75t_R _26619_ (.A(_03846_),
    .B(_03849_),
    .Y(_03850_));
 AOI21x1_ASAP7_75t_R _26620_ (.A1(_03843_),
    .A2(_03850_),
    .B(_03823_),
    .Y(_03851_));
 AOI21x1_ASAP7_75t_R _26621_ (.A1(_03838_),
    .A2(_03851_),
    .B(_03789_),
    .Y(_03852_));
 NAND2x1_ASAP7_75t_R _26622_ (.A(_03824_),
    .B(_03852_),
    .Y(_03853_));
 NAND2x1_ASAP7_75t_R _26623_ (.A(_03792_),
    .B(_03853_),
    .Y(_00112_));
 NOR2x1_ASAP7_75t_R _26624_ (.A(net512),
    .B(_03655_),
    .Y(_03854_));
 OAI21x1_ASAP7_75t_R _26625_ (.A1(net833),
    .A2(_15989_),
    .B(_03771_),
    .Y(_03855_));
 BUFx6f_ASAP7_75t_R _26626_ (.A(_03825_),
    .Y(_03856_));
 OAI21x1_ASAP7_75t_R _26627_ (.A1(_03854_),
    .A2(_03855_),
    .B(_03856_),
    .Y(_03857_));
 AO21x2_ASAP7_75t_R _26628_ (.A1(_03758_),
    .A2(_03744_),
    .B(_03771_),
    .Y(_03858_));
 NOR2x1_ASAP7_75t_R _26629_ (.A(_03666_),
    .B(_03858_),
    .Y(_03859_));
 BUFx10_ASAP7_75t_R _26630_ (.A(_03713_),
    .Y(_03860_));
 OAI21x1_ASAP7_75t_R _26631_ (.A1(_03857_),
    .A2(_03859_),
    .B(_03860_),
    .Y(_03861_));
 BUFx10_ASAP7_75t_R _26632_ (.A(_03799_),
    .Y(_03862_));
 INVx3_ASAP7_75t_R _26633_ (.A(_03808_),
    .Y(_03863_));
 NAND2x2_ASAP7_75t_R _26634_ (.A(_03693_),
    .B(_03863_),
    .Y(_03864_));
 OAI21x1_ASAP7_75t_R _26635_ (.A1(_03862_),
    .A2(_03773_),
    .B(_03864_),
    .Y(_03865_));
 OAI21x1_ASAP7_75t_R _26636_ (.A1(_03673_),
    .A2(_03698_),
    .B(_03687_),
    .Y(_03866_));
 NAND2x2_ASAP7_75t_R _26637_ (.A(_15981_),
    .B(_15989_),
    .Y(_03867_));
 NOR2x2_ASAP7_75t_R _26638_ (.A(_03862_),
    .B(_03867_),
    .Y(_03868_));
 NOR3x1_ASAP7_75t_R _26639_ (.A(_03865_),
    .B(_03866_),
    .C(_03868_),
    .Y(_03869_));
 AOI21x1_ASAP7_75t_R _26640_ (.A1(_03727_),
    .A2(_03726_),
    .B(_01231_),
    .Y(_03870_));
 NOR2x2_ASAP7_75t_R _26641_ (.A(_01234_),
    .B(net923),
    .Y(_03871_));
 OAI21x1_ASAP7_75t_R _26642_ (.A1(_03870_),
    .A2(_03871_),
    .B(_03828_),
    .Y(_03872_));
 INVx4_ASAP7_75t_R _26643_ (.A(_03690_),
    .Y(_03873_));
 AOI21x1_ASAP7_75t_R _26644_ (.A1(_03768_),
    .A2(_15989_),
    .B(_03673_),
    .Y(_03874_));
 AOI21x1_ASAP7_75t_R _26645_ (.A1(_03873_),
    .A2(_03874_),
    .B(_03762_),
    .Y(_03875_));
 NAND2x1_ASAP7_75t_R _26646_ (.A(_03872_),
    .B(_03875_),
    .Y(_03876_));
 NAND2x1_ASAP7_75t_R _26647_ (.A(net915),
    .B(_03750_),
    .Y(_03877_));
 OA21x2_ASAP7_75t_R _26648_ (.A1(_03677_),
    .A2(_03737_),
    .B(_03825_),
    .Y(_03878_));
 AOI21x1_ASAP7_75t_R _26649_ (.A1(_03877_),
    .A2(_03878_),
    .B(_03741_),
    .Y(_03879_));
 NAND2x1_ASAP7_75t_R _26650_ (.A(_03876_),
    .B(_03879_),
    .Y(_03880_));
 OAI21x1_ASAP7_75t_R _26651_ (.A1(_03861_),
    .A2(_03869_),
    .B(_03880_),
    .Y(_03881_));
 NAND2x2_ASAP7_75t_R _26652_ (.A(net588),
    .B(net923),
    .Y(_03882_));
 AO21x1_ASAP7_75t_R _26653_ (.A1(_03734_),
    .A2(_03882_),
    .B(_03712_),
    .Y(_03883_));
 OAI21x1_ASAP7_75t_R _26654_ (.A1(_03666_),
    .A2(_03858_),
    .B(_03688_),
    .Y(_03884_));
 NOR2x1_ASAP7_75t_R _26655_ (.A(_03883_),
    .B(_03884_),
    .Y(_03885_));
 AOI21x1_ASAP7_75t_R _26656_ (.A1(_03760_),
    .A2(_03755_),
    .B(_03673_),
    .Y(_03886_));
 NOR2x1_ASAP7_75t_R _26657_ (.A(_03627_),
    .B(net924),
    .Y(_03887_));
 OAI21x1_ASAP7_75t_R _26658_ (.A1(net513),
    .A2(_15986_),
    .B(_03805_),
    .Y(_03888_));
 NOR2x1_ASAP7_75t_R _26659_ (.A(_03825_),
    .B(_03752_),
    .Y(_03889_));
 OAI21x1_ASAP7_75t_R _26660_ (.A1(_03887_),
    .A2(_03888_),
    .B(_03889_),
    .Y(_03890_));
 AOI21x1_ASAP7_75t_R _26661_ (.A1(net916),
    .A2(_03886_),
    .B(_03890_),
    .Y(_03891_));
 NAND3x2_ASAP7_75t_R _26662_ (.B(_03811_),
    .C(_03771_),
    .Y(_03892_),
    .A(net916));
 INVx1_ASAP7_75t_R _26663_ (.A(_03892_),
    .Y(_03893_));
 INVx1_ASAP7_75t_R _26664_ (.A(_00601_),
    .Y(_03894_));
 BUFx6f_ASAP7_75t_R _26665_ (.A(_03693_),
    .Y(_03895_));
 NAND2x1_ASAP7_75t_R _26666_ (.A(_03895_),
    .B(_03752_),
    .Y(_03896_));
 OAI21x1_ASAP7_75t_R _26667_ (.A1(_03894_),
    .A2(_03896_),
    .B(_03739_),
    .Y(_03897_));
 BUFx10_ASAP7_75t_R _26668_ (.A(_03720_),
    .Y(_03898_));
 OAI21x1_ASAP7_75t_R _26669_ (.A1(_03893_),
    .A2(_03897_),
    .B(_03898_),
    .Y(_03899_));
 NOR3x1_ASAP7_75t_R _26670_ (.A(_03885_),
    .B(_03891_),
    .C(_03899_),
    .Y(_03900_));
 AOI21x1_ASAP7_75t_R _26671_ (.A1(_03823_),
    .A2(_03881_),
    .B(_03900_),
    .Y(_03901_));
 NOR2x2_ASAP7_75t_R _26672_ (.A(_03768_),
    .B(_03670_),
    .Y(_03902_));
 NAND2x1_ASAP7_75t_R _26673_ (.A(_15986_),
    .B(_03902_),
    .Y(_03903_));
 AOI21x1_ASAP7_75t_R _26674_ (.A1(_03781_),
    .A2(_03756_),
    .B(_03762_),
    .Y(_03904_));
 NAND2x1_ASAP7_75t_R _26675_ (.A(_03903_),
    .B(_03904_),
    .Y(_03905_));
 NAND2x1_ASAP7_75t_R _26676_ (.A(_03873_),
    .B(_03874_),
    .Y(_03906_));
 NAND2x1_ASAP7_75t_R _26677_ (.A(_03802_),
    .B(_03665_),
    .Y(_03907_));
 OA21x2_ASAP7_75t_R _26678_ (.A1(_03907_),
    .A2(_15989_),
    .B(_03825_),
    .Y(_03908_));
 AOI21x1_ASAP7_75t_R _26679_ (.A1(_03906_),
    .A2(_03908_),
    .B(_03753_),
    .Y(_03909_));
 AOI21x1_ASAP7_75t_R _26680_ (.A1(_03905_),
    .A2(_03909_),
    .B(_03765_),
    .Y(_03910_));
 BUFx10_ASAP7_75t_R _26681_ (.A(_03762_),
    .Y(_03911_));
 OAI21x1_ASAP7_75t_R _26682_ (.A1(net833),
    .A2(_15986_),
    .B(_03771_),
    .Y(_03912_));
 INVx2_ASAP7_75t_R _26683_ (.A(_03698_),
    .Y(_03913_));
 OA22x2_ASAP7_75t_R _26684_ (.A1(_03796_),
    .A2(_03804_),
    .B1(_03912_),
    .B2(_03913_),
    .Y(_03914_));
 NAND2x1_ASAP7_75t_R _26685_ (.A(_15981_),
    .B(net46),
    .Y(_03915_));
 AOI21x1_ASAP7_75t_R _26686_ (.A1(_03915_),
    .A2(_03767_),
    .B(_03813_),
    .Y(_03916_));
 AO21x1_ASAP7_75t_R _26687_ (.A1(_03736_),
    .A2(_03671_),
    .B(_03694_),
    .Y(_03917_));
 AOI21x1_ASAP7_75t_R _26688_ (.A1(_03916_),
    .A2(_03917_),
    .B(_03741_),
    .Y(_03918_));
 OAI21x1_ASAP7_75t_R _26689_ (.A1(_03911_),
    .A2(_03914_),
    .B(_03918_),
    .Y(_03919_));
 NAND2x1_ASAP7_75t_R _26690_ (.A(_03910_),
    .B(_03919_),
    .Y(_03920_));
 OA21x2_ASAP7_75t_R _26691_ (.A1(_03803_),
    .A2(_03799_),
    .B(_03775_),
    .Y(_03921_));
 NOR2x2_ASAP7_75t_R _26692_ (.A(net587),
    .B(net924),
    .Y(_03922_));
 NAND2x1_ASAP7_75t_R _26693_ (.A(_03816_),
    .B(_03922_),
    .Y(_03923_));
 NAND2x1_ASAP7_75t_R _26694_ (.A(_00602_),
    .B(_03895_),
    .Y(_03924_));
 NAND3x1_ASAP7_75t_R _26695_ (.A(_03921_),
    .B(_03923_),
    .C(_03924_),
    .Y(_03925_));
 OAI21x1_ASAP7_75t_R _26696_ (.A1(_03871_),
    .A2(_03863_),
    .B(_03694_),
    .Y(_03926_));
 NAND2x1_ASAP7_75t_R _26697_ (.A(_03803_),
    .B(_03829_),
    .Y(_03927_));
 AOI21x1_ASAP7_75t_R _26698_ (.A1(_03816_),
    .A2(_03927_),
    .B(_03749_),
    .Y(_03928_));
 AOI21x1_ASAP7_75t_R _26699_ (.A1(_03926_),
    .A2(_03928_),
    .B(_03741_),
    .Y(_03929_));
 NAND2x1_ASAP7_75t_R _26700_ (.A(_03925_),
    .B(_03929_),
    .Y(_03930_));
 NAND2x1_ASAP7_75t_R _26701_ (.A(net901),
    .B(_03767_),
    .Y(_03931_));
 AOI21x1_ASAP7_75t_R _26702_ (.A1(_03744_),
    .A2(_03758_),
    .B(_03693_),
    .Y(_03932_));
 AOI21x1_ASAP7_75t_R _26703_ (.A1(_03867_),
    .A2(_03932_),
    .B(_03739_),
    .Y(_03933_));
 NAND2x1_ASAP7_75t_R _26704_ (.A(_03931_),
    .B(_03933_),
    .Y(_03934_));
 AOI21x1_ASAP7_75t_R _26705_ (.A1(_03862_),
    .A2(_03746_),
    .B(_03688_),
    .Y(_03935_));
 NAND2x1_ASAP7_75t_R _26706_ (.A(_03733_),
    .B(_03809_),
    .Y(_03936_));
 AOI21x1_ASAP7_75t_R _26707_ (.A1(_03935_),
    .A2(_03936_),
    .B(_03753_),
    .Y(_03937_));
 AOI21x1_ASAP7_75t_R _26708_ (.A1(_03934_),
    .A2(_03937_),
    .B(_03823_),
    .Y(_03938_));
 AOI21x1_ASAP7_75t_R _26709_ (.A1(_03930_),
    .A2(_03938_),
    .B(_03789_),
    .Y(_03939_));
 NAND2x1_ASAP7_75t_R _26710_ (.A(_03920_),
    .B(_03939_),
    .Y(_03940_));
 OAI21x1_ASAP7_75t_R _26711_ (.A1(_03790_),
    .A2(_03901_),
    .B(_03940_),
    .Y(_00113_));
 AOI21x1_ASAP7_75t_R _26712_ (.A1(_03803_),
    .A2(_03736_),
    .B(_03828_),
    .Y(_03941_));
 AOI21x1_ASAP7_75t_R _26713_ (.A1(_03674_),
    .A2(_03675_),
    .B(net884),
    .Y(_03942_));
 AOI21x1_ASAP7_75t_R _26714_ (.A1(_03727_),
    .A2(_03726_),
    .B(_01234_),
    .Y(_03943_));
 OA21x2_ASAP7_75t_R _26715_ (.A1(_03942_),
    .A2(net902),
    .B(_03828_),
    .Y(_03944_));
 BUFx6f_ASAP7_75t_R _26716_ (.A(_03749_),
    .Y(_03945_));
 OAI21x1_ASAP7_75t_R _26717_ (.A1(_03941_),
    .A2(_03944_),
    .B(_03945_),
    .Y(_03946_));
 AOI21x1_ASAP7_75t_R _26718_ (.A1(_03744_),
    .A2(_03755_),
    .B(_03673_),
    .Y(_03947_));
 NAND2x1_ASAP7_75t_R _26719_ (.A(_03781_),
    .B(_03947_),
    .Y(_03948_));
 AO21x1_ASAP7_75t_R _26720_ (.A1(_03798_),
    .A2(_03803_),
    .B(_03670_),
    .Y(_03949_));
 AO21x1_ASAP7_75t_R _26721_ (.A1(_03948_),
    .A2(_03949_),
    .B(_03945_),
    .Y(_03950_));
 AOI21x1_ASAP7_75t_R _26722_ (.A1(_03946_),
    .A2(_03950_),
    .B(_03860_),
    .Y(_03951_));
 NOR2x1_ASAP7_75t_R _26723_ (.A(_03863_),
    .B(_03796_),
    .Y(_03952_));
 OAI21x1_ASAP7_75t_R _26724_ (.A1(_03797_),
    .A2(_03655_),
    .B(_03665_),
    .Y(_03953_));
 NOR2x1_ASAP7_75t_R _26725_ (.A(_03887_),
    .B(_03953_),
    .Y(_03954_));
 OAI21x1_ASAP7_75t_R _26726_ (.A1(_03952_),
    .A2(_03954_),
    .B(_03911_),
    .Y(_03955_));
 AO21x1_ASAP7_75t_R _26727_ (.A1(_15989_),
    .A2(net46),
    .B(_03737_),
    .Y(_03956_));
 INVx1_ASAP7_75t_R _26728_ (.A(_03943_),
    .Y(_03957_));
 AOI21x1_ASAP7_75t_R _26729_ (.A1(_03957_),
    .A2(_03734_),
    .B(_03739_),
    .Y(_03958_));
 OAI21x1_ASAP7_75t_R _26730_ (.A1(_03942_),
    .A2(_03956_),
    .B(_03958_),
    .Y(_03959_));
 AOI21x1_ASAP7_75t_R _26731_ (.A1(_03955_),
    .A2(_03959_),
    .B(_03821_),
    .Y(_03960_));
 NOR3x1_ASAP7_75t_R _26732_ (.A(_03951_),
    .B(_03960_),
    .C(_03765_),
    .Y(_03961_));
 AOI21x1_ASAP7_75t_R _26733_ (.A1(net46),
    .A2(_15989_),
    .B(_03799_),
    .Y(_03962_));
 AOI21x1_ASAP7_75t_R _26734_ (.A1(_15981_),
    .A2(_15986_),
    .B(_03805_),
    .Y(_03963_));
 INVx2_ASAP7_75t_R _26735_ (.A(_03870_),
    .Y(_03964_));
 AOI22x1_ASAP7_75t_R _26736_ (.A1(_03962_),
    .A2(_03873_),
    .B1(_03963_),
    .B2(_03964_),
    .Y(_03965_));
 NAND2x1_ASAP7_75t_R _26737_ (.A(_03779_),
    .B(_03874_),
    .Y(_03966_));
 NOR2x1_ASAP7_75t_R _26738_ (.A(_03813_),
    .B(_03761_),
    .Y(_03967_));
 AOI21x1_ASAP7_75t_R _26739_ (.A1(_03966_),
    .A2(_03967_),
    .B(_03753_),
    .Y(_03968_));
 OAI21x1_ASAP7_75t_R _26740_ (.A1(_03911_),
    .A2(_03965_),
    .B(_03968_),
    .Y(_03969_));
 NAND2x2_ASAP7_75t_R _26741_ (.A(net590),
    .B(_03758_),
    .Y(_03970_));
 NAND2x2_ASAP7_75t_R _26742_ (.A(_03970_),
    .B(_03886_),
    .Y(_03971_));
 AO21x2_ASAP7_75t_R _26743_ (.A1(_03726_),
    .A2(_03727_),
    .B(_03778_),
    .Y(_03972_));
 NAND2x2_ASAP7_75t_R _26744_ (.A(_03972_),
    .B(_03932_),
    .Y(_03973_));
 AOI21x1_ASAP7_75t_R _26745_ (.A1(_03971_),
    .A2(_03973_),
    .B(_03856_),
    .Y(_03974_));
 INVx2_ASAP7_75t_R _26746_ (.A(_03810_),
    .Y(_03975_));
 OAI21x1_ASAP7_75t_R _26747_ (.A1(_03828_),
    .A2(_03927_),
    .B(_03739_),
    .Y(_03976_));
 NOR2x1_ASAP7_75t_R _26748_ (.A(_03975_),
    .B(_03976_),
    .Y(_03977_));
 OAI21x1_ASAP7_75t_R _26749_ (.A1(_03974_),
    .A2(_03977_),
    .B(_03821_),
    .Y(_03978_));
 NAND2x1_ASAP7_75t_R _26750_ (.A(_03969_),
    .B(_03978_),
    .Y(_03979_));
 OAI21x1_ASAP7_75t_R _26751_ (.A1(_03823_),
    .A2(_03979_),
    .B(_03789_),
    .Y(_03980_));
 NAND2x1_ASAP7_75t_R _26752_ (.A(_00601_),
    .B(_03805_),
    .Y(_03981_));
 AOI21x1_ASAP7_75t_R _26753_ (.A1(net588),
    .A2(_03758_),
    .B(_03673_),
    .Y(_03982_));
 AOI21x1_ASAP7_75t_R _26754_ (.A1(_03733_),
    .A2(_03982_),
    .B(_03775_),
    .Y(_03983_));
 AOI21x1_ASAP7_75t_R _26755_ (.A1(_03981_),
    .A2(_03983_),
    .B(_03741_),
    .Y(_03984_));
 NAND2x1_ASAP7_75t_R _26756_ (.A(_03808_),
    .B(_03799_),
    .Y(_03985_));
 NOR2x1_ASAP7_75t_R _26757_ (.A(_03724_),
    .B(_03985_),
    .Y(_03986_));
 INVx1_ASAP7_75t_R _26758_ (.A(_03809_),
    .Y(_03987_));
 NOR2x1_ASAP7_75t_R _26759_ (.A(_03692_),
    .B(_03987_),
    .Y(_03988_));
 OAI21x1_ASAP7_75t_R _26760_ (.A1(_03988_),
    .A2(_03986_),
    .B(_03945_),
    .Y(_03989_));
 NAND2x1_ASAP7_75t_R _26761_ (.A(_03984_),
    .B(_03989_),
    .Y(_03990_));
 NAND2x1_ASAP7_75t_R _26762_ (.A(_03840_),
    .B(_03828_),
    .Y(_03991_));
 AO21x1_ASAP7_75t_R _26763_ (.A1(net600),
    .A2(_03829_),
    .B(_03816_),
    .Y(_03992_));
 AOI21x1_ASAP7_75t_R _26764_ (.A1(_03991_),
    .A2(_03992_),
    .B(_03945_),
    .Y(_03993_));
 NAND2x2_ASAP7_75t_R _26765_ (.A(_15976_),
    .B(_03755_),
    .Y(_03994_));
 NAND2x2_ASAP7_75t_R _26766_ (.A(_03994_),
    .B(_03812_),
    .Y(_03995_));
 AOI21x1_ASAP7_75t_R _26767_ (.A1(_03995_),
    .A2(_03810_),
    .B(_03856_),
    .Y(_03996_));
 OAI21x1_ASAP7_75t_R _26768_ (.A1(_03993_),
    .A2(_03996_),
    .B(_03860_),
    .Y(_03997_));
 NAND2x1_ASAP7_75t_R _26769_ (.A(_03997_),
    .B(_03990_),
    .Y(_03998_));
 AOI21x1_ASAP7_75t_R _26770_ (.A1(_03844_),
    .A2(_03758_),
    .B(_03673_),
    .Y(_03999_));
 NAND2x1_ASAP7_75t_R _26771_ (.A(_03728_),
    .B(_03999_),
    .Y(_04000_));
 NAND2x1_ASAP7_75t_R _26772_ (.A(_03892_),
    .B(_04000_),
    .Y(_04001_));
 INVx1_ASAP7_75t_R _26773_ (.A(_03700_),
    .Y(_04002_));
 OAI21x1_ASAP7_75t_R _26774_ (.A1(_03804_),
    .A2(_03690_),
    .B(_03862_),
    .Y(_04003_));
 AOI21x1_ASAP7_75t_R _26775_ (.A1(_04002_),
    .A2(_04003_),
    .B(_03753_),
    .Y(_04004_));
 OAI21x1_ASAP7_75t_R _26776_ (.A1(_03911_),
    .A2(_04001_),
    .B(_04004_),
    .Y(_04005_));
 AND2x2_ASAP7_75t_R _26777_ (.A(_03670_),
    .B(_00603_),
    .Y(_04006_));
 NOR2x1_ASAP7_75t_R _26778_ (.A(_04006_),
    .B(_03761_),
    .Y(_04007_));
 NAND2x1_ASAP7_75t_R _26779_ (.A(_03856_),
    .B(_04007_),
    .Y(_04008_));
 OA21x2_ASAP7_75t_R _26780_ (.A1(_01238_),
    .A2(_03694_),
    .B(_03813_),
    .Y(_04009_));
 AOI21x1_ASAP7_75t_R _26781_ (.A1(_04009_),
    .A2(_03971_),
    .B(_03741_),
    .Y(_04010_));
 AOI21x1_ASAP7_75t_R _26782_ (.A1(_04008_),
    .A2(_04010_),
    .B(_03823_),
    .Y(_04011_));
 AOI21x1_ASAP7_75t_R _26783_ (.A1(_04005_),
    .A2(_04011_),
    .B(_03789_),
    .Y(_04012_));
 OAI21x1_ASAP7_75t_R _26784_ (.A1(_03765_),
    .A2(_03998_),
    .B(_04012_),
    .Y(_04013_));
 OAI21x1_ASAP7_75t_R _26785_ (.A1(_03961_),
    .A2(_03980_),
    .B(_04013_),
    .Y(_00114_));
 OAI21x1_ASAP7_75t_R _26786_ (.A1(net46),
    .A2(_15989_),
    .B(_03752_),
    .Y(_04014_));
 NAND2x2_ASAP7_75t_R _26787_ (.A(_03737_),
    .B(_03811_),
    .Y(_04015_));
 OAI22x1_ASAP7_75t_R _26788_ (.A1(_04014_),
    .A2(_04015_),
    .B1(_03678_),
    .B2(_03752_),
    .Y(_04016_));
 NOR2x1_ASAP7_75t_R _26789_ (.A(_03825_),
    .B(_03831_),
    .Y(_04017_));
 OAI21x1_ASAP7_75t_R _26790_ (.A1(_03671_),
    .A2(_03896_),
    .B(_04017_),
    .Y(_04018_));
 OAI21x1_ASAP7_75t_R _26791_ (.A1(_04016_),
    .A2(_04018_),
    .B(_03898_),
    .Y(_04019_));
 NAND2x1_ASAP7_75t_R _26792_ (.A(net901),
    .B(_03750_),
    .Y(_04020_));
 AOI21x1_ASAP7_75t_R _26793_ (.A1(_03972_),
    .A2(_03999_),
    .B(_03712_),
    .Y(_04021_));
 NAND2x1_ASAP7_75t_R _26794_ (.A(_04020_),
    .B(_04021_),
    .Y(_04022_));
 AO21x1_ASAP7_75t_R _26795_ (.A1(_03942_),
    .A2(_03670_),
    .B(_03711_),
    .Y(_04023_));
 OR2x2_ASAP7_75t_R _26796_ (.A(_04023_),
    .B(_03954_),
    .Y(_04024_));
 AOI21x1_ASAP7_75t_R _26797_ (.A1(_04022_),
    .A2(_04024_),
    .B(_03945_),
    .Y(_04025_));
 NOR2x1_ASAP7_75t_R _26798_ (.A(_04019_),
    .B(_04025_),
    .Y(_04026_));
 OAI21x1_ASAP7_75t_R _26799_ (.A1(net902),
    .A2(_03855_),
    .B(_03813_),
    .Y(_04027_));
 NAND2x1_ASAP7_75t_R _26800_ (.A(_03752_),
    .B(_04027_),
    .Y(_04028_));
 NOR2x1_ASAP7_75t_R _26801_ (.A(net884),
    .B(_15986_),
    .Y(_04029_));
 NOR2x2_ASAP7_75t_R _26802_ (.A(_03844_),
    .B(_03755_),
    .Y(_04030_));
 OAI21x1_ASAP7_75t_R _26803_ (.A1(_04029_),
    .A2(_04030_),
    .B(_03747_),
    .Y(_04031_));
 AOI21x1_ASAP7_75t_R _26804_ (.A1(_03892_),
    .A2(_04031_),
    .B(_03839_),
    .Y(_04032_));
 OAI21x1_ASAP7_75t_R _26805_ (.A1(_04028_),
    .A2(_04032_),
    .B(_03721_),
    .Y(_04033_));
 NAND2x1_ASAP7_75t_R _26806_ (.A(_03972_),
    .B(_03729_),
    .Y(_04034_));
 OAI21x1_ASAP7_75t_R _26807_ (.A1(_15981_),
    .A2(_15986_),
    .B(_03798_),
    .Y(_04035_));
 AOI21x1_ASAP7_75t_R _26808_ (.A1(_03747_),
    .A2(_04035_),
    .B(_03762_),
    .Y(_04036_));
 NAND2x1_ASAP7_75t_R _26809_ (.A(_04036_),
    .B(_04034_),
    .Y(_04037_));
 NAND2x1_ASAP7_75t_R _26810_ (.A(_03936_),
    .B(_03849_),
    .Y(_04038_));
 AOI21x1_ASAP7_75t_R _26811_ (.A1(_04037_),
    .A2(_04038_),
    .B(_03821_),
    .Y(_04039_));
 NOR2x1_ASAP7_75t_R _26812_ (.A(_04033_),
    .B(_04039_),
    .Y(_04040_));
 OAI21x1_ASAP7_75t_R _26813_ (.A1(_04026_),
    .A2(_04040_),
    .B(_03789_),
    .Y(_04041_));
 NOR2x1_ASAP7_75t_R _26814_ (.A(_15981_),
    .B(net587),
    .Y(_04042_));
 NOR2x2_ASAP7_75t_R _26815_ (.A(net833),
    .B(_03758_),
    .Y(_04043_));
 OAI21x1_ASAP7_75t_R _26816_ (.A1(_04042_),
    .A2(_04043_),
    .B(_03805_),
    .Y(_04044_));
 OAI21x1_ASAP7_75t_R _26817_ (.A1(_03677_),
    .A2(_03956_),
    .B(_04044_),
    .Y(_04045_));
 AOI21x1_ASAP7_75t_R _26818_ (.A1(_03747_),
    .A2(_03671_),
    .B(_03762_),
    .Y(_04046_));
 NAND2x1_ASAP7_75t_R _26819_ (.A(_03759_),
    .B(_03962_),
    .Y(_04047_));
 AOI21x1_ASAP7_75t_R _26820_ (.A1(_04046_),
    .A2(_04047_),
    .B(_03713_),
    .Y(_04048_));
 OAI21x1_ASAP7_75t_R _26821_ (.A1(_03945_),
    .A2(_04045_),
    .B(_04048_),
    .Y(_04049_));
 NOR2x1_ASAP7_75t_R _26822_ (.A(_03724_),
    .B(_03912_),
    .Y(_04050_));
 OAI21x1_ASAP7_75t_R _26823_ (.A1(_03913_),
    .A2(_03672_),
    .B(_03813_),
    .Y(_04051_));
 NOR2x1_ASAP7_75t_R _26824_ (.A(_04050_),
    .B(_04051_),
    .Y(_04052_));
 NAND2x1_ASAP7_75t_R _26825_ (.A(_03779_),
    .B(_03947_),
    .Y(_04053_));
 NAND2x1_ASAP7_75t_R _26826_ (.A(_03873_),
    .B(_03962_),
    .Y(_04054_));
 AOI21x1_ASAP7_75t_R _26827_ (.A1(_04053_),
    .A2(_04054_),
    .B(_03839_),
    .Y(_04055_));
 OAI21x1_ASAP7_75t_R _26828_ (.A1(_04052_),
    .A2(_04055_),
    .B(_03860_),
    .Y(_04056_));
 AOI21x1_ASAP7_75t_R _26829_ (.A1(_04049_),
    .A2(_04056_),
    .B(_03823_),
    .Y(_04057_));
 OAI21x1_ASAP7_75t_R _26830_ (.A1(_03724_),
    .A2(_03746_),
    .B(_03747_),
    .Y(_04058_));
 OA21x2_ASAP7_75t_R _26831_ (.A1(_03647_),
    .A2(_03640_),
    .B(_00599_),
    .Y(_04059_));
 OAI21x1_ASAP7_75t_R _26832_ (.A1(_03863_),
    .A2(_04059_),
    .B(_03828_),
    .Y(_04060_));
 AOI21x1_ASAP7_75t_R _26833_ (.A1(_04058_),
    .A2(_04060_),
    .B(_03839_),
    .Y(_04061_));
 AO21x1_ASAP7_75t_R _26834_ (.A1(_03795_),
    .A2(_03696_),
    .B(_03895_),
    .Y(_04062_));
 NOR2x1_ASAP7_75t_R _26835_ (.A(_15981_),
    .B(net46),
    .Y(_04063_));
 OAI21x1_ASAP7_75t_R _26836_ (.A1(_04063_),
    .A2(_04043_),
    .B(_03862_),
    .Y(_04064_));
 AOI21x1_ASAP7_75t_R _26837_ (.A1(_04062_),
    .A2(_04064_),
    .B(_03856_),
    .Y(_04065_));
 OAI21x1_ASAP7_75t_R _26838_ (.A1(_04061_),
    .A2(_04065_),
    .B(_03860_),
    .Y(_04066_));
 INVx1_ASAP7_75t_R _26839_ (.A(_03886_),
    .Y(_04067_));
 AOI21x1_ASAP7_75t_R _26840_ (.A1(_04067_),
    .A2(_04044_),
    .B(_03839_),
    .Y(_04068_));
 NAND2x1_ASAP7_75t_R _26841_ (.A(_03781_),
    .B(_03756_),
    .Y(_04069_));
 AOI21x1_ASAP7_75t_R _26842_ (.A1(net884),
    .A2(_03755_),
    .B(_03693_),
    .Y(_04070_));
 NAND2x1_ASAP7_75t_R _26843_ (.A(_03873_),
    .B(_04070_),
    .Y(_04071_));
 AOI21x1_ASAP7_75t_R _26844_ (.A1(_04069_),
    .A2(_04071_),
    .B(_03856_),
    .Y(_04072_));
 OAI21x1_ASAP7_75t_R _26845_ (.A1(_04068_),
    .A2(_04072_),
    .B(_03821_),
    .Y(_04073_));
 AOI21x1_ASAP7_75t_R _26846_ (.A1(_04066_),
    .A2(_04073_),
    .B(_03765_),
    .Y(_04074_));
 OAI21x1_ASAP7_75t_R _26847_ (.A1(_04057_),
    .A2(_04074_),
    .B(_03790_),
    .Y(_04075_));
 NAND2x1_ASAP7_75t_R _26848_ (.A(_04041_),
    .B(_04075_),
    .Y(_00115_));
 NAND2x1_ASAP7_75t_R _26849_ (.A(_03627_),
    .B(net587),
    .Y(_04076_));
 AOI21x1_ASAP7_75t_R _26850_ (.A1(_04076_),
    .A2(_03781_),
    .B(_03895_),
    .Y(_04077_));
 AOI211x1_ASAP7_75t_R _26851_ (.A1(_03835_),
    .A2(_03736_),
    .B(_04077_),
    .C(_03856_),
    .Y(_04078_));
 NAND2x1_ASAP7_75t_R _26852_ (.A(_03817_),
    .B(_03738_),
    .Y(_04079_));
 OAI21x1_ASAP7_75t_R _26853_ (.A1(_03945_),
    .A2(_04079_),
    .B(_03821_),
    .Y(_04080_));
 NOR2x1_ASAP7_75t_R _26854_ (.A(_03749_),
    .B(_03902_),
    .Y(_04081_));
 AOI21x1_ASAP7_75t_R _26855_ (.A1(_03985_),
    .A2(_04081_),
    .B(_03752_),
    .Y(_04082_));
 OA21x2_ASAP7_75t_R _26856_ (.A1(_03829_),
    .A2(_03799_),
    .B(_03775_),
    .Y(_04083_));
 NAND2x1_ASAP7_75t_R _26857_ (.A(_03781_),
    .B(_03835_),
    .Y(_04084_));
 NAND2x1_ASAP7_75t_R _26858_ (.A(_04083_),
    .B(_04084_),
    .Y(_04085_));
 AOI21x1_ASAP7_75t_R _26859_ (.A1(_04082_),
    .A2(_04085_),
    .B(_03721_),
    .Y(_04086_));
 OAI21x1_ASAP7_75t_R _26860_ (.A1(_04078_),
    .A2(_04080_),
    .B(_04086_),
    .Y(_04087_));
 INVx1_ASAP7_75t_R _26861_ (.A(_03874_),
    .Y(_04088_));
 AO21x1_ASAP7_75t_R _26862_ (.A1(_03726_),
    .A2(_03727_),
    .B(_03772_),
    .Y(_04089_));
 AOI21x1_ASAP7_75t_R _26863_ (.A1(_03805_),
    .A2(_04089_),
    .B(_03762_),
    .Y(_04090_));
 AOI21x1_ASAP7_75t_R _26864_ (.A1(_04088_),
    .A2(_04090_),
    .B(_03753_),
    .Y(_04091_));
 NAND2x1_ASAP7_75t_R _26865_ (.A(_03808_),
    .B(_03932_),
    .Y(_04092_));
 NAND2x1_ASAP7_75t_R _26866_ (.A(_04092_),
    .B(_03793_),
    .Y(_04093_));
 AOI21x1_ASAP7_75t_R _26867_ (.A1(_04091_),
    .A2(_04093_),
    .B(_03765_),
    .Y(_04094_));
 AO21x1_ASAP7_75t_R _26868_ (.A1(_03994_),
    .A2(_03698_),
    .B(_03895_),
    .Y(_04095_));
 OAI21x1_ASAP7_75t_R _26869_ (.A1(_03666_),
    .A2(_03858_),
    .B(_04095_),
    .Y(_04096_));
 NOR2x1_ASAP7_75t_R _26870_ (.A(_03813_),
    .B(_03847_),
    .Y(_04097_));
 NAND2x1_ASAP7_75t_R _26871_ (.A(_03972_),
    .B(_03734_),
    .Y(_04098_));
 AOI21x1_ASAP7_75t_R _26872_ (.A1(_04097_),
    .A2(_04098_),
    .B(_03713_),
    .Y(_04099_));
 OAI21x1_ASAP7_75t_R _26873_ (.A1(_03911_),
    .A2(_04096_),
    .B(_04099_),
    .Y(_04100_));
 AOI21x1_ASAP7_75t_R _26874_ (.A1(_04094_),
    .A2(_04100_),
    .B(_03790_),
    .Y(_04101_));
 NAND2x1_ASAP7_75t_R _26875_ (.A(_04087_),
    .B(_04101_),
    .Y(_04102_));
 NAND2x1_ASAP7_75t_R _26876_ (.A(_03775_),
    .B(_03773_),
    .Y(_04103_));
 OA21x2_ASAP7_75t_R _26877_ (.A1(_03835_),
    .A2(_04103_),
    .B(_03713_),
    .Y(_04104_));
 INVx1_ASAP7_75t_R _26878_ (.A(_03882_),
    .Y(_04105_));
 INVx1_ASAP7_75t_R _26879_ (.A(_03812_),
    .Y(_04106_));
 AOI21x1_ASAP7_75t_R _26880_ (.A1(_03691_),
    .A2(_15989_),
    .B(_03799_),
    .Y(_04107_));
 AOI21x1_ASAP7_75t_R _26881_ (.A1(_03759_),
    .A2(_04107_),
    .B(_03813_),
    .Y(_04108_));
 OAI21x1_ASAP7_75t_R _26882_ (.A1(_04105_),
    .A2(_04106_),
    .B(_04108_),
    .Y(_04109_));
 AOI21x1_ASAP7_75t_R _26883_ (.A1(_04104_),
    .A2(_04109_),
    .B(_03898_),
    .Y(_04110_));
 NAND2x1_ASAP7_75t_R _26884_ (.A(_03882_),
    .B(_03734_),
    .Y(_04111_));
 AOI21x1_ASAP7_75t_R _26885_ (.A1(_04111_),
    .A2(_03983_),
    .B(_03713_),
    .Y(_04112_));
 OA21x2_ASAP7_75t_R _26886_ (.A1(_03854_),
    .A2(_03922_),
    .B(_03895_),
    .Y(_04113_));
 OAI21x1_ASAP7_75t_R _26887_ (.A1(_04077_),
    .A2(_04113_),
    .B(_03839_),
    .Y(_04114_));
 NAND2x1_ASAP7_75t_R _26888_ (.A(_04112_),
    .B(_04114_),
    .Y(_04115_));
 AOI21x1_ASAP7_75t_R _26889_ (.A1(_04110_),
    .A2(_04115_),
    .B(_03789_),
    .Y(_04116_));
 AND2x2_ASAP7_75t_R _26890_ (.A(_03864_),
    .B(_03949_),
    .Y(_04117_));
 OA21x2_ASAP7_75t_R _26891_ (.A1(_03798_),
    .A2(_03816_),
    .B(_03813_),
    .Y(_04118_));
 AO21x1_ASAP7_75t_R _26892_ (.A1(_04117_),
    .A2(_04118_),
    .B(_03753_),
    .Y(_04119_));
 INVx1_ASAP7_75t_R _26893_ (.A(_03871_),
    .Y(_04120_));
 AO21x1_ASAP7_75t_R _26894_ (.A1(_04120_),
    .A2(net600),
    .B(_03694_),
    .Y(_04121_));
 AND3x1_ASAP7_75t_R _26895_ (.A(_04121_),
    .B(_03856_),
    .C(_03836_),
    .Y(_04122_));
 AO21x1_ASAP7_75t_R _26896_ (.A1(_03882_),
    .A2(_03698_),
    .B(_03737_),
    .Y(_04123_));
 AOI21x1_ASAP7_75t_R _26897_ (.A1(_03928_),
    .A2(_04123_),
    .B(_03713_),
    .Y(_04124_));
 AOI21x1_ASAP7_75t_R _26898_ (.A1(_03760_),
    .A2(_03758_),
    .B(_03665_),
    .Y(_04125_));
 NAND2x1_ASAP7_75t_R _26899_ (.A(_03994_),
    .B(_04125_),
    .Y(_04126_));
 NAND3x1_ASAP7_75t_R _26900_ (.A(_03973_),
    .B(_04126_),
    .C(_03688_),
    .Y(_04127_));
 AOI21x1_ASAP7_75t_R _26901_ (.A1(_04124_),
    .A2(_04127_),
    .B(_03823_),
    .Y(_04128_));
 OAI21x1_ASAP7_75t_R _26902_ (.A1(_04122_),
    .A2(_04119_),
    .B(_04128_),
    .Y(_04129_));
 NAND2x1_ASAP7_75t_R _26903_ (.A(_04116_),
    .B(_04129_),
    .Y(_04130_));
 NAND2x1_ASAP7_75t_R _26904_ (.A(_04102_),
    .B(_04130_),
    .Y(_00116_));
 AOI21x1_ASAP7_75t_R _26905_ (.A1(_03757_),
    .A2(_03921_),
    .B(_03721_),
    .Y(_04131_));
 INVx2_ASAP7_75t_R _26906_ (.A(net916),
    .Y(_04132_));
 INVx1_ASAP7_75t_R _26907_ (.A(_03761_),
    .Y(_04133_));
 NOR2x1_ASAP7_75t_R _26908_ (.A(_03749_),
    .B(_03999_),
    .Y(_04134_));
 OAI21x1_ASAP7_75t_R _26909_ (.A1(_04132_),
    .A2(_04133_),
    .B(_04134_),
    .Y(_04135_));
 AOI21x1_ASAP7_75t_R _26910_ (.A1(_04131_),
    .A2(_04135_),
    .B(_03753_),
    .Y(_04136_));
 NAND2x1_ASAP7_75t_R _26911_ (.A(_03694_),
    .B(_15981_),
    .Y(_04137_));
 AOI21x1_ASAP7_75t_R _26912_ (.A1(_04137_),
    .A2(_03735_),
    .B(_03688_),
    .Y(_04138_));
 NAND2x1_ASAP7_75t_R _26913_ (.A(_03781_),
    .B(_04070_),
    .Y(_04139_));
 NAND2x1_ASAP7_75t_R _26914_ (.A(_03795_),
    .B(_03886_),
    .Y(_04140_));
 AOI21x1_ASAP7_75t_R _26915_ (.A1(_04139_),
    .A2(_04140_),
    .B(_03739_),
    .Y(_04141_));
 OAI21x1_ASAP7_75t_R _26916_ (.A1(_04138_),
    .A2(_04141_),
    .B(_03721_),
    .Y(_04142_));
 NAND2x1_ASAP7_75t_R _26917_ (.A(_04136_),
    .B(_04142_),
    .Y(_04143_));
 AOI21x1_ASAP7_75t_R _26918_ (.A1(_03803_),
    .A2(_03736_),
    .B(_03862_),
    .Y(_04144_));
 OAI21x1_ASAP7_75t_R _26919_ (.A1(_03943_),
    .A2(_04059_),
    .B(_03805_),
    .Y(_04145_));
 OA21x2_ASAP7_75t_R _26920_ (.A1(_03696_),
    .A2(_03737_),
    .B(_03749_),
    .Y(_04146_));
 AOI21x1_ASAP7_75t_R _26921_ (.A1(_04145_),
    .A2(_04146_),
    .B(_03898_),
    .Y(_04147_));
 OAI21x1_ASAP7_75t_R _26922_ (.A1(_03794_),
    .A2(_04144_),
    .B(_04147_),
    .Y(_04148_));
 AO21x1_ASAP7_75t_R _26923_ (.A1(_00595_),
    .A2(_03799_),
    .B(_03775_),
    .Y(_04149_));
 NOR2x1_ASAP7_75t_R _26924_ (.A(_03799_),
    .B(_04132_),
    .Y(_04150_));
 OA21x2_ASAP7_75t_R _26925_ (.A1(_04149_),
    .A2(_04150_),
    .B(_03720_),
    .Y(_04151_));
 AO21x1_ASAP7_75t_R _26926_ (.A1(_03957_),
    .A2(_03795_),
    .B(_03895_),
    .Y(_04152_));
 INVx1_ASAP7_75t_R _26927_ (.A(_03796_),
    .Y(_04153_));
 AOI21x1_ASAP7_75t_R _26928_ (.A1(_03811_),
    .A2(_04153_),
    .B(_03762_),
    .Y(_04154_));
 NAND2x1_ASAP7_75t_R _26929_ (.A(_04152_),
    .B(_04154_),
    .Y(_04155_));
 AOI21x1_ASAP7_75t_R _26930_ (.A1(_04151_),
    .A2(_04155_),
    .B(_03741_),
    .Y(_04156_));
 NAND2x1_ASAP7_75t_R _26931_ (.A(_04148_),
    .B(_04156_),
    .Y(_04157_));
 AOI21x1_ASAP7_75t_R _26932_ (.A1(_04143_),
    .A2(_04157_),
    .B(_03790_),
    .Y(_04158_));
 AO21x1_ASAP7_75t_R _26933_ (.A1(net46),
    .A2(_03799_),
    .B(_03775_),
    .Y(_04159_));
 OAI21x1_ASAP7_75t_R _26934_ (.A1(_04159_),
    .A2(_04077_),
    .B(_03898_),
    .Y(_04160_));
 AOI21x1_ASAP7_75t_R _26935_ (.A1(net916),
    .A2(_03811_),
    .B(_03816_),
    .Y(_04161_));
 AOI211x1_ASAP7_75t_R _26936_ (.A1(_03750_),
    .A2(_04076_),
    .B(_04161_),
    .C(_03739_),
    .Y(_04162_));
 OAI21x1_ASAP7_75t_R _26937_ (.A1(_04160_),
    .A2(_04162_),
    .B(_03741_),
    .Y(_04163_));
 NAND2x1_ASAP7_75t_R _26938_ (.A(_03833_),
    .B(_04070_),
    .Y(_04164_));
 INVx1_ASAP7_75t_R _26939_ (.A(_03844_),
    .Y(_04165_));
 AOI21x1_ASAP7_75t_R _26940_ (.A1(_04165_),
    .A2(_03947_),
    .B(_03762_),
    .Y(_04166_));
 NAND2x1_ASAP7_75t_R _26941_ (.A(_04164_),
    .B(_04166_),
    .Y(_04167_));
 OAI21x1_ASAP7_75t_R _26942_ (.A1(_03943_),
    .A2(_03745_),
    .B(_03694_),
    .Y(_04168_));
 NAND3x1_ASAP7_75t_R _26943_ (.A(_03667_),
    .B(_03776_),
    .C(_04168_),
    .Y(_04169_));
 AOI21x1_ASAP7_75t_R _26944_ (.A1(_04167_),
    .A2(_04169_),
    .B(_03898_),
    .Y(_04170_));
 OAI21x1_ASAP7_75t_R _26945_ (.A1(_04163_),
    .A2(_04170_),
    .B(_03790_),
    .Y(_04171_));
 NOR2x1_ASAP7_75t_R _26946_ (.A(_03692_),
    .B(_03796_),
    .Y(_04172_));
 AO21x1_ASAP7_75t_R _26947_ (.A1(_03957_),
    .A2(_03771_),
    .B(_03775_),
    .Y(_04173_));
 OAI21x1_ASAP7_75t_R _26948_ (.A1(_04172_),
    .A2(_04173_),
    .B(_03898_),
    .Y(_04174_));
 AO21x1_ASAP7_75t_R _26949_ (.A1(_03781_),
    .A2(_03964_),
    .B(_03895_),
    .Y(_04175_));
 AOI21x1_ASAP7_75t_R _26950_ (.A1(_03864_),
    .A2(_04175_),
    .B(_03739_),
    .Y(_04176_));
 NOR2x1_ASAP7_75t_R _26951_ (.A(_04174_),
    .B(_04176_),
    .Y(_04177_));
 NAND2x1_ASAP7_75t_R _26952_ (.A(net833),
    .B(net925),
    .Y(_04178_));
 AOI21x1_ASAP7_75t_R _26953_ (.A1(_03798_),
    .A2(_04178_),
    .B(_03771_),
    .Y(_04179_));
 INVx1_ASAP7_75t_R _26954_ (.A(_04179_),
    .Y(_04180_));
 NOR2x1_ASAP7_75t_R _26955_ (.A(_03729_),
    .B(_03749_),
    .Y(_04181_));
 AO21x1_ASAP7_75t_R _26956_ (.A1(_00600_),
    .A2(_03755_),
    .B(_03699_),
    .Y(_04182_));
 NOR2x1_ASAP7_75t_R _26957_ (.A(_03932_),
    .B(_04182_),
    .Y(_04183_));
 AOI21x1_ASAP7_75t_R _26958_ (.A1(_04180_),
    .A2(_04181_),
    .B(_04183_),
    .Y(_04184_));
 OAI21x1_ASAP7_75t_R _26959_ (.A1(_03898_),
    .A2(_04184_),
    .B(_03821_),
    .Y(_04185_));
 NOR2x1_ASAP7_75t_R _26960_ (.A(_04177_),
    .B(_04185_),
    .Y(_04186_));
 NOR2x1_ASAP7_75t_R _26961_ (.A(_04171_),
    .B(_04186_),
    .Y(_04187_));
 NOR2x1_ASAP7_75t_R _26962_ (.A(_04158_),
    .B(_04187_),
    .Y(_00117_));
 AOI211x1_ASAP7_75t_R _26963_ (.A1(_03873_),
    .A2(_03756_),
    .B(_03868_),
    .C(_03911_),
    .Y(_04188_));
 NAND2x1_ASAP7_75t_R _26964_ (.A(_00604_),
    .B(_03747_),
    .Y(_04189_));
 OAI21x1_ASAP7_75t_R _26965_ (.A1(_03922_),
    .A2(_03953_),
    .B(_04189_),
    .Y(_04190_));
 OAI21x1_ASAP7_75t_R _26966_ (.A1(_03945_),
    .A2(_04190_),
    .B(_03860_),
    .Y(_04191_));
 OAI21x1_ASAP7_75t_R _26967_ (.A1(_03922_),
    .A2(_03834_),
    .B(_04015_),
    .Y(_04192_));
 AOI21x1_ASAP7_75t_R _26968_ (.A1(_00600_),
    .A2(_15986_),
    .B(_03805_),
    .Y(_04193_));
 AOI21x1_ASAP7_75t_R _26969_ (.A1(_03803_),
    .A2(_04193_),
    .B(_03839_),
    .Y(_04194_));
 AOI21x1_ASAP7_75t_R _26970_ (.A1(_03945_),
    .A2(_04192_),
    .B(_04194_),
    .Y(_04195_));
 OAI22x1_ASAP7_75t_R _26971_ (.A1(_04188_),
    .A2(_04191_),
    .B1(_04195_),
    .B2(_03860_),
    .Y(_04196_));
 OAI21x1_ASAP7_75t_R _26972_ (.A1(_03823_),
    .A2(_04196_),
    .B(_03789_),
    .Y(_04197_));
 INVx1_ASAP7_75t_R _26973_ (.A(_04063_),
    .Y(_04198_));
 AOI21x1_ASAP7_75t_R _26974_ (.A1(_03736_),
    .A2(_04198_),
    .B(_03828_),
    .Y(_04199_));
 AOI21x1_ASAP7_75t_R _26975_ (.A1(_04178_),
    .A2(_04120_),
    .B(_03862_),
    .Y(_04200_));
 OAI21x1_ASAP7_75t_R _26976_ (.A1(_04199_),
    .A2(_04200_),
    .B(_03945_),
    .Y(_04201_));
 AND2x2_ASAP7_75t_R _26977_ (.A(_03761_),
    .B(_03970_),
    .Y(_04202_));
 OA21x2_ASAP7_75t_R _26978_ (.A1(_04043_),
    .A2(_04042_),
    .B(_03862_),
    .Y(_04203_));
 OAI21x1_ASAP7_75t_R _26979_ (.A1(_04202_),
    .A2(_04203_),
    .B(_03911_),
    .Y(_04204_));
 AOI21x1_ASAP7_75t_R _26980_ (.A1(_04201_),
    .A2(_04204_),
    .B(_03821_),
    .Y(_04205_));
 AND3x2_ASAP7_75t_R _26981_ (.A(_15986_),
    .B(_03676_),
    .C(_03771_),
    .Y(_04206_));
 OAI21x1_ASAP7_75t_R _26982_ (.A1(_04206_),
    .A2(_04179_),
    .B(_03911_),
    .Y(_04207_));
 NAND2x1_ASAP7_75t_R _26983_ (.A(_03759_),
    .B(_03761_),
    .Y(_04208_));
 AO21x1_ASAP7_75t_R _26984_ (.A1(_04208_),
    .A2(_03924_),
    .B(_03856_),
    .Y(_04209_));
 AOI21x1_ASAP7_75t_R _26985_ (.A1(_04207_),
    .A2(_04209_),
    .B(_03860_),
    .Y(_04210_));
 NOR3x2_ASAP7_75t_R _26986_ (.B(_04210_),
    .C(_03765_),
    .Y(_04211_),
    .A(_04205_));
 OAI21x1_ASAP7_75t_R _26987_ (.A1(_03870_),
    .A2(_03942_),
    .B(_03747_),
    .Y(_04212_));
 NAND2x1_ASAP7_75t_R _26988_ (.A(_03816_),
    .B(_03913_),
    .Y(_04213_));
 NAND3x1_ASAP7_75t_R _26989_ (.A(_04212_),
    .B(_04213_),
    .C(_03688_),
    .Y(_04214_));
 AND2x2_ASAP7_75t_R _26990_ (.A(_01235_),
    .B(_01237_),
    .Y(_04215_));
 OA21x2_ASAP7_75t_R _26991_ (.A1(_03895_),
    .A2(_04215_),
    .B(_03825_),
    .Y(_04216_));
 NOR2x1_ASAP7_75t_R _26992_ (.A(net833),
    .B(net46),
    .Y(_04217_));
 OAI21x1_ASAP7_75t_R _26993_ (.A1(_04217_),
    .A2(_03922_),
    .B(_03747_),
    .Y(_04218_));
 AOI21x1_ASAP7_75t_R _26994_ (.A1(_04216_),
    .A2(_04218_),
    .B(_03753_),
    .Y(_04219_));
 AOI21x1_ASAP7_75t_R _26995_ (.A1(_04214_),
    .A2(_04219_),
    .B(_03765_),
    .Y(_04220_));
 OA21x2_ASAP7_75t_R _26996_ (.A1(_03653_),
    .A2(net872),
    .B(_00599_),
    .Y(_04221_));
 OAI21x1_ASAP7_75t_R _26997_ (.A1(_03774_),
    .A2(_04221_),
    .B(_03862_),
    .Y(_04222_));
 NAND2x2_ASAP7_75t_R _26998_ (.A(_03779_),
    .B(_04070_),
    .Y(_04223_));
 AOI21x1_ASAP7_75t_R _26999_ (.A1(_04222_),
    .A2(_04223_),
    .B(_03839_),
    .Y(_04224_));
 NAND2x1_ASAP7_75t_R _27000_ (.A(_03808_),
    .B(_03734_),
    .Y(_04225_));
 OAI21x1_ASAP7_75t_R _27001_ (.A1(_03942_),
    .A2(_03845_),
    .B(_03862_),
    .Y(_04226_));
 AOI21x1_ASAP7_75t_R _27002_ (.A1(_04225_),
    .A2(_04226_),
    .B(_03856_),
    .Y(_04227_));
 OAI21x1_ASAP7_75t_R _27003_ (.A1(_04224_),
    .A2(_04227_),
    .B(_03821_),
    .Y(_04228_));
 AOI21x1_ASAP7_75t_R _27004_ (.A1(_04220_),
    .A2(_04228_),
    .B(_03789_),
    .Y(_04229_));
 INVx1_ASAP7_75t_R _27005_ (.A(_04125_),
    .Y(_04230_));
 OAI21x1_ASAP7_75t_R _27006_ (.A1(_04105_),
    .A2(_04230_),
    .B(_03826_),
    .Y(_04231_));
 INVx1_ASAP7_75t_R _27007_ (.A(_03671_),
    .Y(_04232_));
 OAI21x1_ASAP7_75t_R _27008_ (.A1(_04232_),
    .A2(_04030_),
    .B(_03828_),
    .Y(_04233_));
 AOI21x1_ASAP7_75t_R _27009_ (.A1(_03867_),
    .A2(_04125_),
    .B(_03688_),
    .Y(_04234_));
 NAND2x1_ASAP7_75t_R _27010_ (.A(_04233_),
    .B(_04234_),
    .Y(_04235_));
 AOI21x1_ASAP7_75t_R _27011_ (.A1(_04231_),
    .A2(_04235_),
    .B(_03860_),
    .Y(_04236_));
 AO21x1_ASAP7_75t_R _27012_ (.A1(_03964_),
    .A2(_03795_),
    .B(_03694_),
    .Y(_04237_));
 OAI21x1_ASAP7_75t_R _27013_ (.A1(_03922_),
    .A2(_04067_),
    .B(_04237_),
    .Y(_04238_));
 AO21x1_ASAP7_75t_R _27014_ (.A1(_03677_),
    .A2(_03816_),
    .B(_03825_),
    .Y(_04239_));
 OAI21x1_ASAP7_75t_R _27015_ (.A1(_04239_),
    .A2(_04007_),
    .B(_03741_),
    .Y(_04240_));
 AOI21x1_ASAP7_75t_R _27016_ (.A1(_03911_),
    .A2(_04238_),
    .B(_04240_),
    .Y(_04241_));
 OAI21x1_ASAP7_75t_R _27017_ (.A1(_04236_),
    .A2(_04241_),
    .B(_03765_),
    .Y(_04242_));
 NAND2x1_ASAP7_75t_R _27018_ (.A(_04229_),
    .B(_04242_),
    .Y(_04243_));
 OAI21x1_ASAP7_75t_R _27019_ (.A1(_04197_),
    .A2(_04211_),
    .B(_04243_),
    .Y(_00118_));
 AOI21x1_ASAP7_75t_R _27020_ (.A1(_04020_),
    .A2(_03926_),
    .B(_03739_),
    .Y(_04244_));
 AOI21x1_ASAP7_75t_R _27021_ (.A1(_03995_),
    .A2(_04223_),
    .B(_03688_),
    .Y(_04245_));
 OAI21x1_ASAP7_75t_R _27022_ (.A1(_04244_),
    .A2(_04245_),
    .B(_03821_),
    .Y(_04246_));
 AOI21x1_ASAP7_75t_R _27023_ (.A1(_03816_),
    .A2(_03779_),
    .B(_03749_),
    .Y(_04247_));
 AOI21x1_ASAP7_75t_R _27024_ (.A1(_04247_),
    .A2(_04084_),
    .B(_03752_),
    .Y(_04248_));
 NAND2x1_ASAP7_75t_R _27025_ (.A(_03833_),
    .B(_03750_),
    .Y(_04249_));
 AOI21x1_ASAP7_75t_R _27026_ (.A1(net557),
    .A2(_03847_),
    .B(_03866_),
    .Y(_04250_));
 NAND2x1_ASAP7_75t_R _27027_ (.A(_04249_),
    .B(_04250_),
    .Y(_04251_));
 AOI21x1_ASAP7_75t_R _27028_ (.A1(_04248_),
    .A2(_04251_),
    .B(_03898_),
    .Y(_04252_));
 NAND2x1_ASAP7_75t_R _27029_ (.A(_04252_),
    .B(_04246_),
    .Y(_04253_));
 NOR2x1_ASAP7_75t_R _27030_ (.A(_03670_),
    .B(_15981_),
    .Y(_04254_));
 AO21x1_ASAP7_75t_R _27031_ (.A1(_03812_),
    .A2(_03882_),
    .B(_04254_),
    .Y(_04255_));
 NAND2x1_ASAP7_75t_R _27032_ (.A(_03688_),
    .B(_04255_),
    .Y(_04256_));
 NAND3x1_ASAP7_75t_R _27033_ (.A(_03781_),
    .B(_03728_),
    .C(_03737_),
    .Y(_04257_));
 AOI21x1_ASAP7_75t_R _27034_ (.A1(_03983_),
    .A2(_04257_),
    .B(_03752_),
    .Y(_04258_));
 NAND2x1_ASAP7_75t_R _27035_ (.A(_04256_),
    .B(_04258_),
    .Y(_04259_));
 NOR2x1_ASAP7_75t_R _27036_ (.A(_03768_),
    .B(_03673_),
    .Y(_04260_));
 NAND2x1_ASAP7_75t_R _27037_ (.A(_15986_),
    .B(_04260_),
    .Y(_04261_));
 OA21x2_ASAP7_75t_R _27038_ (.A1(net901),
    .A2(_03895_),
    .B(_03825_),
    .Y(_04262_));
 AOI21x1_ASAP7_75t_R _27039_ (.A1(_04261_),
    .A2(_04262_),
    .B(_03713_),
    .Y(_04263_));
 AOI21x1_ASAP7_75t_R _27040_ (.A1(_03805_),
    .A2(_03728_),
    .B(_04125_),
    .Y(_04264_));
 OAI21x1_ASAP7_75t_R _27041_ (.A1(_04206_),
    .A2(_04264_),
    .B(_03839_),
    .Y(_04265_));
 AOI21x1_ASAP7_75t_R _27042_ (.A1(_04263_),
    .A2(_04265_),
    .B(_03721_),
    .Y(_04266_));
 AOI21x1_ASAP7_75t_R _27043_ (.A1(_04259_),
    .A2(_04266_),
    .B(_03790_),
    .Y(_04267_));
 NAND2x1_ASAP7_75t_R _27044_ (.A(_04267_),
    .B(_04253_),
    .Y(_04268_));
 NAND2x1_ASAP7_75t_R _27045_ (.A(_03728_),
    .B(_03809_),
    .Y(_04269_));
 AND3x1_ASAP7_75t_R _27046_ (.A(_04031_),
    .B(_03839_),
    .C(_04269_),
    .Y(_04270_));
 AO21x1_ASAP7_75t_R _27047_ (.A1(_15989_),
    .A2(_03902_),
    .B(_03700_),
    .Y(_04271_));
 AND3x1_ASAP7_75t_R _27048_ (.A(_03873_),
    .B(_03747_),
    .C(_03811_),
    .Y(_04272_));
 OAI21x1_ASAP7_75t_R _27049_ (.A1(_04271_),
    .A2(_04272_),
    .B(_03823_),
    .Y(_04273_));
 NOR2x1_ASAP7_75t_R _27050_ (.A(_04270_),
    .B(_04273_),
    .Y(_04274_));
 AOI21x1_ASAP7_75t_R _27051_ (.A1(_03816_),
    .A2(_03870_),
    .B(_03813_),
    .Y(_04275_));
 INVx1_ASAP7_75t_R _27052_ (.A(_04275_),
    .Y(_04276_));
 OAI21x1_ASAP7_75t_R _27053_ (.A1(_04260_),
    .A2(_04276_),
    .B(_03765_),
    .Y(_04277_));
 AOI211x1_ASAP7_75t_R _27054_ (.A1(_03828_),
    .A2(_03830_),
    .B(_03884_),
    .C(_03668_),
    .Y(_04278_));
 OAI21x1_ASAP7_75t_R _27055_ (.A1(_04277_),
    .A2(_04278_),
    .B(_03860_),
    .Y(_04279_));
 NAND2x1_ASAP7_75t_R _27056_ (.A(_03907_),
    .B(_04218_),
    .Y(_04280_));
 AOI21x1_ASAP7_75t_R _27057_ (.A1(_03747_),
    .A2(_03666_),
    .B(_03913_),
    .Y(_04281_));
 AOI21x1_ASAP7_75t_R _27058_ (.A1(_04275_),
    .A2(_04281_),
    .B(_03898_),
    .Y(_04282_));
 OAI21x1_ASAP7_75t_R _27059_ (.A1(_03911_),
    .A2(_04280_),
    .B(_04282_),
    .Y(_04283_));
 OA21x2_ASAP7_75t_R _27060_ (.A1(_01237_),
    .A2(_03737_),
    .B(_03825_),
    .Y(_04284_));
 AO21x1_ASAP7_75t_R _27061_ (.A1(_03671_),
    .A2(_03798_),
    .B(_03694_),
    .Y(_04285_));
 AOI21x1_ASAP7_75t_R _27062_ (.A1(_04284_),
    .A2(_04285_),
    .B(_03721_),
    .Y(_04286_));
 AOI21x1_ASAP7_75t_R _27063_ (.A1(_03781_),
    .A2(_03750_),
    .B(_03739_),
    .Y(_04287_));
 OAI21x1_ASAP7_75t_R _27064_ (.A1(_03690_),
    .A2(_03672_),
    .B(_04287_),
    .Y(_04288_));
 AOI21x1_ASAP7_75t_R _27065_ (.A1(_04286_),
    .A2(_04288_),
    .B(_03741_),
    .Y(_04289_));
 AOI21x1_ASAP7_75t_R _27066_ (.A1(_04283_),
    .A2(_04289_),
    .B(_03789_),
    .Y(_04290_));
 OAI21x1_ASAP7_75t_R _27067_ (.A1(_04274_),
    .A2(_04279_),
    .B(_04290_),
    .Y(_04291_));
 NAND2x1_ASAP7_75t_R _27068_ (.A(_04291_),
    .B(_04268_),
    .Y(_00119_));
 NOR2x1_ASAP7_75t_R _27069_ (.A(_12921_),
    .B(_00605_),
    .Y(_04292_));
 XOR2x2_ASAP7_75t_R _27070_ (.A(_13013_),
    .B(_12848_),
    .Y(_04293_));
 XOR2x1_ASAP7_75t_R _27071_ (.A(_12837_),
    .Y(_04294_),
    .B(_04293_));
 XOR2x1_ASAP7_75t_R _27072_ (.A(_01463_),
    .Y(_04295_),
    .B(_12873_));
 NAND2x1_ASAP7_75t_R _27073_ (.A(_04295_),
    .B(_04294_),
    .Y(_04296_));
 XOR2x1_ASAP7_75t_R _27074_ (.A(_12836_),
    .Y(_04297_),
    .B(_04293_));
 XOR2x1_ASAP7_75t_R _27075_ (.A(_12871_),
    .Y(_04298_),
    .B(_01463_));
 NAND2x1_ASAP7_75t_R _27076_ (.A(_04297_),
    .B(_04298_),
    .Y(_04299_));
 AOI21x1_ASAP7_75t_R _27077_ (.A1(_04299_),
    .A2(_04296_),
    .B(_10640_),
    .Y(_04300_));
 OAI21x1_ASAP7_75t_R _27078_ (.A1(_04300_),
    .A2(_04292_),
    .B(_00642_),
    .Y(_04301_));
 AND2x2_ASAP7_75t_R _27079_ (.A(_10643_),
    .B(_00605_),
    .Y(_04302_));
 NAND2x1_ASAP7_75t_R _27080_ (.A(_04297_),
    .B(_04295_),
    .Y(_04303_));
 NAND2x1_ASAP7_75t_R _27081_ (.A(_04294_),
    .B(_04298_),
    .Y(_04304_));
 AOI21x1_ASAP7_75t_R _27082_ (.A1(_04303_),
    .A2(_04304_),
    .B(_10640_),
    .Y(_04305_));
 INVx1_ASAP7_75t_R _27083_ (.A(_00642_),
    .Y(_04306_));
 OAI21x1_ASAP7_75t_R _27084_ (.A1(_04302_),
    .A2(_04305_),
    .B(_04306_),
    .Y(_04307_));
 NAND2x2_ASAP7_75t_R _27085_ (.A(_04301_),
    .B(_04307_),
    .Y(_04308_));
 BUFx16f_ASAP7_75t_R _27086_ (.A(_04308_),
    .Y(_15997_));
 XOR2x1_ASAP7_75t_R _27087_ (.A(net657),
    .Y(_04309_),
    .B(_12834_));
 NAND2x1_ASAP7_75t_R _27088_ (.A(_01702_),
    .B(_04309_),
    .Y(_04310_));
 INVx1_ASAP7_75t_R _27089_ (.A(_04309_),
    .Y(_04311_));
 NAND2x1_ASAP7_75t_R _27090_ (.A(_13011_),
    .B(_04311_),
    .Y(_04312_));
 INVx1_ASAP7_75t_R _27091_ (.A(_04293_),
    .Y(_04313_));
 AOI21x1_ASAP7_75t_R _27092_ (.A1(_04310_),
    .A2(_04312_),
    .B(_04313_),
    .Y(_04314_));
 XOR2x1_ASAP7_75t_R _27093_ (.A(_12834_),
    .Y(_04315_),
    .B(_13011_));
 NAND2x1_ASAP7_75t_R _27094_ (.A(net35),
    .B(_04315_),
    .Y(_04316_));
 INVx1_ASAP7_75t_R _27095_ (.A(_04315_),
    .Y(_04317_));
 NAND2x1_ASAP7_75t_R _27096_ (.A(_01485_),
    .B(_04317_),
    .Y(_04318_));
 AOI21x1_ASAP7_75t_R _27097_ (.A1(_04316_),
    .A2(_04318_),
    .B(_04293_),
    .Y(_04319_));
 OAI21x1_ASAP7_75t_R _27098_ (.A1(_04314_),
    .A2(_04319_),
    .B(_10743_),
    .Y(_04320_));
 INVx2_ASAP7_75t_R _27099_ (.A(_01121_),
    .Y(_04321_));
 NOR2x1_ASAP7_75t_R _27100_ (.A(_12921_),
    .B(_00606_),
    .Y(_04322_));
 INVx3_ASAP7_75t_R _27101_ (.A(_04322_),
    .Y(_04323_));
 NAND3x2_ASAP7_75t_R _27102_ (.B(_04321_),
    .C(_04323_),
    .Y(_04324_),
    .A(_04320_));
 AO21x1_ASAP7_75t_R _27103_ (.A1(_04320_),
    .A2(_04323_),
    .B(_04321_),
    .Y(_04325_));
 NAND2x2_ASAP7_75t_R _27104_ (.A(_04324_),
    .B(_04325_),
    .Y(_04326_));
 BUFx12f_ASAP7_75t_R _27105_ (.A(_04326_),
    .Y(_16000_));
 NOR2x2_ASAP7_75t_R _27106_ (.A(net667),
    .B(_00608_),
    .Y(_04327_));
 INVx4_ASAP7_75t_R _27107_ (.A(_04327_),
    .Y(_04328_));
 XOR2x2_ASAP7_75t_R _27108_ (.A(_12910_),
    .B(_12868_),
    .Y(_04329_));
 XOR2x1_ASAP7_75t_R _27109_ (.A(_04329_),
    .Y(_04330_),
    .B(_12880_));
 NOR2x1_ASAP7_75t_R _27110_ (.A(net878),
    .B(_04330_),
    .Y(_04331_));
 XNOR2x2_ASAP7_75t_R _27111_ (.A(_12831_),
    .B(_12836_),
    .Y(_04332_));
 XOR2x1_ASAP7_75t_R _27112_ (.A(_04329_),
    .Y(_04333_),
    .B(_01496_));
 NOR2x1_ASAP7_75t_R _27113_ (.A(_04332_),
    .B(_04333_),
    .Y(_04334_));
 OAI21x1_ASAP7_75t_R _27114_ (.A1(_04331_),
    .A2(_04334_),
    .B(net767),
    .Y(_04335_));
 INVx2_ASAP7_75t_R _27115_ (.A(_08111_),
    .Y(_04336_));
 AOI21x1_ASAP7_75t_R _27116_ (.A1(_04335_),
    .A2(_04328_),
    .B(_04336_),
    .Y(_04337_));
 NAND2x2_ASAP7_75t_R _27117_ (.A(_00608_),
    .B(_11373_),
    .Y(_04338_));
 NAND2x2_ASAP7_75t_R _27118_ (.A(_12880_),
    .B(_04332_),
    .Y(_04339_));
 NAND2x2_ASAP7_75t_R _27119_ (.A(_01496_),
    .B(net878),
    .Y(_04340_));
 INVx2_ASAP7_75t_R _27120_ (.A(_04329_),
    .Y(_04341_));
 NAND3x2_ASAP7_75t_R _27121_ (.B(_04340_),
    .C(_04341_),
    .Y(_04342_),
    .A(_04339_));
 NOR2x1_ASAP7_75t_R _27122_ (.A(_01496_),
    .B(net878),
    .Y(_04343_));
 NOR2x1_ASAP7_75t_R _27123_ (.A(_12880_),
    .B(_04332_),
    .Y(_04344_));
 OAI21x1_ASAP7_75t_R _27124_ (.A1(_04343_),
    .A2(_04344_),
    .B(_04329_),
    .Y(_04345_));
 NAND3x2_ASAP7_75t_R _27125_ (.B(_10742_),
    .C(_04345_),
    .Y(_04346_),
    .A(_04342_));
 AOI21x1_ASAP7_75t_R _27126_ (.A1(_04338_),
    .A2(_04346_),
    .B(_08111_),
    .Y(_04347_));
 NOR2x2_ASAP7_75t_R _27127_ (.A(_04337_),
    .B(_04347_),
    .Y(_04348_));
 BUFx12f_ASAP7_75t_R _27128_ (.A(_04348_),
    .Y(_04349_));
 BUFx6f_ASAP7_75t_R _27129_ (.A(_04349_),
    .Y(_16008_));
 INVx4_ASAP7_75t_R _27130_ (.A(_04308_),
    .Y(_15995_));
 AOI21x1_ASAP7_75t_R _27131_ (.A1(_04328_),
    .A2(_04335_),
    .B(_08111_),
    .Y(_04350_));
 AOI21x1_ASAP7_75t_R _27132_ (.A1(_04338_),
    .A2(_04346_),
    .B(_04336_),
    .Y(_04351_));
 NOR2x2_ASAP7_75t_R _27133_ (.A(_04350_),
    .B(_04351_),
    .Y(_04352_));
 BUFx10_ASAP7_75t_R _27134_ (.A(_04352_),
    .Y(_16005_));
 XOR2x2_ASAP7_75t_R _27135_ (.A(_01529_),
    .B(_00855_),
    .Y(_04353_));
 XOR2x1_ASAP7_75t_R _27136_ (.A(_00759_),
    .Y(_04354_),
    .B(_00791_));
 XNOR2x1_ASAP7_75t_R _27137_ (.B(_12880_),
    .Y(_04355_),
    .A(_13013_));
 XNOR2x2_ASAP7_75t_R _27138_ (.A(_04354_),
    .B(_04355_),
    .Y(_04356_));
 OAI21x1_ASAP7_75t_R _27139_ (.A1(_04353_),
    .A2(_04356_),
    .B(net867),
    .Y(_04357_));
 AND2x2_ASAP7_75t_R _27140_ (.A(_04356_),
    .B(_04353_),
    .Y(_04358_));
 NAND2x1_ASAP7_75t_R _27141_ (.A(_00710_),
    .B(_11441_),
    .Y(_04359_));
 OAI21x1_ASAP7_75t_R _27142_ (.A1(_04357_),
    .A2(_04358_),
    .B(_04359_),
    .Y(_04360_));
 XOR2x2_ASAP7_75t_R _27143_ (.A(_04360_),
    .B(_08124_),
    .Y(_04361_));
 BUFx6f_ASAP7_75t_R _27144_ (.A(_04361_),
    .Y(_04362_));
 INVx1_ASAP7_75t_R _27145_ (.A(_01239_),
    .Y(_04363_));
 OA21x2_ASAP7_75t_R _27146_ (.A1(_04347_),
    .A2(_04337_),
    .B(_04363_),
    .Y(_04364_));
 NAND2x2_ASAP7_75t_R _27147_ (.A(_04362_),
    .B(_04364_),
    .Y(_04365_));
 OAI21x1_ASAP7_75t_R _27148_ (.A1(_04350_),
    .A2(_04351_),
    .B(_00607_),
    .Y(_04366_));
 OAI21x1_ASAP7_75t_R _27149_ (.A1(net598),
    .A2(_04347_),
    .B(_00612_),
    .Y(_04367_));
 AO21x1_ASAP7_75t_R _27150_ (.A1(_04366_),
    .A2(_04367_),
    .B(_04362_),
    .Y(_04368_));
 XOR2x2_ASAP7_75t_R _27151_ (.A(_13013_),
    .B(_00855_),
    .Y(_04369_));
 XOR2x2_ASAP7_75t_R _27152_ (.A(_12959_),
    .B(_04369_),
    .Y(_04370_));
 XOR2x1_ASAP7_75t_R _27153_ (.A(_04370_),
    .Y(_04371_),
    .B(_01561_));
 NOR2x2_ASAP7_75t_R _27154_ (.A(_10742_),
    .B(_00704_),
    .Y(_04372_));
 AO21x1_ASAP7_75t_R _27155_ (.A1(_04371_),
    .A2(net763),
    .B(_04372_),
    .Y(_04373_));
 BUFx2_ASAP7_75t_R _27156_ (.A(_04373_),
    .Y(_04374_));
 XOR2x2_ASAP7_75t_R _27157_ (.A(_04374_),
    .B(_08133_),
    .Y(_04375_));
 BUFx10_ASAP7_75t_R _27158_ (.A(_04375_),
    .Y(_04376_));
 AOI21x1_ASAP7_75t_R _27159_ (.A1(_04365_),
    .A2(_04368_),
    .B(_04376_),
    .Y(_04377_));
 INVx1_ASAP7_75t_R _27160_ (.A(_04367_),
    .Y(_04378_));
 INVx1_ASAP7_75t_R _27161_ (.A(_01241_),
    .Y(_04379_));
 OA21x2_ASAP7_75t_R _27162_ (.A1(_04351_),
    .A2(_04350_),
    .B(_04379_),
    .Y(_04380_));
 BUFx6f_ASAP7_75t_R _27163_ (.A(_04361_),
    .Y(_04381_));
 OAI21x1_ASAP7_75t_R _27164_ (.A1(_04378_),
    .A2(_04380_),
    .B(_04381_),
    .Y(_04382_));
 BUFx10_ASAP7_75t_R _27165_ (.A(_04361_),
    .Y(_04383_));
 NAND3x2_ASAP7_75t_R _27166_ (.B(_04336_),
    .C(_04328_),
    .Y(_04384_),
    .A(_04335_));
 CKINVDCx5p33_ASAP7_75t_R _27167_ (.A(_04337_),
    .Y(_04385_));
 AO21x2_ASAP7_75t_R _27168_ (.A1(_04384_),
    .A2(_04385_),
    .B(_01239_),
    .Y(_04386_));
 NOR2x2_ASAP7_75t_R _27169_ (.A(_04383_),
    .B(_04386_),
    .Y(_04387_));
 INVx1_ASAP7_75t_R _27170_ (.A(_04387_),
    .Y(_04388_));
 INVx1_ASAP7_75t_R _27171_ (.A(_08133_),
    .Y(_04389_));
 XOR2x2_ASAP7_75t_R _27172_ (.A(_04374_),
    .B(_04389_),
    .Y(_04390_));
 BUFx6f_ASAP7_75t_R _27173_ (.A(_04390_),
    .Y(_04391_));
 AOI21x1_ASAP7_75t_R _27174_ (.A1(_04382_),
    .A2(_04388_),
    .B(_04391_),
    .Y(_04392_));
 NOR2x1_ASAP7_75t_R _27175_ (.A(_10742_),
    .B(_00703_),
    .Y(_04393_));
 INVx2_ASAP7_75t_R _27176_ (.A(_04393_),
    .Y(_04394_));
 XOR2x1_ASAP7_75t_R _27177_ (.A(_12902_),
    .Y(_04395_),
    .B(_00793_));
 NAND2x1_ASAP7_75t_R _27178_ (.A(_12956_),
    .B(_04395_),
    .Y(_04396_));
 NAND2x1_ASAP7_75t_R _27179_ (.A(_12955_),
    .B(_12903_),
    .Y(_04397_));
 INVx1_ASAP7_75t_R _27180_ (.A(_12931_),
    .Y(_04398_));
 AOI21x1_ASAP7_75t_R _27181_ (.A1(_04396_),
    .A2(_04397_),
    .B(_04398_),
    .Y(_04399_));
 NOR2x1_ASAP7_75t_R _27182_ (.A(_12955_),
    .B(_04395_),
    .Y(_04400_));
 NOR2x1_ASAP7_75t_R _27183_ (.A(_12956_),
    .B(_12903_),
    .Y(_04401_));
 OAI21x1_ASAP7_75t_R _27184_ (.A1(_04400_),
    .A2(_04401_),
    .B(_04398_),
    .Y(_04402_));
 INVx1_ASAP7_75t_R _27185_ (.A(_04402_),
    .Y(_04403_));
 OAI21x1_ASAP7_75t_R _27186_ (.A1(_04399_),
    .A2(_04403_),
    .B(net763),
    .Y(_04404_));
 NAND2x1_ASAP7_75t_R _27187_ (.A(_04394_),
    .B(_04404_),
    .Y(_04405_));
 XNOR2x2_ASAP7_75t_R _27188_ (.A(_01095_),
    .B(_04405_),
    .Y(_04406_));
 BUFx6f_ASAP7_75t_R _27189_ (.A(_04406_),
    .Y(_04407_));
 OAI21x1_ASAP7_75t_R _27190_ (.A1(_04377_),
    .A2(_04392_),
    .B(_04407_),
    .Y(_04408_));
 BUFx10_ASAP7_75t_R _27191_ (.A(_04390_),
    .Y(_04409_));
 BUFx6f_ASAP7_75t_R _27192_ (.A(_04383_),
    .Y(_04410_));
 INVx3_ASAP7_75t_R _27193_ (.A(_04350_),
    .Y(_04411_));
 NAND3x2_ASAP7_75t_R _27194_ (.B(_08111_),
    .C(_04328_),
    .Y(_04412_),
    .A(_04335_));
 AOI21x1_ASAP7_75t_R _27195_ (.A1(_04411_),
    .A2(_04412_),
    .B(_00610_),
    .Y(_04413_));
 BUFx4f_ASAP7_75t_R _27196_ (.A(_04361_),
    .Y(_04414_));
 NAND2x1_ASAP7_75t_R _27197_ (.A(_01244_),
    .B(_04414_),
    .Y(_04415_));
 OAI21x1_ASAP7_75t_R _27198_ (.A1(_04410_),
    .A2(net458),
    .B(_04415_),
    .Y(_04416_));
 AOI21x1_ASAP7_75t_R _27199_ (.A1(_04409_),
    .A2(_04416_),
    .B(_04407_),
    .Y(_04417_));
 XOR2x2_ASAP7_75t_R _27200_ (.A(_04360_),
    .B(_08958_),
    .Y(_04418_));
 BUFx6f_ASAP7_75t_R _27201_ (.A(_04418_),
    .Y(_04419_));
 BUFx3_ASAP7_75t_R _27202_ (.A(_01240_),
    .Y(_04420_));
 INVx2_ASAP7_75t_R _27203_ (.A(_04420_),
    .Y(_04421_));
 OAI21x1_ASAP7_75t_R _27204_ (.A1(_04350_),
    .A2(_04351_),
    .B(_04421_),
    .Y(_04422_));
 NAND2x1_ASAP7_75t_R _27205_ (.A(_04367_),
    .B(_04422_),
    .Y(_04423_));
 AOI21x1_ASAP7_75t_R _27206_ (.A1(_04419_),
    .A2(_04423_),
    .B(_04390_),
    .Y(_04424_));
 NAND3x2_ASAP7_75t_R _27207_ (.B(_01121_),
    .C(_04323_),
    .Y(_04425_),
    .A(_04320_));
 AO21x2_ASAP7_75t_R _27208_ (.A1(_04320_),
    .A2(_04323_),
    .B(_01121_),
    .Y(_04426_));
 NAND2x2_ASAP7_75t_R _27209_ (.A(_04426_),
    .B(_04425_),
    .Y(_15994_));
 AOI21x1_ASAP7_75t_R _27210_ (.A1(net48),
    .A2(_04349_),
    .B(_04418_),
    .Y(_04427_));
 NOR2x2_ASAP7_75t_R _27211_ (.A(net467),
    .B(_04348_),
    .Y(_04428_));
 INVx1_ASAP7_75t_R _27212_ (.A(_04428_),
    .Y(_04429_));
 OAI21x1_ASAP7_75t_R _27213_ (.A1(_04350_),
    .A2(_04351_),
    .B(_04363_),
    .Y(_04430_));
 NOR2x2_ASAP7_75t_R _27214_ (.A(_04383_),
    .B(_04430_),
    .Y(_04431_));
 AOI21x1_ASAP7_75t_R _27215_ (.A1(_04427_),
    .A2(_04429_),
    .B(_04431_),
    .Y(_04432_));
 NAND2x1_ASAP7_75t_R _27216_ (.A(_04424_),
    .B(_04432_),
    .Y(_04433_));
 XOR2x1_ASAP7_75t_R _27217_ (.A(_12955_),
    .Y(_04434_),
    .B(_00858_));
 XOR2x1_ASAP7_75t_R _27218_ (.A(_04434_),
    .Y(_04435_),
    .B(_00825_));
 XOR2x1_ASAP7_75t_R _27219_ (.A(_04435_),
    .Y(_04436_),
    .B(_13015_));
 NOR2x1_ASAP7_75t_R _27220_ (.A(_10829_),
    .B(_00702_),
    .Y(_04437_));
 AO21x1_ASAP7_75t_R _27221_ (.A1(_04436_),
    .A2(_11451_),
    .B(_04437_),
    .Y(_04438_));
 XNOR2x2_ASAP7_75t_R _27222_ (.A(_01096_),
    .B(_04438_),
    .Y(_04439_));
 AOI21x1_ASAP7_75t_R _27223_ (.A1(_04417_),
    .A2(_04433_),
    .B(_04439_),
    .Y(_04440_));
 XOR2x1_ASAP7_75t_R _27224_ (.A(_12851_),
    .Y(_04441_),
    .B(_01638_));
 INVx2_ASAP7_75t_R _27225_ (.A(net663),
    .Y(_04442_));
 XOR2x1_ASAP7_75t_R _27226_ (.A(_04441_),
    .Y(_04443_),
    .B(_04442_));
 NOR2x1_ASAP7_75t_R _27227_ (.A(_10786_),
    .B(_00701_),
    .Y(_04444_));
 AO21x1_ASAP7_75t_R _27228_ (.A1(_04443_),
    .A2(_13017_),
    .B(_04444_),
    .Y(_04445_));
 XOR2x2_ASAP7_75t_R _27229_ (.A(_04445_),
    .B(_01097_),
    .Y(_04446_));
 BUFx10_ASAP7_75t_R _27230_ (.A(_04446_),
    .Y(_04447_));
 AOI21x1_ASAP7_75t_R _27231_ (.A1(_04408_),
    .A2(_04440_),
    .B(_04447_),
    .Y(_04448_));
 OAI21x1_ASAP7_75t_R _27232_ (.A1(_16000_),
    .A2(_16005_),
    .B(_04362_),
    .Y(_04449_));
 BUFx6f_ASAP7_75t_R _27233_ (.A(_00611_),
    .Y(_04450_));
 AO21x2_ASAP7_75t_R _27234_ (.A1(_04384_),
    .A2(_04385_),
    .B(_04450_),
    .Y(_04451_));
 INVx1_ASAP7_75t_R _27235_ (.A(_04451_),
    .Y(_04452_));
 OAI21x1_ASAP7_75t_R _27236_ (.A1(_04449_),
    .A2(_04452_),
    .B(_04376_),
    .Y(_04453_));
 BUFx10_ASAP7_75t_R _27237_ (.A(_04352_),
    .Y(_04454_));
 BUFx6f_ASAP7_75t_R _27238_ (.A(_04418_),
    .Y(_04455_));
 AO21x1_ASAP7_75t_R _27239_ (.A1(_04454_),
    .A2(net491),
    .B(_04455_),
    .Y(_04456_));
 AOI21x1_ASAP7_75t_R _27240_ (.A1(_04385_),
    .A2(_04384_),
    .B(_01241_),
    .Y(_04457_));
 INVx2_ASAP7_75t_R _27241_ (.A(_04457_),
    .Y(_04458_));
 OA21x2_ASAP7_75t_R _27242_ (.A1(_04458_),
    .A2(_04414_),
    .B(_04390_),
    .Y(_04459_));
 NAND2x1_ASAP7_75t_R _27243_ (.A(_04456_),
    .B(_04459_),
    .Y(_04460_));
 INVx2_ASAP7_75t_R _27244_ (.A(_04422_),
    .Y(_04461_));
 BUFx6f_ASAP7_75t_R _27245_ (.A(_04418_),
    .Y(_04462_));
 AO21x1_ASAP7_75t_R _27246_ (.A1(_04461_),
    .A2(_04462_),
    .B(_04406_),
    .Y(_04463_));
 AOI21x1_ASAP7_75t_R _27247_ (.A1(_04453_),
    .A2(_04460_),
    .B(_04463_),
    .Y(_04464_));
 BUFx6f_ASAP7_75t_R _27248_ (.A(_04375_),
    .Y(_04465_));
 AOI21x1_ASAP7_75t_R _27249_ (.A1(_04420_),
    .A2(_04454_),
    .B(_04418_),
    .Y(_04466_));
 NOR2x1_ASAP7_75t_R _27250_ (.A(_04465_),
    .B(_04466_),
    .Y(_04467_));
 OAI21x1_ASAP7_75t_R _27251_ (.A1(_04350_),
    .A2(_04351_),
    .B(net467),
    .Y(_04468_));
 AO21x1_ASAP7_75t_R _27252_ (.A1(_04386_),
    .A2(_04468_),
    .B(_04414_),
    .Y(_04469_));
 NAND2x1_ASAP7_75t_R _27253_ (.A(_04467_),
    .B(_04469_),
    .Y(_04470_));
 INVx3_ASAP7_75t_R _27254_ (.A(_04413_),
    .Y(_04471_));
 AOI21x1_ASAP7_75t_R _27255_ (.A1(_15997_),
    .A2(_04352_),
    .B(_04361_),
    .Y(_04472_));
 AOI21x1_ASAP7_75t_R _27256_ (.A1(_04471_),
    .A2(_04472_),
    .B(_04391_),
    .Y(_04473_));
 NAND2x2_ASAP7_75t_R _27257_ (.A(_04326_),
    .B(_04352_),
    .Y(_04474_));
 BUFx6f_ASAP7_75t_R _27258_ (.A(_04418_),
    .Y(_04475_));
 AO21x1_ASAP7_75t_R _27259_ (.A1(_04474_),
    .A2(_04366_),
    .B(_04475_),
    .Y(_04476_));
 NAND2x1_ASAP7_75t_R _27260_ (.A(_04473_),
    .B(_04476_),
    .Y(_04477_));
 NAND3x2_ASAP7_75t_R _27261_ (.B(_01095_),
    .C(_04394_),
    .Y(_04478_),
    .A(_04404_));
 AO21x1_ASAP7_75t_R _27262_ (.A1(_04404_),
    .A2(_04394_),
    .B(_01095_),
    .Y(_04479_));
 NAND2x2_ASAP7_75t_R _27263_ (.A(_04478_),
    .B(_04479_),
    .Y(_04480_));
 BUFx10_ASAP7_75t_R _27264_ (.A(_04480_),
    .Y(_04481_));
 BUFx6f_ASAP7_75t_R _27265_ (.A(_04481_),
    .Y(_04482_));
 AOI21x1_ASAP7_75t_R _27266_ (.A1(_04470_),
    .A2(_04477_),
    .B(_04482_),
    .Y(_04483_));
 BUFx10_ASAP7_75t_R _27267_ (.A(_04439_),
    .Y(_04484_));
 OAI21x1_ASAP7_75t_R _27268_ (.A1(_04464_),
    .A2(_04483_),
    .B(_04484_),
    .Y(_04485_));
 NAND2x1_ASAP7_75t_R _27269_ (.A(_04448_),
    .B(_04485_),
    .Y(_04486_));
 BUFx6f_ASAP7_75t_R _27270_ (.A(_04475_),
    .Y(_04487_));
 INVx4_ASAP7_75t_R _27271_ (.A(net490),
    .Y(_04488_));
 AOI21x1_ASAP7_75t_R _27272_ (.A1(_04385_),
    .A2(_04384_),
    .B(_04488_),
    .Y(_04489_));
 INVx4_ASAP7_75t_R _27273_ (.A(_04489_),
    .Y(_04490_));
 NAND2x2_ASAP7_75t_R _27274_ (.A(_04348_),
    .B(net36),
    .Y(_04491_));
 NAND2x1_ASAP7_75t_R _27275_ (.A(_04490_),
    .B(_04491_),
    .Y(_04492_));
 AOI21x1_ASAP7_75t_R _27276_ (.A1(_04411_),
    .A2(_04412_),
    .B(_04488_),
    .Y(_04493_));
 OAI21x1_ASAP7_75t_R _27277_ (.A1(_04419_),
    .A2(net740),
    .B(_04391_),
    .Y(_04494_));
 AOI21x1_ASAP7_75t_R _27278_ (.A1(_04487_),
    .A2(_04492_),
    .B(_04494_),
    .Y(_04495_));
 OAI21x1_ASAP7_75t_R _27279_ (.A1(net598),
    .A2(_04347_),
    .B(_04488_),
    .Y(_04496_));
 BUFx6f_ASAP7_75t_R _27280_ (.A(_04496_),
    .Y(_04497_));
 AO21x1_ASAP7_75t_R _27281_ (.A1(_04468_),
    .A2(_04497_),
    .B(_04475_),
    .Y(_04498_));
 OAI21x1_ASAP7_75t_R _27282_ (.A1(net598),
    .A2(_04347_),
    .B(net468),
    .Y(_04499_));
 AO21x1_ASAP7_75t_R _27283_ (.A1(_04499_),
    .A2(_04366_),
    .B(_04381_),
    .Y(_04500_));
 AOI21x1_ASAP7_75t_R _27284_ (.A1(_04498_),
    .A2(_04500_),
    .B(_04409_),
    .Y(_04501_));
 OAI21x1_ASAP7_75t_R _27285_ (.A1(_04495_),
    .A2(_04501_),
    .B(_04482_),
    .Y(_04502_));
 OAI21x1_ASAP7_75t_R _27286_ (.A1(_04350_),
    .A2(_04351_),
    .B(_04450_),
    .Y(_04503_));
 AO21x1_ASAP7_75t_R _27287_ (.A1(_04497_),
    .A2(_04503_),
    .B(_04381_),
    .Y(_04504_));
 INVx1_ASAP7_75t_R _27288_ (.A(_04468_),
    .Y(_04505_));
 OA21x2_ASAP7_75t_R _27289_ (.A1(_04347_),
    .A2(net599),
    .B(_00607_),
    .Y(_04506_));
 BUFx10_ASAP7_75t_R _27290_ (.A(_04383_),
    .Y(_04507_));
 OAI21x1_ASAP7_75t_R _27291_ (.A1(_04505_),
    .A2(_04506_),
    .B(_04507_),
    .Y(_04508_));
 AOI21x1_ASAP7_75t_R _27292_ (.A1(_04504_),
    .A2(_04508_),
    .B(_04409_),
    .Y(_04509_));
 NAND2x2_ASAP7_75t_R _27293_ (.A(_15994_),
    .B(net36),
    .Y(_04510_));
 AOI21x1_ASAP7_75t_R _27294_ (.A1(_04326_),
    .A2(_04352_),
    .B(_04361_),
    .Y(_04511_));
 NAND2x1_ASAP7_75t_R _27295_ (.A(_04510_),
    .B(_04511_),
    .Y(_04512_));
 NOR2x2_ASAP7_75t_R _27296_ (.A(_15997_),
    .B(_16000_),
    .Y(_04513_));
 NOR2x2_ASAP7_75t_R _27297_ (.A(_15994_),
    .B(_04349_),
    .Y(_04514_));
 OAI21x1_ASAP7_75t_R _27298_ (.A1(_04513_),
    .A2(_04514_),
    .B(_04507_),
    .Y(_04515_));
 BUFx10_ASAP7_75t_R _27299_ (.A(_04375_),
    .Y(_04516_));
 AOI21x1_ASAP7_75t_R _27300_ (.A1(_04512_),
    .A2(_04515_),
    .B(_04516_),
    .Y(_04517_));
 BUFx10_ASAP7_75t_R _27301_ (.A(_04407_),
    .Y(_04518_));
 OAI21x1_ASAP7_75t_R _27302_ (.A1(_04509_),
    .A2(_04517_),
    .B(_04518_),
    .Y(_04519_));
 AOI21x1_ASAP7_75t_R _27303_ (.A1(_04502_),
    .A2(_04519_),
    .B(_04484_),
    .Y(_04520_));
 INVx1_ASAP7_75t_R _27304_ (.A(_01242_),
    .Y(_04521_));
 AO21x2_ASAP7_75t_R _27305_ (.A1(_04412_),
    .A2(_04411_),
    .B(_04521_),
    .Y(_04522_));
 INVx1_ASAP7_75t_R _27306_ (.A(_04522_),
    .Y(_04523_));
 NAND2x2_ASAP7_75t_R _27307_ (.A(net48),
    .B(_04454_),
    .Y(_04524_));
 INVx3_ASAP7_75t_R _27308_ (.A(net741),
    .Y(_04525_));
 AOI21x1_ASAP7_75t_R _27309_ (.A1(_04525_),
    .A2(_04349_),
    .B(_04383_),
    .Y(_04526_));
 NAND2x2_ASAP7_75t_R _27310_ (.A(_04524_),
    .B(_04526_),
    .Y(_04527_));
 OAI21x1_ASAP7_75t_R _27311_ (.A1(_04456_),
    .A2(_04523_),
    .B(_04527_),
    .Y(_04528_));
 NOR2x1_ASAP7_75t_R _27312_ (.A(_08133_),
    .B(_04374_),
    .Y(_04529_));
 XOR2x1_ASAP7_75t_R _27313_ (.A(_04370_),
    .Y(_04530_),
    .B(_01565_));
 NOR2x1_ASAP7_75t_R _27314_ (.A(_12161_),
    .B(_04530_),
    .Y(_04531_));
 OAI21x1_ASAP7_75t_R _27315_ (.A1(_04372_),
    .A2(_04531_),
    .B(_08133_),
    .Y(_04532_));
 INVx1_ASAP7_75t_R _27316_ (.A(_04532_),
    .Y(_04533_));
 OAI21x1_ASAP7_75t_R _27317_ (.A1(_04529_),
    .A2(_04533_),
    .B(_04406_),
    .Y(_04534_));
 INVx3_ASAP7_75t_R _27318_ (.A(_04534_),
    .Y(_04535_));
 AOI21x1_ASAP7_75t_R _27319_ (.A1(net48),
    .A2(_04349_),
    .B(_04361_),
    .Y(_04536_));
 INVx1_ASAP7_75t_R _27320_ (.A(_04536_),
    .Y(_04537_));
 AO21x1_ASAP7_75t_R _27321_ (.A1(_04412_),
    .A2(_04411_),
    .B(net742),
    .Y(_04538_));
 NAND2x1_ASAP7_75t_R _27322_ (.A(_04538_),
    .B(_04466_),
    .Y(_04539_));
 NOR2x1_ASAP7_75t_R _27323_ (.A(_04389_),
    .B(_04374_),
    .Y(_04540_));
 AND2x2_ASAP7_75t_R _27324_ (.A(_04374_),
    .B(_04389_),
    .Y(_04541_));
 OAI21x1_ASAP7_75t_R _27325_ (.A1(_04540_),
    .A2(_04541_),
    .B(_04406_),
    .Y(_04542_));
 AOI21x1_ASAP7_75t_R _27326_ (.A1(_04537_),
    .A2(_04539_),
    .B(_04542_),
    .Y(_04543_));
 AOI21x1_ASAP7_75t_R _27327_ (.A1(_04528_),
    .A2(_04535_),
    .B(_04543_),
    .Y(_04544_));
 NAND2x1_ASAP7_75t_R _27328_ (.A(_04451_),
    .B(_04427_),
    .Y(_04545_));
 NOR2x2_ASAP7_75t_R _27329_ (.A(_15997_),
    .B(_04454_),
    .Y(_04546_));
 BUFx6f_ASAP7_75t_R _27330_ (.A(_04455_),
    .Y(_04547_));
 OAI21x1_ASAP7_75t_R _27331_ (.A1(_04364_),
    .A2(_04546_),
    .B(_04547_),
    .Y(_04548_));
 AOI21x1_ASAP7_75t_R _27332_ (.A1(_04545_),
    .A2(_04548_),
    .B(_04409_),
    .Y(_04549_));
 AO21x2_ASAP7_75t_R _27333_ (.A1(_04384_),
    .A2(_04385_),
    .B(_04521_),
    .Y(_04550_));
 NAND2x1_ASAP7_75t_R _27334_ (.A(_04550_),
    .B(_04427_),
    .Y(_04551_));
 NOR2x2_ASAP7_75t_R _27335_ (.A(_04525_),
    .B(_04454_),
    .Y(_04552_));
 AOI22x1_ASAP7_75t_R _27336_ (.A1(_04384_),
    .A2(_04385_),
    .B1(_04301_),
    .B2(_04307_),
    .Y(_04553_));
 OAI21x1_ASAP7_75t_R _27337_ (.A1(_04552_),
    .A2(_04553_),
    .B(_04547_),
    .Y(_04554_));
 BUFx6f_ASAP7_75t_R _27338_ (.A(_04375_),
    .Y(_04555_));
 AOI21x1_ASAP7_75t_R _27339_ (.A1(_04551_),
    .A2(_04554_),
    .B(_04555_),
    .Y(_04556_));
 BUFx10_ASAP7_75t_R _27340_ (.A(_04481_),
    .Y(_04557_));
 OAI21x1_ASAP7_75t_R _27341_ (.A1(_04549_),
    .A2(_04556_),
    .B(_04557_),
    .Y(_04558_));
 INVx6_ASAP7_75t_R _27342_ (.A(_04439_),
    .Y(_04559_));
 BUFx10_ASAP7_75t_R _27343_ (.A(_04559_),
    .Y(_04560_));
 AOI21x1_ASAP7_75t_R _27344_ (.A1(_04544_),
    .A2(_04558_),
    .B(_04560_),
    .Y(_04561_));
 OAI21x1_ASAP7_75t_R _27345_ (.A1(_04520_),
    .A2(_04561_),
    .B(_04447_),
    .Y(_04562_));
 NAND2x1_ASAP7_75t_R _27346_ (.A(_04486_),
    .B(_04562_),
    .Y(_00120_));
 NAND2x2_ASAP7_75t_R _27347_ (.A(_04308_),
    .B(_04349_),
    .Y(_04563_));
 AO21x1_ASAP7_75t_R _27348_ (.A1(_04511_),
    .A2(_04563_),
    .B(_04406_),
    .Y(_04564_));
 AO21x1_ASAP7_75t_R _27349_ (.A1(_04466_),
    .A2(_04491_),
    .B(_04465_),
    .Y(_04565_));
 OAI21x1_ASAP7_75t_R _27350_ (.A1(_04564_),
    .A2(_04565_),
    .B(_04559_),
    .Y(_04566_));
 INVx1_ASAP7_75t_R _27351_ (.A(_04524_),
    .Y(_04567_));
 INVx1_ASAP7_75t_R _27352_ (.A(net467),
    .Y(_04568_));
 AO21x1_ASAP7_75t_R _27353_ (.A1(_16008_),
    .A2(_04568_),
    .B(_04362_),
    .Y(_04569_));
 OAI21x1_ASAP7_75t_R _27354_ (.A1(_04567_),
    .A2(_04569_),
    .B(_04535_),
    .Y(_04570_));
 AOI21x1_ASAP7_75t_R _27355_ (.A1(_04525_),
    .A2(_04349_),
    .B(_04418_),
    .Y(_04571_));
 AND2x2_ASAP7_75t_R _27356_ (.A(_04571_),
    .B(_04451_),
    .Y(_04572_));
 INVx1_ASAP7_75t_R _27357_ (.A(_00613_),
    .Y(_04573_));
 NAND2x1_ASAP7_75t_R _27358_ (.A(_04362_),
    .B(_04481_),
    .Y(_04574_));
 NOR2x1_ASAP7_75t_R _27359_ (.A(_04573_),
    .B(_04574_),
    .Y(_04575_));
 NOR2x1_ASAP7_75t_R _27360_ (.A(_00607_),
    .B(_16005_),
    .Y(_04576_));
 OAI21x1_ASAP7_75t_R _27361_ (.A1(_04450_),
    .A2(_04349_),
    .B(_04418_),
    .Y(_04577_));
 OAI21x1_ASAP7_75t_R _27362_ (.A1(_04576_),
    .A2(_04577_),
    .B(_04376_),
    .Y(_04578_));
 OAI22x1_ASAP7_75t_R _27363_ (.A1(_04570_),
    .A2(_04572_),
    .B1(_04575_),
    .B2(_04578_),
    .Y(_04579_));
 NOR2x1_ASAP7_75t_R _27364_ (.A(_04566_),
    .B(_04579_),
    .Y(_04580_));
 BUFx6f_ASAP7_75t_R _27365_ (.A(_04465_),
    .Y(_04581_));
 INVx2_ASAP7_75t_R _27366_ (.A(_04550_),
    .Y(_04582_));
 BUFx6f_ASAP7_75t_R _27367_ (.A(_04348_),
    .Y(_04583_));
 AO21x2_ASAP7_75t_R _27368_ (.A1(_04583_),
    .A2(_01239_),
    .B(_04414_),
    .Y(_04584_));
 INVx1_ASAP7_75t_R _27369_ (.A(_04450_),
    .Y(_04585_));
 AOI21x1_ASAP7_75t_R _27370_ (.A1(_04585_),
    .A2(_04583_),
    .B(_04455_),
    .Y(_04586_));
 NAND2x2_ASAP7_75t_R _27371_ (.A(_04497_),
    .B(_04586_),
    .Y(_04587_));
 OAI21x1_ASAP7_75t_R _27372_ (.A1(_04582_),
    .A2(_04584_),
    .B(_04587_),
    .Y(_04588_));
 NAND2x1_ASAP7_75t_R _27373_ (.A(_04451_),
    .B(_04536_),
    .Y(_04589_));
 OA21x2_ASAP7_75t_R _27374_ (.A1(_04475_),
    .A2(_04489_),
    .B(_04375_),
    .Y(_04590_));
 AOI21x1_ASAP7_75t_R _27375_ (.A1(_04589_),
    .A2(_04590_),
    .B(_04407_),
    .Y(_04591_));
 OAI21x1_ASAP7_75t_R _27376_ (.A1(_04581_),
    .A2(_04588_),
    .B(_04591_),
    .Y(_04592_));
 AOI21x1_ASAP7_75t_R _27377_ (.A1(_04419_),
    .A2(_04364_),
    .B(_04465_),
    .Y(_04593_));
 NOR2x2_ASAP7_75t_R _27378_ (.A(_15994_),
    .B(_04352_),
    .Y(_04594_));
 NAND2x1_ASAP7_75t_R _27379_ (.A(_04475_),
    .B(_04594_),
    .Y(_04595_));
 AOI21x1_ASAP7_75t_R _27380_ (.A1(_04385_),
    .A2(_04384_),
    .B(_04568_),
    .Y(_04596_));
 OAI21x1_ASAP7_75t_R _27381_ (.A1(_04596_),
    .A2(net458),
    .B(_04381_),
    .Y(_04597_));
 NAND3x1_ASAP7_75t_R _27382_ (.A(_04593_),
    .B(_04595_),
    .C(_04597_),
    .Y(_04598_));
 NAND2x1_ASAP7_75t_R _27383_ (.A(_04491_),
    .B(_04466_),
    .Y(_04599_));
 AO21x1_ASAP7_75t_R _27384_ (.A1(_04412_),
    .A2(_04411_),
    .B(net467),
    .Y(_04600_));
 AOI21x1_ASAP7_75t_R _27385_ (.A1(_04600_),
    .A2(_04511_),
    .B(_04391_),
    .Y(_04601_));
 AOI21x1_ASAP7_75t_R _27386_ (.A1(_04599_),
    .A2(_04601_),
    .B(_04481_),
    .Y(_04602_));
 NAND2x1_ASAP7_75t_R _27387_ (.A(_04598_),
    .B(_04602_),
    .Y(_04603_));
 AOI21x1_ASAP7_75t_R _27388_ (.A1(_04592_),
    .A2(_04603_),
    .B(_04560_),
    .Y(_04604_));
 OAI21x1_ASAP7_75t_R _27389_ (.A1(_04580_),
    .A2(_04604_),
    .B(_04447_),
    .Y(_04605_));
 NOR2x2_ASAP7_75t_R _27390_ (.A(_04308_),
    .B(_04349_),
    .Y(_04606_));
 NAND2x1_ASAP7_75t_R _27391_ (.A(_04419_),
    .B(_04606_),
    .Y(_04607_));
 NOR2x2_ASAP7_75t_R _27392_ (.A(_04420_),
    .B(_04383_),
    .Y(_04608_));
 INVx1_ASAP7_75t_R _27393_ (.A(_00614_),
    .Y(_04609_));
 NOR2x1_ASAP7_75t_R _27394_ (.A(_04609_),
    .B(_04455_),
    .Y(_04610_));
 AOI21x1_ASAP7_75t_R _27395_ (.A1(_16008_),
    .A2(_04608_),
    .B(_04610_),
    .Y(_04611_));
 AOI21x1_ASAP7_75t_R _27396_ (.A1(_04607_),
    .A2(_04611_),
    .B(_04376_),
    .Y(_04612_));
 AO21x1_ASAP7_75t_R _27397_ (.A1(_04422_),
    .A2(_04367_),
    .B(_04362_),
    .Y(_04613_));
 OA21x2_ASAP7_75t_R _27398_ (.A1(_04347_),
    .A2(net599),
    .B(_04521_),
    .Y(_04614_));
 OAI21x1_ASAP7_75t_R _27399_ (.A1(_04413_),
    .A2(_04614_),
    .B(_04410_),
    .Y(_04615_));
 AOI21x1_ASAP7_75t_R _27400_ (.A1(_04613_),
    .A2(_04615_),
    .B(_04409_),
    .Y(_04616_));
 OAI21x1_ASAP7_75t_R _27401_ (.A1(_04612_),
    .A2(_04616_),
    .B(_04482_),
    .Y(_04617_));
 NAND2x1_ASAP7_75t_R _27402_ (.A(_04410_),
    .B(_04552_),
    .Y(_04618_));
 NAND2x1_ASAP7_75t_R _27403_ (.A(_04510_),
    .B(_04472_),
    .Y(_04619_));
 AOI21x1_ASAP7_75t_R _27404_ (.A1(_04618_),
    .A2(_04619_),
    .B(_04409_),
    .Y(_04620_));
 NAND2x1_ASAP7_75t_R _27405_ (.A(_04490_),
    .B(_04427_),
    .Y(_04621_));
 AO21x2_ASAP7_75t_R _27406_ (.A1(_04384_),
    .A2(_04385_),
    .B(_04421_),
    .Y(_04622_));
 AOI21x1_ASAP7_75t_R _27407_ (.A1(_16000_),
    .A2(_04583_),
    .B(_04383_),
    .Y(_04623_));
 NAND2x1_ASAP7_75t_R _27408_ (.A(_04622_),
    .B(_04623_),
    .Y(_04624_));
 AOI21x1_ASAP7_75t_R _27409_ (.A1(_04621_),
    .A2(_04624_),
    .B(_04516_),
    .Y(_04625_));
 OAI21x1_ASAP7_75t_R _27410_ (.A1(_04620_),
    .A2(_04625_),
    .B(_04518_),
    .Y(_04626_));
 AOI21x1_ASAP7_75t_R _27411_ (.A1(_04617_),
    .A2(_04626_),
    .B(_04484_),
    .Y(_04627_));
 AO21x2_ASAP7_75t_R _27412_ (.A1(_04583_),
    .A2(_01242_),
    .B(_04455_),
    .Y(_04628_));
 BUFx6f_ASAP7_75t_R _27413_ (.A(_04414_),
    .Y(_04629_));
 OAI21x1_ASAP7_75t_R _27414_ (.A1(net599),
    .A2(_04347_),
    .B(_04450_),
    .Y(_04630_));
 OAI22x1_ASAP7_75t_R _27415_ (.A1(_04628_),
    .A2(_04606_),
    .B1(_04629_),
    .B2(_04630_),
    .Y(_04631_));
 AOI21x1_ASAP7_75t_R _27416_ (.A1(_16005_),
    .A2(_04608_),
    .B(_04391_),
    .Y(_04632_));
 AOI21x1_ASAP7_75t_R _27417_ (.A1(_04632_),
    .A2(_04587_),
    .B(_04481_),
    .Y(_04633_));
 OAI21x1_ASAP7_75t_R _27418_ (.A1(_04581_),
    .A2(_04631_),
    .B(_04633_),
    .Y(_04634_));
 OAI21x1_ASAP7_75t_R _27419_ (.A1(net8),
    .A2(_04461_),
    .B(_04507_),
    .Y(_04635_));
 OAI21x1_ASAP7_75t_R _27420_ (.A1(_04596_),
    .A2(_04594_),
    .B(_04547_),
    .Y(_04636_));
 AOI21x1_ASAP7_75t_R _27421_ (.A1(_04635_),
    .A2(_04636_),
    .B(_04516_),
    .Y(_04637_));
 NAND2x1_ASAP7_75t_R _27422_ (.A(_16000_),
    .B(net36),
    .Y(_04638_));
 NAND2x1_ASAP7_75t_R _27423_ (.A(_04638_),
    .B(_04427_),
    .Y(_04639_));
 OAI21x1_ASAP7_75t_R _27424_ (.A1(net740),
    .A2(_04514_),
    .B(_04547_),
    .Y(_04640_));
 AOI21x1_ASAP7_75t_R _27425_ (.A1(_04639_),
    .A2(_04640_),
    .B(_04409_),
    .Y(_04641_));
 OAI21x1_ASAP7_75t_R _27426_ (.A1(_04637_),
    .A2(_04641_),
    .B(_04482_),
    .Y(_04642_));
 AOI21x1_ASAP7_75t_R _27427_ (.A1(_04634_),
    .A2(_04642_),
    .B(_04560_),
    .Y(_04643_));
 INVx8_ASAP7_75t_R _27428_ (.A(_04446_),
    .Y(_04644_));
 OAI21x1_ASAP7_75t_R _27429_ (.A1(_04627_),
    .A2(_04643_),
    .B(_04644_),
    .Y(_04645_));
 NAND2x1_ASAP7_75t_R _27430_ (.A(_04605_),
    .B(_04645_),
    .Y(_00121_));
 AO21x2_ASAP7_75t_R _27431_ (.A1(_04412_),
    .A2(_04411_),
    .B(_01242_),
    .Y(_04646_));
 BUFx6f_ASAP7_75t_R _27432_ (.A(_04383_),
    .Y(_04647_));
 AOI21x1_ASAP7_75t_R _27433_ (.A1(_04458_),
    .A2(_04646_),
    .B(_04647_),
    .Y(_04648_));
 BUFx6f_ASAP7_75t_R _27434_ (.A(_04455_),
    .Y(_04649_));
 AOI21x1_ASAP7_75t_R _27435_ (.A1(_04422_),
    .A2(_04474_),
    .B(_04649_),
    .Y(_04650_));
 BUFx10_ASAP7_75t_R _27436_ (.A(_04390_),
    .Y(_04651_));
 OAI21x1_ASAP7_75t_R _27437_ (.A1(_04648_),
    .A2(_04650_),
    .B(_04651_),
    .Y(_04652_));
 AO21x1_ASAP7_75t_R _27438_ (.A1(_04583_),
    .A2(_04420_),
    .B(_04455_),
    .Y(_04653_));
 OAI21x1_ASAP7_75t_R _27439_ (.A1(net811),
    .A2(_04461_),
    .B(_04419_),
    .Y(_04654_));
 OAI21x1_ASAP7_75t_R _27440_ (.A1(_04606_),
    .A2(_04653_),
    .B(_04654_),
    .Y(_04655_));
 NAND2x1_ASAP7_75t_R _27441_ (.A(_04555_),
    .B(_04655_),
    .Y(_04656_));
 AOI21x1_ASAP7_75t_R _27442_ (.A1(_04652_),
    .A2(_04656_),
    .B(_04518_),
    .Y(_04657_));
 INVx2_ASAP7_75t_R _27443_ (.A(_04493_),
    .Y(_04658_));
 AOI21x1_ASAP7_75t_R _27444_ (.A1(net37),
    .A2(_04658_),
    .B(_04649_),
    .Y(_04659_));
 AO21x1_ASAP7_75t_R _27445_ (.A1(_04412_),
    .A2(_04411_),
    .B(_01241_),
    .Y(_04660_));
 AOI21x1_ASAP7_75t_R _27446_ (.A1(_04660_),
    .A2(_04474_),
    .B(_04647_),
    .Y(_04661_));
 OAI21x1_ASAP7_75t_R _27447_ (.A1(_04659_),
    .A2(_04661_),
    .B(_04555_),
    .Y(_04662_));
 AO21x1_ASAP7_75t_R _27448_ (.A1(net36),
    .A2(_16008_),
    .B(_04462_),
    .Y(_04663_));
 AOI21x1_ASAP7_75t_R _27449_ (.A1(_04646_),
    .A2(_04511_),
    .B(_04376_),
    .Y(_04664_));
 OAI21x1_ASAP7_75t_R _27450_ (.A1(net810),
    .A2(_04663_),
    .B(_04664_),
    .Y(_04665_));
 AOI21x1_ASAP7_75t_R _27451_ (.A1(_04662_),
    .A2(_04665_),
    .B(_04557_),
    .Y(_04666_));
 NOR3x2_ASAP7_75t_R _27452_ (.B(_04560_),
    .C(_04666_),
    .Y(_04667_),
    .A(_04657_));
 INVx1_ASAP7_75t_R _27453_ (.A(_04430_),
    .Y(_04668_));
 NOR2x1_ASAP7_75t_R _27454_ (.A(_04668_),
    .B(_04514_),
    .Y(_04669_));
 AOI21x1_ASAP7_75t_R _27455_ (.A1(_04563_),
    .A2(_04490_),
    .B(_04410_),
    .Y(_04670_));
 AOI21x1_ASAP7_75t_R _27456_ (.A1(_04629_),
    .A2(_04669_),
    .B(_04670_),
    .Y(_04671_));
 INVx1_ASAP7_75t_R _27457_ (.A(_04586_),
    .Y(_04672_));
 NOR2x1_ASAP7_75t_R _27458_ (.A(_04526_),
    .B(_04542_),
    .Y(_04673_));
 OAI21x1_ASAP7_75t_R _27459_ (.A1(_04582_),
    .A2(_04672_),
    .B(_04673_),
    .Y(_04674_));
 OAI21x1_ASAP7_75t_R _27460_ (.A1(_04534_),
    .A2(_04671_),
    .B(_04674_),
    .Y(_04675_));
 NAND2x1_ASAP7_75t_R _27461_ (.A(_15997_),
    .B(_04454_),
    .Y(_04676_));
 NAND2x1_ASAP7_75t_R _27462_ (.A(_04676_),
    .B(_04571_),
    .Y(_04677_));
 NOR2x2_ASAP7_75t_R _27463_ (.A(_01242_),
    .B(_04454_),
    .Y(_04678_));
 NOR2x1_ASAP7_75t_R _27464_ (.A(_04420_),
    .B(_04583_),
    .Y(_04679_));
 OAI21x1_ASAP7_75t_R _27465_ (.A1(_04678_),
    .A2(_04679_),
    .B(_04462_),
    .Y(_04680_));
 AOI21x1_ASAP7_75t_R _27466_ (.A1(_04677_),
    .A2(_04680_),
    .B(_04516_),
    .Y(_04681_));
 NAND2x2_ASAP7_75t_R _27467_ (.A(_04472_),
    .B(_04471_),
    .Y(_04682_));
 INVx2_ASAP7_75t_R _27468_ (.A(_04682_),
    .Y(_04683_));
 OAI21x1_ASAP7_75t_R _27469_ (.A1(_04419_),
    .A2(_04423_),
    .B(_04465_),
    .Y(_04684_));
 OAI21x1_ASAP7_75t_R _27470_ (.A1(_04683_),
    .A2(_04684_),
    .B(_04481_),
    .Y(_04685_));
 NOR2x1_ASAP7_75t_R _27471_ (.A(_04681_),
    .B(_04685_),
    .Y(_04686_));
 OAI21x1_ASAP7_75t_R _27472_ (.A1(_04686_),
    .A2(_04675_),
    .B(_04560_),
    .Y(_04687_));
 NAND2x1_ASAP7_75t_R _27473_ (.A(_04447_),
    .B(_04687_),
    .Y(_04688_));
 OA21x2_ASAP7_75t_R _27474_ (.A1(_01246_),
    .A2(_04362_),
    .B(_04390_),
    .Y(_04689_));
 NAND2x1_ASAP7_75t_R _27475_ (.A(_04677_),
    .B(_04689_),
    .Y(_04690_));
 AND2x2_ASAP7_75t_R _27476_ (.A(_04361_),
    .B(_00615_),
    .Y(_04691_));
 NOR2x2_ASAP7_75t_R _27477_ (.A(_04691_),
    .B(_04526_),
    .Y(_04692_));
 AOI21x1_ASAP7_75t_R _27478_ (.A1(_04516_),
    .A2(_04692_),
    .B(_04407_),
    .Y(_04693_));
 NAND2x1_ASAP7_75t_R _27479_ (.A(_04690_),
    .B(_04693_),
    .Y(_04694_));
 NOR2x1_ASAP7_75t_R _27480_ (.A(_04383_),
    .B(_04499_),
    .Y(_04695_));
 INVx1_ASAP7_75t_R _27481_ (.A(_04695_),
    .Y(_04696_));
 AO21x1_ASAP7_75t_R _27482_ (.A1(_04497_),
    .A2(_04422_),
    .B(_04475_),
    .Y(_04697_));
 AOI21x1_ASAP7_75t_R _27483_ (.A1(_04696_),
    .A2(_04697_),
    .B(_04542_),
    .Y(_04698_));
 AOI21x1_ASAP7_75t_R _27484_ (.A1(_04366_),
    .A2(_04630_),
    .B(_04414_),
    .Y(_04699_));
 AND2x2_ASAP7_75t_R _27485_ (.A(_01239_),
    .B(_04420_),
    .Y(_04700_));
 INVx2_ASAP7_75t_R _27486_ (.A(_04700_),
    .Y(_04701_));
 OAI21x1_ASAP7_75t_R _27487_ (.A1(net599),
    .A2(_04347_),
    .B(_04701_),
    .Y(_04702_));
 AOI21x1_ASAP7_75t_R _27488_ (.A1(_04503_),
    .A2(_04702_),
    .B(_04475_),
    .Y(_04703_));
 OAI21x1_ASAP7_75t_R _27489_ (.A1(_04699_),
    .A2(_04703_),
    .B(_04535_),
    .Y(_04704_));
 NAND2x1_ASAP7_75t_R _27490_ (.A(_04559_),
    .B(_04704_),
    .Y(_04705_));
 NOR2x1_ASAP7_75t_R _27491_ (.A(_04698_),
    .B(_04705_),
    .Y(_04706_));
 AOI21x1_ASAP7_75t_R _27492_ (.A1(_04694_),
    .A2(_04706_),
    .B(_04447_),
    .Y(_04707_));
 AOI21x1_ASAP7_75t_R _27493_ (.A1(_15997_),
    .A2(_04454_),
    .B(_04455_),
    .Y(_04708_));
 NOR2x1_ASAP7_75t_R _27494_ (.A(_04573_),
    .B(_04414_),
    .Y(_04709_));
 AOI21x1_ASAP7_75t_R _27495_ (.A1(_04510_),
    .A2(_04708_),
    .B(_04709_),
    .Y(_04710_));
 AOI21x1_ASAP7_75t_R _27496_ (.A1(_04516_),
    .A2(_04710_),
    .B(_04407_),
    .Y(_04711_));
 AND2x2_ASAP7_75t_R _27497_ (.A(_04472_),
    .B(_04468_),
    .Y(_04712_));
 AO21x1_ASAP7_75t_R _27498_ (.A1(_04583_),
    .A2(_04488_),
    .B(_04418_),
    .Y(_04713_));
 NOR2x1_ASAP7_75t_R _27499_ (.A(_04506_),
    .B(_04713_),
    .Y(_04714_));
 OAI21x1_ASAP7_75t_R _27500_ (.A1(_04712_),
    .A2(_04714_),
    .B(_04409_),
    .Y(_04715_));
 NAND2x1_ASAP7_75t_R _27501_ (.A(_04711_),
    .B(_04715_),
    .Y(_04716_));
 AOI21x1_ASAP7_75t_R _27502_ (.A1(net48),
    .A2(_04454_),
    .B(_04455_),
    .Y(_04717_));
 NAND2x2_ASAP7_75t_R _27503_ (.A(_04491_),
    .B(_04717_),
    .Y(_04718_));
 AOI21x1_ASAP7_75t_R _27504_ (.A1(_04682_),
    .A2(_04718_),
    .B(_04534_),
    .Y(_04719_));
 OR2x2_ASAP7_75t_R _27505_ (.A(_01244_),
    .B(_04383_),
    .Y(_04720_));
 OAI21x1_ASAP7_75t_R _27506_ (.A1(net458),
    .A2(_04378_),
    .B(_04410_),
    .Y(_04721_));
 AOI21x1_ASAP7_75t_R _27507_ (.A1(_04720_),
    .A2(_04721_),
    .B(_04542_),
    .Y(_04722_));
 NOR3x1_ASAP7_75t_R _27508_ (.A(_04719_),
    .B(_04722_),
    .C(_04559_),
    .Y(_04723_));
 NAND2x1_ASAP7_75t_R _27509_ (.A(_04716_),
    .B(_04723_),
    .Y(_04724_));
 NAND2x1_ASAP7_75t_R _27510_ (.A(_04707_),
    .B(_04724_),
    .Y(_04725_));
 OAI21x1_ASAP7_75t_R _27511_ (.A1(_04667_),
    .A2(_04688_),
    .B(_04725_),
    .Y(_00122_));
 AND3x1_ASAP7_75t_R _27512_ (.A(_04489_),
    .B(_04406_),
    .C(_04419_),
    .Y(_04726_));
 OAI21x1_ASAP7_75t_R _27513_ (.A1(_04658_),
    .A2(_04574_),
    .B(_04365_),
    .Y(_04727_));
 NOR2x1_ASAP7_75t_R _27514_ (.A(_04726_),
    .B(_04727_),
    .Y(_04728_));
 INVx1_ASAP7_75t_R _27515_ (.A(_00607_),
    .Y(_04729_));
 AO21x1_ASAP7_75t_R _27516_ (.A1(_16008_),
    .A2(_04729_),
    .B(_04414_),
    .Y(_04730_));
 OR3x1_ASAP7_75t_R _27517_ (.A(_04730_),
    .B(_04407_),
    .C(_04553_),
    .Y(_04731_));
 AOI21x1_ASAP7_75t_R _27518_ (.A1(_04728_),
    .A2(_04731_),
    .B(_04581_),
    .Y(_04732_));
 NOR2x2_ASAP7_75t_R _27519_ (.A(_04701_),
    .B(_04583_),
    .Y(_04733_));
 NAND2x2_ASAP7_75t_R _27520_ (.A(_04536_),
    .B(_04490_),
    .Y(_04734_));
 OA21x2_ASAP7_75t_R _27521_ (.A1(_04628_),
    .A2(_04733_),
    .B(_04734_),
    .Y(_04735_));
 NOR2x2_ASAP7_75t_R _27522_ (.A(_04406_),
    .B(_04390_),
    .Y(_04736_));
 INVx3_ASAP7_75t_R _27523_ (.A(_04736_),
    .Y(_04737_));
 NOR2x2_ASAP7_75t_R _27524_ (.A(_04481_),
    .B(_04390_),
    .Y(_04738_));
 AO21x2_ASAP7_75t_R _27525_ (.A1(_04583_),
    .A2(_01241_),
    .B(_04414_),
    .Y(_04739_));
 NAND2x1_ASAP7_75t_R _27526_ (.A(_04410_),
    .B(_04457_),
    .Y(_04740_));
 OAI21x1_ASAP7_75t_R _27527_ (.A1(_04567_),
    .A2(_04739_),
    .B(_04740_),
    .Y(_04741_));
 AOI21x1_ASAP7_75t_R _27528_ (.A1(_04738_),
    .A2(_04741_),
    .B(_04484_),
    .Y(_04742_));
 OAI21x1_ASAP7_75t_R _27529_ (.A1(_04735_),
    .A2(_04737_),
    .B(_04742_),
    .Y(_04743_));
 NOR2x1_ASAP7_75t_R _27530_ (.A(_04732_),
    .B(_04743_),
    .Y(_04744_));
 NAND2x1_ASAP7_75t_R _27531_ (.A(_04646_),
    .B(_04511_),
    .Y(_04745_));
 OAI21x1_ASAP7_75t_R _27532_ (.A1(_04581_),
    .A2(_04745_),
    .B(_04482_),
    .Y(_04746_));
 OAI21x1_ASAP7_75t_R _27533_ (.A1(_04379_),
    .A2(_16005_),
    .B(_04381_),
    .Y(_04747_));
 NOR2x1_ASAP7_75t_R _27534_ (.A(_04733_),
    .B(_04747_),
    .Y(_04748_));
 NOR2x1_ASAP7_75t_R _27535_ (.A(_04748_),
    .B(_04578_),
    .Y(_04749_));
 OAI21x1_ASAP7_75t_R _27536_ (.A1(_04746_),
    .A2(_04749_),
    .B(_04484_),
    .Y(_04750_));
 AOI21x1_ASAP7_75t_R _27537_ (.A1(net37),
    .A2(_04646_),
    .B(_04629_),
    .Y(_04751_));
 NAND2x1_ASAP7_75t_R _27538_ (.A(net48),
    .B(_16008_),
    .Y(_04752_));
 AOI21x1_ASAP7_75t_R _27539_ (.A1(_04458_),
    .A2(_04752_),
    .B(_04649_),
    .Y(_04753_));
 OAI21x1_ASAP7_75t_R _27540_ (.A1(_04751_),
    .A2(_04753_),
    .B(_04651_),
    .Y(_04754_));
 NOR2x1_ASAP7_75t_R _27541_ (.A(_04428_),
    .B(_04449_),
    .Y(_04755_));
 INVx1_ASAP7_75t_R _27542_ (.A(_04619_),
    .Y(_04756_));
 OAI21x1_ASAP7_75t_R _27543_ (.A1(_04755_),
    .A2(_04756_),
    .B(_04581_),
    .Y(_04757_));
 AOI21x1_ASAP7_75t_R _27544_ (.A1(_04754_),
    .A2(_04757_),
    .B(_04557_),
    .Y(_04758_));
 OAI21x1_ASAP7_75t_R _27545_ (.A1(_04750_),
    .A2(_04758_),
    .B(_04447_),
    .Y(_04759_));
 NAND2x2_ASAP7_75t_R _27546_ (.A(_16000_),
    .B(_04583_),
    .Y(_04760_));
 AOI21x1_ASAP7_75t_R _27547_ (.A1(_04760_),
    .A2(_04510_),
    .B(_04647_),
    .Y(_04761_));
 OAI21x1_ASAP7_75t_R _27548_ (.A1(_04571_),
    .A2(_04761_),
    .B(_04581_),
    .Y(_04762_));
 NOR2x1_ASAP7_75t_R _27549_ (.A(_04606_),
    .B(_04628_),
    .Y(_04763_));
 INVx1_ASAP7_75t_R _27550_ (.A(_04496_),
    .Y(_04764_));
 NOR2x1_ASAP7_75t_R _27551_ (.A(_04764_),
    .B(_04739_),
    .Y(_04765_));
 OAI21x1_ASAP7_75t_R _27552_ (.A1(_04763_),
    .A2(_04765_),
    .B(_04651_),
    .Y(_04766_));
 AOI21x1_ASAP7_75t_R _27553_ (.A1(_04762_),
    .A2(_04766_),
    .B(_04518_),
    .Y(_04767_));
 INVx3_ASAP7_75t_R _27554_ (.A(_04577_),
    .Y(_04768_));
 NAND2x1_ASAP7_75t_R _27555_ (.A(_04658_),
    .B(_04768_),
    .Y(_04769_));
 OAI21x1_ASAP7_75t_R _27556_ (.A1(_04506_),
    .A2(_04552_),
    .B(_04647_),
    .Y(_04770_));
 AO21x1_ASAP7_75t_R _27557_ (.A1(_04769_),
    .A2(_04770_),
    .B(_04542_),
    .Y(_04771_));
 NOR2x1_ASAP7_75t_R _27558_ (.A(_04381_),
    .B(_04489_),
    .Y(_04772_));
 AOI21x1_ASAP7_75t_R _27559_ (.A1(_04366_),
    .A2(_04772_),
    .B(_04481_),
    .Y(_04773_));
 AOI22x1_ASAP7_75t_R _27560_ (.A1(_04426_),
    .A2(_04425_),
    .B1(_04301_),
    .B2(_04307_),
    .Y(_04774_));
 NOR2x1_ASAP7_75t_R _27561_ (.A(_04774_),
    .B(_04594_),
    .Y(_04775_));
 AOI21x1_ASAP7_75t_R _27562_ (.A1(_04629_),
    .A2(_04775_),
    .B(_04516_),
    .Y(_04776_));
 AOI21x1_ASAP7_75t_R _27563_ (.A1(_04773_),
    .A2(_04776_),
    .B(_04559_),
    .Y(_04777_));
 NAND2x1_ASAP7_75t_R _27564_ (.A(_04771_),
    .B(_04777_),
    .Y(_04778_));
 NOR2x1_ASAP7_75t_R _27565_ (.A(_04767_),
    .B(_04778_),
    .Y(_04779_));
 NOR2x1_ASAP7_75t_R _27566_ (.A(_04651_),
    .B(_04761_),
    .Y(_04780_));
 AO21x1_ASAP7_75t_R _27567_ (.A1(_04563_),
    .A2(net37),
    .B(_04487_),
    .Y(_04781_));
 AOI21x1_ASAP7_75t_R _27568_ (.A1(_04474_),
    .A2(_04563_),
    .B(_04629_),
    .Y(_04782_));
 OAI21x1_ASAP7_75t_R _27569_ (.A1(_04494_),
    .A2(_04782_),
    .B(_04482_),
    .Y(_04783_));
 AOI21x1_ASAP7_75t_R _27570_ (.A1(_04780_),
    .A2(_04781_),
    .B(_04783_),
    .Y(_04784_));
 NOR2x1_ASAP7_75t_R _27571_ (.A(_04582_),
    .B(_04653_),
    .Y(_04785_));
 OAI21x1_ASAP7_75t_R _27572_ (.A1(_04670_),
    .A2(_04785_),
    .B(_04738_),
    .Y(_04786_));
 INVx1_ASAP7_75t_R _27573_ (.A(_04506_),
    .Y(_04787_));
 AOI21x1_ASAP7_75t_R _27574_ (.A1(_04787_),
    .A2(_04623_),
    .B(_04534_),
    .Y(_04788_));
 OR3x1_ASAP7_75t_R _27575_ (.A(_04596_),
    .B(net740),
    .C(_04462_),
    .Y(_04789_));
 AOI21x1_ASAP7_75t_R _27576_ (.A1(_04788_),
    .A2(_04789_),
    .B(_04439_),
    .Y(_04790_));
 NAND2x1_ASAP7_75t_R _27577_ (.A(_04790_),
    .B(_04786_),
    .Y(_04791_));
 OAI21x1_ASAP7_75t_R _27578_ (.A1(_04784_),
    .A2(_04791_),
    .B(_04644_),
    .Y(_04792_));
 OAI22x1_ASAP7_75t_R _27579_ (.A1(_04744_),
    .A2(_04759_),
    .B1(_04779_),
    .B2(_04792_),
    .Y(_00123_));
 NAND2x2_ASAP7_75t_R _27580_ (.A(_04352_),
    .B(_15995_),
    .Y(_04793_));
 NAND2x1_ASAP7_75t_R _27581_ (.A(_15997_),
    .B(_16000_),
    .Y(_04794_));
 AO21x1_ASAP7_75t_R _27582_ (.A1(_04793_),
    .A2(_04794_),
    .B(_04410_),
    .Y(_04795_));
 NAND2x1_ASAP7_75t_R _27583_ (.A(_04468_),
    .B(_04708_),
    .Y(_04796_));
 AO21x1_ASAP7_75t_R _27584_ (.A1(_04795_),
    .A2(_04796_),
    .B(_04581_),
    .Y(_04797_));
 OAI21x1_ASAP7_75t_R _27585_ (.A1(_16008_),
    .A2(net36),
    .B(_04410_),
    .Y(_04798_));
 OAI21x1_ASAP7_75t_R _27586_ (.A1(_04513_),
    .A2(_04798_),
    .B(_04376_),
    .Y(_04799_));
 AND2x2_ASAP7_75t_R _27587_ (.A(_04511_),
    .B(_04563_),
    .Y(_04800_));
 OA21x2_ASAP7_75t_R _27588_ (.A1(_04799_),
    .A2(_04800_),
    .B(_04482_),
    .Y(_04801_));
 AO21x1_ASAP7_75t_R _27589_ (.A1(_04747_),
    .A2(_04386_),
    .B(_04555_),
    .Y(_04802_));
 AOI21x1_ASAP7_75t_R _27590_ (.A1(_04468_),
    .A2(_04474_),
    .B(_04629_),
    .Y(_04803_));
 AOI21x1_ASAP7_75t_R _27591_ (.A1(_04474_),
    .A2(_04491_),
    .B(_04487_),
    .Y(_04804_));
 OAI21x1_ASAP7_75t_R _27592_ (.A1(_04803_),
    .A2(_04804_),
    .B(_04581_),
    .Y(_04805_));
 AOI21x1_ASAP7_75t_R _27593_ (.A1(_04802_),
    .A2(_04805_),
    .B(_04557_),
    .Y(_04806_));
 AOI211x1_ASAP7_75t_R _27594_ (.A1(_04797_),
    .A2(_04801_),
    .B(_04806_),
    .C(_04560_),
    .Y(_04807_));
 AO21x1_ASAP7_75t_R _27595_ (.A1(_04563_),
    .A2(_04499_),
    .B(_04462_),
    .Y(_04808_));
 AO21x1_ASAP7_75t_R _27596_ (.A1(_04808_),
    .A2(_04424_),
    .B(_04407_),
    .Y(_04809_));
 AOI21x1_ASAP7_75t_R _27597_ (.A1(_04525_),
    .A2(_04454_),
    .B(_04455_),
    .Y(_04810_));
 NAND2x1_ASAP7_75t_R _27598_ (.A(_04491_),
    .B(_04810_),
    .Y(_04811_));
 AND3x1_ASAP7_75t_R _27599_ (.A(_04680_),
    .B(_04651_),
    .C(_04811_),
    .Y(_04812_));
 OAI21x1_ASAP7_75t_R _27600_ (.A1(_04413_),
    .A2(net811),
    .B(_04647_),
    .Y(_04813_));
 AOI21x1_ASAP7_75t_R _27601_ (.A1(_04813_),
    .A2(_04654_),
    .B(_04555_),
    .Y(_04814_));
 OAI21x1_ASAP7_75t_R _27602_ (.A1(net458),
    .A2(_04614_),
    .B(_04649_),
    .Y(_04815_));
 AOI21x1_ASAP7_75t_R _27603_ (.A1(_04815_),
    .A2(_04382_),
    .B(_04651_),
    .Y(_04816_));
 OAI21x1_ASAP7_75t_R _27604_ (.A1(_04814_),
    .A2(_04816_),
    .B(_04518_),
    .Y(_04817_));
 OAI21x1_ASAP7_75t_R _27605_ (.A1(_04809_),
    .A2(_04812_),
    .B(_04817_),
    .Y(_04818_));
 OAI21x1_ASAP7_75t_R _27606_ (.A1(_04484_),
    .A2(_04818_),
    .B(_04644_),
    .Y(_04819_));
 OA21x2_ASAP7_75t_R _27607_ (.A1(_16005_),
    .A2(_04419_),
    .B(_04465_),
    .Y(_04820_));
 NAND2x1_ASAP7_75t_R _27608_ (.A(_04522_),
    .B(_04511_),
    .Y(_04821_));
 AO21x1_ASAP7_75t_R _27609_ (.A1(_04820_),
    .A2(_04821_),
    .B(_04559_),
    .Y(_04822_));
 AND3x1_ASAP7_75t_R _27610_ (.A(_04429_),
    .B(_04547_),
    .C(_04563_),
    .Y(_04823_));
 NOR2x1_ASAP7_75t_R _27611_ (.A(_04565_),
    .B(_04823_),
    .Y(_04824_));
 OAI21x1_ASAP7_75t_R _27612_ (.A1(_04822_),
    .A2(_04824_),
    .B(_04557_),
    .Y(_04825_));
 AO21x1_ASAP7_75t_R _27613_ (.A1(_04469_),
    .A2(_04515_),
    .B(_04651_),
    .Y(_04826_));
 AOI21x1_ASAP7_75t_R _27614_ (.A1(_01241_),
    .A2(_04349_),
    .B(_04418_),
    .Y(_04827_));
 NAND2x1_ASAP7_75t_R _27615_ (.A(_04474_),
    .B(_04827_),
    .Y(_04828_));
 AO21x1_ASAP7_75t_R _27616_ (.A1(_04795_),
    .A2(_04828_),
    .B(_04581_),
    .Y(_04829_));
 AOI21x1_ASAP7_75t_R _27617_ (.A1(_04826_),
    .A2(_04829_),
    .B(_04484_),
    .Y(_04830_));
 AND3x1_ASAP7_75t_R _27618_ (.A(_04622_),
    .B(_04471_),
    .C(_04649_),
    .Y(_04831_));
 AO21x1_ASAP7_75t_R _27619_ (.A1(_04412_),
    .A2(_04411_),
    .B(_04363_),
    .Y(_04832_));
 AOI21x1_ASAP7_75t_R _27620_ (.A1(_04649_),
    .A2(_04832_),
    .B(_04376_),
    .Y(_04833_));
 AOI21x1_ASAP7_75t_R _27621_ (.A1(_04672_),
    .A2(_04833_),
    .B(_04559_),
    .Y(_04834_));
 OAI21x1_ASAP7_75t_R _27622_ (.A1(_04453_),
    .A2(_04831_),
    .B(_04834_),
    .Y(_04835_));
 NAND2x2_ASAP7_75t_R _27623_ (.A(_04793_),
    .B(_04827_),
    .Y(_04836_));
 OA21x2_ASAP7_75t_R _27624_ (.A1(_04381_),
    .A2(_04367_),
    .B(_04391_),
    .Y(_04837_));
 NAND2x1_ASAP7_75t_R _27625_ (.A(_04836_),
    .B(_04837_),
    .Y(_04838_));
 AOI21x1_ASAP7_75t_R _27626_ (.A1(_04450_),
    .A2(_04649_),
    .B(_04391_),
    .Y(_04839_));
 AOI21x1_ASAP7_75t_R _27627_ (.A1(_04713_),
    .A2(_04839_),
    .B(_04439_),
    .Y(_04840_));
 AOI21x1_ASAP7_75t_R _27628_ (.A1(_04838_),
    .A2(_04840_),
    .B(_04557_),
    .Y(_04841_));
 AOI21x1_ASAP7_75t_R _27629_ (.A1(_04835_),
    .A2(_04841_),
    .B(_04644_),
    .Y(_04842_));
 OAI21x1_ASAP7_75t_R _27630_ (.A1(_04825_),
    .A2(_04830_),
    .B(_04842_),
    .Y(_04843_));
 OAI21x1_ASAP7_75t_R _27631_ (.A1(_04807_),
    .A2(_04819_),
    .B(_04843_),
    .Y(_00124_));
 AOI21x1_ASAP7_75t_R _27632_ (.A1(_04468_),
    .A2(_04490_),
    .B(_04649_),
    .Y(_04844_));
 AOI211x1_ASAP7_75t_R _27633_ (.A1(_04487_),
    .A2(_04678_),
    .B(_04844_),
    .C(_04737_),
    .Y(_04845_));
 NOR2x1_ASAP7_75t_R _27634_ (.A(_04553_),
    .B(_04584_),
    .Y(_04846_));
 OAI21x1_ASAP7_75t_R _27635_ (.A1(_04533_),
    .A2(_04529_),
    .B(_04480_),
    .Y(_04847_));
 AO21x1_ASAP7_75t_R _27636_ (.A1(_04647_),
    .A2(_04413_),
    .B(_04847_),
    .Y(_04848_));
 OAI21x1_ASAP7_75t_R _27637_ (.A1(_04846_),
    .A2(_04848_),
    .B(_04644_),
    .Y(_04849_));
 NOR2x1_ASAP7_75t_R _27638_ (.A(_04845_),
    .B(_04849_),
    .Y(_04850_));
 NAND2x1_ASAP7_75t_R _27639_ (.A(_04794_),
    .B(_04536_),
    .Y(_04851_));
 OA21x2_ASAP7_75t_R _27640_ (.A1(_16008_),
    .A2(_04585_),
    .B(_04362_),
    .Y(_04852_));
 AOI21x1_ASAP7_75t_R _27641_ (.A1(_04366_),
    .A2(_04852_),
    .B(_04516_),
    .Y(_04853_));
 NAND2x1_ASAP7_75t_R _27642_ (.A(_04851_),
    .B(_04853_),
    .Y(_04854_));
 OA21x2_ASAP7_75t_R _27643_ (.A1(_15997_),
    .A2(_04547_),
    .B(_04376_),
    .Y(_04855_));
 AOI21x1_ASAP7_75t_R _27644_ (.A1(_04855_),
    .A2(_04795_),
    .B(_04482_),
    .Y(_04856_));
 NAND2x1_ASAP7_75t_R _27645_ (.A(_04854_),
    .B(_04856_),
    .Y(_04857_));
 AOI21x1_ASAP7_75t_R _27646_ (.A1(_04850_),
    .A2(_04857_),
    .B(_04484_),
    .Y(_04858_));
 OAI21x1_ASAP7_75t_R _27647_ (.A1(_04649_),
    .A2(_04733_),
    .B(_04376_),
    .Y(_04859_));
 AOI21x1_ASAP7_75t_R _27648_ (.A1(_04538_),
    .A2(_04768_),
    .B(_04859_),
    .Y(_04860_));
 INVx1_ASAP7_75t_R _27649_ (.A(_04628_),
    .Y(_04861_));
 AOI211x1_ASAP7_75t_R _27650_ (.A1(_16008_),
    .A2(_04608_),
    .B(_04861_),
    .C(_04555_),
    .Y(_04862_));
 OAI21x1_ASAP7_75t_R _27651_ (.A1(_04860_),
    .A2(_04862_),
    .B(_04518_),
    .Y(_04863_));
 AO21x1_ASAP7_75t_R _27652_ (.A1(net37),
    .A2(_04366_),
    .B(_04487_),
    .Y(_04864_));
 AND3x1_ASAP7_75t_R _27653_ (.A(_04522_),
    .B(_04462_),
    .C(net37),
    .Y(_04865_));
 NOR2x1_ASAP7_75t_R _27654_ (.A(_04847_),
    .B(_04865_),
    .Y(_04866_));
 OAI21x1_ASAP7_75t_R _27655_ (.A1(_04729_),
    .A2(_04487_),
    .B(_04736_),
    .Y(_04867_));
 OAI21x1_ASAP7_75t_R _27656_ (.A1(_04768_),
    .A2(_04867_),
    .B(_04447_),
    .Y(_04868_));
 AOI21x1_ASAP7_75t_R _27657_ (.A1(_04864_),
    .A2(_04866_),
    .B(_04868_),
    .Y(_04869_));
 NAND2x1_ASAP7_75t_R _27658_ (.A(_04863_),
    .B(_04869_),
    .Y(_04870_));
 AOI21x1_ASAP7_75t_R _27659_ (.A1(_04622_),
    .A2(_04861_),
    .B(_04482_),
    .Y(_04871_));
 OAI21x1_ASAP7_75t_R _27660_ (.A1(_04629_),
    .A2(_04491_),
    .B(_04516_),
    .Y(_04872_));
 NOR2x1_ASAP7_75t_R _27661_ (.A(_04387_),
    .B(_04872_),
    .Y(_04873_));
 AOI21x1_ASAP7_75t_R _27662_ (.A1(_04871_),
    .A2(_04873_),
    .B(_04447_),
    .Y(_04874_));
 AOI211x1_ASAP7_75t_R _27663_ (.A1(_04622_),
    .A2(_04487_),
    .B(_04552_),
    .C(_04555_),
    .Y(_04875_));
 OAI21x1_ASAP7_75t_R _27664_ (.A1(_04507_),
    .A2(net8),
    .B(_04465_),
    .Y(_04876_));
 NOR2x1_ASAP7_75t_R _27665_ (.A(_04876_),
    .B(_04753_),
    .Y(_04877_));
 OAI21x1_ASAP7_75t_R _27666_ (.A1(_04875_),
    .A2(_04877_),
    .B(_04557_),
    .Y(_04878_));
 AO21x1_ASAP7_75t_R _27667_ (.A1(_04660_),
    .A2(_04367_),
    .B(_04629_),
    .Y(_04879_));
 OA21x2_ASAP7_75t_R _27668_ (.A1(_04653_),
    .A2(_04700_),
    .B(_04535_),
    .Y(_04880_));
 NAND2x1_ASAP7_75t_R _27669_ (.A(_04879_),
    .B(_04880_),
    .Y(_04881_));
 NAND3x1_ASAP7_75t_R _27670_ (.A(_04874_),
    .B(_04878_),
    .C(_04881_),
    .Y(_04882_));
 INVx1_ASAP7_75t_R _27671_ (.A(_04512_),
    .Y(_04883_));
 NAND2x1_ASAP7_75t_R _27672_ (.A(_04381_),
    .B(_16000_),
    .Y(_04884_));
 NAND2x1_ASAP7_75t_R _27673_ (.A(_04884_),
    .B(_04738_),
    .Y(_04885_));
 OAI21x1_ASAP7_75t_R _27674_ (.A1(_04883_),
    .A2(_04885_),
    .B(_04446_),
    .Y(_04886_));
 AND2x4_ASAP7_75t_R _27675_ (.A(_04571_),
    .B(_04490_),
    .Y(_04887_));
 OAI21x1_ASAP7_75t_R _27676_ (.A1(_04606_),
    .A2(_04739_),
    .B(_04535_),
    .Y(_04888_));
 NOR2x2_ASAP7_75t_R _27677_ (.A(_04887_),
    .B(_04888_),
    .Y(_04889_));
 NOR2x1_ASAP7_75t_R _27678_ (.A(_04886_),
    .B(_04889_),
    .Y(_04890_));
 INVx1_ASAP7_75t_R _27679_ (.A(_04366_),
    .Y(_04891_));
 AO21x1_ASAP7_75t_R _27680_ (.A1(_04891_),
    .A2(_04647_),
    .B(_04465_),
    .Y(_04892_));
 AOI21x1_ASAP7_75t_R _27681_ (.A1(_04522_),
    .A2(_04768_),
    .B(_04892_),
    .Y(_04893_));
 OA21x2_ASAP7_75t_R _27682_ (.A1(_04514_),
    .A2(_04461_),
    .B(_04547_),
    .Y(_04894_));
 NOR2x1_ASAP7_75t_R _27683_ (.A(_04453_),
    .B(_04894_),
    .Y(_04895_));
 OAI21x1_ASAP7_75t_R _27684_ (.A1(_04893_),
    .A2(_04895_),
    .B(_04557_),
    .Y(_04896_));
 AOI21x1_ASAP7_75t_R _27685_ (.A1(_04896_),
    .A2(_04890_),
    .B(_04560_),
    .Y(_04897_));
 AOI22x1_ASAP7_75t_R _27686_ (.A1(_04858_),
    .A2(_04870_),
    .B1(_04882_),
    .B2(_04897_),
    .Y(_00125_));
 INVx1_ASAP7_75t_R _27687_ (.A(_04610_),
    .Y(_04898_));
 AOI21x1_ASAP7_75t_R _27688_ (.A1(_04898_),
    .A2(_04527_),
    .B(_04516_),
    .Y(_04899_));
 NAND2x1_ASAP7_75t_R _27689_ (.A(_04462_),
    .B(_04764_),
    .Y(_04900_));
 NOR2x1_ASAP7_75t_R _27690_ (.A(_16000_),
    .B(_16005_),
    .Y(_04901_));
 OAI21x1_ASAP7_75t_R _27691_ (.A1(net810),
    .A2(_04901_),
    .B(_04507_),
    .Y(_04902_));
 AOI21x1_ASAP7_75t_R _27692_ (.A1(_04900_),
    .A2(_04902_),
    .B(_04409_),
    .Y(_04903_));
 OAI21x1_ASAP7_75t_R _27693_ (.A1(_04899_),
    .A2(_04903_),
    .B(_04557_),
    .Y(_04904_));
 NAND2x1_ASAP7_75t_R _27694_ (.A(_04550_),
    .B(_04623_),
    .Y(_04905_));
 OAI21x1_ASAP7_75t_R _27695_ (.A1(_04774_),
    .A2(_04514_),
    .B(_04647_),
    .Y(_04906_));
 AOI21x1_ASAP7_75t_R _27696_ (.A1(_04905_),
    .A2(_04906_),
    .B(_04555_),
    .Y(_04907_));
 OAI21x1_ASAP7_75t_R _27697_ (.A1(_04513_),
    .A2(_04594_),
    .B(_04647_),
    .Y(_04908_));
 OAI21x1_ASAP7_75t_R _27698_ (.A1(_04552_),
    .A2(_04606_),
    .B(_04547_),
    .Y(_04909_));
 AOI21x1_ASAP7_75t_R _27699_ (.A1(_04908_),
    .A2(_04909_),
    .B(_04651_),
    .Y(_04910_));
 OAI21x1_ASAP7_75t_R _27700_ (.A1(_04907_),
    .A2(_04910_),
    .B(_04518_),
    .Y(_04911_));
 NAND2x1_ASAP7_75t_R _27701_ (.A(_04904_),
    .B(_04911_),
    .Y(_04912_));
 INVx1_ASAP7_75t_R _27702_ (.A(_04503_),
    .Y(_04913_));
 OAI21x1_ASAP7_75t_R _27703_ (.A1(_04913_),
    .A2(_04364_),
    .B(_04507_),
    .Y(_04914_));
 OAI21x1_ASAP7_75t_R _27704_ (.A1(_04614_),
    .A2(_04380_),
    .B(_04462_),
    .Y(_04915_));
 AOI21x1_ASAP7_75t_R _27705_ (.A1(_04914_),
    .A2(_04915_),
    .B(_04409_),
    .Y(_04916_));
 NAND2x1_ASAP7_75t_R _27706_ (.A(_04471_),
    .B(_04511_),
    .Y(_04917_));
 NOR2x1_ASAP7_75t_R _27707_ (.A(_04700_),
    .B(_16005_),
    .Y(_04918_));
 OAI21x1_ASAP7_75t_R _27708_ (.A1(_04457_),
    .A2(_04918_),
    .B(_04507_),
    .Y(_04919_));
 AOI21x1_ASAP7_75t_R _27709_ (.A1(_04917_),
    .A2(_04919_),
    .B(_04555_),
    .Y(_04920_));
 OAI21x1_ASAP7_75t_R _27710_ (.A1(_04916_),
    .A2(_04920_),
    .B(_04557_),
    .Y(_04921_));
 NAND2x1_ASAP7_75t_R _27711_ (.A(_15997_),
    .B(net48),
    .Y(_04922_));
 NAND2x2_ASAP7_75t_R _27712_ (.A(_04922_),
    .B(_04491_),
    .Y(_04923_));
 AND2x2_ASAP7_75t_R _27713_ (.A(_01243_),
    .B(_01245_),
    .Y(_04924_));
 OA21x2_ASAP7_75t_R _27714_ (.A1(_04381_),
    .A2(_04924_),
    .B(_04465_),
    .Y(_04925_));
 OAI21x1_ASAP7_75t_R _27715_ (.A1(_04487_),
    .A2(_04923_),
    .B(_04925_),
    .Y(_04926_));
 AOI21x1_ASAP7_75t_R _27716_ (.A1(_04507_),
    .A2(_04457_),
    .B(_04465_),
    .Y(_04927_));
 NOR2x1_ASAP7_75t_R _27717_ (.A(_04475_),
    .B(_04430_),
    .Y(_04928_));
 NOR2x1_ASAP7_75t_R _27718_ (.A(_04695_),
    .B(_04928_),
    .Y(_04929_));
 AOI21x1_ASAP7_75t_R _27719_ (.A1(_04927_),
    .A2(_04929_),
    .B(_04481_),
    .Y(_04930_));
 AOI21x1_ASAP7_75t_R _27720_ (.A1(_04926_),
    .A2(_04930_),
    .B(_04447_),
    .Y(_04931_));
 NAND2x1_ASAP7_75t_R _27721_ (.A(_04921_),
    .B(_04931_),
    .Y(_04932_));
 OAI21x1_ASAP7_75t_R _27722_ (.A1(_04644_),
    .A2(_04912_),
    .B(_04932_),
    .Y(_04933_));
 AO21x1_ASAP7_75t_R _27723_ (.A1(_04384_),
    .A2(_04385_),
    .B(_00612_),
    .Y(_04934_));
 NAND2x1_ASAP7_75t_R _27724_ (.A(_04934_),
    .B(_04563_),
    .Y(_04935_));
 OA21x2_ASAP7_75t_R _27725_ (.A1(_04414_),
    .A2(_04366_),
    .B(_04390_),
    .Y(_04936_));
 OAI21x1_ASAP7_75t_R _27726_ (.A1(_04649_),
    .A2(_04935_),
    .B(_04936_),
    .Y(_04937_));
 AOI21x1_ASAP7_75t_R _27727_ (.A1(_04760_),
    .A2(_04810_),
    .B(_04391_),
    .Y(_04938_));
 AO21x1_ASAP7_75t_R _27728_ (.A1(_04702_),
    .A2(_04658_),
    .B(_04362_),
    .Y(_04939_));
 NAND2x1_ASAP7_75t_R _27729_ (.A(_04938_),
    .B(_04939_),
    .Y(_04940_));
 AOI21x1_ASAP7_75t_R _27730_ (.A1(_04937_),
    .A2(_04940_),
    .B(_04407_),
    .Y(_04941_));
 OAI21x1_ASAP7_75t_R _27731_ (.A1(net8),
    .A2(_04668_),
    .B(_04462_),
    .Y(_04942_));
 NAND2x1_ASAP7_75t_R _27732_ (.A(_04793_),
    .B(_04571_),
    .Y(_04943_));
 AOI21x1_ASAP7_75t_R _27733_ (.A1(_04942_),
    .A2(_04943_),
    .B(_04391_),
    .Y(_04944_));
 AO21x1_ASAP7_75t_R _27734_ (.A1(_04475_),
    .A2(_04489_),
    .B(_04375_),
    .Y(_04945_));
 OAI21x1_ASAP7_75t_R _27735_ (.A1(_04692_),
    .A2(_04945_),
    .B(_04407_),
    .Y(_04946_));
 OAI21x1_ASAP7_75t_R _27736_ (.A1(_04944_),
    .A2(_04946_),
    .B(_04644_),
    .Y(_04947_));
 NOR2x1_ASAP7_75t_R _27737_ (.A(_04947_),
    .B(_04941_),
    .Y(_04948_));
 AOI21x1_ASAP7_75t_R _27738_ (.A1(_04730_),
    .A2(_04836_),
    .B(_04376_),
    .Y(_04949_));
 NAND2x1_ASAP7_75t_R _27739_ (.A(_04481_),
    .B(_04684_),
    .Y(_04950_));
 NOR2x1_ASAP7_75t_R _27740_ (.A(_04949_),
    .B(_04950_),
    .Y(_04951_));
 AO21x1_ASAP7_75t_R _27741_ (.A1(_04676_),
    .A2(_04660_),
    .B(_04362_),
    .Y(_04952_));
 AOI21x1_ASAP7_75t_R _27742_ (.A1(_00616_),
    .A2(_04410_),
    .B(_04542_),
    .Y(_04953_));
 NAND2x1_ASAP7_75t_R _27743_ (.A(_04952_),
    .B(_04953_),
    .Y(_04954_));
 OAI21x1_ASAP7_75t_R _27744_ (.A1(net8),
    .A2(_04678_),
    .B(_04507_),
    .Y(_04955_));
 AOI21x1_ASAP7_75t_R _27745_ (.A1(_04462_),
    .A2(_04594_),
    .B(_04534_),
    .Y(_04956_));
 AOI21x1_ASAP7_75t_R _27746_ (.A1(_04955_),
    .A2(_04956_),
    .B(_04644_),
    .Y(_04957_));
 NAND2x1_ASAP7_75t_R _27747_ (.A(_04954_),
    .B(_04957_),
    .Y(_04958_));
 OAI21x1_ASAP7_75t_R _27748_ (.A1(_04951_),
    .A2(_04958_),
    .B(_04560_),
    .Y(_04959_));
 NOR2x1_ASAP7_75t_R _27749_ (.A(_04959_),
    .B(_04948_),
    .Y(_04960_));
 AOI21x1_ASAP7_75t_R _27750_ (.A1(_04484_),
    .A2(_04933_),
    .B(_04960_),
    .Y(_00126_));
 INVx1_ASAP7_75t_R _27751_ (.A(_01245_),
    .Y(_04961_));
 OA21x2_ASAP7_75t_R _27752_ (.A1(_04493_),
    .A2(net811),
    .B(_04547_),
    .Y(_04962_));
 AOI21x1_ASAP7_75t_R _27753_ (.A1(_04961_),
    .A2(_04629_),
    .B(_04962_),
    .Y(_04963_));
 AO21x1_ASAP7_75t_R _27754_ (.A1(_04490_),
    .A2(_04471_),
    .B(_04487_),
    .Y(_04964_));
 AOI21x1_ASAP7_75t_R _27755_ (.A1(_04793_),
    .A2(_04536_),
    .B(_04847_),
    .Y(_04965_));
 AOI22x1_ASAP7_75t_R _27756_ (.A1(_04963_),
    .A2(_04736_),
    .B1(_04964_),
    .B2(_04965_),
    .Y(_04966_));
 AOI211x1_ASAP7_75t_R _27757_ (.A1(_04450_),
    .A2(_04629_),
    .B(_04431_),
    .C(_04651_),
    .Y(_04967_));
 NAND2x1_ASAP7_75t_R _27758_ (.A(_04547_),
    .B(_04546_),
    .Y(_04968_));
 AND3x1_ASAP7_75t_R _27759_ (.A(_04837_),
    .B(_04599_),
    .C(_04968_),
    .Y(_04969_));
 OAI21x1_ASAP7_75t_R _27760_ (.A1(_04967_),
    .A2(_04969_),
    .B(_04518_),
    .Y(_04970_));
 AOI21x1_ASAP7_75t_R _27761_ (.A1(_04966_),
    .A2(_04970_),
    .B(_04484_),
    .Y(_04971_));
 OAI21x1_ASAP7_75t_R _27762_ (.A1(_04450_),
    .A2(_16005_),
    .B(_04475_),
    .Y(_04972_));
 OAI21x1_ASAP7_75t_R _27763_ (.A1(_04428_),
    .A2(_04972_),
    .B(_04555_),
    .Y(_04973_));
 OA21x2_ASAP7_75t_R _27764_ (.A1(_04891_),
    .A2(net8),
    .B(_04647_),
    .Y(_04974_));
 OAI21x1_ASAP7_75t_R _27765_ (.A1(_04733_),
    .A2(_04747_),
    .B(_04651_),
    .Y(_04975_));
 NOR2x1_ASAP7_75t_R _27766_ (.A(_04553_),
    .B(_04972_),
    .Y(_04976_));
 OAI22x1_ASAP7_75t_R _27767_ (.A1(_04973_),
    .A2(_04974_),
    .B1(_04975_),
    .B2(_04976_),
    .Y(_04977_));
 AO21x1_ASAP7_75t_R _27768_ (.A1(_16008_),
    .A2(_15997_),
    .B(_04419_),
    .Y(_04978_));
 AOI21x1_ASAP7_75t_R _27769_ (.A1(_04584_),
    .A2(_04978_),
    .B(_04428_),
    .Y(_04979_));
 NOR2x1_ASAP7_75t_R _27770_ (.A(_04608_),
    .B(_04847_),
    .Y(_04980_));
 OAI21x1_ASAP7_75t_R _27771_ (.A1(_04487_),
    .A2(_04923_),
    .B(_04980_),
    .Y(_04981_));
 OAI21x1_ASAP7_75t_R _27772_ (.A1(_04737_),
    .A2(_04979_),
    .B(_04981_),
    .Y(_04982_));
 AOI21x1_ASAP7_75t_R _27773_ (.A1(_04518_),
    .A2(_04977_),
    .B(_04982_),
    .Y(_04983_));
 OAI21x1_ASAP7_75t_R _27774_ (.A1(_04560_),
    .A2(_04983_),
    .B(_04644_),
    .Y(_04984_));
 NOR2x1_ASAP7_75t_R _27775_ (.A(_04606_),
    .B(_04972_),
    .Y(_04985_));
 NOR2x1_ASAP7_75t_R _27776_ (.A(_04410_),
    .B(_16000_),
    .Y(_04986_));
 AOI21x1_ASAP7_75t_R _27777_ (.A1(_04563_),
    .A2(_04717_),
    .B(_04986_),
    .Y(_04987_));
 OAI22x1_ASAP7_75t_R _27778_ (.A1(_04799_),
    .A2(_04985_),
    .B1(_04581_),
    .B2(_04987_),
    .Y(_04988_));
 OAI21x1_ASAP7_75t_R _27779_ (.A1(_04852_),
    .A2(_04876_),
    .B(_04482_),
    .Y(_04989_));
 INVx1_ASAP7_75t_R _27780_ (.A(_04810_),
    .Y(_04990_));
 OAI21x1_ASAP7_75t_R _27781_ (.A1(_04507_),
    .A2(_04497_),
    .B(_04391_),
    .Y(_04991_));
 AOI21x1_ASAP7_75t_R _27782_ (.A1(_04972_),
    .A2(_04990_),
    .B(_04991_),
    .Y(_04992_));
 OAI21x1_ASAP7_75t_R _27783_ (.A1(_04989_),
    .A2(_04992_),
    .B(_04559_),
    .Y(_04993_));
 AOI21x1_ASAP7_75t_R _27784_ (.A1(_04518_),
    .A2(_04988_),
    .B(_04993_),
    .Y(_04994_));
 AOI21x1_ASAP7_75t_R _27785_ (.A1(_04615_),
    .A2(_04734_),
    .B(_04847_),
    .Y(_04995_));
 AO21x1_ASAP7_75t_R _27786_ (.A1(_16005_),
    .A2(_01242_),
    .B(_04381_),
    .Y(_04996_));
 AOI21x1_ASAP7_75t_R _27787_ (.A1(_04996_),
    .A2(_04836_),
    .B(_04542_),
    .Y(_04997_));
 NOR2x1_ASAP7_75t_R _27788_ (.A(_04997_),
    .B(_04995_),
    .Y(_04998_));
 AO21x1_ASAP7_75t_R _27789_ (.A1(_04503_),
    .A2(_04499_),
    .B(_04419_),
    .Y(_04999_));
 NAND2x1_ASAP7_75t_R _27790_ (.A(_04934_),
    .B(_04536_),
    .Y(_05000_));
 AOI21x1_ASAP7_75t_R _27791_ (.A1(_04999_),
    .A2(_05000_),
    .B(_04534_),
    .Y(_05001_));
 AOI21x1_ASAP7_75t_R _27792_ (.A1(_04915_),
    .A2(_04718_),
    .B(_04737_),
    .Y(_05002_));
 NOR2x1_ASAP7_75t_R _27793_ (.A(_05001_),
    .B(_05002_),
    .Y(_05003_));
 AOI21x1_ASAP7_75t_R _27794_ (.A1(_04998_),
    .A2(_05003_),
    .B(_04560_),
    .Y(_05004_));
 OAI21x1_ASAP7_75t_R _27795_ (.A1(_04994_),
    .A2(_05004_),
    .B(_04447_),
    .Y(_05005_));
 OAI21x1_ASAP7_75t_R _27796_ (.A1(_04971_),
    .A2(_04984_),
    .B(_05005_),
    .Y(_00127_));
 NOR2x2_ASAP7_75t_R _27797_ (.A(_10733_),
    .B(_00617_),
    .Y(_05006_));
 XOR2x1_ASAP7_75t_R _27798_ (.A(net781),
    .Y(_05007_),
    .B(_10628_));
 XOR2x1_ASAP7_75t_R _27799_ (.A(_10677_),
    .Y(_05008_),
    .B(_02211_));
 NAND2x1_ASAP7_75t_R _27800_ (.A(_05007_),
    .B(_05008_),
    .Y(_05009_));
 XNOR2x1_ASAP7_75t_R _27801_ (.B(_10628_),
    .Y(_05010_),
    .A(net781));
 XOR2x1_ASAP7_75t_R _27802_ (.A(_02211_),
    .Y(_05011_),
    .B(_10679_));
 NAND2x1_ASAP7_75t_R _27803_ (.A(_05011_),
    .B(_05010_),
    .Y(_05012_));
 AOI21x1_ASAP7_75t_R _27804_ (.A1(_05009_),
    .A2(_05012_),
    .B(_11374_),
    .Y(_05013_));
 OAI21x1_ASAP7_75t_R _27805_ (.A1(_05006_),
    .A2(_05013_),
    .B(_08023_),
    .Y(_05014_));
 AND2x2_ASAP7_75t_R _27806_ (.A(_11441_),
    .B(_00617_),
    .Y(_05015_));
 NAND2x1_ASAP7_75t_R _27807_ (.A(_05007_),
    .B(_05011_),
    .Y(_05016_));
 NAND2x1_ASAP7_75t_R _27808_ (.A(_05008_),
    .B(_05010_),
    .Y(_05017_));
 AOI21x1_ASAP7_75t_R _27809_ (.A1(_05016_),
    .A2(_05017_),
    .B(_11374_),
    .Y(_05018_));
 INVx1_ASAP7_75t_R _27810_ (.A(_08023_),
    .Y(_05019_));
 OAI21x1_ASAP7_75t_R _27811_ (.A1(_05015_),
    .A2(_05018_),
    .B(_05019_),
    .Y(_05020_));
 NAND2x2_ASAP7_75t_R _27812_ (.A(_05014_),
    .B(_05020_),
    .Y(_05021_));
 BUFx12_ASAP7_75t_R _27813_ (.A(_05021_),
    .Y(_16016_));
 OR2x2_ASAP7_75t_R _27814_ (.A(_10723_),
    .B(_00618_),
    .Y(_05022_));
 NOR2x1_ASAP7_75t_R _27815_ (.A(_10823_),
    .B(_10663_),
    .Y(_05023_));
 NOR2x1_ASAP7_75t_R _27816_ (.A(net683),
    .B(_10659_),
    .Y(_05024_));
 OAI21x1_ASAP7_75t_R _27817_ (.A1(_05023_),
    .A2(_05024_),
    .B(net601),
    .Y(_05025_));
 INVx1_ASAP7_75t_R _27818_ (.A(_05025_),
    .Y(_05026_));
 NAND2x2_ASAP7_75t_R _27819_ (.A(net683),
    .B(_10659_),
    .Y(_05027_));
 NAND2x2_ASAP7_75t_R _27820_ (.A(_10823_),
    .B(_10663_),
    .Y(_05028_));
 NAND3x2_ASAP7_75t_R _27821_ (.B(_05028_),
    .C(net785),
    .Y(_05029_),
    .A(_05027_));
 INVx1_ASAP7_75t_R _27822_ (.A(_05029_),
    .Y(_05030_));
 OAI21x1_ASAP7_75t_R _27823_ (.A1(_05026_),
    .A2(_05030_),
    .B(_11356_),
    .Y(_05031_));
 AOI21x1_ASAP7_75t_R _27824_ (.A1(_05022_),
    .A2(_05031_),
    .B(net617),
    .Y(_05032_));
 NAND2x1_ASAP7_75t_R _27825_ (.A(_00618_),
    .B(_12160_),
    .Y(_05033_));
 NAND3x2_ASAP7_75t_R _27826_ (.B(_10733_),
    .C(_05025_),
    .Y(_05034_),
    .A(_05029_));
 INVx1_ASAP7_75t_R _27827_ (.A(net617),
    .Y(_05035_));
 AOI21x1_ASAP7_75t_R _27828_ (.A1(_05033_),
    .A2(_05034_),
    .B(_05035_),
    .Y(_05036_));
 NOR2x2_ASAP7_75t_R _27829_ (.A(_05032_),
    .B(_05036_),
    .Y(_05037_));
 BUFx10_ASAP7_75t_R _27830_ (.A(_05037_),
    .Y(_16018_));
 XOR2x1_ASAP7_75t_R _27831_ (.A(net52),
    .Y(_05038_),
    .B(_10681_));
 NAND2x1_ASAP7_75t_R _27832_ (.A(_10632_),
    .B(_05038_),
    .Y(_05039_));
 XNOR2x2_ASAP7_75t_R _27833_ (.A(_10676_),
    .B(_10681_),
    .Y(_05040_));
 NAND2x1_ASAP7_75t_R _27834_ (.A(_10624_),
    .B(_05040_),
    .Y(_05041_));
 AOI21x1_ASAP7_75t_R _27835_ (.A1(_05039_),
    .A2(_05041_),
    .B(_02258_),
    .Y(_05042_));
 XOR2x1_ASAP7_75t_R _27836_ (.A(_10681_),
    .Y(_05043_),
    .B(_10624_));
 NAND2x1_ASAP7_75t_R _27837_ (.A(net52),
    .B(_05043_),
    .Y(_05044_));
 XNOR2x2_ASAP7_75t_R _27838_ (.A(_10681_),
    .B(_00829_),
    .Y(_05045_));
 NAND2x1_ASAP7_75t_R _27839_ (.A(_13569_),
    .B(_05045_),
    .Y(_05046_));
 AOI21x1_ASAP7_75t_R _27840_ (.A1(_05044_),
    .A2(_05046_),
    .B(_02246_),
    .Y(_05047_));
 OAI21x1_ASAP7_75t_R _27841_ (.A1(_05042_),
    .A2(_05047_),
    .B(net680),
    .Y(_05048_));
 NOR2x2_ASAP7_75t_R _27842_ (.A(_10619_),
    .B(_00620_),
    .Y(_05049_));
 INVx3_ASAP7_75t_R _27843_ (.A(_05049_),
    .Y(_05050_));
 NAND3x2_ASAP7_75t_R _27844_ (.B(_08031_),
    .C(_05050_),
    .Y(_05051_),
    .A(_05048_));
 AO21x1_ASAP7_75t_R _27845_ (.A1(_05048_),
    .A2(_05050_),
    .B(_08031_),
    .Y(_05052_));
 BUFx4f_ASAP7_75t_R _27846_ (.A(_05052_),
    .Y(_05053_));
 NAND2x2_ASAP7_75t_R _27847_ (.A(_05051_),
    .B(_05053_),
    .Y(_05054_));
 BUFx6f_ASAP7_75t_R _27848_ (.A(_05054_),
    .Y(_16026_));
 AOI21x1_ASAP7_75t_R _27849_ (.A1(_05022_),
    .A2(_05031_),
    .B(_05035_),
    .Y(_05055_));
 AOI21x1_ASAP7_75t_R _27850_ (.A1(_05033_),
    .A2(_05034_),
    .B(net617),
    .Y(_05056_));
 NOR2x2_ASAP7_75t_R _27851_ (.A(_05055_),
    .B(_05056_),
    .Y(_05057_));
 BUFx6f_ASAP7_75t_R rebuffer312 (.A(_05057_),
    .Y(net765));
 INVx3_ASAP7_75t_R _27853_ (.A(_08031_),
    .Y(_05058_));
 NAND3x2_ASAP7_75t_R _27854_ (.B(_05058_),
    .C(_05050_),
    .Y(_05059_),
    .A(_05048_));
 AO21x1_ASAP7_75t_R _27855_ (.A1(_05048_),
    .A2(_05050_),
    .B(_05058_),
    .Y(_05060_));
 BUFx4f_ASAP7_75t_R _27856_ (.A(_05060_),
    .Y(_05061_));
 NAND2x2_ASAP7_75t_R _27857_ (.A(_05059_),
    .B(_05061_),
    .Y(_05062_));
 BUFx12_ASAP7_75t_R _27858_ (.A(_05062_),
    .Y(_05063_));
 BUFx10_ASAP7_75t_R _27859_ (.A(_05063_),
    .Y(_16023_));
 BUFx6f_ASAP7_75t_R _27860_ (.A(_05057_),
    .Y(_05064_));
 NOR2x1_ASAP7_75t_R _27861_ (.A(_16026_),
    .B(_05064_),
    .Y(_05065_));
 INVx1_ASAP7_75t_R _27862_ (.A(_00619_),
    .Y(_05066_));
 AO21x2_ASAP7_75t_R _27863_ (.A1(_05053_),
    .A2(_05051_),
    .B(_05066_),
    .Y(_05067_));
 INVx2_ASAP7_75t_R _27864_ (.A(_05067_),
    .Y(_05068_));
 XNOR2x1_ASAP7_75t_R _27865_ (.B(_10712_),
    .Y(_05069_),
    .A(_10714_));
 NOR2x1_ASAP7_75t_R _27866_ (.A(_05069_),
    .B(_02277_),
    .Y(_05070_));
 XOR2x1_ASAP7_75t_R _27867_ (.A(_10712_),
    .Y(_05071_),
    .B(_10714_));
 OAI21x1_ASAP7_75t_R _27868_ (.A1(_05071_),
    .A2(_02280_),
    .B(_12921_),
    .Y(_05072_));
 NAND2x1_ASAP7_75t_R _27869_ (.A(_00645_),
    .B(net849),
    .Y(_05073_));
 OAI21x1_ASAP7_75t_R _27870_ (.A1(_05070_),
    .A2(_05072_),
    .B(_05073_),
    .Y(_05074_));
 XOR2x2_ASAP7_75t_R _27871_ (.A(_05074_),
    .B(_01020_),
    .Y(_05075_));
 BUFx6f_ASAP7_75t_R _27872_ (.A(_05075_),
    .Y(_05076_));
 BUFx6f_ASAP7_75t_R _27873_ (.A(_05076_),
    .Y(_05077_));
 OA21x2_ASAP7_75t_R _27874_ (.A1(_05065_),
    .A2(_05068_),
    .B(_05077_),
    .Y(_05078_));
 OAI21x1_ASAP7_75t_R _27875_ (.A1(_05013_),
    .A2(_05006_),
    .B(_05019_),
    .Y(_05079_));
 OAI21x1_ASAP7_75t_R _27876_ (.A1(_05015_),
    .A2(_05018_),
    .B(_08023_),
    .Y(_05080_));
 NAND2x2_ASAP7_75t_R _27877_ (.A(_05079_),
    .B(_05080_),
    .Y(_05081_));
 BUFx6f_ASAP7_75t_R _27878_ (.A(_05081_),
    .Y(_16014_));
 BUFx6f_ASAP7_75t_R _27879_ (.A(_05062_),
    .Y(_05082_));
 INVx4_ASAP7_75t_R _27880_ (.A(net473),
    .Y(_05083_));
 AOI21x1_ASAP7_75t_R _27881_ (.A1(_05051_),
    .A2(_05053_),
    .B(_05083_),
    .Y(_05084_));
 AO21x1_ASAP7_75t_R _27882_ (.A1(net43),
    .A2(_05082_),
    .B(net764),
    .Y(_05085_));
 XNOR2x2_ASAP7_75t_R _27883_ (.A(_01020_),
    .B(_05074_),
    .Y(_05086_));
 BUFx10_ASAP7_75t_R _27884_ (.A(_05086_),
    .Y(_05087_));
 BUFx6f_ASAP7_75t_R _27885_ (.A(_05087_),
    .Y(_05088_));
 XNOR2x1_ASAP7_75t_R _27886_ (.B(_10738_),
    .Y(_05089_),
    .A(_00800_));
 XNOR2x1_ASAP7_75t_R _27887_ (.B(_02294_),
    .Y(_05090_),
    .A(_10757_));
 NOR2x1_ASAP7_75t_R _27888_ (.A(_05089_),
    .B(_05090_),
    .Y(_05091_));
 AO21x1_ASAP7_75t_R _27889_ (.A1(_05090_),
    .A2(_05089_),
    .B(_12160_),
    .Y(_05092_));
 NAND2x1_ASAP7_75t_R _27890_ (.A(_00724_),
    .B(_12095_),
    .Y(_05093_));
 OAI21x1_ASAP7_75t_R _27891_ (.A1(_05091_),
    .A2(_05092_),
    .B(_05093_),
    .Y(_05094_));
 XOR2x2_ASAP7_75t_R _27892_ (.A(_05094_),
    .B(_01021_),
    .Y(_05095_));
 BUFx6f_ASAP7_75t_R _27893_ (.A(_05095_),
    .Y(_05096_));
 AO21x1_ASAP7_75t_R _27894_ (.A1(_05085_),
    .A2(_05088_),
    .B(_05096_),
    .Y(_05097_));
 XNOR2x2_ASAP7_75t_R _27895_ (.A(_01021_),
    .B(_05094_),
    .Y(_05098_));
 BUFx6f_ASAP7_75t_R _27896_ (.A(_05098_),
    .Y(_05099_));
 AOI21x1_ASAP7_75t_R _27897_ (.A1(net766),
    .A2(_05082_),
    .B(_05087_),
    .Y(_05100_));
 NOR2x1_ASAP7_75t_R _27898_ (.A(_05099_),
    .B(_05100_),
    .Y(_05101_));
 NOR2x2_ASAP7_75t_R _27899_ (.A(_01247_),
    .B(_05054_),
    .Y(_05102_));
 INVx1_ASAP7_75t_R _27900_ (.A(_00621_),
    .Y(_05103_));
 AO21x2_ASAP7_75t_R _27901_ (.A1(_05053_),
    .A2(_05051_),
    .B(_05103_),
    .Y(_05104_));
 INVx1_ASAP7_75t_R _27902_ (.A(_05104_),
    .Y(_05105_));
 BUFx10_ASAP7_75t_R _27903_ (.A(_05087_),
    .Y(_05106_));
 OAI21x1_ASAP7_75t_R _27904_ (.A1(_05102_),
    .A2(_05105_),
    .B(_05106_),
    .Y(_05107_));
 NOR2x1_ASAP7_75t_R _27905_ (.A(_11450_),
    .B(_00723_),
    .Y(_05108_));
 INVx1_ASAP7_75t_R _27906_ (.A(_05108_),
    .Y(_05109_));
 XOR2x1_ASAP7_75t_R _27907_ (.A(_10756_),
    .Y(_05110_),
    .B(_10783_));
 INVx1_ASAP7_75t_R _27908_ (.A(_05110_),
    .Y(_05111_));
 XOR2x1_ASAP7_75t_R _27909_ (.A(_10755_),
    .Y(_05112_),
    .B(_13671_));
 NAND2x1_ASAP7_75t_R _27910_ (.A(_05111_),
    .B(_05112_),
    .Y(_05113_));
 XOR2x1_ASAP7_75t_R _27911_ (.A(_10755_),
    .Y(_05114_),
    .B(_00832_));
 NAND2x1_ASAP7_75t_R _27912_ (.A(_05110_),
    .B(_05114_),
    .Y(_05115_));
 AO21x1_ASAP7_75t_R _27913_ (.A1(_05113_),
    .A2(_05115_),
    .B(_12092_),
    .Y(_05116_));
 AOI21x1_ASAP7_75t_R _27914_ (.A1(_05109_),
    .A2(_05116_),
    .B(_01022_),
    .Y(_05117_));
 NAND2x1_ASAP7_75t_R _27915_ (.A(_05113_),
    .B(_05115_),
    .Y(_05118_));
 INVx1_ASAP7_75t_R _27916_ (.A(_01022_),
    .Y(_05119_));
 AOI211x1_ASAP7_75t_R _27917_ (.A1(_05118_),
    .A2(_10829_),
    .B(_05108_),
    .C(_05119_),
    .Y(_05120_));
 NOR2x2_ASAP7_75t_R _27918_ (.A(_05117_),
    .B(_05120_),
    .Y(_05121_));
 INVx4_ASAP7_75t_R _27919_ (.A(_05121_),
    .Y(_05122_));
 BUFx10_ASAP7_75t_R _27920_ (.A(_05122_),
    .Y(_05123_));
 AOI21x1_ASAP7_75t_R _27921_ (.A1(_05101_),
    .A2(_05107_),
    .B(_05123_),
    .Y(_05124_));
 OAI21x1_ASAP7_75t_R _27922_ (.A1(_05078_),
    .A2(_05097_),
    .B(_05124_),
    .Y(_05125_));
 OAI21x1_ASAP7_75t_R _27923_ (.A1(_05083_),
    .A2(_05054_),
    .B(_05075_),
    .Y(_05126_));
 BUFx10_ASAP7_75t_R _27924_ (.A(_05086_),
    .Y(_05127_));
 BUFx6f_ASAP7_75t_R _27925_ (.A(_05127_),
    .Y(_05128_));
 NOR2x1_ASAP7_75t_R _27926_ (.A(_10632_),
    .B(_05038_),
    .Y(_05129_));
 NOR2x1_ASAP7_75t_R _27927_ (.A(_10624_),
    .B(_05040_),
    .Y(_05130_));
 OAI21x1_ASAP7_75t_R _27928_ (.A1(_05129_),
    .A2(_05130_),
    .B(_02246_),
    .Y(_05131_));
 NOR2x1_ASAP7_75t_R _27929_ (.A(net52),
    .B(_05043_),
    .Y(_05132_));
 NOR2x1_ASAP7_75t_R _27930_ (.A(_13569_),
    .B(_05045_),
    .Y(_05133_));
 OAI21x1_ASAP7_75t_R _27931_ (.A1(_05132_),
    .A2(_05133_),
    .B(_02258_),
    .Y(_05134_));
 AOI21x1_ASAP7_75t_R _27932_ (.A1(_05131_),
    .A2(_05134_),
    .B(_12161_),
    .Y(_05135_));
 NOR3x2_ASAP7_75t_R _27933_ (.B(_05058_),
    .C(_05049_),
    .Y(_05136_),
    .A(_05135_));
 OA21x2_ASAP7_75t_R _27934_ (.A1(_05135_),
    .A2(_05049_),
    .B(_05058_),
    .Y(_05137_));
 INVx3_ASAP7_75t_R _27935_ (.A(_01248_),
    .Y(_05138_));
 OAI21x1_ASAP7_75t_R _27936_ (.A1(_05136_),
    .A2(_05137_),
    .B(_05138_),
    .Y(_05139_));
 OA21x2_ASAP7_75t_R _27937_ (.A1(_05135_),
    .A2(_05049_),
    .B(_08031_),
    .Y(_05140_));
 INVx1_ASAP7_75t_R _27938_ (.A(_05059_),
    .Y(_05141_));
 INVx1_ASAP7_75t_R _27939_ (.A(_01249_),
    .Y(_05142_));
 OAI21x1_ASAP7_75t_R _27940_ (.A1(_05140_),
    .A2(_05141_),
    .B(_05142_),
    .Y(_05143_));
 NAND2x2_ASAP7_75t_R _27941_ (.A(_05139_),
    .B(_05143_),
    .Y(_05144_));
 AOI21x1_ASAP7_75t_R _27942_ (.A1(_05128_),
    .A2(_05144_),
    .B(_05099_),
    .Y(_05145_));
 NAND2x1_ASAP7_75t_R _27943_ (.A(_05126_),
    .B(_05145_),
    .Y(_05146_));
 BUFx6f_ASAP7_75t_R _27944_ (.A(_05075_),
    .Y(_05147_));
 BUFx6f_ASAP7_75t_R _27945_ (.A(_05098_),
    .Y(_05148_));
 OA21x2_ASAP7_75t_R _27946_ (.A1(net906),
    .A2(_05147_),
    .B(_05148_),
    .Y(_05149_));
 BUFx12_ASAP7_75t_R _27947_ (.A(_05021_),
    .Y(_05150_));
 BUFx10_ASAP7_75t_R _27948_ (.A(_05037_),
    .Y(_05151_));
 NAND2x2_ASAP7_75t_R _27949_ (.A(_05150_),
    .B(_05151_),
    .Y(_05152_));
 AOI21x1_ASAP7_75t_R _27950_ (.A1(_05054_),
    .A2(_05057_),
    .B(_05127_),
    .Y(_05153_));
 OAI21x1_ASAP7_75t_R _27951_ (.A1(_16026_),
    .A2(_05152_),
    .B(_05153_),
    .Y(_05154_));
 BUFx10_ASAP7_75t_R _27952_ (.A(_05121_),
    .Y(_05155_));
 AOI21x1_ASAP7_75t_R _27953_ (.A1(_05149_),
    .A2(_05154_),
    .B(_05155_),
    .Y(_05156_));
 NAND2x1_ASAP7_75t_R _27954_ (.A(_05146_),
    .B(_05156_),
    .Y(_05157_));
 XOR2x1_ASAP7_75t_R _27955_ (.A(_10783_),
    .Y(_05158_),
    .B(_00738_));
 XOR2x1_ASAP7_75t_R _27956_ (.A(_05158_),
    .Y(_05159_),
    .B(_13714_));
 XOR2x1_ASAP7_75t_R _27957_ (.A(_05159_),
    .Y(_05160_),
    .B(_10781_));
 NOR2x1_ASAP7_75t_R _27958_ (.A(_10761_),
    .B(_00722_),
    .Y(_05161_));
 AO21x1_ASAP7_75t_R _27959_ (.A1(_05160_),
    .A2(_10734_),
    .B(_05161_),
    .Y(_05162_));
 XOR2x2_ASAP7_75t_R _27960_ (.A(_05162_),
    .B(_01023_),
    .Y(_05163_));
 BUFx10_ASAP7_75t_R _27961_ (.A(_05163_),
    .Y(_05164_));
 AOI21x1_ASAP7_75t_R _27962_ (.A1(_05125_),
    .A2(_05157_),
    .B(_05164_),
    .Y(_05165_));
 BUFx6f_ASAP7_75t_R _27963_ (.A(_05095_),
    .Y(_05166_));
 BUFx10_ASAP7_75t_R _27964_ (.A(_05166_),
    .Y(_05167_));
 BUFx6f_ASAP7_75t_R _27965_ (.A(_05127_),
    .Y(_05168_));
 NAND2x1_ASAP7_75t_R _27966_ (.A(_05168_),
    .B(_05102_),
    .Y(_05169_));
 NAND2x2_ASAP7_75t_R _27967_ (.A(_05062_),
    .B(_05150_),
    .Y(_05170_));
 BUFx6f_ASAP7_75t_R _27968_ (.A(_05054_),
    .Y(_05171_));
 AOI21x1_ASAP7_75t_R _27969_ (.A1(net919),
    .A2(_05171_),
    .B(_05127_),
    .Y(_05172_));
 OAI21x1_ASAP7_75t_R _27970_ (.A1(_16018_),
    .A2(_05170_),
    .B(_05172_),
    .Y(_05173_));
 NAND2x1_ASAP7_75t_R _27971_ (.A(_05169_),
    .B(_05173_),
    .Y(_05174_));
 AOI21x1_ASAP7_75t_R _27972_ (.A1(_05066_),
    .A2(_05171_),
    .B(_05076_),
    .Y(_05175_));
 OAI21x1_ASAP7_75t_R _27973_ (.A1(_16018_),
    .A2(_05170_),
    .B(_05175_),
    .Y(_05176_));
 AO21x2_ASAP7_75t_R _27974_ (.A1(_05061_),
    .A2(_05059_),
    .B(_01247_),
    .Y(_05177_));
 OA21x2_ASAP7_75t_R _27975_ (.A1(_05177_),
    .A2(_05168_),
    .B(_05166_),
    .Y(_05178_));
 BUFx6f_ASAP7_75t_R _27976_ (.A(_05122_),
    .Y(_05179_));
 AOI21x1_ASAP7_75t_R _27977_ (.A1(_05176_),
    .A2(_05178_),
    .B(_05179_),
    .Y(_05180_));
 OAI21x1_ASAP7_75t_R _27978_ (.A1(_05167_),
    .A2(_05174_),
    .B(_05180_),
    .Y(_05181_));
 INVx2_ASAP7_75t_R _27979_ (.A(_01247_),
    .Y(_05182_));
 AND3x1_ASAP7_75t_R _27980_ (.A(_05087_),
    .B(_05171_),
    .C(_05182_),
    .Y(_05183_));
 AOI21x1_ASAP7_75t_R _27981_ (.A1(_05059_),
    .A2(_05061_),
    .B(_05103_),
    .Y(_05184_));
 AOI21x1_ASAP7_75t_R _27982_ (.A1(_05076_),
    .A2(_05184_),
    .B(_05095_),
    .Y(_05185_));
 INVx1_ASAP7_75t_R _27983_ (.A(_05185_),
    .Y(_05186_));
 NOR2x1_ASAP7_75t_R _27984_ (.A(_05183_),
    .B(_05186_),
    .Y(_05187_));
 INVx1_ASAP7_75t_R _27985_ (.A(_05187_),
    .Y(_05188_));
 OR3x1_ASAP7_75t_R _27986_ (.A(net44),
    .B(_16023_),
    .C(_05168_),
    .Y(_05189_));
 NOR2x2_ASAP7_75t_R _27987_ (.A(_05171_),
    .B(_05150_),
    .Y(_05190_));
 OAI21x1_ASAP7_75t_R _27988_ (.A1(_05171_),
    .A2(_05064_),
    .B(_05139_),
    .Y(_05191_));
 OAI21x1_ASAP7_75t_R _27989_ (.A1(_05190_),
    .A2(_05191_),
    .B(_05128_),
    .Y(_05192_));
 NAND2x1_ASAP7_75t_R _27990_ (.A(_05189_),
    .B(_05192_),
    .Y(_05193_));
 BUFx6f_ASAP7_75t_R _27991_ (.A(_05095_),
    .Y(_05194_));
 INVx1_ASAP7_75t_R _27992_ (.A(_01252_),
    .Y(_05195_));
 OAI21x1_ASAP7_75t_R _27993_ (.A1(net472),
    .A2(_05063_),
    .B(_05087_),
    .Y(_05196_));
 OAI21x1_ASAP7_75t_R _27994_ (.A1(_05195_),
    .A2(_05106_),
    .B(_05196_),
    .Y(_05197_));
 AOI21x1_ASAP7_75t_R _27995_ (.A1(_05194_),
    .A2(_05197_),
    .B(_05155_),
    .Y(_05198_));
 OAI21x1_ASAP7_75t_R _27996_ (.A1(_05188_),
    .A2(_05193_),
    .B(_05198_),
    .Y(_05199_));
 CKINVDCx5p33_ASAP7_75t_R _27997_ (.A(_05163_),
    .Y(_05200_));
 BUFx10_ASAP7_75t_R _27998_ (.A(_05200_),
    .Y(_05201_));
 AOI21x1_ASAP7_75t_R _27999_ (.A1(_05181_),
    .A2(_05199_),
    .B(_05201_),
    .Y(_05202_));
 XOR2x1_ASAP7_75t_R _28000_ (.A(_00738_),
    .Y(_05203_),
    .B(net50));
 XOR2x1_ASAP7_75t_R _28001_ (.A(_05203_),
    .Y(_05204_),
    .B(_00834_));
 XOR2x1_ASAP7_75t_R _28002_ (.A(_05204_),
    .Y(_05205_),
    .B(_10827_));
 NOR2x1_ASAP7_75t_R _28003_ (.A(_11451_),
    .B(_00721_),
    .Y(_05206_));
 AO21x1_ASAP7_75t_R _28004_ (.A1(_05205_),
    .A2(_10831_),
    .B(_05206_),
    .Y(_05207_));
 XOR2x2_ASAP7_75t_R _28005_ (.A(_05207_),
    .B(_01024_),
    .Y(_05208_));
 INVx6_ASAP7_75t_R _28006_ (.A(_05208_),
    .Y(_05209_));
 OAI21x1_ASAP7_75t_R _28007_ (.A1(_05165_),
    .A2(_05202_),
    .B(_05209_),
    .Y(_05210_));
 INVx2_ASAP7_75t_R _28008_ (.A(_01250_),
    .Y(_05211_));
 AO21x2_ASAP7_75t_R _28009_ (.A1(_05061_),
    .A2(_05059_),
    .B(_05211_),
    .Y(_05212_));
 AOI21x1_ASAP7_75t_R _28010_ (.A1(_05212_),
    .A2(_05153_),
    .B(_05099_),
    .Y(_05213_));
 NOR2x2_ASAP7_75t_R _28011_ (.A(_05054_),
    .B(net762),
    .Y(_05214_));
 AOI21x1_ASAP7_75t_R _28012_ (.A1(_16016_),
    .A2(_05064_),
    .B(_05082_),
    .Y(_05215_));
 OAI21x1_ASAP7_75t_R _28013_ (.A1(_05214_),
    .A2(_05215_),
    .B(_05106_),
    .Y(_05216_));
 NAND2x1_ASAP7_75t_R _28014_ (.A(_05213_),
    .B(_05216_),
    .Y(_05217_));
 BUFx6f_ASAP7_75t_R _28015_ (.A(_05075_),
    .Y(_05218_));
 OAI21x1_ASAP7_75t_R _28016_ (.A1(_05218_),
    .A2(_05177_),
    .B(_05148_),
    .Y(_05219_));
 NAND2x2_ASAP7_75t_R _28017_ (.A(_05054_),
    .B(net762),
    .Y(_05220_));
 NOR2x1_ASAP7_75t_R _28018_ (.A(_05076_),
    .B(_05220_),
    .Y(_05221_));
 NOR2x1_ASAP7_75t_R _28019_ (.A(_05219_),
    .B(_05221_),
    .Y(_05222_));
 BUFx10_ASAP7_75t_R _28020_ (.A(_05121_),
    .Y(_05223_));
 AOI21x1_ASAP7_75t_R _28021_ (.A1(_05154_),
    .A2(_05222_),
    .B(_05223_),
    .Y(_05224_));
 NAND2x1_ASAP7_75t_R _28022_ (.A(_05217_),
    .B(_05224_),
    .Y(_05225_));
 NAND2x2_ASAP7_75t_R _28023_ (.A(_05054_),
    .B(_05150_),
    .Y(_05226_));
 OAI21x1_ASAP7_75t_R _28024_ (.A1(_16018_),
    .A2(_05226_),
    .B(_05100_),
    .Y(_05227_));
 AOI21x1_ASAP7_75t_R _28025_ (.A1(_05171_),
    .A2(_05064_),
    .B(_05076_),
    .Y(_05228_));
 NOR2x1_ASAP7_75t_R _28026_ (.A(_05166_),
    .B(_05228_),
    .Y(_05229_));
 AOI21x1_ASAP7_75t_R _28027_ (.A1(_05227_),
    .A2(_05229_),
    .B(_05123_),
    .Y(_05230_));
 AOI21x1_ASAP7_75t_R _28028_ (.A1(_05059_),
    .A2(_05061_),
    .B(_05083_),
    .Y(_05231_));
 AOI21x1_ASAP7_75t_R _28029_ (.A1(_01250_),
    .A2(_05171_),
    .B(_05087_),
    .Y(_05232_));
 INVx2_ASAP7_75t_R _28030_ (.A(_05232_),
    .Y(_05233_));
 NAND2x2_ASAP7_75t_R _28031_ (.A(_05150_),
    .B(net552),
    .Y(_05234_));
 AOI21x1_ASAP7_75t_R _28032_ (.A1(_05082_),
    .A2(_05064_),
    .B(_05218_),
    .Y(_05235_));
 AOI21x1_ASAP7_75t_R _28033_ (.A1(_05234_),
    .A2(_05235_),
    .B(_05099_),
    .Y(_05236_));
 OAI21x1_ASAP7_75t_R _28034_ (.A1(_05231_),
    .A2(_05233_),
    .B(_05236_),
    .Y(_05237_));
 AOI21x1_ASAP7_75t_R _28035_ (.A1(_05230_),
    .A2(_05237_),
    .B(_05163_),
    .Y(_05238_));
 AOI21x1_ASAP7_75t_R _28036_ (.A1(_05225_),
    .A2(_05238_),
    .B(_05209_),
    .Y(_05239_));
 AO21x1_ASAP7_75t_R _28037_ (.A1(_05061_),
    .A2(_05059_),
    .B(_00622_),
    .Y(_05240_));
 BUFx4f_ASAP7_75t_R _28038_ (.A(_05240_),
    .Y(_05241_));
 BUFx6f_ASAP7_75t_R _28039_ (.A(_05127_),
    .Y(_05242_));
 AO21x1_ASAP7_75t_R _28040_ (.A1(_05104_),
    .A2(_05241_),
    .B(_05242_),
    .Y(_05243_));
 NAND2x1_ASAP7_75t_R _28041_ (.A(_05127_),
    .B(_05184_),
    .Y(_05244_));
 OA21x2_ASAP7_75t_R _28042_ (.A1(_05218_),
    .A2(_05067_),
    .B(_05244_),
    .Y(_05245_));
 AOI21x1_ASAP7_75t_R _28043_ (.A1(_05243_),
    .A2(_05245_),
    .B(_05096_),
    .Y(_05246_));
 NAND2x1_ASAP7_75t_R _28044_ (.A(_05127_),
    .B(_05231_),
    .Y(_05247_));
 AND2x2_ASAP7_75t_R _28045_ (.A(_05247_),
    .B(_05095_),
    .Y(_05248_));
 INVx2_ASAP7_75t_R _28046_ (.A(_05248_),
    .Y(_05249_));
 INVx1_ASAP7_75t_R _28047_ (.A(_05220_),
    .Y(_05250_));
 NOR2x2_ASAP7_75t_R _28048_ (.A(_05127_),
    .B(_05084_),
    .Y(_05251_));
 AO21x1_ASAP7_75t_R _28049_ (.A1(_05250_),
    .A2(_05242_),
    .B(_05251_),
    .Y(_05252_));
 OAI21x1_ASAP7_75t_R _28050_ (.A1(_05249_),
    .A2(_05252_),
    .B(_05123_),
    .Y(_05253_));
 NOR2x1_ASAP7_75t_R _28051_ (.A(_05246_),
    .B(_05253_),
    .Y(_05254_));
 NAND2x2_ASAP7_75t_R _28052_ (.A(net43),
    .B(net551),
    .Y(_05255_));
 AOI21x1_ASAP7_75t_R _28053_ (.A1(_05082_),
    .A2(_05151_),
    .B(_05076_),
    .Y(_05256_));
 NAND2x2_ASAP7_75t_R _28054_ (.A(_05255_),
    .B(_05256_),
    .Y(_05257_));
 AOI21x1_ASAP7_75t_R _28055_ (.A1(_16016_),
    .A2(net765),
    .B(_05168_),
    .Y(_05258_));
 NOR2x2_ASAP7_75t_R _28056_ (.A(_05063_),
    .B(net551),
    .Y(_05259_));
 INVx1_ASAP7_75t_R _28057_ (.A(_05259_),
    .Y(_05260_));
 AOI21x1_ASAP7_75t_R _28058_ (.A1(_05258_),
    .A2(_05260_),
    .B(_05099_),
    .Y(_05261_));
 NAND2x1_ASAP7_75t_R _28059_ (.A(_05257_),
    .B(_05261_),
    .Y(_05262_));
 AO21x1_ASAP7_75t_R _28060_ (.A1(_05061_),
    .A2(_05059_),
    .B(_05066_),
    .Y(_05263_));
 INVx1_ASAP7_75t_R _28061_ (.A(_05263_),
    .Y(_05264_));
 BUFx6f_ASAP7_75t_R _28062_ (.A(_05076_),
    .Y(_05265_));
 OAI21x1_ASAP7_75t_R _28063_ (.A1(_05105_),
    .A2(_05264_),
    .B(_05265_),
    .Y(_05266_));
 NOR2x1_ASAP7_75t_R _28064_ (.A(_05218_),
    .B(_05231_),
    .Y(_05267_));
 OAI21x1_ASAP7_75t_R _28065_ (.A1(net44),
    .A2(_05226_),
    .B(_05267_),
    .Y(_05268_));
 BUFx6f_ASAP7_75t_R _28066_ (.A(_05148_),
    .Y(_05269_));
 NAND3x1_ASAP7_75t_R _28067_ (.A(_05266_),
    .B(_05268_),
    .C(_05269_),
    .Y(_05270_));
 BUFx10_ASAP7_75t_R _28068_ (.A(_05122_),
    .Y(_05271_));
 AOI21x1_ASAP7_75t_R _28069_ (.A1(_05262_),
    .A2(_05270_),
    .B(_05271_),
    .Y(_05272_));
 OAI21x1_ASAP7_75t_R _28070_ (.A1(_05272_),
    .A2(_05254_),
    .B(_05164_),
    .Y(_05273_));
 NAND2x1_ASAP7_75t_R _28071_ (.A(_05239_),
    .B(_05273_),
    .Y(_05274_));
 NAND2x1_ASAP7_75t_R _28072_ (.A(_05210_),
    .B(_05274_),
    .Y(_00128_));
 NAND2x1_ASAP7_75t_R _28073_ (.A(_05226_),
    .B(_05256_),
    .Y(_05275_));
 NAND2x1_ASAP7_75t_R _28074_ (.A(_05220_),
    .B(_05100_),
    .Y(_05276_));
 AND3x1_ASAP7_75t_R _28075_ (.A(_05275_),
    .B(_05123_),
    .C(_05276_),
    .Y(_05277_));
 AO21x2_ASAP7_75t_R _28076_ (.A1(_05053_),
    .A2(_05051_),
    .B(_00621_),
    .Y(_05278_));
 AO21x1_ASAP7_75t_R _28077_ (.A1(_05235_),
    .A2(_05278_),
    .B(_05122_),
    .Y(_05279_));
 AOI21x1_ASAP7_75t_R _28078_ (.A1(_05150_),
    .A2(_05151_),
    .B(_05171_),
    .Y(_05280_));
 OA21x2_ASAP7_75t_R _28079_ (.A1(_05280_),
    .A2(_05215_),
    .B(_05077_),
    .Y(_05281_));
 OAI21x1_ASAP7_75t_R _28080_ (.A1(_05279_),
    .A2(_05281_),
    .B(_05167_),
    .Y(_05282_));
 BUFx6f_ASAP7_75t_R _28081_ (.A(_05148_),
    .Y(_05283_));
 NAND2x1_ASAP7_75t_R _28082_ (.A(_00623_),
    .B(_05265_),
    .Y(_05284_));
 NAND2x1_ASAP7_75t_R _28083_ (.A(_05151_),
    .B(_05214_),
    .Y(_05285_));
 NAND2x1_ASAP7_75t_R _28084_ (.A(_05175_),
    .B(_05285_),
    .Y(_05286_));
 OAI21x1_ASAP7_75t_R _28085_ (.A1(_05223_),
    .A2(_05284_),
    .B(_05286_),
    .Y(_05287_));
 AOI21x1_ASAP7_75t_R _28086_ (.A1(_05283_),
    .A2(_05287_),
    .B(_05200_),
    .Y(_05288_));
 OAI21x1_ASAP7_75t_R _28087_ (.A1(_05277_),
    .A2(_05282_),
    .B(_05288_),
    .Y(_05289_));
 AOI21x1_ASAP7_75t_R _28088_ (.A1(_05128_),
    .A2(_05259_),
    .B(_05148_),
    .Y(_05290_));
 INVx2_ASAP7_75t_R _28089_ (.A(_05290_),
    .Y(_05291_));
 NOR2x2_ASAP7_75t_R _28090_ (.A(_05063_),
    .B(_05127_),
    .Y(_05292_));
 NAND2x1_ASAP7_75t_R _28091_ (.A(_05083_),
    .B(_05292_),
    .Y(_05293_));
 NAND2x1_ASAP7_75t_R _28092_ (.A(_05147_),
    .B(_05184_),
    .Y(_05294_));
 NAND3x1_ASAP7_75t_R _28093_ (.A(_05293_),
    .B(_05169_),
    .C(_05294_),
    .Y(_05295_));
 NAND2x1_ASAP7_75t_R _28094_ (.A(_05278_),
    .B(_05256_),
    .Y(_05296_));
 BUFx6f_ASAP7_75t_R _28095_ (.A(_05095_),
    .Y(_05297_));
 AOI21x1_ASAP7_75t_R _28096_ (.A1(_05220_),
    .A2(_05100_),
    .B(_05297_),
    .Y(_05298_));
 AOI21x1_ASAP7_75t_R _28097_ (.A1(_05296_),
    .A2(_05298_),
    .B(_05123_),
    .Y(_05299_));
 OAI21x1_ASAP7_75t_R _28098_ (.A1(_05291_),
    .A2(_05295_),
    .B(_05299_),
    .Y(_05300_));
 INVx2_ASAP7_75t_R _28099_ (.A(_05126_),
    .Y(_05301_));
 NOR2x1_ASAP7_75t_R _28100_ (.A(_05166_),
    .B(_05301_),
    .Y(_05302_));
 OAI21x1_ASAP7_75t_R _28101_ (.A1(_16026_),
    .A2(_05152_),
    .B(_05228_),
    .Y(_05303_));
 AOI21x1_ASAP7_75t_R _28102_ (.A1(_05302_),
    .A2(_05303_),
    .B(_05223_),
    .Y(_05304_));
 INVx4_ASAP7_75t_R _28103_ (.A(_05241_),
    .Y(_05305_));
 NOR2x2_ASAP7_75t_R _28104_ (.A(_05063_),
    .B(_16014_),
    .Y(_05306_));
 AO21x2_ASAP7_75t_R _28105_ (.A1(_05306_),
    .A2(_05151_),
    .B(_05168_),
    .Y(_05307_));
 AO21x2_ASAP7_75t_R _28106_ (.A1(_05053_),
    .A2(_05051_),
    .B(_05182_),
    .Y(_05308_));
 AOI21x1_ASAP7_75t_R _28107_ (.A1(_01250_),
    .A2(_05082_),
    .B(_05076_),
    .Y(_05309_));
 BUFx6f_ASAP7_75t_R _28108_ (.A(_05098_),
    .Y(_05310_));
 AOI21x1_ASAP7_75t_R _28109_ (.A1(_05308_),
    .A2(_05309_),
    .B(_05310_),
    .Y(_05311_));
 OAI21x1_ASAP7_75t_R _28110_ (.A1(_05305_),
    .A2(_05307_),
    .B(_05311_),
    .Y(_05312_));
 AOI21x1_ASAP7_75t_R _28111_ (.A1(_05304_),
    .A2(_05312_),
    .B(_05163_),
    .Y(_05313_));
 AOI21x1_ASAP7_75t_R _28112_ (.A1(_05300_),
    .A2(_05313_),
    .B(_05209_),
    .Y(_05314_));
 NAND2x1_ASAP7_75t_R _28113_ (.A(_05289_),
    .B(_05314_),
    .Y(_05315_));
 OAI21x1_ASAP7_75t_R _28114_ (.A1(_16023_),
    .A2(_05064_),
    .B(_05168_),
    .Y(_05316_));
 INVx2_ASAP7_75t_R _28115_ (.A(_05139_),
    .Y(_05317_));
 OAI22x1_ASAP7_75t_R _28116_ (.A1(_05316_),
    .A2(_05184_),
    .B1(_05126_),
    .B2(_05317_),
    .Y(_05318_));
 AND2x2_ASAP7_75t_R _28117_ (.A(_05318_),
    .B(_05194_),
    .Y(_05319_));
 NAND2x1_ASAP7_75t_R _28118_ (.A(net43),
    .B(_05151_),
    .Y(_05320_));
 INVx1_ASAP7_75t_R _28119_ (.A(_05196_),
    .Y(_05321_));
 NAND2x2_ASAP7_75t_R _28120_ (.A(_05063_),
    .B(net552),
    .Y(_05322_));
 AOI22x1_ASAP7_75t_R _28121_ (.A1(_05153_),
    .A2(_05320_),
    .B1(_05321_),
    .B2(_05322_),
    .Y(_05323_));
 BUFx6f_ASAP7_75t_R _28122_ (.A(_05121_),
    .Y(_05324_));
 AO21x1_ASAP7_75t_R _28123_ (.A1(_05323_),
    .A2(_05283_),
    .B(_05324_),
    .Y(_05325_));
 NAND2x1_ASAP7_75t_R _28124_ (.A(_05128_),
    .B(_05280_),
    .Y(_05326_));
 NAND2x2_ASAP7_75t_R _28125_ (.A(_05063_),
    .B(_16014_),
    .Y(_05327_));
 AOI21x1_ASAP7_75t_R _28126_ (.A1(_05327_),
    .A2(_05232_),
    .B(_05099_),
    .Y(_05328_));
 AOI21x1_ASAP7_75t_R _28127_ (.A1(_05326_),
    .A2(_05328_),
    .B(_05123_),
    .Y(_05329_));
 OAI21x1_ASAP7_75t_R _28128_ (.A1(_05140_),
    .A2(_05141_),
    .B(_05138_),
    .Y(_05330_));
 OA21x2_ASAP7_75t_R _28129_ (.A1(_05330_),
    .A2(_05147_),
    .B(_05148_),
    .Y(_05331_));
 OAI21x1_ASAP7_75t_R _28130_ (.A1(_05305_),
    .A2(_05307_),
    .B(_05331_),
    .Y(_05332_));
 AOI21x1_ASAP7_75t_R _28131_ (.A1(_05329_),
    .A2(_05332_),
    .B(_05163_),
    .Y(_05333_));
 OAI21x1_ASAP7_75t_R _28132_ (.A1(_05319_),
    .A2(_05325_),
    .B(_05333_),
    .Y(_05334_));
 OA21x2_ASAP7_75t_R _28133_ (.A1(net906),
    .A2(_05218_),
    .B(_05095_),
    .Y(_05335_));
 AOI21x1_ASAP7_75t_R _28134_ (.A1(_05054_),
    .A2(_05150_),
    .B(_05127_),
    .Y(_05336_));
 NOR2x1_ASAP7_75t_R _28135_ (.A(_05190_),
    .B(_05336_),
    .Y(_05337_));
 AOI21x1_ASAP7_75t_R _28136_ (.A1(_05335_),
    .A2(_05337_),
    .B(_05223_),
    .Y(_05338_));
 AOI21x1_ASAP7_75t_R _28137_ (.A1(_05212_),
    .A2(_05251_),
    .B(_05297_),
    .Y(_05339_));
 NAND2x1_ASAP7_75t_R _28138_ (.A(_05192_),
    .B(_05339_),
    .Y(_05340_));
 AOI21x1_ASAP7_75t_R _28139_ (.A1(_05338_),
    .A2(_05340_),
    .B(_05200_),
    .Y(_05341_));
 AOI21x1_ASAP7_75t_R _28140_ (.A1(_05226_),
    .A2(_05320_),
    .B(_05147_),
    .Y(_05342_));
 AO21x1_ASAP7_75t_R _28141_ (.A1(_05292_),
    .A2(_05234_),
    .B(_05342_),
    .Y(_05343_));
 INVx3_ASAP7_75t_R _28142_ (.A(_05231_),
    .Y(_05344_));
 AOI21x1_ASAP7_75t_R _28143_ (.A1(_05344_),
    .A2(_05153_),
    .B(_05310_),
    .Y(_05345_));
 NAND2x1_ASAP7_75t_R _28144_ (.A(_05171_),
    .B(_05064_),
    .Y(_05346_));
 BUFx6f_ASAP7_75t_R _28145_ (.A(_05075_),
    .Y(_05347_));
 AO21x1_ASAP7_75t_R _28146_ (.A1(_05346_),
    .A2(_05330_),
    .B(_05347_),
    .Y(_05348_));
 AOI21x1_ASAP7_75t_R _28147_ (.A1(_05345_),
    .A2(_05348_),
    .B(_05179_),
    .Y(_05349_));
 OAI21x1_ASAP7_75t_R _28148_ (.A1(_05167_),
    .A2(_05343_),
    .B(_05349_),
    .Y(_05350_));
 AOI21x1_ASAP7_75t_R _28149_ (.A1(_05341_),
    .A2(_05350_),
    .B(_05208_),
    .Y(_05351_));
 NAND2x1_ASAP7_75t_R _28150_ (.A(_05334_),
    .B(_05351_),
    .Y(_05352_));
 NAND2x1_ASAP7_75t_R _28151_ (.A(_05315_),
    .B(_05352_),
    .Y(_00129_));
 NAND2x1_ASAP7_75t_R _28152_ (.A(_00623_),
    .B(_05128_),
    .Y(_05353_));
 AOI21x1_ASAP7_75t_R _28153_ (.A1(_05082_),
    .A2(_16016_),
    .B(_05087_),
    .Y(_05354_));
 AOI21x1_ASAP7_75t_R _28154_ (.A1(_05255_),
    .A2(_05354_),
    .B(_05095_),
    .Y(_05355_));
 AOI21x1_ASAP7_75t_R _28155_ (.A1(_05353_),
    .A2(_05355_),
    .B(_05223_),
    .Y(_05356_));
 AO21x1_ASAP7_75t_R _28156_ (.A1(_05053_),
    .A2(_05051_),
    .B(net473),
    .Y(_05357_));
 INVx1_ASAP7_75t_R _28157_ (.A(_05357_),
    .Y(_05358_));
 NAND2x1_ASAP7_75t_R _28158_ (.A(_05076_),
    .B(_05263_),
    .Y(_05359_));
 NOR2x1_ASAP7_75t_R _28159_ (.A(_05358_),
    .B(_05359_),
    .Y(_05360_));
 AND3x1_ASAP7_75t_R _28160_ (.A(_05170_),
    .B(_05168_),
    .C(_05104_),
    .Y(_05361_));
 OAI21x1_ASAP7_75t_R _28161_ (.A1(_05360_),
    .A2(_05361_),
    .B(_05096_),
    .Y(_05362_));
 NAND2x1_ASAP7_75t_R _28162_ (.A(_05356_),
    .B(_05362_),
    .Y(_05363_));
 OAI21x1_ASAP7_75t_R _28163_ (.A1(_05063_),
    .A2(_05150_),
    .B(_05075_),
    .Y(_05364_));
 INVx2_ASAP7_75t_R _28164_ (.A(_05364_),
    .Y(_05365_));
 NAND2x1_ASAP7_75t_R _28165_ (.A(_05322_),
    .B(_05365_),
    .Y(_05366_));
 AOI21x1_ASAP7_75t_R _28166_ (.A1(_05128_),
    .A2(_05085_),
    .B(_05099_),
    .Y(_05367_));
 NAND2x1_ASAP7_75t_R _28167_ (.A(_05366_),
    .B(_05367_),
    .Y(_05368_));
 OA21x2_ASAP7_75t_R _28168_ (.A1(_01252_),
    .A2(_05218_),
    .B(_05148_),
    .Y(_05369_));
 NAND2x2_ASAP7_75t_R _28169_ (.A(_05064_),
    .B(_05214_),
    .Y(_05370_));
 NAND2x1_ASAP7_75t_R _28170_ (.A(_05370_),
    .B(_05251_),
    .Y(_05371_));
 AOI21x1_ASAP7_75t_R _28171_ (.A1(_05371_),
    .A2(_05369_),
    .B(_05122_),
    .Y(_05372_));
 AOI21x1_ASAP7_75t_R _28172_ (.A1(_05368_),
    .A2(_05372_),
    .B(_05163_),
    .Y(_05373_));
 NAND2x1_ASAP7_75t_R _28173_ (.A(_05363_),
    .B(_05373_),
    .Y(_05374_));
 AOI21x1_ASAP7_75t_R _28174_ (.A1(_05150_),
    .A2(_05151_),
    .B(_05082_),
    .Y(_05375_));
 AOI21x1_ASAP7_75t_R _28175_ (.A1(_01247_),
    .A2(_01248_),
    .B(_16026_),
    .Y(_05376_));
 OA21x2_ASAP7_75t_R _28176_ (.A1(_05375_),
    .A2(_05376_),
    .B(_05077_),
    .Y(_05377_));
 AO21x1_ASAP7_75t_R _28177_ (.A1(_05285_),
    .A2(_05175_),
    .B(_05310_),
    .Y(_05378_));
 AO21x1_ASAP7_75t_R _28178_ (.A1(_05241_),
    .A2(net906),
    .B(_05242_),
    .Y(_05379_));
 INVx1_ASAP7_75t_R _28179_ (.A(_05244_),
    .Y(_05380_));
 NOR2x1_ASAP7_75t_R _28180_ (.A(_05166_),
    .B(_05380_),
    .Y(_05381_));
 AOI21x1_ASAP7_75t_R _28181_ (.A1(_05379_),
    .A2(_05381_),
    .B(_05123_),
    .Y(_05382_));
 OAI21x1_ASAP7_75t_R _28182_ (.A1(_05377_),
    .A2(_05378_),
    .B(_05382_),
    .Y(_05383_));
 OA21x2_ASAP7_75t_R _28183_ (.A1(_01254_),
    .A2(_05147_),
    .B(_05166_),
    .Y(_05384_));
 OAI21x1_ASAP7_75t_R _28184_ (.A1(_16023_),
    .A2(_05064_),
    .B(_16016_),
    .Y(_05385_));
 NAND2x1_ASAP7_75t_R _28185_ (.A(_05347_),
    .B(_05385_),
    .Y(_05386_));
 AOI21x1_ASAP7_75t_R _28186_ (.A1(_05384_),
    .A2(_05386_),
    .B(_05223_),
    .Y(_05387_));
 OAI21x1_ASAP7_75t_R _28187_ (.A1(_16018_),
    .A2(_05226_),
    .B(_05128_),
    .Y(_05388_));
 NAND2x2_ASAP7_75t_R _28188_ (.A(_00624_),
    .B(_05147_),
    .Y(_05389_));
 NAND3x1_ASAP7_75t_R _28189_ (.A(_05388_),
    .B(_05269_),
    .C(_05389_),
    .Y(_05390_));
 AOI21x1_ASAP7_75t_R _28190_ (.A1(_05387_),
    .A2(_05390_),
    .B(_05200_),
    .Y(_05391_));
 AOI21x1_ASAP7_75t_R _28191_ (.A1(_05383_),
    .A2(_05391_),
    .B(_05208_),
    .Y(_05392_));
 NAND2x1_ASAP7_75t_R _28192_ (.A(_05392_),
    .B(_05374_),
    .Y(_05393_));
 INVx3_ASAP7_75t_R _28193_ (.A(_05143_),
    .Y(_05394_));
 OAI21x1_ASAP7_75t_R _28194_ (.A1(_05136_),
    .A2(_05137_),
    .B(_05211_),
    .Y(_05395_));
 NAND2x2_ASAP7_75t_R _28195_ (.A(_05087_),
    .B(_05395_),
    .Y(_05396_));
 NOR2x1_ASAP7_75t_R _28196_ (.A(_05394_),
    .B(_05396_),
    .Y(_05397_));
 NOR2x2_ASAP7_75t_R _28197_ (.A(_05242_),
    .B(_05191_),
    .Y(_05398_));
 OAI21x1_ASAP7_75t_R _28198_ (.A1(_05397_),
    .A2(_05398_),
    .B(_05096_),
    .Y(_05399_));
 OAI21x1_ASAP7_75t_R _28199_ (.A1(_05317_),
    .A2(_05214_),
    .B(_05265_),
    .Y(_05400_));
 AOI21x1_ASAP7_75t_R _28200_ (.A1(_05106_),
    .A2(_05144_),
    .B(_05297_),
    .Y(_05401_));
 AOI21x1_ASAP7_75t_R _28201_ (.A1(_05400_),
    .A2(_05401_),
    .B(_05223_),
    .Y(_05402_));
 NAND2x1_ASAP7_75t_R _28202_ (.A(_05399_),
    .B(_05402_),
    .Y(_05403_));
 AOI21x1_ASAP7_75t_R _28203_ (.A1(net920),
    .A2(_05171_),
    .B(_05075_),
    .Y(_05404_));
 NAND2x1_ASAP7_75t_R _28204_ (.A(_05322_),
    .B(_05404_),
    .Y(_05405_));
 INVx2_ASAP7_75t_R _28205_ (.A(_05084_),
    .Y(_05406_));
 AO21x1_ASAP7_75t_R _28206_ (.A1(_05241_),
    .A2(_05406_),
    .B(_05128_),
    .Y(_05407_));
 AOI21x1_ASAP7_75t_R _28207_ (.A1(_05405_),
    .A2(_05407_),
    .B(_05194_),
    .Y(_05408_));
 NOR2x1_ASAP7_75t_R _28208_ (.A(_05394_),
    .B(_05364_),
    .Y(_05409_));
 INVx1_ASAP7_75t_R _28209_ (.A(_05395_),
    .Y(_05410_));
 OAI21x1_ASAP7_75t_R _28210_ (.A1(_16026_),
    .A2(_05064_),
    .B(_05168_),
    .Y(_05411_));
 OAI21x1_ASAP7_75t_R _28211_ (.A1(_05410_),
    .A2(_05411_),
    .B(_05297_),
    .Y(_05412_));
 NOR2x1_ASAP7_75t_R _28212_ (.A(_05409_),
    .B(_05412_),
    .Y(_05413_));
 OAI21x1_ASAP7_75t_R _28213_ (.A1(_05408_),
    .A2(_05413_),
    .B(_05324_),
    .Y(_05414_));
 AOI21x1_ASAP7_75t_R _28214_ (.A1(_05403_),
    .A2(_05414_),
    .B(_05164_),
    .Y(_05415_));
 AO21x1_ASAP7_75t_R _28215_ (.A1(_05170_),
    .A2(_05357_),
    .B(_05218_),
    .Y(_05416_));
 OAI21x1_ASAP7_75t_R _28216_ (.A1(_05190_),
    .A2(_05191_),
    .B(_05347_),
    .Y(_05417_));
 AOI21x1_ASAP7_75t_R _28217_ (.A1(_05416_),
    .A2(_05417_),
    .B(_05096_),
    .Y(_05418_));
 AOI21x1_ASAP7_75t_R _28218_ (.A1(_05395_),
    .A2(_05330_),
    .B(_05218_),
    .Y(_05419_));
 AOI21x1_ASAP7_75t_R _28219_ (.A1(_05347_),
    .A2(_05385_),
    .B(_05419_),
    .Y(_05420_));
 OAI21x1_ASAP7_75t_R _28220_ (.A1(_05269_),
    .A2(_05420_),
    .B(_05123_),
    .Y(_05421_));
 NOR2x1_ASAP7_75t_R _28221_ (.A(_05418_),
    .B(_05421_),
    .Y(_05422_));
 NOR2x2_ASAP7_75t_R _28222_ (.A(_01247_),
    .B(_05082_),
    .Y(_05423_));
 OAI21x1_ASAP7_75t_R _28223_ (.A1(_16026_),
    .A2(_05057_),
    .B(_05218_),
    .Y(_05424_));
 NOR2x1_ASAP7_75t_R _28224_ (.A(_05423_),
    .B(_05424_),
    .Y(_05425_));
 OAI21x1_ASAP7_75t_R _28225_ (.A1(_05063_),
    .A2(_05150_),
    .B(_05087_),
    .Y(_05426_));
 OAI21x1_ASAP7_75t_R _28226_ (.A1(_05305_),
    .A2(_05426_),
    .B(_05297_),
    .Y(_05427_));
 OAI21x1_ASAP7_75t_R _28227_ (.A1(_05425_),
    .A2(_05427_),
    .B(_05155_),
    .Y(_05428_));
 NOR2x1_ASAP7_75t_R _28228_ (.A(_01250_),
    .B(_16026_),
    .Y(_05429_));
 OAI21x1_ASAP7_75t_R _28229_ (.A1(_05429_),
    .A2(_05375_),
    .B(_05077_),
    .Y(_05430_));
 AOI21x1_ASAP7_75t_R _28230_ (.A1(_05388_),
    .A2(_05430_),
    .B(_05194_),
    .Y(_05431_));
 OAI21x1_ASAP7_75t_R _28231_ (.A1(_05428_),
    .A2(_05431_),
    .B(_05163_),
    .Y(_05432_));
 NOR2x1_ASAP7_75t_R _28232_ (.A(_05422_),
    .B(_05432_),
    .Y(_05433_));
 OAI21x1_ASAP7_75t_R _28233_ (.A1(_05415_),
    .A2(_05433_),
    .B(_05208_),
    .Y(_05434_));
 NAND2x1_ASAP7_75t_R _28234_ (.A(_05434_),
    .B(_05393_),
    .Y(_00130_));
 AND2x2_ASAP7_75t_R _28235_ (.A(_05412_),
    .B(_05179_),
    .Y(_05435_));
 NOR2x1_ASAP7_75t_R _28236_ (.A(net918),
    .B(_16023_),
    .Y(_05436_));
 OAI21x1_ASAP7_75t_R _28237_ (.A1(_05436_),
    .A2(_05376_),
    .B(_05265_),
    .Y(_05437_));
 AO21x1_ASAP7_75t_R _28238_ (.A1(_05286_),
    .A2(_05437_),
    .B(_05167_),
    .Y(_05438_));
 NAND2x1_ASAP7_75t_R _28239_ (.A(_05435_),
    .B(_05438_),
    .Y(_05439_));
 AO21x2_ASAP7_75t_R _28240_ (.A1(_05053_),
    .A2(_05051_),
    .B(_05211_),
    .Y(_05440_));
 AO21x1_ASAP7_75t_R _28241_ (.A1(_05267_),
    .A2(_05440_),
    .B(_05269_),
    .Y(_05441_));
 NOR2x1_ASAP7_75t_R _28242_ (.A(_16023_),
    .B(_05151_),
    .Y(_05442_));
 OAI21x1_ASAP7_75t_R _28243_ (.A1(_05394_),
    .A2(_05442_),
    .B(_05347_),
    .Y(_05443_));
 INVx1_ASAP7_75t_R _28244_ (.A(_05443_),
    .Y(_05444_));
 NAND2x1_ASAP7_75t_R _28245_ (.A(_05076_),
    .B(_05151_),
    .Y(_05445_));
 OAI21x1_ASAP7_75t_R _28246_ (.A1(_16023_),
    .A2(_05445_),
    .B(_05185_),
    .Y(_05446_));
 OAI22x1_ASAP7_75t_R _28247_ (.A1(_05441_),
    .A2(_05444_),
    .B1(_05446_),
    .B2(_05342_),
    .Y(_05447_));
 AOI21x1_ASAP7_75t_R _28248_ (.A1(_05324_),
    .A2(_05447_),
    .B(_05164_),
    .Y(_05448_));
 NAND2x1_ASAP7_75t_R _28249_ (.A(_05347_),
    .B(net764),
    .Y(_05449_));
 NAND2x1_ASAP7_75t_R _28250_ (.A(_05170_),
    .B(_05175_),
    .Y(_05450_));
 AOI21x1_ASAP7_75t_R _28251_ (.A1(_05449_),
    .A2(_05450_),
    .B(_05155_),
    .Y(_05451_));
 OAI21x1_ASAP7_75t_R _28252_ (.A1(_05179_),
    .A2(_05247_),
    .B(_05178_),
    .Y(_05452_));
 OAI21x1_ASAP7_75t_R _28253_ (.A1(_05451_),
    .A2(_05452_),
    .B(_05163_),
    .Y(_05453_));
 OA21x2_ASAP7_75t_R _28254_ (.A1(_05143_),
    .A2(_05242_),
    .B(_05121_),
    .Y(_05454_));
 NAND2x1_ASAP7_75t_R _28255_ (.A(_05405_),
    .B(_05454_),
    .Y(_05455_));
 AO21x2_ASAP7_75t_R _28256_ (.A1(_05061_),
    .A2(_05059_),
    .B(_05138_),
    .Y(_05456_));
 OAI21x1_ASAP7_75t_R _28257_ (.A1(_05182_),
    .A2(_05456_),
    .B(_05232_),
    .Y(_05457_));
 AOI21x1_ASAP7_75t_R _28258_ (.A1(_05344_),
    .A2(_05228_),
    .B(_05121_),
    .Y(_05458_));
 NAND2x1_ASAP7_75t_R _28259_ (.A(_05457_),
    .B(_05458_),
    .Y(_05459_));
 AOI21x1_ASAP7_75t_R _28260_ (.A1(_05455_),
    .A2(_05459_),
    .B(_05167_),
    .Y(_05460_));
 NOR2x1_ASAP7_75t_R _28261_ (.A(_05453_),
    .B(_05460_),
    .Y(_05461_));
 AOI21x1_ASAP7_75t_R _28262_ (.A1(_05439_),
    .A2(_05448_),
    .B(_05461_),
    .Y(_05462_));
 NAND2x1_ASAP7_75t_R _28263_ (.A(_05241_),
    .B(_05404_),
    .Y(_05463_));
 NAND2x1_ASAP7_75t_R _28264_ (.A(_05463_),
    .B(_05328_),
    .Y(_05464_));
 NAND2x1_ASAP7_75t_R _28265_ (.A(_16023_),
    .B(_05077_),
    .Y(_05465_));
 OAI21x1_ASAP7_75t_R _28266_ (.A1(_16016_),
    .A2(_05151_),
    .B(_05148_),
    .Y(_05466_));
 NOR2x2_ASAP7_75t_R _28267_ (.A(_05259_),
    .B(_05466_),
    .Y(_05467_));
 AOI21x1_ASAP7_75t_R _28268_ (.A1(_05465_),
    .A2(_05467_),
    .B(_05155_),
    .Y(_05468_));
 AOI21x1_ASAP7_75t_R _28269_ (.A1(_05464_),
    .A2(_05468_),
    .B(_05164_),
    .Y(_05469_));
 NOR2x1_ASAP7_75t_R _28270_ (.A(_05215_),
    .B(_05359_),
    .Y(_05470_));
 OAI21x1_ASAP7_75t_R _28271_ (.A1(_05196_),
    .A2(_05280_),
    .B(_05310_),
    .Y(_05471_));
 NOR2x1_ASAP7_75t_R _28272_ (.A(_05470_),
    .B(_05471_),
    .Y(_05472_));
 AO21x1_ASAP7_75t_R _28273_ (.A1(_05067_),
    .A2(_05344_),
    .B(_05347_),
    .Y(_05473_));
 NOR2x2_ASAP7_75t_R _28274_ (.A(_16014_),
    .B(_05037_),
    .Y(_05474_));
 BUFx6f_ASAP7_75t_R _28275_ (.A(_05218_),
    .Y(_05475_));
 OAI21x1_ASAP7_75t_R _28276_ (.A1(_05259_),
    .A2(_05474_),
    .B(_05475_),
    .Y(_05476_));
 AOI21x1_ASAP7_75t_R _28277_ (.A1(_05473_),
    .A2(_05476_),
    .B(_05283_),
    .Y(_05477_));
 OAI21x1_ASAP7_75t_R _28278_ (.A1(_05472_),
    .A2(_05477_),
    .B(_05324_),
    .Y(_05478_));
 AOI21x1_ASAP7_75t_R _28279_ (.A1(_05469_),
    .A2(_05478_),
    .B(_05208_),
    .Y(_05479_));
 AO21x1_ASAP7_75t_R _28280_ (.A1(_05211_),
    .A2(_16023_),
    .B(_05317_),
    .Y(_05480_));
 OAI21x1_ASAP7_75t_R _28281_ (.A1(_05305_),
    .A2(_05426_),
    .B(_05121_),
    .Y(_05481_));
 AO21x1_ASAP7_75t_R _28282_ (.A1(_05480_),
    .A2(_05077_),
    .B(_05481_),
    .Y(_05482_));
 NAND2x1_ASAP7_75t_R _28283_ (.A(_05234_),
    .B(_05256_),
    .Y(_05483_));
 OA21x2_ASAP7_75t_R _28284_ (.A1(_05364_),
    .A2(_05231_),
    .B(_05122_),
    .Y(_05484_));
 AOI21x1_ASAP7_75t_R _28285_ (.A1(_05483_),
    .A2(_05484_),
    .B(_05194_),
    .Y(_05485_));
 NAND2x1_ASAP7_75t_R _28286_ (.A(_05482_),
    .B(_05485_),
    .Y(_05486_));
 OA21x2_ASAP7_75t_R _28287_ (.A1(_05103_),
    .A2(_16026_),
    .B(_05251_),
    .Y(_05487_));
 OAI21x1_ASAP7_75t_R _28288_ (.A1(_05264_),
    .A2(_05316_),
    .B(_05223_),
    .Y(_05488_));
 AOI21x1_ASAP7_75t_R _28289_ (.A1(_05147_),
    .A2(_05084_),
    .B(_05121_),
    .Y(_05489_));
 OAI21x1_ASAP7_75t_R _28290_ (.A1(_05411_),
    .A2(_05306_),
    .B(_05489_),
    .Y(_05490_));
 OAI21x1_ASAP7_75t_R _28291_ (.A1(_05488_),
    .A2(_05487_),
    .B(_05490_),
    .Y(_05491_));
 AOI21x1_ASAP7_75t_R _28292_ (.A1(_05491_),
    .A2(_05167_),
    .B(_05201_),
    .Y(_05492_));
 NAND2x1_ASAP7_75t_R _28293_ (.A(_05486_),
    .B(_05492_),
    .Y(_05493_));
 NAND2x1_ASAP7_75t_R _28294_ (.A(_05493_),
    .B(_05479_),
    .Y(_05494_));
 OAI21x1_ASAP7_75t_R _28295_ (.A1(_05209_),
    .A2(_05462_),
    .B(_05494_),
    .Y(_00131_));
 AOI211x1_ASAP7_75t_R _28296_ (.A1(_05370_),
    .A2(_05365_),
    .B(_05419_),
    .C(_05283_),
    .Y(_05495_));
 OA21x2_ASAP7_75t_R _28297_ (.A1(_05128_),
    .A2(_05226_),
    .B(_05185_),
    .Y(_05496_));
 AO21x1_ASAP7_75t_R _28298_ (.A1(_05496_),
    .A2(_05192_),
    .B(_05324_),
    .Y(_05497_));
 NOR2x1_ASAP7_75t_R _28299_ (.A(_05495_),
    .B(_05497_),
    .Y(_05498_));
 NAND2x1_ASAP7_75t_R _28300_ (.A(_05406_),
    .B(_05309_),
    .Y(_05499_));
 NAND3x1_ASAP7_75t_R _28301_ (.A(_05173_),
    .B(_05283_),
    .C(_05499_),
    .Y(_05500_));
 AO21x1_ASAP7_75t_R _28302_ (.A1(_05357_),
    .A2(_05143_),
    .B(_05106_),
    .Y(_05501_));
 AOI21x1_ASAP7_75t_R _28303_ (.A1(_05501_),
    .A2(_05145_),
    .B(_05271_),
    .Y(_05502_));
 AO21x1_ASAP7_75t_R _28304_ (.A1(_05500_),
    .A2(_05502_),
    .B(_05201_),
    .Y(_05503_));
 NAND2x1_ASAP7_75t_R _28305_ (.A(_05095_),
    .B(_05177_),
    .Y(_05504_));
 OA21x2_ASAP7_75t_R _28306_ (.A1(_05504_),
    .A2(_05172_),
    .B(_05223_),
    .Y(_05505_));
 NAND2x1_ASAP7_75t_R _28307_ (.A(_05322_),
    .B(_05336_),
    .Y(_05506_));
 AOI21x1_ASAP7_75t_R _28308_ (.A1(_05278_),
    .A2(_05235_),
    .B(_05297_),
    .Y(_05507_));
 NAND2x1_ASAP7_75t_R _28309_ (.A(_05506_),
    .B(_05507_),
    .Y(_05508_));
 AOI21x1_ASAP7_75t_R _28310_ (.A1(_05505_),
    .A2(_05508_),
    .B(_05163_),
    .Y(_05509_));
 AND3x1_ASAP7_75t_R _28311_ (.A(_05327_),
    .B(_05265_),
    .C(_05278_),
    .Y(_05510_));
 AO21x1_ASAP7_75t_R _28312_ (.A1(_05234_),
    .A2(_05220_),
    .B(_05347_),
    .Y(_05511_));
 NAND2x1_ASAP7_75t_R _28313_ (.A(_05096_),
    .B(_05511_),
    .Y(_05512_));
 AOI21x1_ASAP7_75t_R _28314_ (.A1(_05275_),
    .A2(_05355_),
    .B(_05155_),
    .Y(_05513_));
 OAI21x1_ASAP7_75t_R _28315_ (.A1(_05510_),
    .A2(_05512_),
    .B(_05513_),
    .Y(_05514_));
 AOI21x1_ASAP7_75t_R _28316_ (.A1(_05509_),
    .A2(_05514_),
    .B(_05208_),
    .Y(_05515_));
 OAI21x1_ASAP7_75t_R _28317_ (.A1(_05498_),
    .A2(_05503_),
    .B(_05515_),
    .Y(_05516_));
 NAND2x2_ASAP7_75t_R _28318_ (.A(_05063_),
    .B(_05037_),
    .Y(_05517_));
 AOI21x1_ASAP7_75t_R _28319_ (.A1(_05517_),
    .A2(_05255_),
    .B(_05168_),
    .Y(_05518_));
 INVx1_ASAP7_75t_R _28320_ (.A(_05518_),
    .Y(_05519_));
 NAND2x1_ASAP7_75t_R _28321_ (.A(_05177_),
    .B(_05104_),
    .Y(_05520_));
 AOI21x1_ASAP7_75t_R _28322_ (.A1(_05128_),
    .A2(_05520_),
    .B(_05166_),
    .Y(_05521_));
 AOI21x1_ASAP7_75t_R _28323_ (.A1(_05519_),
    .A2(_05521_),
    .B(_05223_),
    .Y(_05522_));
 OAI21x1_ASAP7_75t_R _28324_ (.A1(_05474_),
    .A2(_05426_),
    .B(_05166_),
    .Y(_05523_));
 AO21x1_ASAP7_75t_R _28325_ (.A1(_05517_),
    .A2(_05172_),
    .B(_05523_),
    .Y(_05524_));
 NAND2x1_ASAP7_75t_R _28326_ (.A(_05522_),
    .B(_05524_),
    .Y(_05525_));
 INVx1_ASAP7_75t_R _28327_ (.A(_00625_),
    .Y(_05526_));
 NAND2x1_ASAP7_75t_R _28328_ (.A(_05526_),
    .B(_05242_),
    .Y(_05527_));
 AO21x1_ASAP7_75t_R _28329_ (.A1(_05293_),
    .A2(_05527_),
    .B(_05096_),
    .Y(_05528_));
 NAND2x2_ASAP7_75t_R _28330_ (.A(_05327_),
    .B(_05172_),
    .Y(_05529_));
 NAND2x1_ASAP7_75t_R _28331_ (.A(_05082_),
    .B(_05087_),
    .Y(_05530_));
 OA21x2_ASAP7_75t_R _28332_ (.A1(_05474_),
    .A2(_05530_),
    .B(_05166_),
    .Y(_05531_));
 AOI21x1_ASAP7_75t_R _28333_ (.A1(_05529_),
    .A2(_05531_),
    .B(_05123_),
    .Y(_05532_));
 AOI21x1_ASAP7_75t_R _28334_ (.A1(_05528_),
    .A2(_05532_),
    .B(_05200_),
    .Y(_05533_));
 NAND2x1_ASAP7_75t_R _28335_ (.A(_05525_),
    .B(_05533_),
    .Y(_05534_));
 AOI21x1_ASAP7_75t_R _28336_ (.A1(_05100_),
    .A2(_05220_),
    .B(_05380_),
    .Y(_05535_));
 NOR2x1_ASAP7_75t_R _28337_ (.A(_05099_),
    .B(_05221_),
    .Y(_05536_));
 NAND2x1_ASAP7_75t_R _28338_ (.A(_05535_),
    .B(_05536_),
    .Y(_05537_));
 AOI21x1_ASAP7_75t_R _28339_ (.A1(_05440_),
    .A2(_05256_),
    .B(_05292_),
    .Y(_05538_));
 AOI21x1_ASAP7_75t_R _28340_ (.A1(_05269_),
    .A2(_05538_),
    .B(_05155_),
    .Y(_05539_));
 AOI21x1_ASAP7_75t_R _28341_ (.A1(_05537_),
    .A2(_05539_),
    .B(_05163_),
    .Y(_05540_));
 AO21x1_ASAP7_75t_R _28342_ (.A1(_05330_),
    .A2(_05406_),
    .B(_05147_),
    .Y(_05541_));
 AOI21x1_ASAP7_75t_R _28343_ (.A1(_05541_),
    .A2(_05154_),
    .B(_05194_),
    .Y(_05542_));
 NAND2x2_ASAP7_75t_R _28344_ (.A(_05242_),
    .B(_05308_),
    .Y(_05543_));
 AOI21x1_ASAP7_75t_R _28345_ (.A1(_05543_),
    .A2(_05307_),
    .B(_05269_),
    .Y(_05544_));
 OAI21x1_ASAP7_75t_R _28346_ (.A1(_05544_),
    .A2(_05542_),
    .B(_05324_),
    .Y(_05545_));
 AOI21x1_ASAP7_75t_R _28347_ (.A1(_05545_),
    .A2(_05540_),
    .B(_05209_),
    .Y(_05546_));
 NAND2x1_ASAP7_75t_R _28348_ (.A(_05546_),
    .B(_05534_),
    .Y(_05547_));
 NAND2x1_ASAP7_75t_R _28349_ (.A(_05516_),
    .B(_05547_),
    .Y(_00132_));
 AND2x2_ASAP7_75t_R _28350_ (.A(_05445_),
    .B(_05148_),
    .Y(_05548_));
 AO21x1_ASAP7_75t_R _28351_ (.A1(_05548_),
    .A2(_05257_),
    .B(_05179_),
    .Y(_05549_));
 NAND2x1_ASAP7_75t_R _28352_ (.A(net44),
    .B(_05306_),
    .Y(_05550_));
 AO21x1_ASAP7_75t_R _28353_ (.A1(_05404_),
    .A2(_05327_),
    .B(_05310_),
    .Y(_05551_));
 AOI21x1_ASAP7_75t_R _28354_ (.A1(_05301_),
    .A2(_05550_),
    .B(_05551_),
    .Y(_05552_));
 OAI21x1_ASAP7_75t_R _28355_ (.A1(_05549_),
    .A2(_05552_),
    .B(_05201_),
    .Y(_05553_));
 AO21x1_ASAP7_75t_R _28356_ (.A1(_05068_),
    .A2(_05077_),
    .B(_05310_),
    .Y(_05554_));
 OA21x2_ASAP7_75t_R _28357_ (.A1(_05280_),
    .A2(_05410_),
    .B(_05088_),
    .Y(_05555_));
 OAI21x1_ASAP7_75t_R _28358_ (.A1(_05554_),
    .A2(_05555_),
    .B(_05271_),
    .Y(_05556_));
 NAND2x1_ASAP7_75t_R _28359_ (.A(_05106_),
    .B(_05191_),
    .Y(_05557_));
 AND3x1_ASAP7_75t_R _28360_ (.A(_05154_),
    .B(_05269_),
    .C(_05557_),
    .Y(_05558_));
 NOR2x1_ASAP7_75t_R _28361_ (.A(_05556_),
    .B(_05558_),
    .Y(_05559_));
 NOR2x1_ASAP7_75t_R _28362_ (.A(_05553_),
    .B(_05559_),
    .Y(_05560_));
 AO21x1_ASAP7_75t_R _28363_ (.A1(_00619_),
    .A2(_05077_),
    .B(_05096_),
    .Y(_05561_));
 AOI21x1_ASAP7_75t_R _28364_ (.A1(_16018_),
    .A2(_05214_),
    .B(_05475_),
    .Y(_05562_));
 OAI21x1_ASAP7_75t_R _28365_ (.A1(_05561_),
    .A2(_05562_),
    .B(_05271_),
    .Y(_05563_));
 OA21x2_ASAP7_75t_R _28366_ (.A1(_05068_),
    .A2(_05305_),
    .B(_05077_),
    .Y(_05564_));
 NAND2x1_ASAP7_75t_R _28367_ (.A(_05106_),
    .B(_05440_),
    .Y(_05565_));
 OAI21x1_ASAP7_75t_R _28368_ (.A1(_05305_),
    .A2(_05565_),
    .B(_05194_),
    .Y(_05566_));
 NOR2x1_ASAP7_75t_R _28369_ (.A(_05564_),
    .B(_05566_),
    .Y(_05567_));
 OAI21x1_ASAP7_75t_R _28370_ (.A1(_05563_),
    .A2(_05567_),
    .B(_05164_),
    .Y(_05568_));
 OR3x2_ASAP7_75t_R _28371_ (.A(_16026_),
    .B(_05182_),
    .C(_05138_),
    .Y(_05569_));
 AOI21x1_ASAP7_75t_R _28372_ (.A1(_05475_),
    .A2(_05569_),
    .B(_05167_),
    .Y(_05570_));
 AO21x1_ASAP7_75t_R _28373_ (.A1(_16018_),
    .A2(_05214_),
    .B(_05388_),
    .Y(_05571_));
 AO21x1_ASAP7_75t_R _28374_ (.A1(_05335_),
    .A2(_05233_),
    .B(_05179_),
    .Y(_05572_));
 AOI21x1_ASAP7_75t_R _28375_ (.A1(_05570_),
    .A2(_05571_),
    .B(_05572_),
    .Y(_05573_));
 OAI21x1_ASAP7_75t_R _28376_ (.A1(_05568_),
    .A2(_05573_),
    .B(_05208_),
    .Y(_05574_));
 AOI221x1_ASAP7_75t_R _28377_ (.A1(_05088_),
    .A2(_05456_),
    .B1(_05292_),
    .B2(_05234_),
    .C(_05283_),
    .Y(_05575_));
 AO21x1_ASAP7_75t_R _28378_ (.A1(_05168_),
    .A2(_05344_),
    .B(_05095_),
    .Y(_05576_));
 OAI21x1_ASAP7_75t_R _28379_ (.A1(_05576_),
    .A2(_05444_),
    .B(_05271_),
    .Y(_05577_));
 OAI21x1_ASAP7_75t_R _28380_ (.A1(_05575_),
    .A2(_05577_),
    .B(_05201_),
    .Y(_05578_));
 OA21x2_ASAP7_75t_R _28381_ (.A1(_05102_),
    .A2(_05138_),
    .B(_05265_),
    .Y(_05579_));
 AOI211x1_ASAP7_75t_R _28382_ (.A1(_05370_),
    .A2(_05404_),
    .B(_05579_),
    .C(_05283_),
    .Y(_05580_));
 AND2x2_ASAP7_75t_R _28383_ (.A(_05232_),
    .B(_05456_),
    .Y(_05581_));
 INVx1_ASAP7_75t_R _28384_ (.A(_05222_),
    .Y(_05582_));
 OAI21x1_ASAP7_75t_R _28385_ (.A1(_05581_),
    .A2(_05582_),
    .B(_05324_),
    .Y(_05583_));
 NOR2x1_ASAP7_75t_R _28386_ (.A(_05580_),
    .B(_05583_),
    .Y(_05584_));
 NOR2x1_ASAP7_75t_R _28387_ (.A(_05578_),
    .B(_05584_),
    .Y(_05585_));
 NAND2x1_ASAP7_75t_R _28388_ (.A(_05104_),
    .B(_05301_),
    .Y(_05586_));
 AOI21x1_ASAP7_75t_R _28389_ (.A1(_05396_),
    .A2(_05586_),
    .B(_05167_),
    .Y(_05587_));
 NOR2x1_ASAP7_75t_R _28390_ (.A(_05214_),
    .B(_05543_),
    .Y(_05588_));
 AO21x1_ASAP7_75t_R _28391_ (.A1(_05292_),
    .A2(_05083_),
    .B(_05269_),
    .Y(_05589_));
 OAI21x1_ASAP7_75t_R _28392_ (.A1(_05588_),
    .A2(_05589_),
    .B(_05271_),
    .Y(_05590_));
 OAI21x1_ASAP7_75t_R _28393_ (.A1(_05587_),
    .A2(_05590_),
    .B(_05164_),
    .Y(_05591_));
 OA21x2_ASAP7_75t_R _28394_ (.A1(_16016_),
    .A2(_05088_),
    .B(_05269_),
    .Y(_05592_));
 OAI21x1_ASAP7_75t_R _28395_ (.A1(_05474_),
    .A2(_05426_),
    .B(_05592_),
    .Y(_05593_));
 INVx1_ASAP7_75t_R _28396_ (.A(_05280_),
    .Y(_05594_));
 NAND2x1_ASAP7_75t_R _28397_ (.A(_05067_),
    .B(_05594_),
    .Y(_05595_));
 AOI21x1_ASAP7_75t_R _28398_ (.A1(_05152_),
    .A2(_05228_),
    .B(_05283_),
    .Y(_05596_));
 OAI21x1_ASAP7_75t_R _28399_ (.A1(_05088_),
    .A2(_05595_),
    .B(_05596_),
    .Y(_05597_));
 AOI21x1_ASAP7_75t_R _28400_ (.A1(_05593_),
    .A2(_05597_),
    .B(_05271_),
    .Y(_05598_));
 OAI21x1_ASAP7_75t_R _28401_ (.A1(_05591_),
    .A2(_05598_),
    .B(_05209_),
    .Y(_05599_));
 OAI22x1_ASAP7_75t_R _28402_ (.A1(_05560_),
    .A2(_05574_),
    .B1(_05585_),
    .B2(_05599_),
    .Y(_00133_));
 NAND2x1_ASAP7_75t_R _28403_ (.A(_05389_),
    .B(_05388_),
    .Y(_05600_));
 AOI21x1_ASAP7_75t_R _28404_ (.A1(_05600_),
    .A2(_05248_),
    .B(_05200_),
    .Y(_05601_));
 INVx1_ASAP7_75t_R _28405_ (.A(_05543_),
    .Y(_05602_));
 OA21x2_ASAP7_75t_R _28406_ (.A1(_05215_),
    .A2(_05214_),
    .B(_05475_),
    .Y(_05603_));
 OA21x2_ASAP7_75t_R _28407_ (.A1(_05241_),
    .A2(_05147_),
    .B(_05099_),
    .Y(_05604_));
 OAI21x1_ASAP7_75t_R _28408_ (.A1(_05602_),
    .A2(_05603_),
    .B(_05604_),
    .Y(_05605_));
 NAND2x1_ASAP7_75t_R _28409_ (.A(_05605_),
    .B(_05601_),
    .Y(_05606_));
 OAI21x1_ASAP7_75t_R _28410_ (.A1(_05394_),
    .A2(_05423_),
    .B(_05475_),
    .Y(_05607_));
 AND3x1_ASAP7_75t_R _28411_ (.A(_05607_),
    .B(_05194_),
    .C(_05244_),
    .Y(_05608_));
 NAND2x1_ASAP7_75t_R _28412_ (.A(_05234_),
    .B(_05365_),
    .Y(_05609_));
 AO21x1_ASAP7_75t_R _28413_ (.A1(_01253_),
    .A2(_01251_),
    .B(_05265_),
    .Y(_05610_));
 AND3x1_ASAP7_75t_R _28414_ (.A(_05609_),
    .B(_05283_),
    .C(_05610_),
    .Y(_05611_));
 OAI21x1_ASAP7_75t_R _28415_ (.A1(_05608_),
    .A2(_05611_),
    .B(_05201_),
    .Y(_05612_));
 AOI21x1_ASAP7_75t_R _28416_ (.A1(_05612_),
    .A2(_05606_),
    .B(_05271_),
    .Y(_05613_));
 OAI21x1_ASAP7_75t_R _28417_ (.A1(_05423_),
    .A2(_05144_),
    .B(_05475_),
    .Y(_05614_));
 OA21x2_ASAP7_75t_R _28418_ (.A1(_05065_),
    .A2(_05196_),
    .B(_05614_),
    .Y(_05615_));
 AO21x1_ASAP7_75t_R _28419_ (.A1(_05404_),
    .A2(_05212_),
    .B(_05297_),
    .Y(_05616_));
 OA21x2_ASAP7_75t_R _28420_ (.A1(_05375_),
    .A2(_05102_),
    .B(_05475_),
    .Y(_05617_));
 OAI21x1_ASAP7_75t_R _28421_ (.A1(_05616_),
    .A2(_05617_),
    .B(_05201_),
    .Y(_05618_));
 AOI21x1_ASAP7_75t_R _28422_ (.A1(_05167_),
    .A2(_05615_),
    .B(_05618_),
    .Y(_05619_));
 AO21x1_ASAP7_75t_R _28423_ (.A1(_05292_),
    .A2(net44),
    .B(_05096_),
    .Y(_05620_));
 AOI211x1_ASAP7_75t_R _28424_ (.A1(_05569_),
    .A2(_05321_),
    .B(_05620_),
    .C(_05518_),
    .Y(_05621_));
 AO21x1_ASAP7_75t_R _28425_ (.A1(_05517_),
    .A2(_16016_),
    .B(_05088_),
    .Y(_05622_));
 OA21x2_ASAP7_75t_R _28426_ (.A1(_05067_),
    .A2(_05265_),
    .B(_05297_),
    .Y(_05623_));
 AO21x1_ASAP7_75t_R _28427_ (.A1(_05622_),
    .A2(_05623_),
    .B(_05200_),
    .Y(_05624_));
 OAI21x1_ASAP7_75t_R _28428_ (.A1(_05621_),
    .A2(_05624_),
    .B(_05271_),
    .Y(_05625_));
 OAI21x1_ASAP7_75t_R _28429_ (.A1(_05619_),
    .A2(_05625_),
    .B(_05209_),
    .Y(_05626_));
 NOR2x1_ASAP7_75t_R _28430_ (.A(_05305_),
    .B(_05233_),
    .Y(_05627_));
 AOI21x1_ASAP7_75t_R _28431_ (.A1(_00626_),
    .A2(_05475_),
    .B(_05096_),
    .Y(_05628_));
 NAND2x1_ASAP7_75t_R _28432_ (.A(_05327_),
    .B(_05404_),
    .Y(_05629_));
 AOI21x1_ASAP7_75t_R _28433_ (.A1(_05628_),
    .A2(_05629_),
    .B(_05179_),
    .Y(_05630_));
 OAI21x1_ASAP7_75t_R _28434_ (.A1(_05291_),
    .A2(_05627_),
    .B(_05630_),
    .Y(_05631_));
 NAND2x1_ASAP7_75t_R _28435_ (.A(_05327_),
    .B(_05398_),
    .Y(_05632_));
 NOR2x1_ASAP7_75t_R _28436_ (.A(_05310_),
    .B(_05175_),
    .Y(_05633_));
 AOI21x1_ASAP7_75t_R _28437_ (.A1(_05529_),
    .A2(_05633_),
    .B(_05324_),
    .Y(_05634_));
 OAI21x1_ASAP7_75t_R _28438_ (.A1(_05167_),
    .A2(_05632_),
    .B(_05634_),
    .Y(_05635_));
 AOI21x1_ASAP7_75t_R _28439_ (.A1(_05631_),
    .A2(_05635_),
    .B(_05201_),
    .Y(_05636_));
 INVx1_ASAP7_75t_R _28440_ (.A(_05336_),
    .Y(_05637_));
 NAND2x1_ASAP7_75t_R _28441_ (.A(_05637_),
    .B(_05236_),
    .Y(_05638_));
 AOI21x1_ASAP7_75t_R _28442_ (.A1(_05604_),
    .A2(_05443_),
    .B(_05324_),
    .Y(_05639_));
 NAND2x1_ASAP7_75t_R _28443_ (.A(_05638_),
    .B(_05639_),
    .Y(_05640_));
 AOI21x1_ASAP7_75t_R _28444_ (.A1(net43),
    .A2(net765),
    .B(_05242_),
    .Y(_05641_));
 OAI21x1_ASAP7_75t_R _28445_ (.A1(_05309_),
    .A2(_05641_),
    .B(_05260_),
    .Y(_05642_));
 NAND2x1_ASAP7_75t_R _28446_ (.A(_05194_),
    .B(_05642_),
    .Y(_05643_));
 NAND2x1_ASAP7_75t_R _28447_ (.A(_05088_),
    .B(net43),
    .Y(_05644_));
 AOI21x1_ASAP7_75t_R _28448_ (.A1(_05644_),
    .A2(_05467_),
    .B(_05179_),
    .Y(_05645_));
 NAND2x1_ASAP7_75t_R _28449_ (.A(_05643_),
    .B(_05645_),
    .Y(_05646_));
 AOI21x1_ASAP7_75t_R _28450_ (.A1(_05640_),
    .A2(_05646_),
    .B(_05164_),
    .Y(_05647_));
 OAI21x1_ASAP7_75t_R _28451_ (.A1(_05636_),
    .A2(_05647_),
    .B(_05208_),
    .Y(_05648_));
 OAI21x1_ASAP7_75t_R _28452_ (.A1(_05626_),
    .A2(_05613_),
    .B(_05648_),
    .Y(_00134_));
 NOR2x1_ASAP7_75t_R _28453_ (.A(_05184_),
    .B(_05375_),
    .Y(_05649_));
 NOR2x1_ASAP7_75t_R _28454_ (.A(_05088_),
    .B(_05649_),
    .Y(_05650_));
 AO21x1_ASAP7_75t_R _28455_ (.A1(_16016_),
    .A2(net44),
    .B(_05530_),
    .Y(_05651_));
 NAND2x1_ASAP7_75t_R _28456_ (.A(_05290_),
    .B(_05651_),
    .Y(_05652_));
 NOR2x1_ASAP7_75t_R _28457_ (.A(_05297_),
    .B(_05309_),
    .Y(_05653_));
 AOI21x1_ASAP7_75t_R _28458_ (.A1(_05529_),
    .A2(_05653_),
    .B(_05123_),
    .Y(_05654_));
 OAI21x1_ASAP7_75t_R _28459_ (.A1(_05650_),
    .A2(_05652_),
    .B(_05654_),
    .Y(_05655_));
 INVx1_ASAP7_75t_R _28460_ (.A(_05366_),
    .Y(_05656_));
 AOI21x1_ASAP7_75t_R _28461_ (.A1(_05212_),
    .A2(_05251_),
    .B(_05310_),
    .Y(_05657_));
 NAND2x1_ASAP7_75t_R _28462_ (.A(_05344_),
    .B(_05228_),
    .Y(_05658_));
 AOI21x1_ASAP7_75t_R _28463_ (.A1(_05657_),
    .A2(_05658_),
    .B(_05155_),
    .Y(_05659_));
 OAI21x1_ASAP7_75t_R _28464_ (.A1(_05656_),
    .A2(_05616_),
    .B(_05659_),
    .Y(_05660_));
 AOI21x1_ASAP7_75t_R _28465_ (.A1(_05655_),
    .A2(_05660_),
    .B(_05164_),
    .Y(_05661_));
 AOI21x1_ASAP7_75t_R _28466_ (.A1(_05475_),
    .A2(_05594_),
    .B(_05576_),
    .Y(_05662_));
 OAI21x1_ASAP7_75t_R _28467_ (.A1(net44),
    .A2(_05226_),
    .B(_05106_),
    .Y(_05663_));
 OAI21x1_ASAP7_75t_R _28468_ (.A1(_16018_),
    .A2(_05170_),
    .B(_05077_),
    .Y(_05664_));
 OAI21x1_ASAP7_75t_R _28469_ (.A1(_05265_),
    .A2(_05241_),
    .B(_05297_),
    .Y(_05665_));
 AOI21x1_ASAP7_75t_R _28470_ (.A1(_05663_),
    .A2(_05664_),
    .B(_05665_),
    .Y(_05666_));
 OAI21x1_ASAP7_75t_R _28471_ (.A1(_05662_),
    .A2(_05666_),
    .B(_05271_),
    .Y(_05667_));
 NOR2x1_ASAP7_75t_R _28472_ (.A(_05347_),
    .B(_16018_),
    .Y(_05668_));
 INVx1_ASAP7_75t_R _28473_ (.A(_05506_),
    .Y(_05669_));
 OAI21x1_ASAP7_75t_R _28474_ (.A1(_05668_),
    .A2(_05669_),
    .B(_05194_),
    .Y(_05670_));
 OAI21x1_ASAP7_75t_R _28475_ (.A1(_05214_),
    .A2(_05375_),
    .B(_05106_),
    .Y(_05671_));
 AOI21x1_ASAP7_75t_R _28476_ (.A1(_05355_),
    .A2(_05671_),
    .B(_05179_),
    .Y(_05672_));
 NAND2x1_ASAP7_75t_R _28477_ (.A(_05670_),
    .B(_05672_),
    .Y(_05673_));
 AOI21x1_ASAP7_75t_R _28478_ (.A1(_05667_),
    .A2(_05673_),
    .B(_05201_),
    .Y(_05674_));
 OAI21x1_ASAP7_75t_R _28479_ (.A1(_05661_),
    .A2(_05674_),
    .B(_05208_),
    .Y(_05675_));
 AND3x1_ASAP7_75t_R _28480_ (.A(_05241_),
    .B(_05265_),
    .C(_05406_),
    .Y(_05676_));
 AO21x1_ASAP7_75t_R _28481_ (.A1(_05228_),
    .A2(_05327_),
    .B(_05310_),
    .Y(_05677_));
 OA21x2_ASAP7_75t_R _28482_ (.A1(_01253_),
    .A2(_05242_),
    .B(_05148_),
    .Y(_05678_));
 AO21x1_ASAP7_75t_R _28483_ (.A1(_05406_),
    .A2(_05143_),
    .B(_05347_),
    .Y(_05679_));
 AOI21x1_ASAP7_75t_R _28484_ (.A1(_05678_),
    .A2(_05679_),
    .B(_05155_),
    .Y(_05680_));
 OAI21x1_ASAP7_75t_R _28485_ (.A1(_05676_),
    .A2(_05677_),
    .B(_05680_),
    .Y(_05681_));
 AO21x1_ASAP7_75t_R _28486_ (.A1(_05100_),
    .A2(_05220_),
    .B(_05269_),
    .Y(_05682_));
 OA21x2_ASAP7_75t_R _28487_ (.A1(_05065_),
    .A2(net43),
    .B(_05088_),
    .Y(_05683_));
 OA21x2_ASAP7_75t_R _28488_ (.A1(_05526_),
    .A2(_05242_),
    .B(_05099_),
    .Y(_05684_));
 INVx1_ASAP7_75t_R _28489_ (.A(_05183_),
    .Y(_05685_));
 AOI21x1_ASAP7_75t_R _28490_ (.A1(_05684_),
    .A2(_05685_),
    .B(_05179_),
    .Y(_05686_));
 OAI21x1_ASAP7_75t_R _28491_ (.A1(_05682_),
    .A2(_05683_),
    .B(_05686_),
    .Y(_05687_));
 AOI21x1_ASAP7_75t_R _28492_ (.A1(_05681_),
    .A2(_05687_),
    .B(_05201_),
    .Y(_05688_));
 AO21x1_ASAP7_75t_R _28493_ (.A1(_05475_),
    .A2(_05250_),
    .B(_05380_),
    .Y(_05689_));
 OA21x2_ASAP7_75t_R _28494_ (.A1(_01248_),
    .A2(_05147_),
    .B(_05166_),
    .Y(_05690_));
 AOI21x1_ASAP7_75t_R _28495_ (.A1(_05690_),
    .A2(_05609_),
    .B(_05155_),
    .Y(_05691_));
 OAI21x1_ASAP7_75t_R _28496_ (.A1(_05188_),
    .A2(_05689_),
    .B(_05691_),
    .Y(_05692_));
 OAI21x1_ASAP7_75t_R _28497_ (.A1(_05068_),
    .A2(_05126_),
    .B(_05310_),
    .Y(_05693_));
 AOI21x1_ASAP7_75t_R _28498_ (.A1(_05088_),
    .A2(_05649_),
    .B(_05693_),
    .Y(_05694_));
 OAI21x1_ASAP7_75t_R _28499_ (.A1(_16023_),
    .A2(_16018_),
    .B(_16016_),
    .Y(_05695_));
 NAND2x1_ASAP7_75t_R _28500_ (.A(_05106_),
    .B(_05695_),
    .Y(_05696_));
 AOI21x1_ASAP7_75t_R _28501_ (.A1(_05437_),
    .A2(_05696_),
    .B(_05283_),
    .Y(_05697_));
 OAI21x1_ASAP7_75t_R _28502_ (.A1(_05694_),
    .A2(_05697_),
    .B(_05324_),
    .Y(_05698_));
 AOI21x1_ASAP7_75t_R _28503_ (.A1(_05692_),
    .A2(_05698_),
    .B(_05164_),
    .Y(_05699_));
 OAI21x1_ASAP7_75t_R _28504_ (.A1(_05688_),
    .A2(_05699_),
    .B(_05209_),
    .Y(_05700_));
 NAND2x1_ASAP7_75t_R _28505_ (.A(_05700_),
    .B(_05675_),
    .Y(_00135_));
 NOR2x1_ASAP7_75t_R _28506_ (.A(_10733_),
    .B(_00627_),
    .Y(_05701_));
 XOR2x1_ASAP7_75t_R _28507_ (.A(_11364_),
    .Y(_05702_),
    .B(_11365_));
 XOR2x1_ASAP7_75t_R _28508_ (.A(_11405_),
    .Y(_05703_),
    .B(_02909_));
 NAND2x1_ASAP7_75t_R _28509_ (.A(_05702_),
    .B(_05703_),
    .Y(_05704_));
 XNOR2x1_ASAP7_75t_R _28510_ (.B(_11365_),
    .Y(_05705_),
    .A(_11364_));
 XOR2x1_ASAP7_75t_R _28511_ (.A(_02909_),
    .Y(_05706_),
    .B(_11407_));
 NAND2x1_ASAP7_75t_R _28512_ (.A(_05706_),
    .B(_05705_),
    .Y(_05707_));
 AOI21x1_ASAP7_75t_R _28513_ (.A1(_05707_),
    .A2(_05704_),
    .B(_11374_),
    .Y(_05708_));
 OAI21x1_ASAP7_75t_R _28514_ (.A1(_05701_),
    .A2(_05708_),
    .B(_08024_),
    .Y(_05709_));
 AND2x2_ASAP7_75t_R _28515_ (.A(_11441_),
    .B(_00627_),
    .Y(_05710_));
 NAND2x1_ASAP7_75t_R _28516_ (.A(_05706_),
    .B(_05702_),
    .Y(_05711_));
 NAND2x1_ASAP7_75t_R _28517_ (.A(_05705_),
    .B(_05703_),
    .Y(_05712_));
 AOI21x1_ASAP7_75t_R _28518_ (.A1(_05712_),
    .A2(_05711_),
    .B(_11374_),
    .Y(_05713_));
 INVx1_ASAP7_75t_R _28519_ (.A(_08024_),
    .Y(_05714_));
 OAI21x1_ASAP7_75t_R _28520_ (.A1(_05710_),
    .A2(_05713_),
    .B(_05714_),
    .Y(_05715_));
 NAND2x2_ASAP7_75t_R _28521_ (.A(_05709_),
    .B(_05715_),
    .Y(_05716_));
 BUFx12_ASAP7_75t_R _28522_ (.A(_05716_),
    .Y(_16033_));
 OR2x2_ASAP7_75t_R _28523_ (.A(_10723_),
    .B(_00628_),
    .Y(_05717_));
 NOR2x2_ASAP7_75t_R _28524_ (.A(_11537_),
    .B(_11393_),
    .Y(_05718_));
 NOR2x2_ASAP7_75t_R _28525_ (.A(_11536_),
    .B(_11389_),
    .Y(_05719_));
 OAI21x1_ASAP7_75t_R _28526_ (.A1(_05718_),
    .A2(_05719_),
    .B(net625),
    .Y(_05720_));
 INVx1_ASAP7_75t_R _28527_ (.A(_05720_),
    .Y(_05721_));
 NOR3x1_ASAP7_75t_R _28528_ (.A(_05719_),
    .B(_05718_),
    .C(net626),
    .Y(_05722_));
 OAI21x1_ASAP7_75t_R _28529_ (.A1(_05721_),
    .A2(_05722_),
    .B(_11356_),
    .Y(_05723_));
 AOI21x1_ASAP7_75t_R _28530_ (.A1(_05717_),
    .A2(_05723_),
    .B(net858),
    .Y(_05724_));
 NAND2x1_ASAP7_75t_R _28531_ (.A(_00628_),
    .B(_12160_),
    .Y(_05725_));
 NAND2x2_ASAP7_75t_R _28532_ (.A(_11537_),
    .B(_11393_),
    .Y(_05726_));
 INVx1_ASAP7_75t_R _28533_ (.A(net625),
    .Y(_05727_));
 NOR2x1_ASAP7_75t_R _28534_ (.A(net705),
    .B(_11388_),
    .Y(_05728_));
 AND2x2_ASAP7_75t_R _28535_ (.A(net705),
    .B(_11388_),
    .Y(_05729_));
 OAI21x1_ASAP7_75t_R _28536_ (.A1(_05728_),
    .A2(_05729_),
    .B(_11536_),
    .Y(_05730_));
 NAND3x2_ASAP7_75t_R _28537_ (.B(_05726_),
    .C(_05730_),
    .Y(_05731_),
    .A(_05727_));
 NAND3x2_ASAP7_75t_R _28538_ (.B(_05731_),
    .C(_05720_),
    .Y(_05732_),
    .A(_10733_));
 INVx1_ASAP7_75t_R _28539_ (.A(net858),
    .Y(_05733_));
 AOI21x1_ASAP7_75t_R _28540_ (.A1(_05725_),
    .A2(_05732_),
    .B(_05733_),
    .Y(_05734_));
 NOR2x2_ASAP7_75t_R _28541_ (.A(_05724_),
    .B(_05734_),
    .Y(_05735_));
 BUFx12_ASAP7_75t_R _28542_ (.A(_05735_),
    .Y(_16035_));
 NOR2x1_ASAP7_75t_R _28543_ (.A(net680),
    .B(_00630_),
    .Y(_05736_));
 INVx3_ASAP7_75t_R _28544_ (.A(_05736_),
    .Y(_05737_));
 XOR2x1_ASAP7_75t_R _28545_ (.A(net789),
    .Y(_05738_),
    .B(_11409_));
 NAND2x1_ASAP7_75t_R _28546_ (.A(_02910_),
    .B(_05738_),
    .Y(_05739_));
 XNOR2x1_ASAP7_75t_R _28547_ (.B(_11409_),
    .Y(_05740_),
    .A(net789));
 NAND2x1_ASAP7_75t_R _28548_ (.A(net700),
    .B(_05740_),
    .Y(_05741_));
 AOI21x1_ASAP7_75t_R _28549_ (.A1(_05739_),
    .A2(_05741_),
    .B(_02960_),
    .Y(_05742_));
 XOR2x1_ASAP7_75t_R _28550_ (.A(_11409_),
    .Y(_05743_),
    .B(net702));
 NAND2x1_ASAP7_75t_R _28551_ (.A(net789),
    .B(_05743_),
    .Y(_05744_));
 XNOR2x1_ASAP7_75t_R _28552_ (.B(net702),
    .Y(_05745_),
    .A(_11409_));
 NAND2x1_ASAP7_75t_R _28553_ (.A(_14315_),
    .B(_05745_),
    .Y(_05746_));
 AOI21x1_ASAP7_75t_R _28554_ (.A1(_05744_),
    .A2(_05746_),
    .B(_02950_),
    .Y(_05747_));
 OAI21x1_ASAP7_75t_R _28555_ (.A1(_05742_),
    .A2(_05747_),
    .B(net767),
    .Y(_05748_));
 AOI21x1_ASAP7_75t_R _28556_ (.A1(_05737_),
    .A2(_05748_),
    .B(_08033_),
    .Y(_05749_));
 INVx4_ASAP7_75t_R _28557_ (.A(_05749_),
    .Y(_05750_));
 NAND3x2_ASAP7_75t_R _28558_ (.B(_08033_),
    .C(_05737_),
    .Y(_05751_),
    .A(_05748_));
 NAND2x2_ASAP7_75t_R _28559_ (.A(_05750_),
    .B(_05751_),
    .Y(_05752_));
 BUFx10_ASAP7_75t_R _28560_ (.A(_05752_),
    .Y(_16043_));
 AOI21x1_ASAP7_75t_R _28561_ (.A1(_05717_),
    .A2(_05723_),
    .B(_05733_),
    .Y(_05753_));
 AOI21x1_ASAP7_75t_R _28562_ (.A1(_05732_),
    .A2(_05725_),
    .B(net860),
    .Y(_05754_));
 NOR2x2_ASAP7_75t_R _28563_ (.A(_05753_),
    .B(_05754_),
    .Y(_05755_));
 BUFx6f_ASAP7_75t_R _28564_ (.A(_05755_),
    .Y(_16030_));
 INVx2_ASAP7_75t_R _28565_ (.A(_08033_),
    .Y(_05756_));
 NAND3x2_ASAP7_75t_R _28566_ (.B(_05756_),
    .C(_05737_),
    .Y(_05757_),
    .A(_05748_));
 AO21x1_ASAP7_75t_R _28567_ (.A1(_05748_),
    .A2(_05737_),
    .B(_05756_),
    .Y(_05758_));
 BUFx4f_ASAP7_75t_R _28568_ (.A(_05758_),
    .Y(_05759_));
 NAND2x2_ASAP7_75t_R _28569_ (.A(_05757_),
    .B(_05759_),
    .Y(_05760_));
 BUFx10_ASAP7_75t_R _28570_ (.A(_05760_),
    .Y(_16040_));
 XNOR2x1_ASAP7_75t_R _28571_ (.B(_11434_),
    .Y(_05761_),
    .A(_00807_));
 XOR2x1_ASAP7_75t_R _28572_ (.A(_02976_),
    .Y(_05762_),
    .B(_02975_));
 NOR2x1_ASAP7_75t_R _28573_ (.A(_05761_),
    .B(_05762_),
    .Y(_05763_));
 XOR2x1_ASAP7_75t_R _28574_ (.A(_11434_),
    .Y(_05764_),
    .B(_00807_));
 OAI21x1_ASAP7_75t_R _28575_ (.A1(_05764_),
    .A2(_02977_),
    .B(net867),
    .Y(_05765_));
 NAND2x1_ASAP7_75t_R _28576_ (.A(_00667_),
    .B(_10689_),
    .Y(_05766_));
 OAI21x1_ASAP7_75t_R _28577_ (.A1(_05763_),
    .A2(_05765_),
    .B(_05766_),
    .Y(_05767_));
 XOR2x2_ASAP7_75t_R _28578_ (.A(_05767_),
    .B(_08262_),
    .Y(_05768_));
 BUFx10_ASAP7_75t_R _28579_ (.A(_05768_),
    .Y(_05769_));
 BUFx6f_ASAP7_75t_R _28580_ (.A(_05769_),
    .Y(_05770_));
 INVx1_ASAP7_75t_R _28581_ (.A(_00631_),
    .Y(_05771_));
 AO21x2_ASAP7_75t_R _28582_ (.A1(_05759_),
    .A2(_05757_),
    .B(_05771_),
    .Y(_05772_));
 INVx2_ASAP7_75t_R _28583_ (.A(_05772_),
    .Y(_05773_));
 XNOR2x1_ASAP7_75t_R _28584_ (.B(_11463_),
    .Y(_05774_),
    .A(_00808_));
 XOR2x2_ASAP7_75t_R _28585_ (.A(_05774_),
    .B(_02987_),
    .Y(_05775_));
 NOR2x1_ASAP7_75t_R _28586_ (.A(_10743_),
    .B(_00666_),
    .Y(_05776_));
 AOI21x1_ASAP7_75t_R _28587_ (.A1(_10734_),
    .A2(_05775_),
    .B(_05776_),
    .Y(_05777_));
 XOR2x2_ASAP7_75t_R _28588_ (.A(_05777_),
    .B(_01053_),
    .Y(_05778_));
 BUFx6f_ASAP7_75t_R _28589_ (.A(_05778_),
    .Y(_05779_));
 AOI21x1_ASAP7_75t_R _28590_ (.A1(_05770_),
    .A2(_05773_),
    .B(_05779_),
    .Y(_05780_));
 BUFx4f_ASAP7_75t_R _28591_ (.A(_05751_),
    .Y(_05781_));
 BUFx4f_ASAP7_75t_R _28592_ (.A(_05750_),
    .Y(_05782_));
 AO21x2_ASAP7_75t_R _28593_ (.A1(_05781_),
    .A2(_05782_),
    .B(_00631_),
    .Y(_05783_));
 INVx1_ASAP7_75t_R _28594_ (.A(_00632_),
    .Y(_05784_));
 AOI21x1_ASAP7_75t_R _28595_ (.A1(_05757_),
    .A2(_05759_),
    .B(_05784_),
    .Y(_05785_));
 NOR2x2_ASAP7_75t_R _28596_ (.A(_05768_),
    .B(_05785_),
    .Y(_05786_));
 NAND2x1_ASAP7_75t_R _28597_ (.A(_05783_),
    .B(_05786_),
    .Y(_05787_));
 INVx3_ASAP7_75t_R _28598_ (.A(_00629_),
    .Y(_05788_));
 AO21x2_ASAP7_75t_R _28599_ (.A1(_05781_),
    .A2(_05782_),
    .B(_05788_),
    .Y(_05789_));
 INVx1_ASAP7_75t_R _28600_ (.A(_05789_),
    .Y(_05790_));
 NAND2x1_ASAP7_75t_R _28601_ (.A(_05770_),
    .B(_05790_),
    .Y(_05791_));
 AND3x1_ASAP7_75t_R _28602_ (.A(_05780_),
    .B(_05787_),
    .C(_05791_),
    .Y(_05792_));
 XOR2x2_ASAP7_75t_R _28603_ (.A(_05777_),
    .B(_08058_),
    .Y(_05793_));
 BUFx6f_ASAP7_75t_R _28604_ (.A(_05793_),
    .Y(_05794_));
 BUFx6f_ASAP7_75t_R _28605_ (.A(_05794_),
    .Y(_05795_));
 BUFx10_ASAP7_75t_R _28606_ (.A(_05752_),
    .Y(_05796_));
 BUFx12_ASAP7_75t_R _28607_ (.A(_05716_),
    .Y(_05797_));
 NAND2x2_ASAP7_75t_R _28608_ (.A(_05796_),
    .B(_05797_),
    .Y(_05798_));
 AO21x2_ASAP7_75t_R _28609_ (.A1(_05759_),
    .A2(_05757_),
    .B(_00632_),
    .Y(_05799_));
 NAND2x1_ASAP7_75t_R _28610_ (.A(_05769_),
    .B(_05799_),
    .Y(_05800_));
 INVx1_ASAP7_75t_R _28611_ (.A(_05800_),
    .Y(_05801_));
 AOI21x1_ASAP7_75t_R _28612_ (.A1(_05750_),
    .A2(_05751_),
    .B(_05784_),
    .Y(_05802_));
 NOR2x2_ASAP7_75t_R _28613_ (.A(_05802_),
    .B(_05769_),
    .Y(_05803_));
 AOI21x1_ASAP7_75t_R _28614_ (.A1(_05798_),
    .A2(_05801_),
    .B(_05803_),
    .Y(_05804_));
 NOR2x2_ASAP7_75t_R _28615_ (.A(net585),
    .B(_00665_),
    .Y(_05805_));
 INVx1_ASAP7_75t_R _28616_ (.A(_05805_),
    .Y(_05806_));
 XOR2x1_ASAP7_75t_R _28617_ (.A(_00744_),
    .Y(_05807_),
    .B(_00745_));
 XOR2x1_ASAP7_75t_R _28618_ (.A(_11487_),
    .Y(_05808_),
    .B(_00840_));
 NAND2x1_ASAP7_75t_R _28619_ (.A(_05807_),
    .B(_05808_),
    .Y(_05809_));
 INVx1_ASAP7_75t_R _28620_ (.A(_05807_),
    .Y(_05810_));
 XNOR2x1_ASAP7_75t_R _28621_ (.B(_11487_),
    .Y(_05811_),
    .A(_00840_));
 NAND2x1_ASAP7_75t_R _28622_ (.A(_05810_),
    .B(_05811_),
    .Y(_05812_));
 AOI21x1_ASAP7_75t_R _28623_ (.A1(_05809_),
    .A2(_05812_),
    .B(_12095_),
    .Y(_05813_));
 INVx1_ASAP7_75t_R _28624_ (.A(_05813_),
    .Y(_05814_));
 AOI21x1_ASAP7_75t_R _28625_ (.A1(_05806_),
    .A2(_05814_),
    .B(_01054_),
    .Y(_05815_));
 NOR3x2_ASAP7_75t_R _28626_ (.B(_08066_),
    .C(_05805_),
    .Y(_05816_),
    .A(_05813_));
 NOR2x2_ASAP7_75t_R _28627_ (.A(_05815_),
    .B(_05816_),
    .Y(_05817_));
 INVx3_ASAP7_75t_R _28628_ (.A(_05817_),
    .Y(_05818_));
 BUFx10_ASAP7_75t_R _28629_ (.A(_05818_),
    .Y(_05819_));
 OAI21x1_ASAP7_75t_R _28630_ (.A1(_05795_),
    .A2(_05804_),
    .B(_05819_),
    .Y(_05820_));
 OAI21x1_ASAP7_75t_R _28631_ (.A1(_05701_),
    .A2(_05708_),
    .B(_05714_),
    .Y(_05821_));
 OAI21x1_ASAP7_75t_R _28632_ (.A1(_05713_),
    .A2(_05710_),
    .B(_08024_),
    .Y(_05822_));
 NAND2x2_ASAP7_75t_R _28633_ (.A(_05821_),
    .B(_05822_),
    .Y(_05823_));
 BUFx6f_ASAP7_75t_R _28634_ (.A(_05823_),
    .Y(_16031_));
 NAND2x2_ASAP7_75t_R _28635_ (.A(_05752_),
    .B(_05735_),
    .Y(_05824_));
 XOR2x2_ASAP7_75t_R _28636_ (.A(_05767_),
    .B(_01052_),
    .Y(_05825_));
 NOR2x2_ASAP7_75t_R _28637_ (.A(_05825_),
    .B(net459),
    .Y(_05826_));
 OAI21x1_ASAP7_75t_R _28638_ (.A1(net29),
    .A2(_05824_),
    .B(_05826_),
    .Y(_05827_));
 BUFx6f_ASAP7_75t_R _28639_ (.A(_05825_),
    .Y(_05828_));
 BUFx6f_ASAP7_75t_R _28640_ (.A(_05828_),
    .Y(_05829_));
 INVx1_ASAP7_75t_R _28641_ (.A(_05781_),
    .Y(_05830_));
 OAI21x1_ASAP7_75t_R _28642_ (.A1(_05749_),
    .A2(_05830_),
    .B(_00631_),
    .Y(_05831_));
 OAI21x1_ASAP7_75t_R _28643_ (.A1(_05788_),
    .A2(_16043_),
    .B(_05831_),
    .Y(_05832_));
 AOI21x1_ASAP7_75t_R _28644_ (.A1(_05829_),
    .A2(_05832_),
    .B(_05779_),
    .Y(_05833_));
 NAND2x1_ASAP7_75t_R _28645_ (.A(_05827_),
    .B(_05833_),
    .Y(_05834_));
 NAND2x2_ASAP7_75t_R _28646_ (.A(_16030_),
    .B(net29),
    .Y(_05835_));
 BUFx6f_ASAP7_75t_R _28647_ (.A(_05760_),
    .Y(_05836_));
 AOI21x1_ASAP7_75t_R _28648_ (.A1(_05836_),
    .A2(_16035_),
    .B(_05828_),
    .Y(_05837_));
 NAND2x2_ASAP7_75t_R _28649_ (.A(_05835_),
    .B(_05837_),
    .Y(_05838_));
 AOI21x1_ASAP7_75t_R _28650_ (.A1(_16030_),
    .A2(_05797_),
    .B(_05769_),
    .Y(_05839_));
 AOI21x1_ASAP7_75t_R _28651_ (.A1(_05824_),
    .A2(_05839_),
    .B(_05794_),
    .Y(_05840_));
 BUFx6f_ASAP7_75t_R _28652_ (.A(_05818_),
    .Y(_05841_));
 AOI21x1_ASAP7_75t_R _28653_ (.A1(_05838_),
    .A2(_05840_),
    .B(_05841_),
    .Y(_05842_));
 XOR2x1_ASAP7_75t_R _28654_ (.A(_00745_),
    .Y(_05843_),
    .B(_00746_));
 XOR2x1_ASAP7_75t_R _28655_ (.A(_05843_),
    .Y(_05844_),
    .B(_11485_));
 XOR2x2_ASAP7_75t_R _28656_ (.A(_05844_),
    .B(_11497_),
    .Y(_05845_));
 NOR2x1_ASAP7_75t_R _28657_ (.A(_10787_),
    .B(_00663_),
    .Y(_05846_));
 AO21x1_ASAP7_75t_R _28658_ (.A1(_05845_),
    .A2(_10786_),
    .B(_05846_),
    .Y(_05847_));
 XOR2x2_ASAP7_75t_R _28659_ (.A(_05847_),
    .B(_01055_),
    .Y(_05848_));
 INVx2_ASAP7_75t_R _28660_ (.A(_05848_),
    .Y(_05849_));
 AOI21x1_ASAP7_75t_R _28661_ (.A1(_05834_),
    .A2(_05842_),
    .B(_05849_),
    .Y(_05850_));
 OAI21x1_ASAP7_75t_R _28662_ (.A1(_05792_),
    .A2(_05820_),
    .B(_05850_),
    .Y(_05851_));
 INVx2_ASAP7_75t_R _28663_ (.A(_01258_),
    .Y(_05852_));
 AO21x1_ASAP7_75t_R _28664_ (.A1(_05781_),
    .A2(_05782_),
    .B(_05852_),
    .Y(_05853_));
 BUFx4f_ASAP7_75t_R _28665_ (.A(_05853_),
    .Y(_05854_));
 BUFx6f_ASAP7_75t_R _28666_ (.A(_05793_),
    .Y(_05855_));
 AOI21x1_ASAP7_75t_R _28667_ (.A1(_05854_),
    .A2(_05786_),
    .B(_05855_),
    .Y(_05856_));
 NOR2x2_ASAP7_75t_R _28668_ (.A(_05828_),
    .B(_05797_),
    .Y(_05857_));
 AOI21x1_ASAP7_75t_R _28669_ (.A1(_05752_),
    .A2(net522),
    .B(_05825_),
    .Y(_05858_));
 NAND2x2_ASAP7_75t_R _28670_ (.A(_05760_),
    .B(net522),
    .Y(_05859_));
 OAI21x1_ASAP7_75t_R _28671_ (.A1(_05857_),
    .A2(_05858_),
    .B(_05859_),
    .Y(_05860_));
 NAND2x1_ASAP7_75t_R _28672_ (.A(_05856_),
    .B(_05860_),
    .Y(_05861_));
 NOR2x1_ASAP7_75t_R _28673_ (.A(_05779_),
    .B(_05858_),
    .Y(_05862_));
 NAND2x2_ASAP7_75t_R _28674_ (.A(_05752_),
    .B(net523),
    .Y(_05863_));
 INVx2_ASAP7_75t_R _28675_ (.A(_01256_),
    .Y(_05864_));
 AOI21x1_ASAP7_75t_R _28676_ (.A1(_05757_),
    .A2(_05759_),
    .B(_05864_),
    .Y(_05865_));
 NOR2x2_ASAP7_75t_R _28677_ (.A(_05769_),
    .B(_05865_),
    .Y(_05866_));
 OAI21x1_ASAP7_75t_R _28678_ (.A1(net29),
    .A2(_05863_),
    .B(_05866_),
    .Y(_05867_));
 AOI21x1_ASAP7_75t_R _28679_ (.A1(_05862_),
    .A2(_05867_),
    .B(_05841_),
    .Y(_05868_));
 BUFx10_ASAP7_75t_R _28680_ (.A(_05848_),
    .Y(_05869_));
 AOI21x1_ASAP7_75t_R _28681_ (.A1(_05861_),
    .A2(_05868_),
    .B(_05869_),
    .Y(_05870_));
 AOI21x1_ASAP7_75t_R _28682_ (.A1(_05757_),
    .A2(_05759_),
    .B(_05852_),
    .Y(_05871_));
 AOI21x1_ASAP7_75t_R _28683_ (.A1(net30),
    .A2(_16043_),
    .B(_05871_),
    .Y(_05872_));
 OAI21x1_ASAP7_75t_R _28684_ (.A1(_05770_),
    .A2(_05872_),
    .B(_05779_),
    .Y(_05873_));
 BUFx10_ASAP7_75t_R _28685_ (.A(_05768_),
    .Y(_05874_));
 OAI21x1_ASAP7_75t_R _28686_ (.A1(_05796_),
    .A2(_16031_),
    .B(_05874_),
    .Y(_05875_));
 NAND2x2_ASAP7_75t_R _28687_ (.A(_05752_),
    .B(net515),
    .Y(_05876_));
 NAND2x1_ASAP7_75t_R _28688_ (.A(_05824_),
    .B(_05876_),
    .Y(_05877_));
 NOR2x1_ASAP7_75t_R _28689_ (.A(_05875_),
    .B(_05877_),
    .Y(_05878_));
 NOR2x1_ASAP7_75t_R _28690_ (.A(_05873_),
    .B(_05878_),
    .Y(_05879_));
 INVx2_ASAP7_75t_R _28691_ (.A(_01255_),
    .Y(_05880_));
 NAND3x2_ASAP7_75t_R _28692_ (.B(_05750_),
    .C(_05880_),
    .Y(_05881_),
    .A(_05751_));
 OAI21x1_ASAP7_75t_R _28693_ (.A1(_16033_),
    .A2(_16040_),
    .B(_05881_),
    .Y(_05882_));
 NAND2x1_ASAP7_75t_R _28694_ (.A(_05770_),
    .B(_05882_),
    .Y(_05883_));
 AOI21x1_ASAP7_75t_R _28695_ (.A1(_05796_),
    .A2(_16030_),
    .B(_05769_),
    .Y(_05884_));
 NAND3x2_ASAP7_75t_R _28696_ (.B(_16035_),
    .C(_05836_),
    .Y(_05885_),
    .A(_05797_));
 NAND2x1_ASAP7_75t_R _28697_ (.A(_05884_),
    .B(_05885_),
    .Y(_05886_));
 BUFx6f_ASAP7_75t_R _28698_ (.A(_05778_),
    .Y(_05887_));
 BUFx6f_ASAP7_75t_R _28699_ (.A(_05887_),
    .Y(_05888_));
 AOI21x1_ASAP7_75t_R _28700_ (.A1(_05883_),
    .A2(_05886_),
    .B(_05888_),
    .Y(_05889_));
 OAI21x1_ASAP7_75t_R _28701_ (.A1(_05879_),
    .A2(_05889_),
    .B(_05819_),
    .Y(_05890_));
 XOR2x1_ASAP7_75t_R _28702_ (.A(_00746_),
    .Y(_05891_),
    .B(_11363_));
 XOR2x1_ASAP7_75t_R _28703_ (.A(_05891_),
    .Y(_05892_),
    .B(_00842_));
 XOR2x1_ASAP7_75t_R _28704_ (.A(_05892_),
    .Y(_05893_),
    .B(_11540_));
 NOR2x1_ASAP7_75t_R _28705_ (.A(_13017_),
    .B(_00662_),
    .Y(_05894_));
 AO21x1_ASAP7_75t_R _28706_ (.A1(_05893_),
    .A2(_10831_),
    .B(_05894_),
    .Y(_05895_));
 XOR2x2_ASAP7_75t_R _28707_ (.A(_05895_),
    .B(_01056_),
    .Y(_05896_));
 CKINVDCx8_ASAP7_75t_R _28708_ (.A(_05896_),
    .Y(_05897_));
 AOI21x1_ASAP7_75t_R _28709_ (.A1(_05870_),
    .A2(_05890_),
    .B(_05897_),
    .Y(_05898_));
 NAND2x1_ASAP7_75t_R _28710_ (.A(_05851_),
    .B(_05898_),
    .Y(_05899_));
 BUFx6f_ASAP7_75t_R _28711_ (.A(_05778_),
    .Y(_05900_));
 BUFx10_ASAP7_75t_R _28712_ (.A(_05900_),
    .Y(_05901_));
 NOR2x2_ASAP7_75t_R _28713_ (.A(net29),
    .B(_05859_),
    .Y(_05902_));
 INVx1_ASAP7_75t_R _28714_ (.A(_01257_),
    .Y(_05903_));
 OA21x2_ASAP7_75t_R _28715_ (.A1(_05836_),
    .A2(_05903_),
    .B(_05828_),
    .Y(_05904_));
 INVx1_ASAP7_75t_R _28716_ (.A(_05904_),
    .Y(_05905_));
 INVx2_ASAP7_75t_R _28717_ (.A(_05881_),
    .Y(_05906_));
 NAND2x1_ASAP7_75t_R _28718_ (.A(_05770_),
    .B(_05906_),
    .Y(_05907_));
 OAI21x1_ASAP7_75t_R _28719_ (.A1(_05902_),
    .A2(_05905_),
    .B(_05907_),
    .Y(_05908_));
 NAND2x2_ASAP7_75t_R _28720_ (.A(net522),
    .B(_05716_),
    .Y(_05909_));
 BUFx6f_ASAP7_75t_R _28721_ (.A(_05825_),
    .Y(_05910_));
 AOI21x1_ASAP7_75t_R _28722_ (.A1(_05788_),
    .A2(_05796_),
    .B(_05910_),
    .Y(_05911_));
 OAI21x1_ASAP7_75t_R _28723_ (.A1(_16043_),
    .A2(_05909_),
    .B(_05911_),
    .Y(_05912_));
 BUFx6f_ASAP7_75t_R _28724_ (.A(_05769_),
    .Y(_05913_));
 OA21x2_ASAP7_75t_R _28725_ (.A1(_05881_),
    .A2(_05913_),
    .B(_05887_),
    .Y(_05914_));
 BUFx6f_ASAP7_75t_R _28726_ (.A(_05818_),
    .Y(_05915_));
 AOI21x1_ASAP7_75t_R _28727_ (.A1(_05912_),
    .A2(_05914_),
    .B(_05915_),
    .Y(_05916_));
 OAI21x1_ASAP7_75t_R _28728_ (.A1(_05901_),
    .A2(_05908_),
    .B(_05916_),
    .Y(_05917_));
 AOI21x1_ASAP7_75t_R _28729_ (.A1(_05782_),
    .A2(_05751_),
    .B(_01256_),
    .Y(_05918_));
 INVx1_ASAP7_75t_R _28730_ (.A(_05918_),
    .Y(_05919_));
 OA21x2_ASAP7_75t_R _28731_ (.A1(net514),
    .A2(_16035_),
    .B(_05836_),
    .Y(_05920_));
 INVx1_ASAP7_75t_R _28732_ (.A(_05920_),
    .Y(_05921_));
 BUFx6f_ASAP7_75t_R _28733_ (.A(_05910_),
    .Y(_05922_));
 AOI21x1_ASAP7_75t_R _28734_ (.A1(_05919_),
    .A2(_05921_),
    .B(_05922_),
    .Y(_05923_));
 NOR2x1_ASAP7_75t_R _28735_ (.A(_01255_),
    .B(_05760_),
    .Y(_05924_));
 AOI21x1_ASAP7_75t_R _28736_ (.A1(_05770_),
    .A2(_05924_),
    .B(_05779_),
    .Y(_05925_));
 AO21x2_ASAP7_75t_R _28737_ (.A1(_05759_),
    .A2(_05757_),
    .B(_00631_),
    .Y(_05926_));
 NAND2x1_ASAP7_75t_R _28738_ (.A(_05926_),
    .B(_05884_),
    .Y(_05927_));
 NAND2x1_ASAP7_75t_R _28739_ (.A(_05925_),
    .B(_05927_),
    .Y(_05928_));
 BUFx6f_ASAP7_75t_R _28740_ (.A(_05887_),
    .Y(_05929_));
 INVx1_ASAP7_75t_R _28741_ (.A(_01260_),
    .Y(_05930_));
 BUFx6f_ASAP7_75t_R _28742_ (.A(_05874_),
    .Y(_05931_));
 AOI21x1_ASAP7_75t_R _28743_ (.A1(_05750_),
    .A2(_05751_),
    .B(net496),
    .Y(_05932_));
 NOR2x2_ASAP7_75t_R _28744_ (.A(_05825_),
    .B(net595),
    .Y(_05933_));
 INVx2_ASAP7_75t_R _28745_ (.A(_05933_),
    .Y(_05934_));
 OAI21x1_ASAP7_75t_R _28746_ (.A1(_05930_),
    .A2(_05931_),
    .B(_05934_),
    .Y(_05935_));
 BUFx10_ASAP7_75t_R _28747_ (.A(_05817_),
    .Y(_05936_));
 AOI21x1_ASAP7_75t_R _28748_ (.A1(_05929_),
    .A2(_05935_),
    .B(_05936_),
    .Y(_05937_));
 OAI21x1_ASAP7_75t_R _28749_ (.A1(_05923_),
    .A2(_05928_),
    .B(_05937_),
    .Y(_05938_));
 BUFx10_ASAP7_75t_R _28750_ (.A(_05849_),
    .Y(_05939_));
 AOI21x1_ASAP7_75t_R _28751_ (.A1(_05917_),
    .A2(_05938_),
    .B(_05939_),
    .Y(_05940_));
 NOR2x2_ASAP7_75t_R _28752_ (.A(_01257_),
    .B(_05796_),
    .Y(_05941_));
 BUFx6f_ASAP7_75t_R _28753_ (.A(_05769_),
    .Y(_05942_));
 OAI21x1_ASAP7_75t_R _28754_ (.A1(_05918_),
    .A2(_05941_),
    .B(_05942_),
    .Y(_05943_));
 INVx3_ASAP7_75t_R _28755_ (.A(_05786_),
    .Y(_05944_));
 NAND3x1_ASAP7_75t_R _28756_ (.A(_05944_),
    .B(_05900_),
    .C(_05943_),
    .Y(_05945_));
 NAND2x1_ASAP7_75t_R _28757_ (.A(_05769_),
    .B(_05918_),
    .Y(_05946_));
 AND2x2_ASAP7_75t_R _28758_ (.A(_05946_),
    .B(_05794_),
    .Y(_05947_));
 AOI21x1_ASAP7_75t_R _28759_ (.A1(_05947_),
    .A2(_05886_),
    .B(_05936_),
    .Y(_05948_));
 NAND2x1_ASAP7_75t_R _28760_ (.A(_05945_),
    .B(_05948_),
    .Y(_05949_));
 BUFx6f_ASAP7_75t_R _28761_ (.A(_05817_),
    .Y(_05950_));
 BUFx10_ASAP7_75t_R _28762_ (.A(_05950_),
    .Y(_05951_));
 NAND2x2_ASAP7_75t_R _28763_ (.A(_05760_),
    .B(_05735_),
    .Y(_05952_));
 AO21x1_ASAP7_75t_R _28764_ (.A1(_05952_),
    .A2(_05789_),
    .B(_05942_),
    .Y(_05953_));
 INVx2_ASAP7_75t_R _28765_ (.A(net595),
    .Y(_05954_));
 AOI21x1_ASAP7_75t_R _28766_ (.A1(_16040_),
    .A2(_05797_),
    .B(_05910_),
    .Y(_05955_));
 AOI21x1_ASAP7_75t_R _28767_ (.A1(_05954_),
    .A2(_05955_),
    .B(_05900_),
    .Y(_05956_));
 OAI21x1_ASAP7_75t_R _28768_ (.A1(_05874_),
    .A2(_05865_),
    .B(_05887_),
    .Y(_05957_));
 AOI21x1_ASAP7_75t_R _28769_ (.A1(_05831_),
    .A2(_05881_),
    .B(_05910_),
    .Y(_05958_));
 NOR2x1_ASAP7_75t_R _28770_ (.A(_05957_),
    .B(_05958_),
    .Y(_05959_));
 AOI21x1_ASAP7_75t_R _28771_ (.A1(_05953_),
    .A2(_05956_),
    .B(_05959_),
    .Y(_05960_));
 NAND2x1_ASAP7_75t_R _28772_ (.A(_05951_),
    .B(_05960_),
    .Y(_05961_));
 BUFx10_ASAP7_75t_R _28773_ (.A(_05848_),
    .Y(_05962_));
 AOI21x1_ASAP7_75t_R _28774_ (.A1(_05949_),
    .A2(_05961_),
    .B(_05962_),
    .Y(_05963_));
 OAI21x1_ASAP7_75t_R _28775_ (.A1(_05940_),
    .A2(_05963_),
    .B(_05897_),
    .Y(_05964_));
 NAND2x1_ASAP7_75t_R _28776_ (.A(_05899_),
    .B(_05964_),
    .Y(_00136_));
 NOR2x2_ASAP7_75t_R _28777_ (.A(_16040_),
    .B(net29),
    .Y(_05965_));
 OAI21x1_ASAP7_75t_R _28778_ (.A1(_16043_),
    .A2(net30),
    .B(_05913_),
    .Y(_05966_));
 NOR2x1_ASAP7_75t_R _28779_ (.A(_05965_),
    .B(_05966_),
    .Y(_05967_));
 BUFx6f_ASAP7_75t_R _28780_ (.A(_05817_),
    .Y(_05968_));
 AOI211x1_ASAP7_75t_R _28781_ (.A1(_05866_),
    .A2(_05876_),
    .B(_05967_),
    .C(_05968_),
    .Y(_05969_));
 INVx2_ASAP7_75t_R _28782_ (.A(_05859_),
    .Y(_05970_));
 NAND2x1_ASAP7_75t_R _28783_ (.A(_05942_),
    .B(_05783_),
    .Y(_05971_));
 OAI21x1_ASAP7_75t_R _28784_ (.A1(_05970_),
    .A2(_05971_),
    .B(_05968_),
    .Y(_05972_));
 AOI21x1_ASAP7_75t_R _28785_ (.A1(_16035_),
    .A2(_05716_),
    .B(_05752_),
    .Y(_05973_));
 INVx2_ASAP7_75t_R _28786_ (.A(_05973_),
    .Y(_05974_));
 AO21x1_ASAP7_75t_R _28787_ (.A1(_05797_),
    .A2(net30),
    .B(_05836_),
    .Y(_05975_));
 BUFx6f_ASAP7_75t_R _28788_ (.A(_05874_),
    .Y(_05976_));
 AOI21x1_ASAP7_75t_R _28789_ (.A1(_05974_),
    .A2(_05975_),
    .B(_05976_),
    .Y(_05977_));
 OAI21x1_ASAP7_75t_R _28790_ (.A1(_05972_),
    .A2(_05977_),
    .B(_05901_),
    .Y(_05978_));
 NOR2x1_ASAP7_75t_R _28791_ (.A(_05969_),
    .B(_05978_),
    .Y(_05979_));
 INVx1_ASAP7_75t_R _28792_ (.A(_00633_),
    .Y(_05980_));
 OR3x1_ASAP7_75t_R _28793_ (.A(_05950_),
    .B(_05980_),
    .C(_05942_),
    .Y(_05981_));
 NAND2x2_ASAP7_75t_R _28794_ (.A(_16035_),
    .B(_05797_),
    .Y(_05982_));
 OAI21x1_ASAP7_75t_R _28795_ (.A1(_16043_),
    .A2(_05982_),
    .B(_05911_),
    .Y(_05983_));
 AO21x1_ASAP7_75t_R _28796_ (.A1(_05981_),
    .A2(_05983_),
    .B(_05929_),
    .Y(_05984_));
 NAND2x1_ASAP7_75t_R _28797_ (.A(_05869_),
    .B(_05984_),
    .Y(_05985_));
 OAI21x1_ASAP7_75t_R _28798_ (.A1(_05979_),
    .A2(_05985_),
    .B(_05896_),
    .Y(_05986_));
 AOI221x1_ASAP7_75t_R _28799_ (.A1(_05876_),
    .A2(_05866_),
    .B1(_05783_),
    .B2(_05837_),
    .C(_05819_),
    .Y(_05987_));
 INVx4_ASAP7_75t_R _28800_ (.A(net459),
    .Y(_05988_));
 BUFx6f_ASAP7_75t_R _28801_ (.A(_05828_),
    .Y(_05989_));
 AO21x1_ASAP7_75t_R _28802_ (.A1(_05988_),
    .A2(_05989_),
    .B(_05950_),
    .Y(_05990_));
 OA21x2_ASAP7_75t_R _28803_ (.A1(_16043_),
    .A2(_05982_),
    .B(_05858_),
    .Y(_05991_));
 OAI21x1_ASAP7_75t_R _28804_ (.A1(_05990_),
    .A2(_05991_),
    .B(_05795_),
    .Y(_05992_));
 OAI21x1_ASAP7_75t_R _28805_ (.A1(_05987_),
    .A2(_05992_),
    .B(_05939_),
    .Y(_05993_));
 NAND2x1_ASAP7_75t_R _28806_ (.A(_05926_),
    .B(_05803_),
    .Y(_05994_));
 NOR2x2_ASAP7_75t_R _28807_ (.A(_05760_),
    .B(net524),
    .Y(_05995_));
 AO21x1_ASAP7_75t_R _28808_ (.A1(_05906_),
    .A2(_05931_),
    .B(_05841_),
    .Y(_05996_));
 AOI21x1_ASAP7_75t_R _28809_ (.A1(_05976_),
    .A2(_05995_),
    .B(_05996_),
    .Y(_05997_));
 NOR2x2_ASAP7_75t_R _28810_ (.A(_05910_),
    .B(_05871_),
    .Y(_05998_));
 AO21x2_ASAP7_75t_R _28811_ (.A1(_05781_),
    .A2(_05782_),
    .B(_05880_),
    .Y(_05999_));
 AO21x1_ASAP7_75t_R _28812_ (.A1(_05998_),
    .A2(_05999_),
    .B(_05950_),
    .Y(_06000_));
 AO21x2_ASAP7_75t_R _28813_ (.A1(_05797_),
    .A2(_16035_),
    .B(_16040_),
    .Y(_06001_));
 AOI21x1_ASAP7_75t_R _28814_ (.A1(_05988_),
    .A2(_06001_),
    .B(_05931_),
    .Y(_06002_));
 OAI21x1_ASAP7_75t_R _28815_ (.A1(_06000_),
    .A2(_06002_),
    .B(_05901_),
    .Y(_06003_));
 AOI21x1_ASAP7_75t_R _28816_ (.A1(_05994_),
    .A2(_05997_),
    .B(_06003_),
    .Y(_06004_));
 NOR2x1_ASAP7_75t_R _28817_ (.A(_05993_),
    .B(_06004_),
    .Y(_06005_));
 INVx2_ASAP7_75t_R _28818_ (.A(_05871_),
    .Y(_06006_));
 AO21x1_ASAP7_75t_R _28819_ (.A1(_05803_),
    .A2(_06006_),
    .B(_05888_),
    .Y(_06007_));
 AOI21x1_ASAP7_75t_R _28820_ (.A1(_05829_),
    .A2(_05798_),
    .B(_05794_),
    .Y(_06008_));
 NAND2x2_ASAP7_75t_R _28821_ (.A(_05760_),
    .B(net514),
    .Y(_06009_));
 BUFx6f_ASAP7_75t_R _28822_ (.A(_06009_),
    .Y(_06010_));
 AND2x2_ASAP7_75t_R _28823_ (.A(_05946_),
    .B(_06010_),
    .Y(_06011_));
 AOI21x1_ASAP7_75t_R _28824_ (.A1(_06008_),
    .A2(_06011_),
    .B(_05968_),
    .Y(_06012_));
 OA21x2_ASAP7_75t_R _28825_ (.A1(_05923_),
    .A2(_06007_),
    .B(_06012_),
    .Y(_06013_));
 BUFx6f_ASAP7_75t_R _28826_ (.A(_05825_),
    .Y(_06014_));
 AO21x1_ASAP7_75t_R _28827_ (.A1(_16040_),
    .A2(net563),
    .B(_06014_),
    .Y(_06015_));
 BUFx6f_ASAP7_75t_R _28828_ (.A(_05793_),
    .Y(_06016_));
 AOI21x1_ASAP7_75t_R _28829_ (.A1(_05863_),
    .A2(_05786_),
    .B(_06016_),
    .Y(_06017_));
 OA21x2_ASAP7_75t_R _28830_ (.A1(_05995_),
    .A2(_06015_),
    .B(_06017_),
    .Y(_06018_));
 NAND2x1_ASAP7_75t_R _28831_ (.A(_05835_),
    .B(_05955_),
    .Y(_06019_));
 INVx1_ASAP7_75t_R _28832_ (.A(_06019_),
    .Y(_06020_));
 NOR2x2_ASAP7_75t_R _28833_ (.A(_05760_),
    .B(_05769_),
    .Y(_06021_));
 AO21x1_ASAP7_75t_R _28834_ (.A1(_05909_),
    .A2(_06021_),
    .B(_05888_),
    .Y(_06022_));
 OAI21x1_ASAP7_75t_R _28835_ (.A1(_06020_),
    .A2(_06022_),
    .B(_05951_),
    .Y(_06023_));
 OAI21x1_ASAP7_75t_R _28836_ (.A1(_06018_),
    .A2(_06023_),
    .B(_05962_),
    .Y(_06024_));
 OAI21x1_ASAP7_75t_R _28837_ (.A1(_06013_),
    .A2(_06024_),
    .B(_05897_),
    .Y(_06025_));
 NOR2x2_ASAP7_75t_R _28838_ (.A(net563),
    .B(_05796_),
    .Y(_06026_));
 AO21x1_ASAP7_75t_R _28839_ (.A1(_06026_),
    .A2(_05931_),
    .B(_05900_),
    .Y(_06027_));
 NOR2x1_ASAP7_75t_R _28840_ (.A(_06027_),
    .B(_06002_),
    .Y(_06028_));
 NOR2x1_ASAP7_75t_R _28841_ (.A(_05922_),
    .B(_05974_),
    .Y(_06029_));
 INVx1_ASAP7_75t_R _28842_ (.A(_06010_),
    .Y(_06030_));
 NAND2x1_ASAP7_75t_R _28843_ (.A(_05829_),
    .B(_05854_),
    .Y(_06031_));
 OAI21x1_ASAP7_75t_R _28844_ (.A1(_06030_),
    .A2(_06031_),
    .B(_05888_),
    .Y(_06032_));
 OAI21x1_ASAP7_75t_R _28845_ (.A1(_06029_),
    .A2(_06032_),
    .B(_05951_),
    .Y(_06033_));
 OAI21x1_ASAP7_75t_R _28846_ (.A1(_06028_),
    .A2(_06033_),
    .B(_05939_),
    .Y(_06034_));
 AO21x1_ASAP7_75t_R _28847_ (.A1(_05933_),
    .A2(_05859_),
    .B(_05900_),
    .Y(_06035_));
 OA21x2_ASAP7_75t_R _28848_ (.A1(_16033_),
    .A2(net30),
    .B(_05884_),
    .Y(_06036_));
 OAI21x1_ASAP7_75t_R _28849_ (.A1(_06035_),
    .A2(_06036_),
    .B(_05819_),
    .Y(_06037_));
 AO21x1_ASAP7_75t_R _28850_ (.A1(_16035_),
    .A2(_05796_),
    .B(_05828_),
    .Y(_06038_));
 NOR2x1_ASAP7_75t_R _28851_ (.A(_05773_),
    .B(_06038_),
    .Y(_06039_));
 NOR2x1p5_ASAP7_75t_R _28852_ (.A(_05918_),
    .B(_05944_),
    .Y(_06040_));
 OA21x2_ASAP7_75t_R _28853_ (.A1(_06040_),
    .A2(_06039_),
    .B(_05929_),
    .Y(_06041_));
 NOR2x1_ASAP7_75t_R _28854_ (.A(_06037_),
    .B(_06041_),
    .Y(_06042_));
 NOR2x1_ASAP7_75t_R _28855_ (.A(_06034_),
    .B(_06042_),
    .Y(_06043_));
 OAI22x1_ASAP7_75t_R _28856_ (.A1(_05986_),
    .A2(_06005_),
    .B1(_06043_),
    .B2(_06025_),
    .Y(_00137_));
 AO21x1_ASAP7_75t_R _28857_ (.A1(_05798_),
    .A2(_05988_),
    .B(_05922_),
    .Y(_06044_));
 INVx1_ASAP7_75t_R _28858_ (.A(_05924_),
    .Y(_06045_));
 NAND3x1_ASAP7_75t_R _28859_ (.A(_06045_),
    .B(_05952_),
    .C(_05922_),
    .Y(_06046_));
 AOI21x1_ASAP7_75t_R _28860_ (.A1(_06044_),
    .A2(_06046_),
    .B(_05795_),
    .Y(_06047_));
 BUFx6f_ASAP7_75t_R _28861_ (.A(_05794_),
    .Y(_06048_));
 NOR2x2_ASAP7_75t_R _28862_ (.A(_05857_),
    .B(_05858_),
    .Y(_06049_));
 NAND2x1_ASAP7_75t_R _28863_ (.A(_06048_),
    .B(_06049_),
    .Y(_06050_));
 AOI211x1_ASAP7_75t_R _28864_ (.A1(_05995_),
    .A2(_16033_),
    .B(_05871_),
    .C(_05976_),
    .Y(_06051_));
 OAI21x1_ASAP7_75t_R _28865_ (.A1(_06050_),
    .A2(_06051_),
    .B(_05951_),
    .Y(_06052_));
 OAI21x1_ASAP7_75t_R _28866_ (.A1(_06047_),
    .A2(_06052_),
    .B(_05962_),
    .Y(_06053_));
 NOR2x1_ASAP7_75t_R _28867_ (.A(_05913_),
    .B(_16033_),
    .Y(_06054_));
 AOI21x1_ASAP7_75t_R _28868_ (.A1(_06021_),
    .A2(_05909_),
    .B(_06054_),
    .Y(_06055_));
 NOR2x2_ASAP7_75t_R _28869_ (.A(_01258_),
    .B(_05836_),
    .Y(_06056_));
 OAI21x1_ASAP7_75t_R _28870_ (.A1(_06026_),
    .A2(_06056_),
    .B(_05931_),
    .Y(_06057_));
 AO21x1_ASAP7_75t_R _28871_ (.A1(_06055_),
    .A2(_06057_),
    .B(_05795_),
    .Y(_06058_));
 NOR2x1_ASAP7_75t_R _28872_ (.A(_05874_),
    .B(_05918_),
    .Y(_06059_));
 AOI21x1_ASAP7_75t_R _28873_ (.A1(_06059_),
    .A2(_05921_),
    .B(_05888_),
    .Y(_06060_));
 OAI21x1_ASAP7_75t_R _28874_ (.A1(net595),
    .A2(_05875_),
    .B(_06060_),
    .Y(_06061_));
 AOI21x1_ASAP7_75t_R _28875_ (.A1(_06058_),
    .A2(_06061_),
    .B(_05951_),
    .Y(_06062_));
 OAI21x1_ASAP7_75t_R _28876_ (.A1(_06053_),
    .A2(_06062_),
    .B(_05896_),
    .Y(_06063_));
 NAND2x1_ASAP7_75t_R _28877_ (.A(_06016_),
    .B(_05943_),
    .Y(_06064_));
 AO21x2_ASAP7_75t_R _28878_ (.A1(_05781_),
    .A2(_05782_),
    .B(_05864_),
    .Y(_06065_));
 AND3x1_ASAP7_75t_R _28879_ (.A(_06010_),
    .B(_05989_),
    .C(_06065_),
    .Y(_06066_));
 OAI21x1_ASAP7_75t_R _28880_ (.A1(_06064_),
    .A2(_06066_),
    .B(_05819_),
    .Y(_06067_));
 AO21x2_ASAP7_75t_R _28881_ (.A1(_05759_),
    .A2(_05757_),
    .B(_01257_),
    .Y(_06068_));
 AO21x2_ASAP7_75t_R _28882_ (.A1(_05781_),
    .A2(_05782_),
    .B(_01258_),
    .Y(_06069_));
 AND3x1_ASAP7_75t_R _28883_ (.A(_06068_),
    .B(_06069_),
    .C(_05942_),
    .Y(_06070_));
 AND2x2_ASAP7_75t_R _28884_ (.A(_06059_),
    .B(_05952_),
    .Y(_06071_));
 OA21x2_ASAP7_75t_R _28885_ (.A1(_06070_),
    .A2(_06071_),
    .B(_05929_),
    .Y(_06072_));
 NOR2x1_ASAP7_75t_R _28886_ (.A(_06067_),
    .B(_06072_),
    .Y(_06073_));
 AOI21x1_ASAP7_75t_R _28887_ (.A1(_06069_),
    .A2(_05952_),
    .B(_05922_),
    .Y(_06074_));
 AOI21x1_ASAP7_75t_R _28888_ (.A1(_06068_),
    .A2(_05876_),
    .B(_05976_),
    .Y(_06075_));
 OAI21x1_ASAP7_75t_R _28889_ (.A1(_06074_),
    .A2(_06075_),
    .B(_05901_),
    .Y(_06076_));
 AOI21x1_ASAP7_75t_R _28890_ (.A1(_01257_),
    .A2(_05796_),
    .B(_05828_),
    .Y(_06077_));
 INVx2_ASAP7_75t_R _28891_ (.A(_06077_),
    .Y(_06078_));
 NOR2x1_ASAP7_75t_R _28892_ (.A(_05970_),
    .B(_06078_),
    .Y(_06079_));
 AND3x1_ASAP7_75t_R _28893_ (.A(_05988_),
    .B(_05954_),
    .C(_05989_),
    .Y(_06080_));
 OAI21x1_ASAP7_75t_R _28894_ (.A1(_06079_),
    .A2(_06080_),
    .B(_05795_),
    .Y(_06081_));
 AOI21x1_ASAP7_75t_R _28895_ (.A1(_06076_),
    .A2(_06081_),
    .B(_05819_),
    .Y(_06082_));
 NOR3x1_ASAP7_75t_R _28896_ (.A(_06082_),
    .B(_06073_),
    .C(_05962_),
    .Y(_06083_));
 AND2x2_ASAP7_75t_R _28897_ (.A(_01256_),
    .B(_01255_),
    .Y(_06084_));
 AO21x2_ASAP7_75t_R _28898_ (.A1(_05759_),
    .A2(_05757_),
    .B(_06084_),
    .Y(_06085_));
 AOI21x1_ASAP7_75t_R _28899_ (.A1(_06085_),
    .A2(_06001_),
    .B(_05976_),
    .Y(_06086_));
 NAND2x1_ASAP7_75t_R _28900_ (.A(_05929_),
    .B(_05983_),
    .Y(_06087_));
 NAND2x1_ASAP7_75t_R _28901_ (.A(_06065_),
    .B(_05786_),
    .Y(_06088_));
 AOI21x1_ASAP7_75t_R _28902_ (.A1(_06088_),
    .A2(_05780_),
    .B(_05915_),
    .Y(_06089_));
 OAI21x1_ASAP7_75t_R _28903_ (.A1(_06086_),
    .A2(_06087_),
    .B(_06089_),
    .Y(_06090_));
 NAND2x1_ASAP7_75t_R _28904_ (.A(_00634_),
    .B(_06014_),
    .Y(_06091_));
 NAND2x1_ASAP7_75t_R _28905_ (.A(_06091_),
    .B(_06049_),
    .Y(_06092_));
 OA21x2_ASAP7_75t_R _28906_ (.A1(_01262_),
    .A2(_05829_),
    .B(_05779_),
    .Y(_06093_));
 AOI21x1_ASAP7_75t_R _28907_ (.A1(_06093_),
    .A2(_06055_),
    .B(_05968_),
    .Y(_06094_));
 OAI21x1_ASAP7_75t_R _28908_ (.A1(_05901_),
    .A2(_06092_),
    .B(_06094_),
    .Y(_06095_));
 AOI21x1_ASAP7_75t_R _28909_ (.A1(_06090_),
    .A2(_06095_),
    .B(_05939_),
    .Y(_06096_));
 OAI21x1_ASAP7_75t_R _28910_ (.A1(_05796_),
    .A2(_16035_),
    .B(_05828_),
    .Y(_06097_));
 INVx1_ASAP7_75t_R _28911_ (.A(_05876_),
    .Y(_06098_));
 NOR2x1_ASAP7_75t_R _28912_ (.A(_06097_),
    .B(_06098_),
    .Y(_06099_));
 AO21x1_ASAP7_75t_R _28913_ (.A1(_05955_),
    .A2(_05954_),
    .B(_06016_),
    .Y(_06100_));
 OA21x2_ASAP7_75t_R _28914_ (.A1(_01260_),
    .A2(_05829_),
    .B(_05855_),
    .Y(_06101_));
 OAI21x1_ASAP7_75t_R _28915_ (.A1(net29),
    .A2(_05859_),
    .B(_05803_),
    .Y(_06102_));
 AOI21x1_ASAP7_75t_R _28916_ (.A1(_06101_),
    .A2(_06102_),
    .B(_05915_),
    .Y(_06103_));
 OAI21x1_ASAP7_75t_R _28917_ (.A1(_06099_),
    .A2(_06100_),
    .B(_06103_),
    .Y(_06104_));
 INVx1_ASAP7_75t_R _28918_ (.A(_05831_),
    .Y(_06105_));
 NOR2x1_ASAP7_75t_R _28919_ (.A(_06105_),
    .B(_05875_),
    .Y(_06106_));
 NOR2x2_ASAP7_75t_R _28920_ (.A(_05788_),
    .B(_16043_),
    .Y(_06107_));
 NOR3x1_ASAP7_75t_R _28921_ (.A(_06107_),
    .B(_05931_),
    .C(net595),
    .Y(_06108_));
 OAI21x1_ASAP7_75t_R _28922_ (.A1(_06106_),
    .A2(_06108_),
    .B(_05929_),
    .Y(_06109_));
 NAND2x2_ASAP7_75t_R _28923_ (.A(_05836_),
    .B(_05797_),
    .Y(_06110_));
 AOI21x1_ASAP7_75t_R _28924_ (.A1(net30),
    .A2(net29),
    .B(_05874_),
    .Y(_06111_));
 NOR2x1_ASAP7_75t_R _28925_ (.A(_05980_),
    .B(_06014_),
    .Y(_06112_));
 AOI21x1_ASAP7_75t_R _28926_ (.A1(_06110_),
    .A2(_06111_),
    .B(_06112_),
    .Y(_06113_));
 AOI21x1_ASAP7_75t_R _28927_ (.A1(_06048_),
    .A2(_06113_),
    .B(_05968_),
    .Y(_06114_));
 NAND2x1_ASAP7_75t_R _28928_ (.A(_06109_),
    .B(_06114_),
    .Y(_06115_));
 AOI21x1_ASAP7_75t_R _28929_ (.A1(_06104_),
    .A2(_06115_),
    .B(_05962_),
    .Y(_06116_));
 OAI21x1_ASAP7_75t_R _28930_ (.A1(_06096_),
    .A2(_06116_),
    .B(_05897_),
    .Y(_06117_));
 OAI21x1_ASAP7_75t_R _28931_ (.A1(_06063_),
    .A2(_06083_),
    .B(_06117_),
    .Y(_00138_));
 NAND2x1_ASAP7_75t_R _28932_ (.A(_16040_),
    .B(_05829_),
    .Y(_06118_));
 AOI21x1_ASAP7_75t_R _28933_ (.A1(_05952_),
    .A2(_05909_),
    .B(_05887_),
    .Y(_06119_));
 AOI21x1_ASAP7_75t_R _28934_ (.A1(_06118_),
    .A2(_06119_),
    .B(_05936_),
    .Y(_06120_));
 NAND2x1_ASAP7_75t_R _28935_ (.A(_05799_),
    .B(_06077_),
    .Y(_06121_));
 OA21x2_ASAP7_75t_R _28936_ (.A1(_05836_),
    .A2(_05852_),
    .B(_05910_),
    .Y(_06122_));
 AOI21x1_ASAP7_75t_R _28937_ (.A1(_06010_),
    .A2(_06122_),
    .B(_05855_),
    .Y(_06123_));
 NAND2x1_ASAP7_75t_R _28938_ (.A(_06121_),
    .B(_06123_),
    .Y(_06124_));
 AOI21x1_ASAP7_75t_R _28939_ (.A1(_06120_),
    .A2(_06124_),
    .B(_05869_),
    .Y(_06125_));
 OAI21x1_ASAP7_75t_R _28940_ (.A1(_05973_),
    .A2(_05934_),
    .B(_05855_),
    .Y(_06126_));
 AO21x1_ASAP7_75t_R _28941_ (.A1(_05836_),
    .A2(_00629_),
    .B(_05874_),
    .Y(_06127_));
 NOR2x1_ASAP7_75t_R _28942_ (.A(_06127_),
    .B(_05877_),
    .Y(_06128_));
 NOR2x1_ASAP7_75t_R _28943_ (.A(_06126_),
    .B(_06128_),
    .Y(_06129_));
 NAND2x1_ASAP7_75t_R _28944_ (.A(_05789_),
    .B(_05826_),
    .Y(_06130_));
 AND2x2_ASAP7_75t_R _28945_ (.A(_05840_),
    .B(_06130_),
    .Y(_06131_));
 OAI21x1_ASAP7_75t_R _28946_ (.A1(_06129_),
    .A2(_06131_),
    .B(_05951_),
    .Y(_06132_));
 NAND2x1_ASAP7_75t_R _28947_ (.A(_06125_),
    .B(_06132_),
    .Y(_06133_));
 AND3x1_ASAP7_75t_R _28948_ (.A(_06065_),
    .B(_06006_),
    .C(_05989_),
    .Y(_06134_));
 AO21x1_ASAP7_75t_R _28949_ (.A1(_05801_),
    .A2(_05876_),
    .B(_05841_),
    .Y(_06135_));
 NAND2x1_ASAP7_75t_R _28950_ (.A(_05876_),
    .B(_05786_),
    .Y(_06136_));
 AOI21x1_ASAP7_75t_R _28951_ (.A1(_05909_),
    .A2(_05837_),
    .B(_05950_),
    .Y(_06137_));
 AOI21x1_ASAP7_75t_R _28952_ (.A1(_06136_),
    .A2(_06137_),
    .B(_05888_),
    .Y(_06138_));
 OAI21x1_ASAP7_75t_R _28953_ (.A1(_06134_),
    .A2(_06135_),
    .B(_06138_),
    .Y(_06139_));
 NOR2x1_ASAP7_75t_R _28954_ (.A(_06107_),
    .B(_06038_),
    .Y(_06140_));
 AO21x1_ASAP7_75t_R _28955_ (.A1(_05803_),
    .A2(_05772_),
    .B(_05818_),
    .Y(_06141_));
 AOI21x1_ASAP7_75t_R _28956_ (.A1(_06014_),
    .A2(net871),
    .B(_05817_),
    .Y(_06142_));
 OAI21x1_ASAP7_75t_R _28957_ (.A1(_05965_),
    .A2(_05966_),
    .B(_06142_),
    .Y(_06143_));
 OAI21x1_ASAP7_75t_R _28958_ (.A1(_06140_),
    .A2(_06141_),
    .B(_06143_),
    .Y(_06144_));
 AOI21x1_ASAP7_75t_R _28959_ (.A1(_05901_),
    .A2(_06144_),
    .B(_05939_),
    .Y(_06145_));
 NAND2x1_ASAP7_75t_R _28960_ (.A(_06139_),
    .B(_06145_),
    .Y(_06146_));
 NAND2x1_ASAP7_75t_R _28961_ (.A(_06133_),
    .B(_06146_),
    .Y(_06147_));
 NAND2x1_ASAP7_75t_R _28962_ (.A(_05829_),
    .B(net871),
    .Y(_06148_));
 NAND2x1_ASAP7_75t_R _28963_ (.A(_06110_),
    .B(_05911_),
    .Y(_06149_));
 AOI21x1_ASAP7_75t_R _28964_ (.A1(_06148_),
    .A2(_06149_),
    .B(_05936_),
    .Y(_06150_));
 NAND2x2_ASAP7_75t_R _28965_ (.A(_05874_),
    .B(net459),
    .Y(_06151_));
 OAI21x1_ASAP7_75t_R _28966_ (.A1(_05841_),
    .A2(_06151_),
    .B(_05914_),
    .Y(_06152_));
 OAI21x1_ASAP7_75t_R _28967_ (.A1(_06150_),
    .A2(_06152_),
    .B(_05869_),
    .Y(_06153_));
 AO21x1_ASAP7_75t_R _28968_ (.A1(_06085_),
    .A2(_06069_),
    .B(_05913_),
    .Y(_06154_));
 AOI21x1_ASAP7_75t_R _28969_ (.A1(_05988_),
    .A2(_05858_),
    .B(_05950_),
    .Y(_06155_));
 NAND2x1_ASAP7_75t_R _28970_ (.A(_06154_),
    .B(_06155_),
    .Y(_06156_));
 OA21x2_ASAP7_75t_R _28971_ (.A1(_06068_),
    .A2(_05942_),
    .B(_05950_),
    .Y(_06157_));
 OAI21x1_ASAP7_75t_R _28972_ (.A1(_05970_),
    .A2(_06078_),
    .B(_06157_),
    .Y(_06158_));
 AOI21x1_ASAP7_75t_R _28973_ (.A1(_06156_),
    .A2(_06158_),
    .B(_05901_),
    .Y(_06159_));
 OAI21x1_ASAP7_75t_R _28974_ (.A1(_06153_),
    .A2(_06159_),
    .B(_05896_),
    .Y(_06160_));
 OA21x2_ASAP7_75t_R _28975_ (.A1(_05966_),
    .A2(_06056_),
    .B(_05900_),
    .Y(_06161_));
 AO21x1_ASAP7_75t_R _28976_ (.A1(_05781_),
    .A2(_05782_),
    .B(_01257_),
    .Y(_06162_));
 AOI21x1_ASAP7_75t_R _28977_ (.A1(_06162_),
    .A2(_06085_),
    .B(_05913_),
    .Y(_06163_));
 INVx1_ASAP7_75t_R _28978_ (.A(_06163_),
    .Y(_06164_));
 AOI21x1_ASAP7_75t_R _28979_ (.A1(_06164_),
    .A2(_05983_),
    .B(_05888_),
    .Y(_06165_));
 OAI21x1_ASAP7_75t_R _28980_ (.A1(_06161_),
    .A2(_06165_),
    .B(_05819_),
    .Y(_06166_));
 NAND2x1_ASAP7_75t_R _28981_ (.A(_05854_),
    .B(_05826_),
    .Y(_06167_));
 AO21x2_ASAP7_75t_R _28982_ (.A1(_05863_),
    .A2(_06068_),
    .B(_05874_),
    .Y(_06168_));
 NAND2x1_ASAP7_75t_R _28983_ (.A(_06167_),
    .B(_06168_),
    .Y(_06169_));
 AOI21x1_ASAP7_75t_R _28984_ (.A1(_05926_),
    .A2(_05884_),
    .B(_05900_),
    .Y(_06170_));
 AOI21x1_ASAP7_75t_R _28985_ (.A1(_06019_),
    .A2(_06170_),
    .B(_05915_),
    .Y(_06171_));
 OAI21x1_ASAP7_75t_R _28986_ (.A1(_05795_),
    .A2(_06169_),
    .B(_06171_),
    .Y(_06172_));
 AOI21x1_ASAP7_75t_R _28987_ (.A1(_06166_),
    .A2(_06172_),
    .B(_05962_),
    .Y(_06173_));
 NOR2x1_ASAP7_75t_R _28988_ (.A(_06160_),
    .B(_06173_),
    .Y(_06174_));
 AOI21x1_ASAP7_75t_R _28989_ (.A1(_05897_),
    .A2(_06147_),
    .B(_06174_),
    .Y(_00139_));
 AO21x1_ASAP7_75t_R _28990_ (.A1(_06111_),
    .A2(_06110_),
    .B(_05900_),
    .Y(_06175_));
 OAI21x1_ASAP7_75t_R _28991_ (.A1(_05967_),
    .A2(_06175_),
    .B(_05819_),
    .Y(_06176_));
 AND3x1_ASAP7_75t_R _28992_ (.A(_05982_),
    .B(_06010_),
    .C(_05931_),
    .Y(_06177_));
 OA21x2_ASAP7_75t_R _28993_ (.A1(_05797_),
    .A2(_05796_),
    .B(_05910_),
    .Y(_06178_));
 AO21x1_ASAP7_75t_R _28994_ (.A1(_06178_),
    .A2(_05783_),
    .B(_06016_),
    .Y(_06179_));
 NOR2x1_ASAP7_75t_R _28995_ (.A(_06177_),
    .B(_06179_),
    .Y(_06180_));
 AO21x1_ASAP7_75t_R _28996_ (.A1(_16033_),
    .A2(_16043_),
    .B(_05913_),
    .Y(_06181_));
 AOI21x1_ASAP7_75t_R _28997_ (.A1(_05971_),
    .A2(_06181_),
    .B(_05970_),
    .Y(_06182_));
 AO21x1_ASAP7_75t_R _28998_ (.A1(_05781_),
    .A2(_05782_),
    .B(_05903_),
    .Y(_06183_));
 AOI21x1_ASAP7_75t_R _28999_ (.A1(_05989_),
    .A2(_06183_),
    .B(_05906_),
    .Y(_06184_));
 AOI21x1_ASAP7_75t_R _29000_ (.A1(_05929_),
    .A2(_06184_),
    .B(_05915_),
    .Y(_06185_));
 OAI21x1_ASAP7_75t_R _29001_ (.A1(_05901_),
    .A2(_06182_),
    .B(_06185_),
    .Y(_06186_));
 OAI21x1_ASAP7_75t_R _29002_ (.A1(_06176_),
    .A2(_06180_),
    .B(_06186_),
    .Y(_06187_));
 OAI21x1_ASAP7_75t_R _29003_ (.A1(_05962_),
    .A2(_06187_),
    .B(_05897_),
    .Y(_06188_));
 INVx1_ASAP7_75t_R _29004_ (.A(_05923_),
    .Y(_06189_));
 NOR2x1_ASAP7_75t_R _29005_ (.A(_05976_),
    .B(_06098_),
    .Y(_06190_));
 NAND2x1_ASAP7_75t_R _29006_ (.A(_05855_),
    .B(_05926_),
    .Y(_06191_));
 OAI21x1_ASAP7_75t_R _29007_ (.A1(_06048_),
    .A2(_05902_),
    .B(_06191_),
    .Y(_06192_));
 OAI21x1_ASAP7_75t_R _29008_ (.A1(_06048_),
    .A2(_06057_),
    .B(_05915_),
    .Y(_06193_));
 AOI21x1_ASAP7_75t_R _29009_ (.A1(_06190_),
    .A2(_06192_),
    .B(_06193_),
    .Y(_06194_));
 OAI21x1_ASAP7_75t_R _29010_ (.A1(_06189_),
    .A2(_05901_),
    .B(_06194_),
    .Y(_06195_));
 AOI21x1_ASAP7_75t_R _29011_ (.A1(_05829_),
    .A2(_05941_),
    .B(_05794_),
    .Y(_06196_));
 NAND2x2_ASAP7_75t_R _29012_ (.A(_05910_),
    .B(net595),
    .Y(_06197_));
 AND3x1_ASAP7_75t_R _29013_ (.A(_05943_),
    .B(_06196_),
    .C(_06197_),
    .Y(_06198_));
 INVx1_ASAP7_75t_R _29014_ (.A(_05802_),
    .Y(_06199_));
 OAI21x1_ASAP7_75t_R _29015_ (.A1(_05902_),
    .A2(_05905_),
    .B(_06048_),
    .Y(_06200_));
 AOI21x1_ASAP7_75t_R _29016_ (.A1(_06199_),
    .A2(_05998_),
    .B(_06200_),
    .Y(_06201_));
 OAI21x1_ASAP7_75t_R _29017_ (.A1(_06198_),
    .A2(_06201_),
    .B(_05951_),
    .Y(_06202_));
 AOI21x1_ASAP7_75t_R _29018_ (.A1(_06195_),
    .A2(_06202_),
    .B(_05939_),
    .Y(_06203_));
 AOI21x1_ASAP7_75t_R _29019_ (.A1(_06010_),
    .A2(_05982_),
    .B(_06014_),
    .Y(_06204_));
 AO21x1_ASAP7_75t_R _29020_ (.A1(_05952_),
    .A2(_05904_),
    .B(_06204_),
    .Y(_06205_));
 NAND2x1_ASAP7_75t_R _29021_ (.A(_05824_),
    .B(_05839_),
    .Y(_06206_));
 NOR2x1_ASAP7_75t_R _29022_ (.A(_05779_),
    .B(_05958_),
    .Y(_06207_));
 AOI21x1_ASAP7_75t_R _29023_ (.A1(_06206_),
    .A2(_06207_),
    .B(_05936_),
    .Y(_06208_));
 OAI21x1_ASAP7_75t_R _29024_ (.A1(_05795_),
    .A2(_06205_),
    .B(_06208_),
    .Y(_06209_));
 OAI21x1_ASAP7_75t_R _29025_ (.A1(_00635_),
    .A2(_05989_),
    .B(_06197_),
    .Y(_06210_));
 AOI21x1_ASAP7_75t_R _29026_ (.A1(_06048_),
    .A2(_06210_),
    .B(_05915_),
    .Y(_06211_));
 NAND2x2_ASAP7_75t_R _29027_ (.A(_06010_),
    .B(_05904_),
    .Y(_06212_));
 AOI21x1_ASAP7_75t_R _29028_ (.A1(_05931_),
    .A2(_05920_),
    .B(_06016_),
    .Y(_06213_));
 NAND2x1_ASAP7_75t_R _29029_ (.A(_06212_),
    .B(_06213_),
    .Y(_06214_));
 AOI21x1_ASAP7_75t_R _29030_ (.A1(_06211_),
    .A2(_06214_),
    .B(_05939_),
    .Y(_06215_));
 NAND2x1_ASAP7_75t_R _29031_ (.A(_06209_),
    .B(_06215_),
    .Y(_06216_));
 AOI21x1_ASAP7_75t_R _29032_ (.A1(_05931_),
    .A2(_05999_),
    .B(_06016_),
    .Y(_06217_));
 AO21x1_ASAP7_75t_R _29033_ (.A1(_05995_),
    .A2(_16033_),
    .B(_05770_),
    .Y(_06218_));
 AOI21x1_ASAP7_75t_R _29034_ (.A1(_06217_),
    .A2(_06218_),
    .B(_05915_),
    .Y(_06219_));
 OR3x1_ASAP7_75t_R _29035_ (.A(_05865_),
    .B(net595),
    .C(_06014_),
    .Y(_06220_));
 AOI21x1_ASAP7_75t_R _29036_ (.A1(_05884_),
    .A2(_05885_),
    .B(_05779_),
    .Y(_06221_));
 NAND2x1_ASAP7_75t_R _29037_ (.A(_06221_),
    .B(_06220_),
    .Y(_06222_));
 NAND2x1_ASAP7_75t_R _29038_ (.A(_06222_),
    .B(_06219_),
    .Y(_06223_));
 AOI21x1_ASAP7_75t_R _29039_ (.A1(_05876_),
    .A2(_05866_),
    .B(_05855_),
    .Y(_06224_));
 AO21x1_ASAP7_75t_R _29040_ (.A1(_05876_),
    .A2(_05772_),
    .B(_05829_),
    .Y(_06225_));
 NAND2x1_ASAP7_75t_R _29041_ (.A(_06224_),
    .B(_06225_),
    .Y(_06226_));
 AOI21x1_ASAP7_75t_R _29042_ (.A1(_05854_),
    .A2(_05837_),
    .B(_06021_),
    .Y(_06227_));
 AOI21x1_ASAP7_75t_R _29043_ (.A1(_06048_),
    .A2(_06227_),
    .B(_05968_),
    .Y(_06228_));
 AOI21x1_ASAP7_75t_R _29044_ (.A1(_06226_),
    .A2(_06228_),
    .B(_05869_),
    .Y(_06229_));
 AOI21x1_ASAP7_75t_R _29045_ (.A1(_06223_),
    .A2(_06229_),
    .B(_05897_),
    .Y(_06230_));
 NAND2x1_ASAP7_75t_R _29046_ (.A(_06230_),
    .B(_06216_),
    .Y(_06231_));
 OAI21x1_ASAP7_75t_R _29047_ (.A1(_06188_),
    .A2(_06203_),
    .B(_06231_),
    .Y(_00140_));
 AO21x1_ASAP7_75t_R _29048_ (.A1(_05801_),
    .A2(_05854_),
    .B(_05950_),
    .Y(_06232_));
 OA21x2_ASAP7_75t_R _29049_ (.A1(_00629_),
    .A2(_16040_),
    .B(_05786_),
    .Y(_06233_));
 NAND2x1_ASAP7_75t_R _29050_ (.A(_05950_),
    .B(_05946_),
    .Y(_06234_));
 OA21x2_ASAP7_75t_R _29051_ (.A1(_06234_),
    .A2(_06122_),
    .B(_05888_),
    .Y(_06235_));
 OA21x2_ASAP7_75t_R _29052_ (.A1(_06232_),
    .A2(_06233_),
    .B(_06235_),
    .Y(_06236_));
 NAND2x1_ASAP7_75t_R _29053_ (.A(_05974_),
    .B(_05975_),
    .Y(_06237_));
 NAND2x1_ASAP7_75t_R _29054_ (.A(_06084_),
    .B(_05836_),
    .Y(_06238_));
 AO21x1_ASAP7_75t_R _29055_ (.A1(_06238_),
    .A2(_06014_),
    .B(_05818_),
    .Y(_06239_));
 AO21x1_ASAP7_75t_R _29056_ (.A1(_06237_),
    .A2(_05976_),
    .B(_06239_),
    .Y(_06240_));
 NOR2x1_ASAP7_75t_R _29057_ (.A(_05825_),
    .B(_16035_),
    .Y(_06241_));
 INVx1_ASAP7_75t_R _29058_ (.A(_06241_),
    .Y(_06242_));
 NAND2x1_ASAP7_75t_R _29059_ (.A(_05875_),
    .B(_06242_),
    .Y(_06243_));
 AO21x1_ASAP7_75t_R _29060_ (.A1(_00629_),
    .A2(_06014_),
    .B(_05817_),
    .Y(_06244_));
 OA21x2_ASAP7_75t_R _29061_ (.A1(_06243_),
    .A2(_06244_),
    .B(_06016_),
    .Y(_06245_));
 AO21x1_ASAP7_75t_R _29062_ (.A1(_06240_),
    .A2(_06245_),
    .B(_05939_),
    .Y(_06246_));
 OA21x2_ASAP7_75t_R _29063_ (.A1(net30),
    .A2(_05913_),
    .B(_05794_),
    .Y(_06247_));
 AOI21x1_ASAP7_75t_R _29064_ (.A1(_06247_),
    .A2(_05838_),
    .B(_05841_),
    .Y(_06248_));
 NOR2x1_ASAP7_75t_R _29065_ (.A(net29),
    .B(_05863_),
    .Y(_06249_));
 AOI21x1_ASAP7_75t_R _29066_ (.A1(_06010_),
    .A2(_06077_),
    .B(_06016_),
    .Y(_06250_));
 OAI21x1_ASAP7_75t_R _29067_ (.A1(_06249_),
    .A2(_05944_),
    .B(_06250_),
    .Y(_06251_));
 AOI21x1_ASAP7_75t_R _29068_ (.A1(_06248_),
    .A2(_06251_),
    .B(_05869_),
    .Y(_06252_));
 INVx1_ASAP7_75t_R _29069_ (.A(_06221_),
    .Y(_06253_));
 AND3x1_ASAP7_75t_R _29070_ (.A(_05859_),
    .B(_05931_),
    .C(_06065_),
    .Y(_06254_));
 OA21x2_ASAP7_75t_R _29071_ (.A1(_05789_),
    .A2(_05913_),
    .B(_05887_),
    .Y(_06255_));
 OAI21x1_ASAP7_75t_R _29072_ (.A1(_06241_),
    .A2(_05955_),
    .B(_05854_),
    .Y(_06256_));
 AOI21x1_ASAP7_75t_R _29073_ (.A1(_06255_),
    .A2(_06256_),
    .B(_05936_),
    .Y(_06257_));
 OAI21x1_ASAP7_75t_R _29074_ (.A1(_06253_),
    .A2(_06254_),
    .B(_06257_),
    .Y(_06258_));
 AOI21x1_ASAP7_75t_R _29075_ (.A1(_06252_),
    .A2(_06258_),
    .B(_05897_),
    .Y(_06259_));
 OAI21x1_ASAP7_75t_R _29076_ (.A1(_06236_),
    .A2(_06246_),
    .B(_06259_),
    .Y(_06260_));
 INVx1_ASAP7_75t_R _29077_ (.A(_05858_),
    .Y(_06261_));
 NOR2x2_ASAP7_75t_R _29078_ (.A(net524),
    .B(net516),
    .Y(_06262_));
 OA21x2_ASAP7_75t_R _29079_ (.A1(_06261_),
    .A2(_06262_),
    .B(_05900_),
    .Y(_06263_));
 OR3x1_ASAP7_75t_R _29080_ (.A(_05973_),
    .B(_05770_),
    .C(_05790_),
    .Y(_06264_));
 NAND2x2_ASAP7_75t_R _29081_ (.A(_05828_),
    .B(net516),
    .Y(_06265_));
 NAND2x1_ASAP7_75t_R _29082_ (.A(_05794_),
    .B(_06265_),
    .Y(_06266_));
 OAI21x1_ASAP7_75t_R _29083_ (.A1(_06266_),
    .A2(_06204_),
    .B(_05936_),
    .Y(_06267_));
 AOI21x1_ASAP7_75t_R _29084_ (.A1(_06263_),
    .A2(_06264_),
    .B(_06267_),
    .Y(_06268_));
 AO21x1_ASAP7_75t_R _29085_ (.A1(_06045_),
    .A2(_06009_),
    .B(_06014_),
    .Y(_06269_));
 NAND2x1_ASAP7_75t_R _29086_ (.A(_06197_),
    .B(_06269_),
    .Y(_06270_));
 AO21x1_ASAP7_75t_R _29087_ (.A1(_06069_),
    .A2(_05913_),
    .B(_05887_),
    .Y(_06271_));
 NOR2x1_ASAP7_75t_R _29088_ (.A(_06105_),
    .B(_05944_),
    .Y(_06272_));
 OAI21x1_ASAP7_75t_R _29089_ (.A1(_06271_),
    .A2(_06272_),
    .B(_05841_),
    .Y(_06273_));
 AOI21x1_ASAP7_75t_R _29090_ (.A1(_05901_),
    .A2(_06270_),
    .B(_06273_),
    .Y(_06274_));
 OAI21x1_ASAP7_75t_R _29091_ (.A1(_06268_),
    .A2(_06274_),
    .B(_05869_),
    .Y(_06275_));
 AOI21x1_ASAP7_75t_R _29092_ (.A1(_06021_),
    .A2(_05909_),
    .B(_05855_),
    .Y(_06276_));
 NAND2x1_ASAP7_75t_R _29093_ (.A(_06015_),
    .B(_06276_),
    .Y(_06277_));
 NOR2x1_ASAP7_75t_R _29094_ (.A(_05779_),
    .B(_05826_),
    .Y(_06278_));
 AOI21x1_ASAP7_75t_R _29095_ (.A1(_06278_),
    .A2(_06168_),
    .B(_05936_),
    .Y(_06279_));
 AOI21x1_ASAP7_75t_R _29096_ (.A1(_06277_),
    .A2(_06279_),
    .B(_05869_),
    .Y(_06280_));
 OAI21x1_ASAP7_75t_R _29097_ (.A1(_06026_),
    .A2(_06056_),
    .B(_05989_),
    .Y(_06281_));
 AOI21x1_ASAP7_75t_R _29098_ (.A1(_05770_),
    .A2(_05882_),
    .B(_05779_),
    .Y(_06282_));
 AOI21x1_ASAP7_75t_R _29099_ (.A1(_06281_),
    .A2(_06282_),
    .B(_05841_),
    .Y(_06283_));
 NOR2x1_ASAP7_75t_R _29100_ (.A(net563),
    .B(_05874_),
    .Y(_06284_));
 AOI211x1_ASAP7_75t_R _29101_ (.A1(_05906_),
    .A2(_05829_),
    .B(_06284_),
    .C(_05855_),
    .Y(_06285_));
 OAI21x1_ASAP7_75t_R _29102_ (.A1(_05902_),
    .A2(_06078_),
    .B(_06285_),
    .Y(_06286_));
 NAND2x1_ASAP7_75t_R _29103_ (.A(_06283_),
    .B(_06286_),
    .Y(_06287_));
 AOI21x1_ASAP7_75t_R _29104_ (.A1(_06280_),
    .A2(_06287_),
    .B(_05896_),
    .Y(_06288_));
 NAND2x1_ASAP7_75t_R _29105_ (.A(_06288_),
    .B(_06275_),
    .Y(_06289_));
 NAND2x1_ASAP7_75t_R _29106_ (.A(_06260_),
    .B(_06289_),
    .Y(_00141_));
 OA21x2_ASAP7_75t_R _29107_ (.A1(_05789_),
    .A2(_05910_),
    .B(_05887_),
    .Y(_06290_));
 AO21x1_ASAP7_75t_R _29108_ (.A1(_05952_),
    .A2(_16033_),
    .B(_05913_),
    .Y(_06291_));
 AOI21x1_ASAP7_75t_R _29109_ (.A1(_06290_),
    .A2(_06291_),
    .B(_05950_),
    .Y(_06292_));
 AOI21x1_ASAP7_75t_R _29110_ (.A1(_06238_),
    .A2(_05933_),
    .B(_05887_),
    .Y(_06293_));
 AO21x1_ASAP7_75t_R _29111_ (.A1(_06097_),
    .A2(_06265_),
    .B(_05995_),
    .Y(_06294_));
 NAND2x1_ASAP7_75t_R _29112_ (.A(_06293_),
    .B(_06294_),
    .Y(_06295_));
 AOI21x1_ASAP7_75t_R _29113_ (.A1(_06292_),
    .A2(_06295_),
    .B(_05849_),
    .Y(_06296_));
 NAND2x1_ASAP7_75t_R _29114_ (.A(_05887_),
    .B(_06151_),
    .Y(_06297_));
 AOI21x1_ASAP7_75t_R _29115_ (.A1(_06091_),
    .A2(_06049_),
    .B(_06297_),
    .Y(_06298_));
 NAND2x2_ASAP7_75t_R _29116_ (.A(_05942_),
    .B(_05999_),
    .Y(_06299_));
 OAI21x1_ASAP7_75t_R _29117_ (.A1(_16040_),
    .A2(_05909_),
    .B(_06178_),
    .Y(_06300_));
 OA21x2_ASAP7_75t_R _29118_ (.A1(_05799_),
    .A2(_05828_),
    .B(_05794_),
    .Y(_06301_));
 INVx1_ASAP7_75t_R _29119_ (.A(_06301_),
    .Y(_06302_));
 AOI21x1_ASAP7_75t_R _29120_ (.A1(_06299_),
    .A2(_06300_),
    .B(_06302_),
    .Y(_06303_));
 OAI21x1_ASAP7_75t_R _29121_ (.A1(_06298_),
    .A2(_06303_),
    .B(_05951_),
    .Y(_06304_));
 NAND2x1_ASAP7_75t_R _29122_ (.A(_06296_),
    .B(_06304_),
    .Y(_06305_));
 AO21x1_ASAP7_75t_R _29123_ (.A1(_06077_),
    .A2(_06006_),
    .B(_05900_),
    .Y(_06306_));
 AOI21x1_ASAP7_75t_R _29124_ (.A1(_05881_),
    .A2(_06001_),
    .B(_05976_),
    .Y(_06307_));
 AO21x1_ASAP7_75t_R _29125_ (.A1(_05781_),
    .A2(_05782_),
    .B(_06084_),
    .Y(_06308_));
 AO21x1_ASAP7_75t_R _29126_ (.A1(_06068_),
    .A2(_06308_),
    .B(_05942_),
    .Y(_06309_));
 AOI21x1_ASAP7_75t_R _29127_ (.A1(_05954_),
    .A2(_05837_),
    .B(_06016_),
    .Y(_06310_));
 AOI21x1_ASAP7_75t_R _29128_ (.A1(_06309_),
    .A2(_06310_),
    .B(_05936_),
    .Y(_06311_));
 OAI21x1_ASAP7_75t_R _29129_ (.A1(_06306_),
    .A2(_06307_),
    .B(_06311_),
    .Y(_06312_));
 NAND2x1_ASAP7_75t_R _29130_ (.A(_05942_),
    .B(_05773_),
    .Y(_06313_));
 NAND2x1_ASAP7_75t_R _29131_ (.A(_05880_),
    .B(_06021_),
    .Y(_06314_));
 NAND3x1_ASAP7_75t_R _29132_ (.A(_06196_),
    .B(_06313_),
    .C(_06314_),
    .Y(_06315_));
 AND2x2_ASAP7_75t_R _29133_ (.A(_01261_),
    .B(_01259_),
    .Y(_06316_));
 OA21x2_ASAP7_75t_R _29134_ (.A1(_06014_),
    .A2(_06316_),
    .B(_05794_),
    .Y(_06317_));
 AO21x1_ASAP7_75t_R _29135_ (.A1(_05982_),
    .A2(_06009_),
    .B(_05942_),
    .Y(_06318_));
 AOI21x1_ASAP7_75t_R _29136_ (.A1(_06317_),
    .A2(_06318_),
    .B(_05841_),
    .Y(_06319_));
 AOI21x1_ASAP7_75t_R _29137_ (.A1(_06315_),
    .A2(_06319_),
    .B(_05869_),
    .Y(_06320_));
 AOI21x1_ASAP7_75t_R _29138_ (.A1(_06312_),
    .A2(_06320_),
    .B(_05896_),
    .Y(_06321_));
 NAND2x1_ASAP7_75t_R _29139_ (.A(_06305_),
    .B(_06321_),
    .Y(_06322_));
 OA21x2_ASAP7_75t_R _29140_ (.A1(_06111_),
    .A2(_05998_),
    .B(_05824_),
    .Y(_06323_));
 INVx1_ASAP7_75t_R _29141_ (.A(_05857_),
    .Y(_06324_));
 AOI21x1_ASAP7_75t_R _29142_ (.A1(_06324_),
    .A2(_06119_),
    .B(_05841_),
    .Y(_06325_));
 OAI21x1_ASAP7_75t_R _29143_ (.A1(_05795_),
    .A2(_06323_),
    .B(_06325_),
    .Y(_06326_));
 NAND2x1_ASAP7_75t_R _29144_ (.A(_06301_),
    .B(_06168_),
    .Y(_06327_));
 AOI21x1_ASAP7_75t_R _29145_ (.A1(_06008_),
    .A2(_05860_),
    .B(_05936_),
    .Y(_06328_));
 NAND2x1_ASAP7_75t_R _29146_ (.A(_06327_),
    .B(_06328_),
    .Y(_06329_));
 AOI21x1_ASAP7_75t_R _29147_ (.A1(_06326_),
    .A2(_06329_),
    .B(_05869_),
    .Y(_06330_));
 OA21x2_ASAP7_75t_R _29148_ (.A1(_05944_),
    .A2(_06056_),
    .B(_06038_),
    .Y(_06331_));
 AND2x2_ASAP7_75t_R _29149_ (.A(_05910_),
    .B(_00636_),
    .Y(_06332_));
 AOI21x1_ASAP7_75t_R _29150_ (.A1(_06010_),
    .A2(_06077_),
    .B(_06332_),
    .Y(_06333_));
 AOI21x1_ASAP7_75t_R _29151_ (.A1(_06048_),
    .A2(_06333_),
    .B(_05915_),
    .Y(_06334_));
 OAI21x1_ASAP7_75t_R _29152_ (.A1(_05795_),
    .A2(_06331_),
    .B(_06334_),
    .Y(_06335_));
 INVx1_ASAP7_75t_R _29153_ (.A(_05911_),
    .Y(_06336_));
 AOI21x1_ASAP7_75t_R _29154_ (.A1(_06336_),
    .A2(_06212_),
    .B(_06048_),
    .Y(_06337_));
 OAI21x1_ASAP7_75t_R _29155_ (.A1(_06060_),
    .A2(_06337_),
    .B(_05819_),
    .Y(_06338_));
 AOI21x1_ASAP7_75t_R _29156_ (.A1(_06335_),
    .A2(_06338_),
    .B(_05939_),
    .Y(_06339_));
 OAI21x1_ASAP7_75t_R _29157_ (.A1(_06330_),
    .A2(_06339_),
    .B(_05896_),
    .Y(_06340_));
 NAND2x1_ASAP7_75t_R _29158_ (.A(_06322_),
    .B(_06340_),
    .Y(_00142_));
 OAI21x1_ASAP7_75t_R _29159_ (.A1(_16040_),
    .A2(_06262_),
    .B(_05772_),
    .Y(_06341_));
 AOI21x1_ASAP7_75t_R _29160_ (.A1(_05789_),
    .A2(_05786_),
    .B(_05888_),
    .Y(_06342_));
 OAI21x1_ASAP7_75t_R _29161_ (.A1(_05922_),
    .A2(_06341_),
    .B(_06342_),
    .Y(_06343_));
 AOI21x1_ASAP7_75t_R _29162_ (.A1(_16033_),
    .A2(_05863_),
    .B(_05922_),
    .Y(_06344_));
 OAI21x1_ASAP7_75t_R _29163_ (.A1(_06163_),
    .A2(_06344_),
    .B(_05929_),
    .Y(_06345_));
 NAND3x1_ASAP7_75t_R _29164_ (.A(_06343_),
    .B(_06345_),
    .C(_05951_),
    .Y(_06346_));
 INVx1_ASAP7_75t_R _29165_ (.A(_06191_),
    .Y(_06347_));
 NAND2x1_ASAP7_75t_R _29166_ (.A(_06299_),
    .B(_06181_),
    .Y(_06348_));
 AOI21x1_ASAP7_75t_R _29167_ (.A1(_06347_),
    .A2(_06348_),
    .B(_05951_),
    .Y(_06349_));
 NAND2x1_ASAP7_75t_R _29168_ (.A(_05864_),
    .B(_05976_),
    .Y(_06350_));
 AO21x1_ASAP7_75t_R _29169_ (.A1(_06318_),
    .A2(_06350_),
    .B(_05795_),
    .Y(_06351_));
 NAND2x1_ASAP7_75t_R _29170_ (.A(_06349_),
    .B(_06351_),
    .Y(_06352_));
 AOI21x1_ASAP7_75t_R _29171_ (.A1(_06346_),
    .A2(_06352_),
    .B(_05962_),
    .Y(_06353_));
 AO21x1_ASAP7_75t_R _29172_ (.A1(_05952_),
    .A2(_16033_),
    .B(_05922_),
    .Y(_06354_));
 NAND2x1_ASAP7_75t_R _29173_ (.A(_00635_),
    .B(_05989_),
    .Y(_06355_));
 AO21x1_ASAP7_75t_R _29174_ (.A1(_05925_),
    .A2(_06355_),
    .B(_05915_),
    .Y(_06356_));
 AOI21x1_ASAP7_75t_R _29175_ (.A1(_06224_),
    .A2(_06354_),
    .B(_06356_),
    .Y(_06357_));
 OA21x2_ASAP7_75t_R _29176_ (.A1(_01261_),
    .A2(_05770_),
    .B(_05855_),
    .Y(_06358_));
 OAI21x1_ASAP7_75t_R _29177_ (.A1(_05802_),
    .A2(_05941_),
    .B(_05976_),
    .Y(_06359_));
 AO21x1_ASAP7_75t_R _29178_ (.A1(_06358_),
    .A2(_06359_),
    .B(_05968_),
    .Y(_06360_));
 AND3x1_ASAP7_75t_R _29179_ (.A(_05799_),
    .B(_05989_),
    .C(_06199_),
    .Y(_06361_));
 AO21x1_ASAP7_75t_R _29180_ (.A1(_05858_),
    .A2(_06010_),
    .B(_06016_),
    .Y(_06362_));
 NOR2x1_ASAP7_75t_R _29181_ (.A(_06361_),
    .B(_06362_),
    .Y(_06363_));
 OAI21x1_ASAP7_75t_R _29182_ (.A1(_06360_),
    .A2(_06363_),
    .B(_05962_),
    .Y(_06364_));
 OAI21x1_ASAP7_75t_R _29183_ (.A1(_06357_),
    .A2(_06364_),
    .B(_05897_),
    .Y(_06365_));
 AOI21x1_ASAP7_75t_R _29184_ (.A1(_06110_),
    .A2(_06001_),
    .B(_05922_),
    .Y(_06366_));
 NOR2x1_ASAP7_75t_R _29185_ (.A(_06366_),
    .B(_06175_),
    .Y(_06367_));
 OAI21x1_ASAP7_75t_R _29186_ (.A1(_05965_),
    .A2(_06097_),
    .B(_06242_),
    .Y(_06368_));
 AO21x1_ASAP7_75t_R _29187_ (.A1(_06368_),
    .A2(_05929_),
    .B(_05819_),
    .Y(_06369_));
 NOR2x1_ASAP7_75t_R _29188_ (.A(_06367_),
    .B(_06369_),
    .Y(_06370_));
 AOI21x1_ASAP7_75t_R _29189_ (.A1(_16043_),
    .A2(_06262_),
    .B(_05800_),
    .Y(_06371_));
 NAND3x1_ASAP7_75t_R _29190_ (.A(_06097_),
    .B(_05888_),
    .C(_06265_),
    .Y(_06372_));
 NOR2x1_ASAP7_75t_R _29191_ (.A(_06371_),
    .B(_06372_),
    .Y(_06373_));
 AND2x2_ASAP7_75t_R _29192_ (.A(_06151_),
    .B(_05855_),
    .Y(_06374_));
 NAND2x1_ASAP7_75t_R _29193_ (.A(_05922_),
    .B(_05973_),
    .Y(_06375_));
 AO21x1_ASAP7_75t_R _29194_ (.A1(_06374_),
    .A2(_06375_),
    .B(_05968_),
    .Y(_06376_));
 OAI21x1_ASAP7_75t_R _29195_ (.A1(_06373_),
    .A2(_06376_),
    .B(_05962_),
    .Y(_06377_));
 OAI21x1_ASAP7_75t_R _29196_ (.A1(_06370_),
    .A2(_06377_),
    .B(_05896_),
    .Y(_06378_));
 AND2x2_ASAP7_75t_R _29197_ (.A(_06341_),
    .B(_05989_),
    .Y(_06379_));
 OAI21x1_ASAP7_75t_R _29198_ (.A1(_06261_),
    .A2(_05902_),
    .B(_05968_),
    .Y(_06380_));
 NAND2x1_ASAP7_75t_R _29199_ (.A(_06006_),
    .B(_05803_),
    .Y(_06381_));
 AOI21x1_ASAP7_75t_R _29200_ (.A1(_06381_),
    .A2(_06155_),
    .B(_06048_),
    .Y(_06382_));
 OA21x2_ASAP7_75t_R _29201_ (.A1(_06379_),
    .A2(_06380_),
    .B(_06382_),
    .Y(_06383_));
 AOI211x1_ASAP7_75t_R _29202_ (.A1(_06006_),
    .A2(_06077_),
    .B(_06099_),
    .C(_05968_),
    .Y(_06384_));
 NOR2x1_ASAP7_75t_R _29203_ (.A(_05818_),
    .B(_05998_),
    .Y(_06385_));
 AO21x1_ASAP7_75t_R _29204_ (.A1(_06212_),
    .A2(_06385_),
    .B(_05929_),
    .Y(_06386_));
 OAI21x1_ASAP7_75t_R _29205_ (.A1(_06384_),
    .A2(_06386_),
    .B(_05939_),
    .Y(_06387_));
 NOR2x1_ASAP7_75t_R _29206_ (.A(_06383_),
    .B(_06387_),
    .Y(_06388_));
 OAI22x1_ASAP7_75t_R _29207_ (.A1(_06353_),
    .A2(_06365_),
    .B1(_06378_),
    .B2(_06388_),
    .Y(_00143_));
 NOR2x2_ASAP7_75t_R _29208_ (.A(net621),
    .B(_00637_),
    .Y(_06389_));
 XOR2x1_ASAP7_75t_R _29209_ (.A(net597),
    .Y(_06390_),
    .B(net850));
 XOR2x1_ASAP7_75t_R _29210_ (.A(net829),
    .Y(_06391_),
    .B(_12128_));
 NAND2x1_ASAP7_75t_R _29211_ (.A(_06390_),
    .B(_06391_),
    .Y(_06392_));
 XNOR2x1_ASAP7_75t_R _29212_ (.B(net597),
    .Y(_06393_),
    .A(net850));
 XOR2x1_ASAP7_75t_R _29213_ (.A(_12130_),
    .Y(_06394_),
    .B(net829));
 NAND2x1_ASAP7_75t_R _29214_ (.A(_06393_),
    .B(_06394_),
    .Y(_06395_));
 AOI21x1_ASAP7_75t_R _29215_ (.A1(_06392_),
    .A2(_06395_),
    .B(_11441_),
    .Y(_06396_));
 OAI21x1_ASAP7_75t_R _29216_ (.A1(_06389_),
    .A2(_06396_),
    .B(_08026_),
    .Y(_06397_));
 AND2x2_ASAP7_75t_R _29217_ (.A(_10643_),
    .B(_00637_),
    .Y(_06398_));
 NAND2x1_ASAP7_75t_R _29218_ (.A(_06390_),
    .B(_06394_),
    .Y(_06399_));
 NAND2x1_ASAP7_75t_R _29219_ (.A(_06393_),
    .B(_06391_),
    .Y(_06400_));
 AOI21x1_ASAP7_75t_R _29220_ (.A1(_06400_),
    .A2(_06399_),
    .B(_11441_),
    .Y(_06401_));
 INVx1_ASAP7_75t_R _29221_ (.A(_08026_),
    .Y(_06402_));
 OAI21x1_ASAP7_75t_R _29222_ (.A1(_06398_),
    .A2(_06401_),
    .B(_06402_),
    .Y(_06403_));
 NAND2x2_ASAP7_75t_R _29223_ (.A(_06403_),
    .B(_06397_),
    .Y(_06404_));
 BUFx12f_ASAP7_75t_R _29224_ (.A(_06404_),
    .Y(_16050_));
 OR2x2_ASAP7_75t_R _29225_ (.A(_10666_),
    .B(_00638_),
    .Y(_06405_));
 NOR2x2_ASAP7_75t_R _29226_ (.A(_12276_),
    .B(_12116_),
    .Y(_06406_));
 NOR2x2_ASAP7_75t_R _29227_ (.A(_12275_),
    .B(_12111_),
    .Y(_06407_));
 OAI21x1_ASAP7_75t_R _29228_ (.A1(_06407_),
    .A2(_06406_),
    .B(net597),
    .Y(_06408_));
 INVx1_ASAP7_75t_R _29229_ (.A(_06408_),
    .Y(_06409_));
 NOR3x1_ASAP7_75t_R _29230_ (.A(_06407_),
    .B(_06406_),
    .C(net591),
    .Y(_06410_));
 OAI21x1_ASAP7_75t_R _29231_ (.A1(_06410_),
    .A2(_06409_),
    .B(_10761_),
    .Y(_06411_));
 AOI21x1_ASAP7_75t_R _29232_ (.A1(_06405_),
    .A2(_06411_),
    .B(net854),
    .Y(_06412_));
 NAND2x1_ASAP7_75t_R _29233_ (.A(_00638_),
    .B(_12095_),
    .Y(_06413_));
 NAND2x2_ASAP7_75t_R _29234_ (.A(_12275_),
    .B(_12111_),
    .Y(_06414_));
 NAND2x2_ASAP7_75t_R _29235_ (.A(_12276_),
    .B(_12116_),
    .Y(_06415_));
 INVx1_ASAP7_75t_R _29236_ (.A(net597),
    .Y(_06416_));
 NAND3x2_ASAP7_75t_R _29237_ (.B(_06415_),
    .C(_06416_),
    .Y(_06417_),
    .A(_06414_));
 NAND3x2_ASAP7_75t_R _29238_ (.B(_11356_),
    .C(_06417_),
    .Y(_06418_),
    .A(_06408_));
 INVx1_ASAP7_75t_R _29239_ (.A(net854),
    .Y(_06419_));
 AOI21x1_ASAP7_75t_R _29240_ (.A1(_06413_),
    .A2(_06418_),
    .B(_06419_),
    .Y(_06420_));
 NOR2x2_ASAP7_75t_R _29241_ (.A(_06420_),
    .B(_06412_),
    .Y(_06421_));
 BUFx12_ASAP7_75t_R _29242_ (.A(_06421_),
    .Y(_16052_));
 XOR2x1_ASAP7_75t_R _29243_ (.A(net59),
    .Y(_06422_),
    .B(_12132_));
 NAND2x1_ASAP7_75t_R _29244_ (.A(_12097_),
    .B(_06422_),
    .Y(_06423_));
 XNOR2x1_ASAP7_75t_R _29245_ (.B(_12132_),
    .Y(_06424_),
    .A(_12127_));
 NAND2x1_ASAP7_75t_R _29246_ (.A(net844),
    .B(_06424_),
    .Y(_06425_));
 AOI21x1_ASAP7_75t_R _29247_ (.A1(_06423_),
    .A2(_06425_),
    .B(_03644_),
    .Y(_06426_));
 XOR2x1_ASAP7_75t_R _29248_ (.A(_12132_),
    .Y(_06427_),
    .B(net844));
 NAND2x1_ASAP7_75t_R _29249_ (.A(net59),
    .B(_06427_),
    .Y(_06428_));
 XNOR2x1_ASAP7_75t_R _29250_ (.B(net844),
    .Y(_06429_),
    .A(_12132_));
 NAND2x1_ASAP7_75t_R _29251_ (.A(_15019_),
    .B(_06429_),
    .Y(_06430_));
 AOI21x1_ASAP7_75t_R _29252_ (.A1(_06428_),
    .A2(_06430_),
    .B(_03634_),
    .Y(_06431_));
 OAI21x1_ASAP7_75t_R _29253_ (.A1(_06426_),
    .A2(_06431_),
    .B(net680),
    .Y(_06432_));
 NOR2x2_ASAP7_75t_R _29254_ (.A(net786),
    .B(_00639_),
    .Y(_06433_));
 INVx3_ASAP7_75t_R _29255_ (.A(_06433_),
    .Y(_06434_));
 NAND3x2_ASAP7_75t_R _29256_ (.B(_08035_),
    .C(_06434_),
    .Y(_06435_),
    .A(_06432_));
 AO21x2_ASAP7_75t_R _29257_ (.A1(_06432_),
    .A2(_06434_),
    .B(_08035_),
    .Y(_06436_));
 NAND2x2_ASAP7_75t_R _29258_ (.A(_06435_),
    .B(_06436_),
    .Y(_06437_));
 BUFx12_ASAP7_75t_R _29259_ (.A(_06437_),
    .Y(_06438_));
 BUFx10_ASAP7_75t_R _29260_ (.A(_06438_),
    .Y(_16060_));
 AOI21x1_ASAP7_75t_R _29261_ (.A1(_06411_),
    .A2(_06405_),
    .B(_06419_),
    .Y(_06439_));
 AOI21x1_ASAP7_75t_R _29262_ (.A1(_06418_),
    .A2(_06413_),
    .B(net855),
    .Y(_06440_));
 NOR2x2_ASAP7_75t_R _29263_ (.A(_06440_),
    .B(_06439_),
    .Y(_06441_));
 BUFx2_ASAP7_75t_R rebuffer354 (.A(_06441_),
    .Y(net807));
 BUFx6f_ASAP7_75t_R _29265_ (.A(_06441_),
    .Y(_16047_));
 NAND3x2_ASAP7_75t_R _29266_ (.B(_08258_),
    .C(_06434_),
    .Y(_06443_),
    .A(_06432_));
 AO21x1_ASAP7_75t_R _29267_ (.A1(_06432_),
    .A2(_06434_),
    .B(_08258_),
    .Y(_06444_));
 BUFx4f_ASAP7_75t_R _29268_ (.A(_06444_),
    .Y(_06445_));
 NAND2x2_ASAP7_75t_R _29269_ (.A(_06443_),
    .B(_06445_),
    .Y(_06446_));
 BUFx10_ASAP7_75t_R _29270_ (.A(_06446_),
    .Y(_16057_));
 XNOR2x1_ASAP7_75t_R _29271_ (.B(_12170_),
    .Y(_06447_),
    .A(_00815_));
 XOR2x1_ASAP7_75t_R _29272_ (.A(_03658_),
    .Y(_06448_),
    .B(_03657_));
 NOR2x1_ASAP7_75t_R _29273_ (.A(_06447_),
    .B(_06448_),
    .Y(_06449_));
 XOR2x1_ASAP7_75t_R _29274_ (.A(_12170_),
    .Y(_06450_),
    .B(_00815_));
 OAI21x1_ASAP7_75t_R _29275_ (.A1(_06450_),
    .A2(_03659_),
    .B(net621),
    .Y(_06451_));
 NAND2x2_ASAP7_75t_R _29276_ (.A(_00690_),
    .B(_10643_),
    .Y(_06452_));
 OAI21x1_ASAP7_75t_R _29277_ (.A1(_06449_),
    .A2(_06451_),
    .B(_06452_),
    .Y(_06453_));
 XOR2x2_ASAP7_75t_R _29278_ (.A(_06453_),
    .B(_08047_),
    .Y(_06454_));
 BUFx6f_ASAP7_75t_R _29279_ (.A(_06454_),
    .Y(_06455_));
 NOR2x1_ASAP7_75t_R _29280_ (.A(_12097_),
    .B(_06422_),
    .Y(_06456_));
 NOR2x1_ASAP7_75t_R _29281_ (.A(net844),
    .B(_06424_),
    .Y(_06457_));
 OAI21x1_ASAP7_75t_R _29282_ (.A1(_06456_),
    .A2(_06457_),
    .B(_03634_),
    .Y(_06458_));
 NOR2x1_ASAP7_75t_R _29283_ (.A(net59),
    .B(_06427_),
    .Y(_06459_));
 NOR2x1_ASAP7_75t_R _29284_ (.A(_15019_),
    .B(_06429_),
    .Y(_06460_));
 OAI21x1_ASAP7_75t_R _29285_ (.A1(_06459_),
    .A2(_06460_),
    .B(_03644_),
    .Y(_06461_));
 AOI21x1_ASAP7_75t_R _29286_ (.A1(_06458_),
    .A2(_06461_),
    .B(_12161_),
    .Y(_06462_));
 NOR3x2_ASAP7_75t_R _29287_ (.B(_08035_),
    .C(_06433_),
    .Y(_06463_),
    .A(_06462_));
 OA21x2_ASAP7_75t_R _29288_ (.A1(_06462_),
    .A2(_06433_),
    .B(_08035_),
    .Y(_06464_));
 INVx2_ASAP7_75t_R _29289_ (.A(_01263_),
    .Y(_06465_));
 OAI21x1_ASAP7_75t_R _29290_ (.A1(_06463_),
    .A2(_06464_),
    .B(_06465_),
    .Y(_06466_));
 XNOR2x1_ASAP7_75t_R _29291_ (.B(_12184_),
    .Y(_06467_),
    .A(_00816_));
 XOR2x1_ASAP7_75t_R _29292_ (.A(_06467_),
    .Y(_06468_),
    .B(_03682_));
 NOR2x1_ASAP7_75t_R _29293_ (.A(_10743_),
    .B(_00689_),
    .Y(_06469_));
 AOI21x1_ASAP7_75t_R _29294_ (.A1(_10734_),
    .A2(_06468_),
    .B(_06469_),
    .Y(_06470_));
 XNOR2x2_ASAP7_75t_R _29295_ (.A(_01085_),
    .B(_06470_),
    .Y(_06471_));
 OAI21x1_ASAP7_75t_R _29296_ (.A1(_06455_),
    .A2(_06466_),
    .B(_06471_),
    .Y(_06472_));
 OAI21x1_ASAP7_75t_R _29297_ (.A1(_06389_),
    .A2(_06396_),
    .B(_06402_),
    .Y(_06473_));
 OAI21x1_ASAP7_75t_R _29298_ (.A1(_06401_),
    .A2(_06398_),
    .B(_08026_),
    .Y(_06474_));
 NAND2x2_ASAP7_75t_R _29299_ (.A(_06474_),
    .B(_06473_),
    .Y(_06475_));
 NOR2x2_ASAP7_75t_R _29300_ (.A(_06437_),
    .B(net627),
    .Y(_06476_));
 INVx1_ASAP7_75t_R _29301_ (.A(_01265_),
    .Y(_06477_));
 BUFx10_ASAP7_75t_R _29302_ (.A(_06446_),
    .Y(_06478_));
 OAI21x1_ASAP7_75t_R _29303_ (.A1(_06477_),
    .A2(_06478_),
    .B(_06454_),
    .Y(_06479_));
 AOI21x1_ASAP7_75t_R _29304_ (.A1(net21),
    .A2(_06476_),
    .B(_06479_),
    .Y(_06480_));
 NOR2x1_ASAP7_75t_R _29305_ (.A(_11450_),
    .B(_00688_),
    .Y(_06481_));
 INVx1_ASAP7_75t_R _29306_ (.A(_06481_),
    .Y(_06482_));
 XOR2x1_ASAP7_75t_R _29307_ (.A(_12258_),
    .Y(_06483_),
    .B(_00848_));
 XNOR2x1_ASAP7_75t_R _29308_ (.B(_00753_),
    .Y(_06484_),
    .A(_00752_));
 XOR2x2_ASAP7_75t_R _29309_ (.A(_06483_),
    .B(_06484_),
    .Y(_06485_));
 NAND2x1_ASAP7_75t_R _29310_ (.A(_10787_),
    .B(_06485_),
    .Y(_06486_));
 AOI21x1_ASAP7_75t_R _29311_ (.A1(_06482_),
    .A2(_06486_),
    .B(_01086_),
    .Y(_06487_));
 INVx1_ASAP7_75t_R _29312_ (.A(_01086_),
    .Y(_06488_));
 AOI211x1_ASAP7_75t_R _29313_ (.A1(_06485_),
    .A2(_10786_),
    .B(_06481_),
    .C(_06488_),
    .Y(_06489_));
 NOR2x2_ASAP7_75t_R _29314_ (.A(_06487_),
    .B(_06489_),
    .Y(_06490_));
 BUFx6f_ASAP7_75t_R _29315_ (.A(_06490_),
    .Y(_06491_));
 OAI21x1_ASAP7_75t_R _29316_ (.A1(_06472_),
    .A2(_06480_),
    .B(_06491_),
    .Y(_06492_));
 NAND2x1_ASAP7_75t_R _29317_ (.A(net21),
    .B(_06476_),
    .Y(_06493_));
 INVx3_ASAP7_75t_R _29318_ (.A(_00408_),
    .Y(_06494_));
 BUFx6f_ASAP7_75t_R _29319_ (.A(_06438_),
    .Y(_06495_));
 BUFx6f_ASAP7_75t_R _29320_ (.A(_06454_),
    .Y(_06496_));
 AOI21x1_ASAP7_75t_R _29321_ (.A1(_06494_),
    .A2(_06495_),
    .B(_06496_),
    .Y(_06497_));
 AOI21x1_ASAP7_75t_R _29322_ (.A1(_06443_),
    .A2(_06445_),
    .B(_01263_),
    .Y(_06498_));
 AO21x2_ASAP7_75t_R _29323_ (.A1(_06496_),
    .A2(_06498_),
    .B(_06471_),
    .Y(_06499_));
 AOI21x1_ASAP7_75t_R _29324_ (.A1(_06493_),
    .A2(_06497_),
    .B(_06499_),
    .Y(_06500_));
 BUFx4f_ASAP7_75t_R _29325_ (.A(_06436_),
    .Y(_06501_));
 BUFx4f_ASAP7_75t_R _29326_ (.A(_06435_),
    .Y(_06502_));
 AND2x2_ASAP7_75t_R _29327_ (.A(_01263_),
    .B(_01264_),
    .Y(_06503_));
 AO21x1_ASAP7_75t_R _29328_ (.A1(_06501_),
    .A2(_06502_),
    .B(_06503_),
    .Y(_06504_));
 BUFx6f_ASAP7_75t_R _29329_ (.A(_06475_),
    .Y(_16048_));
 OAI21x1_ASAP7_75t_R _29330_ (.A1(net26),
    .A2(_16052_),
    .B(_16057_),
    .Y(_06505_));
 BUFx6f_ASAP7_75t_R _29331_ (.A(_06454_),
    .Y(_06506_));
 BUFx6f_ASAP7_75t_R _29332_ (.A(_06506_),
    .Y(_06507_));
 AOI21x1_ASAP7_75t_R _29333_ (.A1(_06504_),
    .A2(_06505_),
    .B(_06507_),
    .Y(_06508_));
 NOR2x2_ASAP7_75t_R _29334_ (.A(net511),
    .B(_06438_),
    .Y(_06509_));
 BUFx6f_ASAP7_75t_R _29335_ (.A(_06455_),
    .Y(_06510_));
 OAI21x1_ASAP7_75t_R _29336_ (.A1(_16057_),
    .A2(_16052_),
    .B(_06510_),
    .Y(_06511_));
 BUFx6f_ASAP7_75t_R _29337_ (.A(_06471_),
    .Y(_06512_));
 OAI21x1_ASAP7_75t_R _29338_ (.A1(_06509_),
    .A2(_06511_),
    .B(_06512_),
    .Y(_06513_));
 XOR2x2_ASAP7_75t_R _29339_ (.A(_06470_),
    .B(_01085_),
    .Y(_06514_));
 BUFx6f_ASAP7_75t_R _29340_ (.A(_06514_),
    .Y(_06515_));
 AOI21x1_ASAP7_75t_R _29341_ (.A1(_06502_),
    .A2(_06501_),
    .B(net484),
    .Y(_06516_));
 NAND2x1_ASAP7_75t_R _29342_ (.A(_06450_),
    .B(_03659_),
    .Y(_06517_));
 AOI21x1_ASAP7_75t_R _29343_ (.A1(_06447_),
    .A2(_06448_),
    .B(_11441_),
    .Y(_06518_));
 NAND2x1_ASAP7_75t_R _29344_ (.A(_06517_),
    .B(_06518_),
    .Y(_06519_));
 AOI21x1_ASAP7_75t_R _29345_ (.A1(_06452_),
    .A2(_06519_),
    .B(_08047_),
    .Y(_06520_));
 INVx1_ASAP7_75t_R _29346_ (.A(_08047_),
    .Y(_06521_));
 NOR2x2_ASAP7_75t_R _29347_ (.A(_06521_),
    .B(_06453_),
    .Y(_06522_));
 OAI21x1_ASAP7_75t_R _29348_ (.A1(_06520_),
    .A2(_06522_),
    .B(_01268_),
    .Y(_06523_));
 OAI21x1_ASAP7_75t_R _29349_ (.A1(_06510_),
    .A2(net482),
    .B(_06523_),
    .Y(_06524_));
 BUFx10_ASAP7_75t_R _29350_ (.A(_06490_),
    .Y(_06525_));
 AOI21x1_ASAP7_75t_R _29351_ (.A1(_06515_),
    .A2(_06524_),
    .B(_06525_),
    .Y(_06526_));
 OAI21x1_ASAP7_75t_R _29352_ (.A1(_06508_),
    .A2(_06513_),
    .B(_06526_),
    .Y(_06527_));
 OAI21x1_ASAP7_75t_R _29353_ (.A1(_06492_),
    .A2(_06500_),
    .B(_06527_),
    .Y(_06528_));
 XOR2x1_ASAP7_75t_R _29354_ (.A(_00753_),
    .Y(_06529_),
    .B(_00754_));
 XOR2x1_ASAP7_75t_R _29355_ (.A(_06529_),
    .Y(_06530_),
    .B(_12260_));
 XOR2x1_ASAP7_75t_R _29356_ (.A(_06530_),
    .Y(_06531_),
    .B(_12220_));
 NOR2x1_ASAP7_75t_R _29357_ (.A(_10761_),
    .B(_00687_),
    .Y(_06532_));
 AO21x1_ASAP7_75t_R _29358_ (.A1(_06531_),
    .A2(_10734_),
    .B(_06532_),
    .Y(_06533_));
 XOR2x2_ASAP7_75t_R _29359_ (.A(_06533_),
    .B(_01087_),
    .Y(_06534_));
 BUFx10_ASAP7_75t_R _29360_ (.A(_06534_),
    .Y(_06535_));
 AO21x1_ASAP7_75t_R _29361_ (.A1(_06501_),
    .A2(_06502_),
    .B(_06494_),
    .Y(_06536_));
 BUFx4f_ASAP7_75t_R _29362_ (.A(_06536_),
    .Y(_06537_));
 NAND2x2_ASAP7_75t_R _29363_ (.A(_06446_),
    .B(_06421_),
    .Y(_06538_));
 NOR2x2_ASAP7_75t_R _29364_ (.A(_06520_),
    .B(_06522_),
    .Y(_06539_));
 BUFx6f_ASAP7_75t_R _29365_ (.A(_06539_),
    .Y(_06540_));
 BUFx6f_ASAP7_75t_R _29366_ (.A(_06540_),
    .Y(_06541_));
 AOI21x1_ASAP7_75t_R _29367_ (.A1(_06537_),
    .A2(_06538_),
    .B(_06541_),
    .Y(_06542_));
 AOI21x1_ASAP7_75t_R _29368_ (.A1(_06478_),
    .A2(_16050_),
    .B(_06496_),
    .Y(_06543_));
 INVx1_ASAP7_75t_R _29369_ (.A(_06543_),
    .Y(_06544_));
 OAI21x1_ASAP7_75t_R _29370_ (.A1(net483),
    .A2(_06544_),
    .B(_06512_),
    .Y(_06545_));
 INVx3_ASAP7_75t_R _29371_ (.A(_00640_),
    .Y(_06546_));
 AOI21x1_ASAP7_75t_R _29372_ (.A1(_06502_),
    .A2(_06501_),
    .B(_06546_),
    .Y(_06547_));
 BUFx6f_ASAP7_75t_R _29373_ (.A(_06539_),
    .Y(_06548_));
 BUFx6f_ASAP7_75t_R _29374_ (.A(_06548_),
    .Y(_06549_));
 OAI21x1_ASAP7_75t_R _29375_ (.A1(_06498_),
    .A2(_06547_),
    .B(_06549_),
    .Y(_06550_));
 OAI21x1_ASAP7_75t_R _29376_ (.A1(_06463_),
    .A2(_06464_),
    .B(net917),
    .Y(_06551_));
 BUFx6f_ASAP7_75t_R _29377_ (.A(_06471_),
    .Y(_06552_));
 AOI21x1_ASAP7_75t_R _29378_ (.A1(_06510_),
    .A2(_06551_),
    .B(_06552_),
    .Y(_06553_));
 CKINVDCx5p33_ASAP7_75t_R _29379_ (.A(_06490_),
    .Y(_06554_));
 AOI21x1_ASAP7_75t_R _29380_ (.A1(_06550_),
    .A2(_06553_),
    .B(_06554_),
    .Y(_06555_));
 OAI21x1_ASAP7_75t_R _29381_ (.A1(_06542_),
    .A2(_06545_),
    .B(_06555_),
    .Y(_06556_));
 BUFx6f_ASAP7_75t_R _29382_ (.A(_06548_),
    .Y(_06557_));
 AOI21x1_ASAP7_75t_R _29383_ (.A1(_06435_),
    .A2(_06436_),
    .B(_01264_),
    .Y(_06558_));
 BUFx6f_ASAP7_75t_R _29384_ (.A(_06514_),
    .Y(_06559_));
 AO21x1_ASAP7_75t_R _29385_ (.A1(_06557_),
    .A2(net593),
    .B(_06559_),
    .Y(_06560_));
 NAND2x2_ASAP7_75t_R _29386_ (.A(net633),
    .B(net891),
    .Y(_06561_));
 AOI21x1_ASAP7_75t_R _29387_ (.A1(_06438_),
    .A2(net807),
    .B(_06548_),
    .Y(_06562_));
 OAI21x1_ASAP7_75t_R _29388_ (.A1(_16060_),
    .A2(_06561_),
    .B(_06562_),
    .Y(_06563_));
 INVx1_ASAP7_75t_R _29389_ (.A(_06563_),
    .Y(_06564_));
 AOI21x1_ASAP7_75t_R _29390_ (.A1(_06443_),
    .A2(_06445_),
    .B(_01265_),
    .Y(_06565_));
 OAI21x1_ASAP7_75t_R _29391_ (.A1(_06558_),
    .A2(net846),
    .B(_06549_),
    .Y(_06566_));
 BUFx6f_ASAP7_75t_R _29392_ (.A(_06455_),
    .Y(_06567_));
 INVx3_ASAP7_75t_R _29393_ (.A(net484),
    .Y(_06568_));
 AOI21x1_ASAP7_75t_R _29394_ (.A1(_06443_),
    .A2(_06445_),
    .B(_06568_),
    .Y(_06569_));
 INVx2_ASAP7_75t_R _29395_ (.A(_06569_),
    .Y(_06570_));
 BUFx6f_ASAP7_75t_R _29396_ (.A(_06570_),
    .Y(_06571_));
 AOI21x1_ASAP7_75t_R _29397_ (.A1(_06567_),
    .A2(_06571_),
    .B(_06552_),
    .Y(_06572_));
 AOI21x1_ASAP7_75t_R _29398_ (.A1(_06566_),
    .A2(_06572_),
    .B(_06525_),
    .Y(_06573_));
 OAI21x1_ASAP7_75t_R _29399_ (.A1(_06560_),
    .A2(_06564_),
    .B(_06573_),
    .Y(_06574_));
 AOI21x1_ASAP7_75t_R _29400_ (.A1(_06574_),
    .A2(_06556_),
    .B(_06535_),
    .Y(_06575_));
 XOR2x1_ASAP7_75t_R _29401_ (.A(_00754_),
    .Y(_06576_),
    .B(_12085_));
 XOR2x1_ASAP7_75t_R _29402_ (.A(_06576_),
    .Y(_06577_),
    .B(_00850_));
 XOR2x1_ASAP7_75t_R _29403_ (.A(_06577_),
    .Y(_06578_),
    .B(_12279_));
 NOR2x1_ASAP7_75t_R _29404_ (.A(_10830_),
    .B(_00686_),
    .Y(_06579_));
 AO21x1_ASAP7_75t_R _29405_ (.A1(_06578_),
    .A2(_10830_),
    .B(_06579_),
    .Y(_06580_));
 XOR2x2_ASAP7_75t_R _29406_ (.A(_06580_),
    .B(_01088_),
    .Y(_06581_));
 BUFx10_ASAP7_75t_R _29407_ (.A(_06581_),
    .Y(_06582_));
 AOI211x1_ASAP7_75t_R _29408_ (.A1(_06528_),
    .A2(_06535_),
    .B(_06575_),
    .C(_06582_),
    .Y(_06583_));
 BUFx6f_ASAP7_75t_R _29409_ (.A(_06514_),
    .Y(_06584_));
 AOI21x1_ASAP7_75t_R _29410_ (.A1(_06495_),
    .A2(net809),
    .B(_06496_),
    .Y(_06585_));
 NOR2x1_ASAP7_75t_R _29411_ (.A(_06584_),
    .B(_06585_),
    .Y(_06586_));
 AO21x2_ASAP7_75t_R _29412_ (.A1(_06445_),
    .A2(_06443_),
    .B(_01264_),
    .Y(_06587_));
 INVx1_ASAP7_75t_R _29413_ (.A(_06587_),
    .Y(_06588_));
 AOI21x1_ASAP7_75t_R _29414_ (.A1(_16050_),
    .A2(net808),
    .B(_06478_),
    .Y(_06589_));
 OAI21x1_ASAP7_75t_R _29415_ (.A1(_06588_),
    .A2(_06589_),
    .B(_06510_),
    .Y(_06590_));
 AOI21x1_ASAP7_75t_R _29416_ (.A1(_06586_),
    .A2(_06590_),
    .B(_06554_),
    .Y(_06591_));
 INVx2_ASAP7_75t_R _29417_ (.A(_06538_),
    .Y(_06592_));
 BUFx6f_ASAP7_75t_R _29418_ (.A(_06548_),
    .Y(_06593_));
 OAI21x1_ASAP7_75t_R _29419_ (.A1(_06589_),
    .A2(_06592_),
    .B(_06593_),
    .Y(_06594_));
 INVx1_ASAP7_75t_R _29420_ (.A(_01266_),
    .Y(_06595_));
 AO21x2_ASAP7_75t_R _29421_ (.A1(_06436_),
    .A2(_06435_),
    .B(_06595_),
    .Y(_06596_));
 AND2x2_ASAP7_75t_R _29422_ (.A(_06596_),
    .B(_06496_),
    .Y(_06597_));
 AOI21x1_ASAP7_75t_R _29423_ (.A1(net22),
    .A2(_06597_),
    .B(_06552_),
    .Y(_06598_));
 NAND2x1_ASAP7_75t_R _29424_ (.A(_06594_),
    .B(_06598_),
    .Y(_06599_));
 NAND2x1_ASAP7_75t_R _29425_ (.A(_06591_),
    .B(_06599_),
    .Y(_06600_));
 NOR2x2_ASAP7_75t_R _29426_ (.A(_06438_),
    .B(net633),
    .Y(_06601_));
 NAND2x2_ASAP7_75t_R _29427_ (.A(_06438_),
    .B(net633),
    .Y(_06602_));
 OAI21x1_ASAP7_75t_R _29428_ (.A1(_16052_),
    .A2(_06602_),
    .B(_06540_),
    .Y(_06603_));
 NOR2x2_ASAP7_75t_R _29429_ (.A(_06595_),
    .B(_06438_),
    .Y(_06604_));
 INVx3_ASAP7_75t_R _29430_ (.A(_06604_),
    .Y(_06605_));
 AOI21x1_ASAP7_75t_R _29431_ (.A1(_06605_),
    .A2(_06562_),
    .B(_06552_),
    .Y(_06606_));
 OAI21x1_ASAP7_75t_R _29432_ (.A1(_06601_),
    .A2(_06603_),
    .B(_06606_),
    .Y(_06607_));
 NAND2x2_ASAP7_75t_R _29433_ (.A(_06438_),
    .B(net628),
    .Y(_06608_));
 INVx1_ASAP7_75t_R _29434_ (.A(_06608_),
    .Y(_06609_));
 AOI21x1_ASAP7_75t_R _29435_ (.A1(_06593_),
    .A2(_06609_),
    .B(_06472_),
    .Y(_06610_));
 AOI21x1_ASAP7_75t_R _29436_ (.A1(_06563_),
    .A2(_06610_),
    .B(_06525_),
    .Y(_06611_));
 NAND2x1_ASAP7_75t_R _29437_ (.A(_06607_),
    .B(_06611_),
    .Y(_06612_));
 AOI21x1_ASAP7_75t_R _29438_ (.A1(_06600_),
    .A2(_06612_),
    .B(_06535_),
    .Y(_06613_));
 AOI21x1_ASAP7_75t_R _29439_ (.A1(_06502_),
    .A2(_06501_),
    .B(_06568_),
    .Y(_06614_));
 INVx2_ASAP7_75t_R _29440_ (.A(_06614_),
    .Y(_06615_));
 BUFx6f_ASAP7_75t_R _29441_ (.A(_06471_),
    .Y(_06616_));
 AO21x1_ASAP7_75t_R _29442_ (.A1(_06615_),
    .A2(_06506_),
    .B(_06616_),
    .Y(_06617_));
 AOI21x1_ASAP7_75t_R _29443_ (.A1(net22),
    .A2(_06608_),
    .B(_06567_),
    .Y(_06618_));
 BUFx6f_ASAP7_75t_R _29444_ (.A(_06554_),
    .Y(_06619_));
 OAI21x1_ASAP7_75t_R _29445_ (.A1(_06617_),
    .A2(_06618_),
    .B(_06619_),
    .Y(_06620_));
 INVx3_ASAP7_75t_R _29446_ (.A(_06509_),
    .Y(_06621_));
 NAND2x1_ASAP7_75t_R _29447_ (.A(_06621_),
    .B(_06497_),
    .Y(_06622_));
 AO21x2_ASAP7_75t_R _29448_ (.A1(_06445_),
    .A2(_06443_),
    .B(net485),
    .Y(_06623_));
 INVx2_ASAP7_75t_R _29449_ (.A(_06547_),
    .Y(_06624_));
 AO21x1_ASAP7_75t_R _29450_ (.A1(_06623_),
    .A2(_06624_),
    .B(_06593_),
    .Y(_06625_));
 AOI21x1_ASAP7_75t_R _29451_ (.A1(_06622_),
    .A2(_06625_),
    .B(_06515_),
    .Y(_06626_));
 BUFx10_ASAP7_75t_R _29452_ (.A(_06534_),
    .Y(_06627_));
 OAI21x1_ASAP7_75t_R _29453_ (.A1(_06620_),
    .A2(_06626_),
    .B(_06627_),
    .Y(_06628_));
 NAND2x2_ASAP7_75t_R _29454_ (.A(_16048_),
    .B(net556),
    .Y(_06629_));
 AOI21x1_ASAP7_75t_R _29455_ (.A1(_06478_),
    .A2(net891),
    .B(_06454_),
    .Y(_06630_));
 NAND2x2_ASAP7_75t_R _29456_ (.A(_06629_),
    .B(_06630_),
    .Y(_06631_));
 NAND2x2_ASAP7_75t_R _29457_ (.A(_06438_),
    .B(net891),
    .Y(_06632_));
 AOI21x1_ASAP7_75t_R _29458_ (.A1(_16050_),
    .A2(net21),
    .B(_06548_),
    .Y(_06633_));
 AOI21x1_ASAP7_75t_R _29459_ (.A1(_06632_),
    .A2(_06633_),
    .B(_06616_),
    .Y(_06634_));
 NAND2x1_ASAP7_75t_R _29460_ (.A(_06631_),
    .B(_06634_),
    .Y(_06635_));
 NOR2x2_ASAP7_75t_R _29461_ (.A(_06496_),
    .B(net821),
    .Y(_06636_));
 OAI21x1_ASAP7_75t_R _29462_ (.A1(net23),
    .A2(_06602_),
    .B(_06636_),
    .Y(_06637_));
 NOR2x2_ASAP7_75t_R _29463_ (.A(_06494_),
    .B(_06495_),
    .Y(_06638_));
 OAI21x1_ASAP7_75t_R _29464_ (.A1(_06547_),
    .A2(_06638_),
    .B(_06510_),
    .Y(_06639_));
 NAND3x1_ASAP7_75t_R _29465_ (.A(_06637_),
    .B(_06512_),
    .C(_06639_),
    .Y(_06640_));
 BUFx6f_ASAP7_75t_R _29466_ (.A(_06554_),
    .Y(_06641_));
 AOI21x1_ASAP7_75t_R _29467_ (.A1(_06635_),
    .A2(_06640_),
    .B(_06641_),
    .Y(_06642_));
 OAI21x1_ASAP7_75t_R _29468_ (.A1(_06642_),
    .A2(_06628_),
    .B(_06582_),
    .Y(_06643_));
 NOR2x1_ASAP7_75t_R _29469_ (.A(_06643_),
    .B(_06613_),
    .Y(_06644_));
 NOR2x1_ASAP7_75t_R _29470_ (.A(_06583_),
    .B(_06644_),
    .Y(_00144_));
 NOR2x2_ASAP7_75t_R _29471_ (.A(_06614_),
    .B(_06548_),
    .Y(_06645_));
 NAND2x1_ASAP7_75t_R _29472_ (.A(_06645_),
    .B(_06621_),
    .Y(_06646_));
 BUFx6f_ASAP7_75t_R _29473_ (.A(_06490_),
    .Y(_06647_));
 NAND2x1_ASAP7_75t_R _29474_ (.A(_06593_),
    .B(_06498_),
    .Y(_06648_));
 NAND3x2_ASAP7_75t_R _29475_ (.B(_06540_),
    .C(_16060_),
    .Y(_06649_),
    .A(_16052_));
 AND4x1_ASAP7_75t_R _29476_ (.A(_06646_),
    .B(_06647_),
    .C(_06648_),
    .D(_06649_),
    .Y(_06650_));
 AOI21x1_ASAP7_75t_R _29477_ (.A1(_16050_),
    .A2(net891),
    .B(_16057_),
    .Y(_06651_));
 OAI21x1_ASAP7_75t_R _29478_ (.A1(_06569_),
    .A2(_06651_),
    .B(_06567_),
    .Y(_06652_));
 AO21x2_ASAP7_75t_R _29479_ (.A1(_06501_),
    .A2(_06502_),
    .B(_06465_),
    .Y(_06653_));
 AOI21x1_ASAP7_75t_R _29480_ (.A1(_01266_),
    .A2(_06478_),
    .B(_06496_),
    .Y(_06654_));
 AOI21x1_ASAP7_75t_R _29481_ (.A1(_06653_),
    .A2(_06654_),
    .B(_06647_),
    .Y(_06655_));
 BUFx6f_ASAP7_75t_R _29482_ (.A(_06616_),
    .Y(_06656_));
 AO21x1_ASAP7_75t_R _29483_ (.A1(_06652_),
    .A2(_06655_),
    .B(_06656_),
    .Y(_06657_));
 OAI21x1_ASAP7_75t_R _29484_ (.A1(_06568_),
    .A2(_06438_),
    .B(_06454_),
    .Y(_06658_));
 INVx1_ASAP7_75t_R _29485_ (.A(_06658_),
    .Y(_06659_));
 NOR2x1_ASAP7_75t_R _29486_ (.A(_06647_),
    .B(_06659_),
    .Y(_06660_));
 OAI21x1_ASAP7_75t_R _29487_ (.A1(_16060_),
    .A2(_06561_),
    .B(_06585_),
    .Y(_06661_));
 AOI21x1_ASAP7_75t_R _29488_ (.A1(_06660_),
    .A2(_06661_),
    .B(_06515_),
    .Y(_06662_));
 NAND2x2_ASAP7_75t_R _29489_ (.A(_06478_),
    .B(net555),
    .Y(_06663_));
 BUFx6f_ASAP7_75t_R _29490_ (.A(_06454_),
    .Y(_06664_));
 AO21x1_ASAP7_75t_R _29491_ (.A1(_06663_),
    .A2(_06624_),
    .B(_06664_),
    .Y(_06665_));
 AND2x2_ASAP7_75t_R _29492_ (.A(_06551_),
    .B(_06496_),
    .Y(_06666_));
 AOI21x1_ASAP7_75t_R _29493_ (.A1(_06608_),
    .A2(_06666_),
    .B(_06554_),
    .Y(_06667_));
 NAND2x1_ASAP7_75t_R _29494_ (.A(_06665_),
    .B(_06667_),
    .Y(_06668_));
 AOI21x1_ASAP7_75t_R _29495_ (.A1(_06662_),
    .A2(_06668_),
    .B(_06534_),
    .Y(_06669_));
 OAI21x1_ASAP7_75t_R _29496_ (.A1(_06650_),
    .A2(_06657_),
    .B(_06669_),
    .Y(_06670_));
 NAND2x2_ASAP7_75t_R _29497_ (.A(_06478_),
    .B(net634),
    .Y(_06671_));
 OAI21x1_ASAP7_75t_R _29498_ (.A1(_16047_),
    .A2(_06671_),
    .B(_06497_),
    .Y(_06672_));
 INVx1_ASAP7_75t_R _29499_ (.A(_00405_),
    .Y(_06673_));
 OR3x1_ASAP7_75t_R _29500_ (.A(_06490_),
    .B(_06673_),
    .C(_06540_),
    .Y(_06674_));
 NAND2x1_ASAP7_75t_R _29501_ (.A(_06672_),
    .B(_06674_),
    .Y(_06675_));
 INVx2_ASAP7_75t_R _29502_ (.A(_06534_),
    .Y(_06676_));
 BUFx6f_ASAP7_75t_R _29503_ (.A(_06676_),
    .Y(_06677_));
 AOI21x1_ASAP7_75t_R _29504_ (.A1(_06656_),
    .A2(_06675_),
    .B(_06677_),
    .Y(_06678_));
 BUFx6f_ASAP7_75t_R _29505_ (.A(_06647_),
    .Y(_06679_));
 AO22x1_ASAP7_75t_R _29506_ (.A1(_06602_),
    .A2(_06630_),
    .B1(_06666_),
    .B2(_06608_),
    .Y(_06680_));
 AOI21x1_ASAP7_75t_R _29507_ (.A1(_16050_),
    .A2(net891),
    .B(_06495_),
    .Y(_06681_));
 OAI21x1_ASAP7_75t_R _29508_ (.A1(_06681_),
    .A2(_06589_),
    .B(_06567_),
    .Y(_06682_));
 OA21x2_ASAP7_75t_R _29509_ (.A1(_16057_),
    .A2(net511),
    .B(_06548_),
    .Y(_06683_));
 AOI21x1_ASAP7_75t_R _29510_ (.A1(_06663_),
    .A2(_06683_),
    .B(_06554_),
    .Y(_06684_));
 AOI21x1_ASAP7_75t_R _29511_ (.A1(_06682_),
    .A2(_06684_),
    .B(_06656_),
    .Y(_06685_));
 OAI21x1_ASAP7_75t_R _29512_ (.A1(_06679_),
    .A2(_06680_),
    .B(_06685_),
    .Y(_06686_));
 INVx5_ASAP7_75t_R _29513_ (.A(_06581_),
    .Y(_06687_));
 AOI21x1_ASAP7_75t_R _29514_ (.A1(_06678_),
    .A2(_06686_),
    .B(_06687_),
    .Y(_06688_));
 NAND2x1_ASAP7_75t_R _29515_ (.A(_06670_),
    .B(_06688_),
    .Y(_06689_));
 OA21x2_ASAP7_75t_R _29516_ (.A1(_06587_),
    .A2(_06507_),
    .B(_06512_),
    .Y(_06690_));
 NAND2x1_ASAP7_75t_R _29517_ (.A(_06541_),
    .B(_06681_),
    .Y(_06691_));
 NAND2x2_ASAP7_75t_R _29518_ (.A(_06478_),
    .B(net26),
    .Y(_06692_));
 AOI21x1_ASAP7_75t_R _29519_ (.A1(_06692_),
    .A2(_06597_),
    .B(_06512_),
    .Y(_06693_));
 AOI221x1_ASAP7_75t_R _29520_ (.A1(_06690_),
    .A2(_06652_),
    .B1(_06691_),
    .B2(_06693_),
    .C(_06641_),
    .Y(_06694_));
 NOR2x2_ASAP7_75t_R _29521_ (.A(_06455_),
    .B(_06516_),
    .Y(_06695_));
 NAND2x1_ASAP7_75t_R _29522_ (.A(_06695_),
    .B(_06663_),
    .Y(_06696_));
 OAI21x1_ASAP7_75t_R _29523_ (.A1(_16050_),
    .A2(net23),
    .B(_06562_),
    .Y(_06697_));
 BUFx6f_ASAP7_75t_R _29524_ (.A(_06514_),
    .Y(_06698_));
 AOI21x1_ASAP7_75t_R _29525_ (.A1(_06696_),
    .A2(_06697_),
    .B(_06698_),
    .Y(_06699_));
 NOR2x1_ASAP7_75t_R _29526_ (.A(_06558_),
    .B(_06658_),
    .Y(_06700_));
 NOR2x2_ASAP7_75t_R _29527_ (.A(_06546_),
    .B(_06495_),
    .Y(_06701_));
 AO21x1_ASAP7_75t_R _29528_ (.A1(_16052_),
    .A2(_06495_),
    .B(_06455_),
    .Y(_06702_));
 OAI21x1_ASAP7_75t_R _29529_ (.A1(_06701_),
    .A2(_06702_),
    .B(_06559_),
    .Y(_06703_));
 NOR2x1_ASAP7_75t_R _29530_ (.A(_06700_),
    .B(_06703_),
    .Y(_06704_));
 OAI21x1_ASAP7_75t_R _29531_ (.A1(_06699_),
    .A2(_06704_),
    .B(_06641_),
    .Y(_06705_));
 NAND2x1_ASAP7_75t_R _29532_ (.A(_06677_),
    .B(_06705_),
    .Y(_06706_));
 AOI21x1_ASAP7_75t_R _29533_ (.A1(_06664_),
    .A2(_06602_),
    .B(_06616_),
    .Y(_06707_));
 AOI21x1_ASAP7_75t_R _29534_ (.A1(_06557_),
    .A2(net593),
    .B(_06601_),
    .Y(_06708_));
 AOI21x1_ASAP7_75t_R _29535_ (.A1(_06707_),
    .A2(_06708_),
    .B(_06525_),
    .Y(_06709_));
 NAND2x2_ASAP7_75t_R _29536_ (.A(net633),
    .B(net807),
    .Y(_06710_));
 AOI21x1_ASAP7_75t_R _29537_ (.A1(_16057_),
    .A2(_06710_),
    .B(net593),
    .Y(_06711_));
 AOI21x1_ASAP7_75t_R _29538_ (.A1(_06645_),
    .A2(_06605_),
    .B(_06559_),
    .Y(_06712_));
 OAI21x1_ASAP7_75t_R _29539_ (.A1(_06507_),
    .A2(_06711_),
    .B(_06712_),
    .Y(_06713_));
 AOI21x1_ASAP7_75t_R _29540_ (.A1(_06709_),
    .A2(_06713_),
    .B(_06677_),
    .Y(_06714_));
 BUFx10_ASAP7_75t_R _29541_ (.A(_06584_),
    .Y(_06715_));
 NOR2x2_ASAP7_75t_R _29542_ (.A(_06478_),
    .B(_06539_),
    .Y(_06716_));
 NAND2x1_ASAP7_75t_R _29543_ (.A(_06716_),
    .B(_06710_),
    .Y(_06717_));
 NAND2x1_ASAP7_75t_R _29544_ (.A(_06629_),
    .B(_06543_),
    .Y(_06718_));
 NAND2x1_ASAP7_75t_R _29545_ (.A(_06717_),
    .B(_06718_),
    .Y(_06719_));
 NOR2x1_ASAP7_75t_R _29546_ (.A(_16057_),
    .B(_16052_),
    .Y(_06720_));
 OAI21x1_ASAP7_75t_R _29547_ (.A1(_06588_),
    .A2(_06720_),
    .B(_06557_),
    .Y(_06721_));
 BUFx6f_ASAP7_75t_R _29548_ (.A(_06471_),
    .Y(_06722_));
 AOI21x1_ASAP7_75t_R _29549_ (.A1(net22),
    .A2(_06562_),
    .B(_06722_),
    .Y(_06723_));
 AOI21x1_ASAP7_75t_R _29550_ (.A1(_06723_),
    .A2(_06721_),
    .B(_06619_),
    .Y(_06724_));
 OAI21x1_ASAP7_75t_R _29551_ (.A1(_06715_),
    .A2(_06719_),
    .B(_06724_),
    .Y(_06725_));
 AOI21x1_ASAP7_75t_R _29552_ (.A1(_06714_),
    .A2(_06725_),
    .B(_06582_),
    .Y(_06726_));
 OAI21x1_ASAP7_75t_R _29553_ (.A1(_06694_),
    .A2(_06706_),
    .B(_06726_),
    .Y(_06727_));
 NAND2x1_ASAP7_75t_R _29554_ (.A(_06689_),
    .B(_06727_),
    .Y(_00145_));
 OA21x2_ASAP7_75t_R _29555_ (.A1(_16060_),
    .A2(_00641_),
    .B(_06540_),
    .Y(_06728_));
 NAND2x1_ASAP7_75t_R _29556_ (.A(_06608_),
    .B(_06728_),
    .Y(_06729_));
 AO21x2_ASAP7_75t_R _29557_ (.A1(_06501_),
    .A2(_06502_),
    .B(_01263_),
    .Y(_06730_));
 NAND3x1_ASAP7_75t_R _29558_ (.A(_06538_),
    .B(_06507_),
    .C(_06730_),
    .Y(_06731_));
 AOI21x1_ASAP7_75t_R _29559_ (.A1(_06729_),
    .A2(_06731_),
    .B(_06656_),
    .Y(_06732_));
 NAND2x1_ASAP7_75t_R _29560_ (.A(_06656_),
    .B(_06603_),
    .Y(_06733_));
 OAI21x1_ASAP7_75t_R _29561_ (.A1(_16047_),
    .A2(_06602_),
    .B(_06567_),
    .Y(_06734_));
 NOR2x1_ASAP7_75t_R _29562_ (.A(_06604_),
    .B(_06734_),
    .Y(_06735_));
 OAI21x1_ASAP7_75t_R _29563_ (.A1(_06733_),
    .A2(_06735_),
    .B(_06679_),
    .Y(_06736_));
 OAI21x1_ASAP7_75t_R _29564_ (.A1(_06732_),
    .A2(_06736_),
    .B(_06535_),
    .Y(_06737_));
 OAI21x1_ASAP7_75t_R _29565_ (.A1(_16057_),
    .A2(net21),
    .B(_16050_),
    .Y(_06738_));
 NAND2x1_ASAP7_75t_R _29566_ (.A(_06567_),
    .B(_06738_),
    .Y(_06739_));
 AO21x2_ASAP7_75t_R _29567_ (.A1(_06501_),
    .A2(_06502_),
    .B(_01266_),
    .Y(_06740_));
 AO21x1_ASAP7_75t_R _29568_ (.A1(_06740_),
    .A2(_06587_),
    .B(_06567_),
    .Y(_06741_));
 AO21x1_ASAP7_75t_R _29569_ (.A1(_06739_),
    .A2(_06741_),
    .B(_06656_),
    .Y(_06742_));
 INVx3_ASAP7_75t_R _29570_ (.A(net482),
    .Y(_06743_));
 NAND2x1_ASAP7_75t_R _29571_ (.A(_06743_),
    .B(_06543_),
    .Y(_06744_));
 AOI21x1_ASAP7_75t_R _29572_ (.A1(_06507_),
    .A2(_06711_),
    .B(_06515_),
    .Y(_06745_));
 NAND2x1_ASAP7_75t_R _29573_ (.A(_06744_),
    .B(_06745_),
    .Y(_06746_));
 AOI21x1_ASAP7_75t_R _29574_ (.A1(_06742_),
    .A2(_06746_),
    .B(_06679_),
    .Y(_06747_));
 OAI21x1_ASAP7_75t_R _29575_ (.A1(_06737_),
    .A2(_06747_),
    .B(_06582_),
    .Y(_06748_));
 AOI21x1_ASAP7_75t_R _29576_ (.A1(_06495_),
    .A2(_16048_),
    .B(_06548_),
    .Y(_06749_));
 INVx2_ASAP7_75t_R _29577_ (.A(_06565_),
    .Y(_06750_));
 AND2x2_ASAP7_75t_R _29578_ (.A(_06749_),
    .B(_06750_),
    .Y(_06751_));
 INVx2_ASAP7_75t_R _29579_ (.A(_06740_),
    .Y(_06752_));
 BUFx6f_ASAP7_75t_R _29580_ (.A(_06539_),
    .Y(_06753_));
 OAI21x1_ASAP7_75t_R _29581_ (.A1(_16060_),
    .A2(net21),
    .B(_06753_),
    .Y(_06754_));
 OAI21x1_ASAP7_75t_R _29582_ (.A1(_06752_),
    .A2(_06754_),
    .B(_06559_),
    .Y(_06755_));
 NOR2x1_ASAP7_75t_R _29583_ (.A(_06751_),
    .B(_06755_),
    .Y(_06756_));
 AOI21x1_ASAP7_75t_R _29584_ (.A1(_01265_),
    .A2(_06495_),
    .B(_06496_),
    .Y(_06757_));
 NAND2x1_ASAP7_75t_R _29585_ (.A(_06663_),
    .B(_06757_),
    .Y(_06758_));
 AO21x1_ASAP7_75t_R _29586_ (.A1(_06623_),
    .A2(_06615_),
    .B(_06549_),
    .Y(_06759_));
 AOI21x1_ASAP7_75t_R _29587_ (.A1(_06758_),
    .A2(_06759_),
    .B(_06698_),
    .Y(_06760_));
 OA21x2_ASAP7_75t_R _29588_ (.A1(_06756_),
    .A2(_06760_),
    .B(_06679_),
    .Y(_06761_));
 INVx1_ASAP7_75t_R _29589_ (.A(_06566_),
    .Y(_06762_));
 INVx3_ASAP7_75t_R _29590_ (.A(_06558_),
    .Y(_06763_));
 AOI21x1_ASAP7_75t_R _29591_ (.A1(_06763_),
    .A2(_06671_),
    .B(_06541_),
    .Y(_06764_));
 OAI21x1_ASAP7_75t_R _29592_ (.A1(_06762_),
    .A2(_06764_),
    .B(_06656_),
    .Y(_06765_));
 AOI21x1_ASAP7_75t_R _29593_ (.A1(_06763_),
    .A2(_06538_),
    .B(_06541_),
    .Y(_06766_));
 OA21x2_ASAP7_75t_R _29594_ (.A1(_06752_),
    .A2(net846),
    .B(_06541_),
    .Y(_06767_));
 OAI21x1_ASAP7_75t_R _29595_ (.A1(_06766_),
    .A2(_06767_),
    .B(_06715_),
    .Y(_06768_));
 AOI21x1_ASAP7_75t_R _29596_ (.A1(_06765_),
    .A2(_06768_),
    .B(_06679_),
    .Y(_06769_));
 NOR3x2_ASAP7_75t_R _29597_ (.B(_06769_),
    .C(_06535_),
    .Y(_06770_),
    .A(_06761_));
 OA21x2_ASAP7_75t_R _29598_ (.A1(net26),
    .A2(_06495_),
    .B(_06455_),
    .Y(_06771_));
 AOI21x1_ASAP7_75t_R _29599_ (.A1(_06629_),
    .A2(_06771_),
    .B(_06584_),
    .Y(_06772_));
 OA21x2_ASAP7_75t_R _29600_ (.A1(_06673_),
    .A2(_06507_),
    .B(_06772_),
    .Y(_06773_));
 NOR2x1_ASAP7_75t_R _29601_ (.A(_06557_),
    .B(_06638_),
    .Y(_06774_));
 AOI22x1_ASAP7_75t_R _29602_ (.A1(_06774_),
    .A2(_06743_),
    .B1(_06543_),
    .B2(_06624_),
    .Y(_06775_));
 OAI21x1_ASAP7_75t_R _29603_ (.A1(_06656_),
    .A2(_06775_),
    .B(_06677_),
    .Y(_06776_));
 NOR2x1_ASAP7_75t_R _29604_ (.A(_06773_),
    .B(_06776_),
    .Y(_06777_));
 NAND2x2_ASAP7_75t_R _29605_ (.A(_00406_),
    .B(_06664_),
    .Y(_06778_));
 AOI21x1_ASAP7_75t_R _29606_ (.A1(_06778_),
    .A2(_06603_),
    .B(_06698_),
    .Y(_06779_));
 OR3x1_ASAP7_75t_R _29607_ (.A(_06522_),
    .B(_06520_),
    .C(_01270_),
    .Y(_06780_));
 AOI21x1_ASAP7_75t_R _29608_ (.A1(_06780_),
    .A2(_06739_),
    .B(_06656_),
    .Y(_06781_));
 OAI21x1_ASAP7_75t_R _29609_ (.A1(_06779_),
    .A2(_06781_),
    .B(_06535_),
    .Y(_06782_));
 NAND2x1_ASAP7_75t_R _29610_ (.A(_06641_),
    .B(_06782_),
    .Y(_06783_));
 AO21x1_ASAP7_75t_R _29611_ (.A1(_06445_),
    .A2(_06443_),
    .B(_06503_),
    .Y(_06784_));
 INVx1_ASAP7_75t_R _29612_ (.A(_06784_),
    .Y(_06785_));
 OA21x2_ASAP7_75t_R _29613_ (.A1(_06651_),
    .A2(_06785_),
    .B(_06507_),
    .Y(_06786_));
 NAND2x1_ASAP7_75t_R _29614_ (.A(_06698_),
    .B(_06672_),
    .Y(_06787_));
 AOI21x1_ASAP7_75t_R _29615_ (.A1(_06541_),
    .A2(_06701_),
    .B(_06559_),
    .Y(_06788_));
 AO21x1_ASAP7_75t_R _29616_ (.A1(_06623_),
    .A2(_06763_),
    .B(_06549_),
    .Y(_06789_));
 AOI21x1_ASAP7_75t_R _29617_ (.A1(_06788_),
    .A2(_06789_),
    .B(_06676_),
    .Y(_06790_));
 OAI21x1_ASAP7_75t_R _29618_ (.A1(_06786_),
    .A2(_06787_),
    .B(_06790_),
    .Y(_06791_));
 NAND2x2_ASAP7_75t_R _29619_ (.A(_06663_),
    .B(_06749_),
    .Y(_06792_));
 AOI21x1_ASAP7_75t_R _29620_ (.A1(_06743_),
    .A2(_06543_),
    .B(_06722_),
    .Y(_06793_));
 NAND2x1_ASAP7_75t_R _29621_ (.A(_06792_),
    .B(_06793_),
    .Y(_06794_));
 OA21x2_ASAP7_75t_R _29622_ (.A1(_01268_),
    .A2(_06510_),
    .B(_06552_),
    .Y(_06795_));
 OAI21x1_ASAP7_75t_R _29623_ (.A1(_16052_),
    .A2(_06671_),
    .B(_06645_),
    .Y(_06796_));
 AOI21x1_ASAP7_75t_R _29624_ (.A1(_06795_),
    .A2(_06796_),
    .B(_06534_),
    .Y(_06797_));
 AOI21x1_ASAP7_75t_R _29625_ (.A1(_06794_),
    .A2(_06797_),
    .B(_06641_),
    .Y(_06798_));
 AOI21x1_ASAP7_75t_R _29626_ (.A1(_06791_),
    .A2(_06798_),
    .B(_06582_),
    .Y(_06799_));
 OAI21x1_ASAP7_75t_R _29627_ (.A1(_06777_),
    .A2(_06783_),
    .B(_06799_),
    .Y(_06800_));
 OAI21x1_ASAP7_75t_R _29628_ (.A1(_06748_),
    .A2(_06770_),
    .B(_06800_),
    .Y(_00146_));
 AO21x1_ASAP7_75t_R _29629_ (.A1(_06445_),
    .A2(_06443_),
    .B(_01266_),
    .Y(_06801_));
 AO21x1_ASAP7_75t_R _29630_ (.A1(_06801_),
    .A2(_06763_),
    .B(_06549_),
    .Y(_06802_));
 AOI21x1_ASAP7_75t_R _29631_ (.A1(_06608_),
    .A2(_06728_),
    .B(_06515_),
    .Y(_06803_));
 AOI21x1_ASAP7_75t_R _29632_ (.A1(_06802_),
    .A2(_06803_),
    .B(_06641_),
    .Y(_06804_));
 OA21x2_ASAP7_75t_R _29633_ (.A1(_06546_),
    .A2(_16060_),
    .B(_06645_),
    .Y(_06805_));
 NOR2x1_ASAP7_75t_R _29634_ (.A(_06638_),
    .B(_06702_),
    .Y(_06806_));
 OAI21x1_ASAP7_75t_R _29635_ (.A1(_06805_),
    .A2(_06806_),
    .B(_06715_),
    .Y(_06807_));
 AO21x1_ASAP7_75t_R _29636_ (.A1(_06804_),
    .A2(_06807_),
    .B(_06677_),
    .Y(_06808_));
 AO21x1_ASAP7_75t_R _29637_ (.A1(_06630_),
    .A2(_06710_),
    .B(_06514_),
    .Y(_06809_));
 AO21x1_ASAP7_75t_R _29638_ (.A1(net22),
    .A2(_06749_),
    .B(_06809_),
    .Y(_06810_));
 NAND2x1_ASAP7_75t_R _29639_ (.A(_06506_),
    .B(net828),
    .Y(_06811_));
 NAND2x2_ASAP7_75t_R _29640_ (.A(_06602_),
    .B(_06630_),
    .Y(_06812_));
 NAND2x1_ASAP7_75t_R _29641_ (.A(_06811_),
    .B(_06812_),
    .Y(_06813_));
 AOI21x1_ASAP7_75t_R _29642_ (.A1(_06715_),
    .A2(_06813_),
    .B(_06491_),
    .Y(_06814_));
 AND2x2_ASAP7_75t_R _29643_ (.A(_06810_),
    .B(_06814_),
    .Y(_06815_));
 NOR2x1_ASAP7_75t_R _29644_ (.A(_06808_),
    .B(_06815_),
    .Y(_06816_));
 OAI21x1_ASAP7_75t_R _29645_ (.A1(_06638_),
    .A2(_06589_),
    .B(_06507_),
    .Y(_06817_));
 OAI21x1_ASAP7_75t_R _29646_ (.A1(_06516_),
    .A2(_06681_),
    .B(_06541_),
    .Y(_06818_));
 AOI21x1_ASAP7_75t_R _29647_ (.A1(_06817_),
    .A2(_06818_),
    .B(_06715_),
    .Y(_06819_));
 NAND2x1_ASAP7_75t_R _29648_ (.A(_06537_),
    .B(_06636_),
    .Y(_06820_));
 AND2x2_ASAP7_75t_R _29649_ (.A(_06634_),
    .B(_06820_),
    .Y(_06821_));
 OA21x2_ASAP7_75t_R _29650_ (.A1(_06819_),
    .A2(_06821_),
    .B(_06679_),
    .Y(_06822_));
 AO21x1_ASAP7_75t_R _29651_ (.A1(_06501_),
    .A2(_06502_),
    .B(_01265_),
    .Y(_06823_));
 AO21x1_ASAP7_75t_R _29652_ (.A1(_06823_),
    .A2(_06571_),
    .B(_06567_),
    .Y(_06824_));
 NAND2x1_ASAP7_75t_R _29653_ (.A(_06693_),
    .B(_06824_),
    .Y(_06825_));
 NAND2x1_ASAP7_75t_R _29654_ (.A(_06632_),
    .B(_06629_),
    .Y(_06826_));
 AO21x1_ASAP7_75t_R _29655_ (.A1(_16057_),
    .A2(_06664_),
    .B(_06584_),
    .Y(_06827_));
 OA21x2_ASAP7_75t_R _29656_ (.A1(_06826_),
    .A2(_06827_),
    .B(_06619_),
    .Y(_06828_));
 AO21x1_ASAP7_75t_R _29657_ (.A1(_06828_),
    .A2(_06825_),
    .B(_06535_),
    .Y(_06829_));
 OAI21x1_ASAP7_75t_R _29658_ (.A1(_06822_),
    .A2(_06829_),
    .B(_06687_),
    .Y(_06830_));
 AOI21x1_ASAP7_75t_R _29659_ (.A1(_06596_),
    .A2(_06636_),
    .B(_06722_),
    .Y(_06831_));
 OAI21x1_ASAP7_75t_R _29660_ (.A1(net846),
    .A2(_06720_),
    .B(_06664_),
    .Y(_06832_));
 NAND2x1_ASAP7_75t_R _29661_ (.A(_06831_),
    .B(_06832_),
    .Y(_06833_));
 AOI21x1_ASAP7_75t_R _29662_ (.A1(_06621_),
    .A2(_06562_),
    .B(_06559_),
    .Y(_06834_));
 NAND2x1_ASAP7_75t_R _29663_ (.A(_06718_),
    .B(_06834_),
    .Y(_06835_));
 AOI21x1_ASAP7_75t_R _29664_ (.A1(_06833_),
    .A2(_06835_),
    .B(_06641_),
    .Y(_06836_));
 NAND2x1_ASAP7_75t_R _29665_ (.A(_06619_),
    .B(_06755_),
    .Y(_06837_));
 AO21x1_ASAP7_75t_R _29666_ (.A1(_06823_),
    .A2(_06784_),
    .B(_06753_),
    .Y(_06838_));
 AOI21x1_ASAP7_75t_R _29667_ (.A1(_06672_),
    .A2(_06838_),
    .B(_06698_),
    .Y(_06839_));
 OAI21x1_ASAP7_75t_R _29668_ (.A1(_06837_),
    .A2(_06839_),
    .B(_06677_),
    .Y(_06840_));
 NOR2x1_ASAP7_75t_R _29669_ (.A(_06840_),
    .B(_06836_),
    .Y(_06841_));
 NOR2x2_ASAP7_75t_R _29670_ (.A(_06540_),
    .B(_06750_),
    .Y(_06842_));
 NOR2x1_ASAP7_75t_R _29671_ (.A(_06554_),
    .B(_06842_),
    .Y(_06843_));
 NAND2x1_ASAP7_75t_R _29672_ (.A(_06758_),
    .B(_06843_),
    .Y(_06844_));
 AO21x1_ASAP7_75t_R _29673_ (.A1(_06740_),
    .A2(_06784_),
    .B(_06593_),
    .Y(_06845_));
 AOI21x1_ASAP7_75t_R _29674_ (.A1(_06571_),
    .A2(_06585_),
    .B(_06647_),
    .Y(_06846_));
 NAND2x1_ASAP7_75t_R _29675_ (.A(_06845_),
    .B(_06846_),
    .Y(_06847_));
 AOI21x1_ASAP7_75t_R _29676_ (.A1(_06844_),
    .A2(_06847_),
    .B(_06715_),
    .Y(_06848_));
 NAND2x1_ASAP7_75t_R _29677_ (.A(_06671_),
    .B(_06497_),
    .Y(_06849_));
 AOI21x1_ASAP7_75t_R _29678_ (.A1(_06811_),
    .A2(_06849_),
    .B(_06491_),
    .Y(_06850_));
 NOR2x1_ASAP7_75t_R _29679_ (.A(_06506_),
    .B(_06570_),
    .Y(_06851_));
 AO21x1_ASAP7_75t_R _29680_ (.A1(_06851_),
    .A2(_06525_),
    .B(_06499_),
    .Y(_06852_));
 OAI21x1_ASAP7_75t_R _29681_ (.A1(_06850_),
    .A2(_06852_),
    .B(_06627_),
    .Y(_06853_));
 NOR2x1_ASAP7_75t_R _29682_ (.A(_06848_),
    .B(_06853_),
    .Y(_06854_));
 OAI21x1_ASAP7_75t_R _29683_ (.A1(_06841_),
    .A2(_06854_),
    .B(_06582_),
    .Y(_06855_));
 OAI21x1_ASAP7_75t_R _29684_ (.A1(_06816_),
    .A2(_06830_),
    .B(_06855_),
    .Y(_00147_));
 AOI21x1_ASAP7_75t_R _29685_ (.A1(_06632_),
    .A2(_06633_),
    .B(_06584_),
    .Y(_06856_));
 NOR2x2_ASAP7_75t_R _29686_ (.A(net26),
    .B(net892),
    .Y(_06857_));
 AO21x2_ASAP7_75t_R _29687_ (.A1(net26),
    .A2(_06495_),
    .B(_06496_),
    .Y(_06858_));
 NOR2x2_ASAP7_75t_R _29688_ (.A(_06857_),
    .B(_06858_),
    .Y(_06859_));
 INVx1_ASAP7_75t_R _29689_ (.A(_06859_),
    .Y(_06860_));
 OA21x2_ASAP7_75t_R _29690_ (.A1(_06592_),
    .A2(_06479_),
    .B(_06698_),
    .Y(_06861_));
 AOI221x1_ASAP7_75t_R _29691_ (.A1(_06550_),
    .A2(_06856_),
    .B1(_06860_),
    .B2(_06861_),
    .C(_06679_),
    .Y(_06862_));
 NOR2x1_ASAP7_75t_R _29692_ (.A(_06601_),
    .B(_06479_),
    .Y(_06863_));
 INVx1_ASAP7_75t_R _29693_ (.A(_06863_),
    .Y(_06864_));
 OAI21x1_ASAP7_75t_R _29694_ (.A1(_06507_),
    .A2(_06505_),
    .B(_06864_),
    .Y(_06865_));
 NAND2x2_ASAP7_75t_R _29695_ (.A(_06455_),
    .B(_06516_),
    .Y(_06866_));
 INVx1_ASAP7_75t_R _29696_ (.A(_00407_),
    .Y(_06867_));
 NAND2x1_ASAP7_75t_R _29697_ (.A(_06867_),
    .B(_06753_),
    .Y(_06868_));
 AND3x1_ASAP7_75t_R _29698_ (.A(_06866_),
    .B(_06722_),
    .C(_06868_),
    .Y(_06869_));
 AOI21x1_ASAP7_75t_R _29699_ (.A1(_06715_),
    .A2(_06865_),
    .B(_06869_),
    .Y(_06870_));
 OAI21x1_ASAP7_75t_R _29700_ (.A1(_06641_),
    .A2(_06870_),
    .B(_06535_),
    .Y(_06871_));
 AND2x2_ASAP7_75t_R _29701_ (.A(_06551_),
    .B(_06548_),
    .Y(_06872_));
 AO21x1_ASAP7_75t_R _29702_ (.A1(_06743_),
    .A2(_06872_),
    .B(_06515_),
    .Y(_06873_));
 AOI21x1_ASAP7_75t_R _29703_ (.A1(_06557_),
    .A2(_06653_),
    .B(_06722_),
    .Y(_06874_));
 AOI21x1_ASAP7_75t_R _29704_ (.A1(_06874_),
    .A2(_06734_),
    .B(_06619_),
    .Y(_06875_));
 OAI21x1_ASAP7_75t_R _29705_ (.A1(_06564_),
    .A2(_06873_),
    .B(_06875_),
    .Y(_06876_));
 NOR2x1_ASAP7_75t_R _29706_ (.A(_06559_),
    .B(_06716_),
    .Y(_06877_));
 NAND2x1_ASAP7_75t_R _29707_ (.A(_06596_),
    .B(_06630_),
    .Y(_06878_));
 AOI21x1_ASAP7_75t_R _29708_ (.A1(_06877_),
    .A2(_06878_),
    .B(_06491_),
    .Y(_06879_));
 OAI21x1_ASAP7_75t_R _29709_ (.A1(_06701_),
    .A2(_06609_),
    .B(_06557_),
    .Y(_06880_));
 AOI21x1_ASAP7_75t_R _29710_ (.A1(_06608_),
    .A2(_06666_),
    .B(_06552_),
    .Y(_06881_));
 NAND2x1_ASAP7_75t_R _29711_ (.A(_06880_),
    .B(_06881_),
    .Y(_06882_));
 AOI21x1_ASAP7_75t_R _29712_ (.A1(_06879_),
    .A2(_06882_),
    .B(_06627_),
    .Y(_06883_));
 AOI21x1_ASAP7_75t_R _29713_ (.A1(_06876_),
    .A2(_06883_),
    .B(_06687_),
    .Y(_06884_));
 OAI21x1_ASAP7_75t_R _29714_ (.A1(_06862_),
    .A2(_06871_),
    .B(_06884_),
    .Y(_06885_));
 AOI21x1_ASAP7_75t_R _29715_ (.A1(_06621_),
    .A2(_06749_),
    .B(_06559_),
    .Y(_06886_));
 OA21x2_ASAP7_75t_R _29716_ (.A1(_06507_),
    .A2(_06711_),
    .B(_06886_),
    .Y(_06887_));
 AO21x1_ASAP7_75t_R _29717_ (.A1(_06505_),
    .A2(_06602_),
    .B(_06549_),
    .Y(_06888_));
 AOI21x1_ASAP7_75t_R _29718_ (.A1(_06596_),
    .A2(_06872_),
    .B(_06722_),
    .Y(_06889_));
 AO21x1_ASAP7_75t_R _29719_ (.A1(_06888_),
    .A2(_06889_),
    .B(_06491_),
    .Y(_06890_));
 AOI211x1_ASAP7_75t_R _29720_ (.A1(_06558_),
    .A2(_06593_),
    .B(net846),
    .C(_06552_),
    .Y(_06891_));
 AOI21x1_ASAP7_75t_R _29721_ (.A1(_06866_),
    .A2(_06891_),
    .B(_06619_),
    .Y(_06892_));
 AOI21x1_ASAP7_75t_R _29722_ (.A1(_06615_),
    .A2(_06654_),
    .B(_06584_),
    .Y(_06893_));
 INVx1_ASAP7_75t_R _29723_ (.A(_06480_),
    .Y(_06894_));
 NAND2x1_ASAP7_75t_R _29724_ (.A(_06893_),
    .B(_06894_),
    .Y(_06895_));
 AOI21x1_ASAP7_75t_R _29725_ (.A1(_06892_),
    .A2(_06895_),
    .B(_06677_),
    .Y(_06896_));
 OAI21x1_ASAP7_75t_R _29726_ (.A1(_06887_),
    .A2(_06890_),
    .B(_06896_),
    .Y(_06897_));
 NAND2x1_ASAP7_75t_R _29727_ (.A(_06466_),
    .B(_06479_),
    .Y(_06898_));
 OA21x2_ASAP7_75t_R _29728_ (.A1(_06898_),
    .A2(_06722_),
    .B(_06647_),
    .Y(_06899_));
 OA21x2_ASAP7_75t_R _29729_ (.A1(net26),
    .A2(_06478_),
    .B(_06455_),
    .Y(_06900_));
 NAND2x1_ASAP7_75t_R _29730_ (.A(_06663_),
    .B(_06900_),
    .Y(_06901_));
 AOI21x1_ASAP7_75t_R _29731_ (.A1(_06663_),
    .A2(_06683_),
    .B(_06559_),
    .Y(_06902_));
 NAND2x1_ASAP7_75t_R _29732_ (.A(_06901_),
    .B(_06902_),
    .Y(_06903_));
 AOI21x1_ASAP7_75t_R _29733_ (.A1(_06899_),
    .A2(_06903_),
    .B(_06627_),
    .Y(_06904_));
 NOR3x1_ASAP7_75t_R _29734_ (.A(_06476_),
    .B(_06549_),
    .C(_06547_),
    .Y(_06905_));
 OAI21x1_ASAP7_75t_R _29735_ (.A1(_06859_),
    .A2(_06905_),
    .B(_06698_),
    .Y(_06906_));
 AOI21x1_ASAP7_75t_R _29736_ (.A1(_06812_),
    .A2(_06772_),
    .B(_06525_),
    .Y(_06907_));
 NAND2x1_ASAP7_75t_R _29737_ (.A(_06906_),
    .B(_06907_),
    .Y(_06908_));
 AOI21x1_ASAP7_75t_R _29738_ (.A1(_06904_),
    .A2(_06908_),
    .B(_06582_),
    .Y(_06909_));
 NAND2x1_ASAP7_75t_R _29739_ (.A(_06897_),
    .B(_06909_),
    .Y(_06910_));
 NAND2x1_ASAP7_75t_R _29740_ (.A(_06910_),
    .B(_06885_),
    .Y(_00148_));
 AO21x1_ASAP7_75t_R _29741_ (.A1(_06537_),
    .A2(_06623_),
    .B(_06593_),
    .Y(_06911_));
 AO21x1_ASAP7_75t_R _29742_ (.A1(_06740_),
    .A2(_06571_),
    .B(_06664_),
    .Y(_06912_));
 AND3x1_ASAP7_75t_R _29743_ (.A(_06912_),
    .B(_06911_),
    .C(_06515_),
    .Y(_06913_));
 AO21x1_ASAP7_75t_R _29744_ (.A1(_06476_),
    .A2(_16052_),
    .B(_06510_),
    .Y(_06914_));
 OA21x2_ASAP7_75t_R _29745_ (.A1(_06494_),
    .A2(_06593_),
    .B(_06552_),
    .Y(_06915_));
 AO21x1_ASAP7_75t_R _29746_ (.A1(_06914_),
    .A2(_06915_),
    .B(_06491_),
    .Y(_06916_));
 AO21x1_ASAP7_75t_R _29747_ (.A1(_06540_),
    .A2(_06558_),
    .B(_06471_),
    .Y(_06917_));
 OA21x2_ASAP7_75t_R _29748_ (.A1(_06917_),
    .A2(_06597_),
    .B(_06647_),
    .Y(_06918_));
 NOR2x1_ASAP7_75t_R _29749_ (.A(net23),
    .B(_06671_),
    .Y(_06919_));
 AND3x1_ASAP7_75t_R _29750_ (.A(_06501_),
    .B(_06502_),
    .C(_06503_),
    .Y(_06920_));
 OA21x2_ASAP7_75t_R _29751_ (.A1(_06920_),
    .A2(_06753_),
    .B(_06616_),
    .Y(_06921_));
 OAI21x1_ASAP7_75t_R _29752_ (.A1(_06919_),
    .A2(_06603_),
    .B(_06921_),
    .Y(_06922_));
 AOI21x1_ASAP7_75t_R _29753_ (.A1(_06918_),
    .A2(_06922_),
    .B(_06677_),
    .Y(_06923_));
 OAI21x1_ASAP7_75t_R _29754_ (.A1(_06916_),
    .A2(_06913_),
    .B(_06923_),
    .Y(_06924_));
 OA21x2_ASAP7_75t_R _29755_ (.A1(net23),
    .A2(_06753_),
    .B(_06616_),
    .Y(_06925_));
 AOI21x1_ASAP7_75t_R _29756_ (.A1(_06925_),
    .A2(_06631_),
    .B(_06619_),
    .Y(_06926_));
 AOI21x1_ASAP7_75t_R _29757_ (.A1(_06692_),
    .A2(_06757_),
    .B(_06552_),
    .Y(_06927_));
 AO21x1_ASAP7_75t_R _29758_ (.A1(_06857_),
    .A2(_16060_),
    .B(_06658_),
    .Y(_06928_));
 NAND2x1_ASAP7_75t_R _29759_ (.A(_06927_),
    .B(_06928_),
    .Y(_06929_));
 AOI21x1_ASAP7_75t_R _29760_ (.A1(_06926_),
    .A2(_06929_),
    .B(_06627_),
    .Y(_06930_));
 AO21x1_ASAP7_75t_R _29761_ (.A1(_06538_),
    .A2(_06763_),
    .B(_06664_),
    .Y(_06931_));
 NAND2x1_ASAP7_75t_R _29762_ (.A(_06563_),
    .B(_06931_),
    .Y(_06932_));
 OA21x2_ASAP7_75t_R _29763_ (.A1(_06537_),
    .A2(_06753_),
    .B(_06584_),
    .Y(_06933_));
 OAI21x1_ASAP7_75t_R _29764_ (.A1(_06752_),
    .A2(_06681_),
    .B(_06557_),
    .Y(_06934_));
 AOI21x1_ASAP7_75t_R _29765_ (.A1(_06933_),
    .A2(_06934_),
    .B(_06525_),
    .Y(_06935_));
 OAI21x1_ASAP7_75t_R _29766_ (.A1(_06715_),
    .A2(_06932_),
    .B(_06935_),
    .Y(_06936_));
 AOI21x1_ASAP7_75t_R _29767_ (.A1(_06930_),
    .A2(_06936_),
    .B(_06687_),
    .Y(_06937_));
 NAND2x1_ASAP7_75t_R _29768_ (.A(_06937_),
    .B(_06924_),
    .Y(_06938_));
 NOR2x1_ASAP7_75t_R _29769_ (.A(_06552_),
    .B(_06872_),
    .Y(_06939_));
 NAND2x1_ASAP7_75t_R _29770_ (.A(_06717_),
    .B(_06939_),
    .Y(_06940_));
 NOR2x1_ASAP7_75t_R _29771_ (.A(_06584_),
    .B(_06636_),
    .Y(_06941_));
 AOI21x1_ASAP7_75t_R _29772_ (.A1(_06941_),
    .A2(_06832_),
    .B(_06534_),
    .Y(_06942_));
 AOI21x1_ASAP7_75t_R _29773_ (.A1(_06940_),
    .A2(_06942_),
    .B(_06491_),
    .Y(_06943_));
 AO21x1_ASAP7_75t_R _29774_ (.A1(_06740_),
    .A2(_06753_),
    .B(_06514_),
    .Y(_06944_));
 AOI21x1_ASAP7_75t_R _29775_ (.A1(_06624_),
    .A2(_06659_),
    .B(_06944_),
    .Y(_06945_));
 AO21x1_ASAP7_75t_R _29776_ (.A1(_06692_),
    .A2(_06730_),
    .B(_06664_),
    .Y(_06946_));
 AOI21x1_ASAP7_75t_R _29777_ (.A1(_06866_),
    .A2(_06946_),
    .B(_06512_),
    .Y(_06947_));
 OAI21x1_ASAP7_75t_R _29778_ (.A1(_06945_),
    .A2(_06947_),
    .B(_06627_),
    .Y(_06948_));
 AOI21x1_ASAP7_75t_R _29779_ (.A1(_06943_),
    .A2(_06948_),
    .B(_06582_),
    .Y(_06949_));
 AO21x1_ASAP7_75t_R _29780_ (.A1(_06740_),
    .A2(_06587_),
    .B(_06540_),
    .Y(_06950_));
 NAND2x1_ASAP7_75t_R _29781_ (.A(_06950_),
    .B(_06610_),
    .Y(_06951_));
 NAND2x1_ASAP7_75t_R _29782_ (.A(_06757_),
    .B(_06493_),
    .Y(_06952_));
 INVx1_ASAP7_75t_R _29783_ (.A(_01264_),
    .Y(_06953_));
 AOI21x1_ASAP7_75t_R _29784_ (.A1(_06953_),
    .A2(_06510_),
    .B(_06499_),
    .Y(_06954_));
 AOI21x1_ASAP7_75t_R _29785_ (.A1(_06952_),
    .A2(_06954_),
    .B(_06534_),
    .Y(_06955_));
 NAND2x1_ASAP7_75t_R _29786_ (.A(_06951_),
    .B(_06955_),
    .Y(_06956_));
 NAND2x1_ASAP7_75t_R _29787_ (.A(_06455_),
    .B(_06537_),
    .Y(_06957_));
 NOR2x1_ASAP7_75t_R _29788_ (.A(_06681_),
    .B(_06957_),
    .Y(_06958_));
 AO21x1_ASAP7_75t_R _29789_ (.A1(_06585_),
    .A2(_06561_),
    .B(_06616_),
    .Y(_06959_));
 OA21x2_ASAP7_75t_R _29790_ (.A1(_16050_),
    .A2(_06548_),
    .B(_06471_),
    .Y(_06960_));
 OAI21x1_ASAP7_75t_R _29791_ (.A1(_06857_),
    .A2(_06858_),
    .B(_06960_),
    .Y(_06961_));
 OAI21x1_ASAP7_75t_R _29792_ (.A1(_06958_),
    .A2(_06959_),
    .B(_06961_),
    .Y(_06962_));
 AOI21x1_ASAP7_75t_R _29793_ (.A1(_06627_),
    .A2(_06962_),
    .B(_06641_),
    .Y(_06963_));
 NAND2x1_ASAP7_75t_R _29794_ (.A(_06956_),
    .B(_06963_),
    .Y(_06964_));
 NAND2x1_ASAP7_75t_R _29795_ (.A(_06949_),
    .B(_06964_),
    .Y(_06965_));
 NAND2x1_ASAP7_75t_R _29796_ (.A(_06938_),
    .B(_06965_),
    .Y(_00149_));
 AO21x1_ASAP7_75t_R _29797_ (.A1(_06540_),
    .A2(net596),
    .B(_06471_),
    .Y(_06966_));
 AOI21x1_ASAP7_75t_R _29798_ (.A1(_06778_),
    .A2(_06603_),
    .B(_06966_),
    .Y(_06967_));
 AO21x1_ASAP7_75t_R _29799_ (.A1(_06730_),
    .A2(_06570_),
    .B(_06506_),
    .Y(_06968_));
 OAI21x1_ASAP7_75t_R _29800_ (.A1(_06476_),
    .A2(_06589_),
    .B(_06510_),
    .Y(_06969_));
 AOI21x1_ASAP7_75t_R _29801_ (.A1(_06968_),
    .A2(_06969_),
    .B(_06515_),
    .Y(_06970_));
 OAI21x1_ASAP7_75t_R _29802_ (.A1(_06967_),
    .A2(_06970_),
    .B(_06491_),
    .Y(_06971_));
 OA21x2_ASAP7_75t_R _29803_ (.A1(_06537_),
    .A2(_06506_),
    .B(_06514_),
    .Y(_06972_));
 NAND2x1_ASAP7_75t_R _29804_ (.A(_06710_),
    .B(_06900_),
    .Y(_06973_));
 AOI21x1_ASAP7_75t_R _29805_ (.A1(_06972_),
    .A2(_06973_),
    .B(_06525_),
    .Y(_06974_));
 INVx1_ASAP7_75t_R _29806_ (.A(_06920_),
    .Y(_06975_));
 AOI22x1_ASAP7_75t_R _29807_ (.A1(_06975_),
    .A2(_06695_),
    .B1(_16047_),
    .B2(_06716_),
    .Y(_06976_));
 NAND2x1_ASAP7_75t_R _29808_ (.A(_06856_),
    .B(_06976_),
    .Y(_06977_));
 AOI21x1_ASAP7_75t_R _29809_ (.A1(_06974_),
    .A2(_06977_),
    .B(_06677_),
    .Y(_06978_));
 NAND2x1_ASAP7_75t_R _29810_ (.A(_06971_),
    .B(_06978_),
    .Y(_06979_));
 AND2x2_ASAP7_75t_R _29811_ (.A(_01267_),
    .B(_01269_),
    .Y(_06980_));
 OA21x2_ASAP7_75t_R _29812_ (.A1(_06506_),
    .A2(_06980_),
    .B(_06647_),
    .Y(_06981_));
 NAND2x1_ASAP7_75t_R _29813_ (.A(_06710_),
    .B(_06749_),
    .Y(_06982_));
 AOI21x1_ASAP7_75t_R _29814_ (.A1(_06981_),
    .A2(_06982_),
    .B(_06515_),
    .Y(_06983_));
 NAND2x2_ASAP7_75t_R _29815_ (.A(_06605_),
    .B(_06757_),
    .Y(_06984_));
 NAND2x1_ASAP7_75t_R _29816_ (.A(_06716_),
    .B(_06561_),
    .Y(_06985_));
 AOI21x1_ASAP7_75t_R _29817_ (.A1(_06664_),
    .A2(_06498_),
    .B(_06647_),
    .Y(_06986_));
 NAND3x1_ASAP7_75t_R _29818_ (.A(_06984_),
    .B(_06985_),
    .C(_06986_),
    .Y(_06987_));
 AOI21x1_ASAP7_75t_R _29819_ (.A1(_06983_),
    .A2(_06987_),
    .B(_06534_),
    .Y(_06988_));
 NAND2x1_ASAP7_75t_R _29820_ (.A(_06695_),
    .B(_06538_),
    .Y(_06989_));
 AO21x1_ASAP7_75t_R _29821_ (.A1(_06763_),
    .A2(_06750_),
    .B(_06593_),
    .Y(_06990_));
 AOI21x1_ASAP7_75t_R _29822_ (.A1(_06989_),
    .A2(_06990_),
    .B(_06525_),
    .Y(_06991_));
 NAND2x1_ASAP7_75t_R _29823_ (.A(_06465_),
    .B(_06716_),
    .Y(_06992_));
 NOR3x1_ASAP7_75t_R _29824_ (.A(_06506_),
    .B(_16060_),
    .C(_06546_),
    .Y(_06993_));
 OAI21x1_ASAP7_75t_R _29825_ (.A1(_06842_),
    .A2(_06993_),
    .B(_06647_),
    .Y(_06994_));
 NAND2x1_ASAP7_75t_R _29826_ (.A(_06992_),
    .B(_06994_),
    .Y(_06995_));
 OAI21x1_ASAP7_75t_R _29827_ (.A1(_06991_),
    .A2(_06995_),
    .B(_06715_),
    .Y(_06996_));
 AOI21x1_ASAP7_75t_R _29828_ (.A1(_06988_),
    .A2(_06996_),
    .B(_06582_),
    .Y(_06997_));
 NAND2x1_ASAP7_75t_R _29829_ (.A(_06979_),
    .B(_06997_),
    .Y(_06998_));
 NAND2x1_ASAP7_75t_R _29830_ (.A(_00409_),
    .B(_06510_),
    .Y(_06999_));
 NAND2x1_ASAP7_75t_R _29831_ (.A(_06692_),
    .B(_06757_),
    .Y(_07000_));
 AOI21x1_ASAP7_75t_R _29832_ (.A1(_06999_),
    .A2(_07000_),
    .B(_06698_),
    .Y(_07001_));
 AO21x1_ASAP7_75t_R _29833_ (.A1(_06740_),
    .A2(_06571_),
    .B(_06593_),
    .Y(_07002_));
 AOI21x1_ASAP7_75t_R _29834_ (.A1(_06649_),
    .A2(_07002_),
    .B(_06512_),
    .Y(_07003_));
 OAI21x1_ASAP7_75t_R _29835_ (.A1(_07001_),
    .A2(_07003_),
    .B(_06627_),
    .Y(_07004_));
 NAND2x1_ASAP7_75t_R _29836_ (.A(_07004_),
    .B(_06679_),
    .Y(_07005_));
 NOR2x1_ASAP7_75t_R _29837_ (.A(_06753_),
    .B(_06826_),
    .Y(_07006_));
 AO21x1_ASAP7_75t_R _29838_ (.A1(_06654_),
    .A2(_06632_),
    .B(_06471_),
    .Y(_07007_));
 OA21x2_ASAP7_75t_R _29839_ (.A1(_07006_),
    .A2(_07007_),
    .B(_06676_),
    .Y(_07008_));
 INVx1_ASAP7_75t_R _29840_ (.A(_06738_),
    .Y(_07009_));
 OAI21x1_ASAP7_75t_R _29841_ (.A1(_07009_),
    .A2(_07006_),
    .B(_06656_),
    .Y(_07010_));
 AND2x2_ASAP7_75t_R _29842_ (.A(_07008_),
    .B(_07010_),
    .Y(_07011_));
 NAND2x1_ASAP7_75t_R _29843_ (.A(_06707_),
    .B(_06594_),
    .Y(_07012_));
 OA21x2_ASAP7_75t_R _29844_ (.A1(_06623_),
    .A2(_06664_),
    .B(_06616_),
    .Y(_07013_));
 AOI21x1_ASAP7_75t_R _29845_ (.A1(_07013_),
    .A2(_06832_),
    .B(_06534_),
    .Y(_07014_));
 AOI21x1_ASAP7_75t_R _29846_ (.A1(_07012_),
    .A2(_07014_),
    .B(_06679_),
    .Y(_07015_));
 OA21x2_ASAP7_75t_R _29847_ (.A1(_06863_),
    .A2(_06497_),
    .B(_06515_),
    .Y(_07016_));
 OAI21x1_ASAP7_75t_R _29848_ (.A1(_06745_),
    .A2(_07016_),
    .B(_06627_),
    .Y(_07017_));
 AOI21x1_ASAP7_75t_R _29849_ (.A1(_07015_),
    .A2(_07017_),
    .B(_06687_),
    .Y(_07018_));
 OAI21x1_ASAP7_75t_R _29850_ (.A1(_07005_),
    .A2(_07011_),
    .B(_07018_),
    .Y(_07019_));
 NAND2x1_ASAP7_75t_R _29851_ (.A(_06998_),
    .B(_07019_),
    .Y(_00150_));
 NOR2x1_ASAP7_75t_R _29852_ (.A(_06559_),
    .B(_06851_),
    .Y(_07020_));
 NAND2x1_ASAP7_75t_R _29853_ (.A(_06567_),
    .B(_06681_),
    .Y(_07021_));
 AO21x1_ASAP7_75t_R _29854_ (.A1(_07020_),
    .A2(_07021_),
    .B(_06491_),
    .Y(_07022_));
 AO21x1_ASAP7_75t_R _29855_ (.A1(_06476_),
    .A2(net23),
    .B(_06549_),
    .Y(_07023_));
 OAI21x1_ASAP7_75t_R _29856_ (.A1(net596),
    .A2(_06651_),
    .B(_06541_),
    .Y(_07024_));
 AND3x1_ASAP7_75t_R _29857_ (.A(_07023_),
    .B(_07024_),
    .C(_06698_),
    .Y(_07025_));
 OAI21x1_ASAP7_75t_R _29858_ (.A1(_07022_),
    .A2(_07025_),
    .B(_06535_),
    .Y(_07026_));
 NOR2x1_ASAP7_75t_R _29859_ (.A(_06455_),
    .B(_16052_),
    .Y(_07027_));
 AO21x1_ASAP7_75t_R _29860_ (.A1(_06900_),
    .A2(_06663_),
    .B(_07027_),
    .Y(_07028_));
 AOI21x1_ASAP7_75t_R _29861_ (.A1(_06698_),
    .A2(_07028_),
    .B(_06619_),
    .Y(_07029_));
 OAI21x1_ASAP7_75t_R _29862_ (.A1(_06476_),
    .A2(_06651_),
    .B(_06557_),
    .Y(_07030_));
 NAND2x1_ASAP7_75t_R _29863_ (.A(_07030_),
    .B(_06772_),
    .Y(_07031_));
 AND2x2_ASAP7_75t_R _29864_ (.A(_07029_),
    .B(_07031_),
    .Y(_07032_));
 NAND2x1_ASAP7_75t_R _29865_ (.A(_06984_),
    .B(_06792_),
    .Y(_07033_));
 NAND2x2_ASAP7_75t_R _29866_ (.A(net22),
    .B(_06585_),
    .Y(_07034_));
 AOI21x1_ASAP7_75t_R _29867_ (.A1(_06645_),
    .A2(_06605_),
    .B(_06722_),
    .Y(_07035_));
 AOI21x1_ASAP7_75t_R _29868_ (.A1(_07034_),
    .A2(_07035_),
    .B(_06525_),
    .Y(_07036_));
 OAI21x1_ASAP7_75t_R _29869_ (.A1(_06715_),
    .A2(_07033_),
    .B(_07036_),
    .Y(_07037_));
 NOR2x1_ASAP7_75t_R _29870_ (.A(_06584_),
    .B(_06654_),
    .Y(_07038_));
 AOI21x1_ASAP7_75t_R _29871_ (.A1(_07038_),
    .A2(_06864_),
    .B(_06619_),
    .Y(_07039_));
 NOR2x1_ASAP7_75t_R _29872_ (.A(_06701_),
    .B(_06651_),
    .Y(_07040_));
 OAI21x1_ASAP7_75t_R _29873_ (.A1(_16060_),
    .A2(_16050_),
    .B(net23),
    .Y(_07041_));
 AOI21x1_ASAP7_75t_R _29874_ (.A1(_06557_),
    .A2(_07041_),
    .B(_06722_),
    .Y(_07042_));
 OAI21x1_ASAP7_75t_R _29875_ (.A1(_06541_),
    .A2(_07040_),
    .B(_07042_),
    .Y(_07043_));
 AOI21x1_ASAP7_75t_R _29876_ (.A1(_07039_),
    .A2(_07043_),
    .B(_06627_),
    .Y(_07044_));
 AOI21x1_ASAP7_75t_R _29877_ (.A1(_07037_),
    .A2(_07044_),
    .B(_06687_),
    .Y(_07045_));
 OAI21x1_ASAP7_75t_R _29878_ (.A1(_07026_),
    .A2(_07032_),
    .B(_07045_),
    .Y(_07046_));
 NAND2x1_ASAP7_75t_R _29879_ (.A(_06561_),
    .B(_06543_),
    .Y(_07047_));
 AOI21x1_ASAP7_75t_R _29880_ (.A1(_07047_),
    .A2(_06838_),
    .B(_06512_),
    .Y(_07048_));
 INVx1_ASAP7_75t_R _29881_ (.A(_06537_),
    .Y(_07049_));
 OAI21x1_ASAP7_75t_R _29882_ (.A1(_07049_),
    .A2(_06658_),
    .B(_06722_),
    .Y(_07050_));
 AOI21x1_ASAP7_75t_R _29883_ (.A1(_06541_),
    .A2(_07040_),
    .B(_07050_),
    .Y(_07051_));
 OAI21x1_ASAP7_75t_R _29884_ (.A1(_07048_),
    .A2(_07051_),
    .B(_06679_),
    .Y(_07052_));
 NAND2x1_ASAP7_75t_R _29885_ (.A(_06953_),
    .B(_06549_),
    .Y(_07053_));
 AOI21x1_ASAP7_75t_R _29886_ (.A1(_07053_),
    .A2(_06982_),
    .B(_06512_),
    .Y(_07054_));
 AND2x2_ASAP7_75t_R _29887_ (.A(_06653_),
    .B(_06540_),
    .Y(_07055_));
 NOR2x1_ASAP7_75t_R _29888_ (.A(_06584_),
    .B(_06509_),
    .Y(_07056_));
 OA21x2_ASAP7_75t_R _29889_ (.A1(_07055_),
    .A2(_06900_),
    .B(_07056_),
    .Y(_07057_));
 OAI21x1_ASAP7_75t_R _29890_ (.A1(_07054_),
    .A2(_07057_),
    .B(_06641_),
    .Y(_07058_));
 NAND2x1_ASAP7_75t_R _29891_ (.A(_07052_),
    .B(_07058_),
    .Y(_07059_));
 AND3x1_ASAP7_75t_R _29892_ (.A(_06623_),
    .B(_06567_),
    .C(_06615_),
    .Y(_07060_));
 AO21x1_ASAP7_75t_R _29893_ (.A1(_06585_),
    .A2(_06692_),
    .B(_06512_),
    .Y(_07061_));
 NAND2x1_ASAP7_75t_R _29894_ (.A(_06549_),
    .B(net828),
    .Y(_07062_));
 NOR2x1_ASAP7_75t_R _29895_ (.A(_06506_),
    .B(_06750_),
    .Y(_07063_));
 OAI21x1_ASAP7_75t_R _29896_ (.A1(_01269_),
    .A2(_06753_),
    .B(_06616_),
    .Y(_07064_));
 NOR2x1_ASAP7_75t_R _29897_ (.A(_07063_),
    .B(_07064_),
    .Y(_07065_));
 AOI21x1_ASAP7_75t_R _29898_ (.A1(_07062_),
    .A2(_07065_),
    .B(_06491_),
    .Y(_07066_));
 OAI21x1_ASAP7_75t_R _29899_ (.A1(_07060_),
    .A2(_07061_),
    .B(_07066_),
    .Y(_07067_));
 OA21x2_ASAP7_75t_R _29900_ (.A1(_06867_),
    .A2(_06753_),
    .B(_06616_),
    .Y(_07068_));
 OR3x1_ASAP7_75t_R _29901_ (.A(_06506_),
    .B(_16057_),
    .C(_01263_),
    .Y(_07069_));
 AOI21x1_ASAP7_75t_R _29902_ (.A1(_07068_),
    .A2(_07069_),
    .B(_06619_),
    .Y(_07070_));
 OAI21x1_ASAP7_75t_R _29903_ (.A1(net26),
    .A2(_06592_),
    .B(_06557_),
    .Y(_07071_));
 NAND2x1_ASAP7_75t_R _29904_ (.A(_07071_),
    .B(_06881_),
    .Y(_07072_));
 AOI21x1_ASAP7_75t_R _29905_ (.A1(_07070_),
    .A2(_07072_),
    .B(_06677_),
    .Y(_07073_));
 AOI21x1_ASAP7_75t_R _29906_ (.A1(_07067_),
    .A2(_07073_),
    .B(_06582_),
    .Y(_07074_));
 OAI21x1_ASAP7_75t_R _29907_ (.A1(_06535_),
    .A2(_07059_),
    .B(_07074_),
    .Y(_07075_));
 NAND2x1_ASAP7_75t_R _29908_ (.A(_07046_),
    .B(_07075_),
    .Y(_00151_));
 NOR2x1_ASAP7_75t_R _29909_ (.A(_10763_),
    .B(_00410_),
    .Y(_07076_));
 XOR2x1_ASAP7_75t_R _29910_ (.A(net619),
    .Y(_07077_),
    .B(_12831_));
 XOR2x1_ASAP7_75t_R _29911_ (.A(net939),
    .Y(_07078_),
    .B(_12871_));
 NAND2x1_ASAP7_75t_R _29912_ (.A(_07078_),
    .B(_07077_),
    .Y(_07079_));
 INVx1_ASAP7_75t_R _29913_ (.A(_12831_),
    .Y(_07080_));
 XOR2x1_ASAP7_75t_R _29914_ (.A(net619),
    .Y(_07081_),
    .B(_07080_));
 XOR2x1_ASAP7_75t_R _29915_ (.A(_12873_),
    .Y(_07082_),
    .B(net939));
 NAND2x1_ASAP7_75t_R _29916_ (.A(_07082_),
    .B(_07081_),
    .Y(_07083_));
 AOI21x1_ASAP7_75t_R _29917_ (.A1(_07083_),
    .A2(_07079_),
    .B(_12095_),
    .Y(_07084_));
 OAI21x1_ASAP7_75t_R _29918_ (.A1(_07084_),
    .A2(_07076_),
    .B(_01102_),
    .Y(_07085_));
 AND2x2_ASAP7_75t_R _29919_ (.A(_10640_),
    .B(_00410_),
    .Y(_07086_));
 NAND2x1_ASAP7_75t_R _29920_ (.A(_07081_),
    .B(_07078_),
    .Y(_07087_));
 NAND2x1_ASAP7_75t_R _29921_ (.A(_07082_),
    .B(_07077_),
    .Y(_07088_));
 AOI21x1_ASAP7_75t_R _29922_ (.A1(_07088_),
    .A2(_07087_),
    .B(_12095_),
    .Y(_07089_));
 INVx1_ASAP7_75t_R _29923_ (.A(_01102_),
    .Y(_07090_));
 OAI21x1_ASAP7_75t_R _29924_ (.A1(_07089_),
    .A2(_07086_),
    .B(_07090_),
    .Y(_07091_));
 NAND2x2_ASAP7_75t_R _29925_ (.A(_07091_),
    .B(_07085_),
    .Y(_07092_));
 BUFx12f_ASAP7_75t_R _29926_ (.A(_07092_),
    .Y(_07093_));
 BUFx16f_ASAP7_75t_R _29927_ (.A(_07093_),
    .Y(_16067_));
 NOR2x1_ASAP7_75t_R _29928_ (.A(_10666_),
    .B(_00411_),
    .Y(_07094_));
 NAND2x1_ASAP7_75t_R _29929_ (.A(net663),
    .B(_12855_),
    .Y(_07095_));
 NAND2x1_ASAP7_75t_R _29930_ (.A(_04442_),
    .B(_12859_),
    .Y(_07096_));
 XNOR2x2_ASAP7_75t_R _29931_ (.A(_00756_),
    .B(_12829_),
    .Y(_07097_));
 AO21x1_ASAP7_75t_R _29932_ (.A1(_07095_),
    .A2(_07096_),
    .B(_07097_),
    .Y(_07098_));
 NAND3x1_ASAP7_75t_R _29933_ (.A(_07095_),
    .B(_07096_),
    .C(_07097_),
    .Y(_07099_));
 AOI21x1_ASAP7_75t_R _29934_ (.A1(_07098_),
    .A2(_07099_),
    .B(_11441_),
    .Y(_07100_));
 INVx1_ASAP7_75t_R _29935_ (.A(_01091_),
    .Y(_07101_));
 OAI21x1_ASAP7_75t_R _29936_ (.A1(_07094_),
    .A2(_07100_),
    .B(_07101_),
    .Y(_07102_));
 AND2x2_ASAP7_75t_R _29937_ (.A(_11373_),
    .B(_00411_),
    .Y(_07103_));
 XOR2x1_ASAP7_75t_R _29938_ (.A(net619),
    .Y(_07104_),
    .B(_12859_));
 NAND2x1_ASAP7_75t_R _29939_ (.A(_04442_),
    .B(_07104_),
    .Y(_07105_));
 XOR2x1_ASAP7_75t_R _29940_ (.A(_07097_),
    .Y(_07106_),
    .B(_12859_));
 NAND2x1_ASAP7_75t_R _29941_ (.A(net663),
    .B(_07106_),
    .Y(_07107_));
 AOI21x1_ASAP7_75t_R _29942_ (.A1(_07105_),
    .A2(_07107_),
    .B(_11441_),
    .Y(_07108_));
 OAI21x1_ASAP7_75t_R _29943_ (.A1(_07103_),
    .A2(_07108_),
    .B(_01091_),
    .Y(_07109_));
 NAND2x2_ASAP7_75t_R _29944_ (.A(_07102_),
    .B(_07109_),
    .Y(_07110_));
 INVx6_ASAP7_75t_R _29945_ (.A(net935),
    .Y(_16069_));
 NOR2x2_ASAP7_75t_R _29946_ (.A(net786),
    .B(_00413_),
    .Y(_07111_));
 XOR2x1_ASAP7_75t_R _29947_ (.A(_12870_),
    .Y(_07112_),
    .B(_12879_));
 NAND2x1_ASAP7_75t_R _29948_ (.A(_12837_),
    .B(_07112_),
    .Y(_07113_));
 XNOR2x1_ASAP7_75t_R _29949_ (.B(_00822_),
    .Y(_07114_),
    .A(_12870_));
 NAND2x1_ASAP7_75t_R _29950_ (.A(_12836_),
    .B(_07114_),
    .Y(_07115_));
 AOI21x1_ASAP7_75t_R _29951_ (.A1(_07113_),
    .A2(_07115_),
    .B(_04341_),
    .Y(_07116_));
 XOR2x1_ASAP7_75t_R _29952_ (.A(_12879_),
    .Y(_07117_),
    .B(_12836_));
 NAND2x1_ASAP7_75t_R _29953_ (.A(_12870_),
    .B(_07117_),
    .Y(_07118_));
 XNOR2x1_ASAP7_75t_R _29954_ (.B(_12836_),
    .Y(_07119_),
    .A(_12879_));
 NAND2x1_ASAP7_75t_R _29955_ (.A(_01456_),
    .B(_07119_),
    .Y(_07120_));
 AOI21x1_ASAP7_75t_R _29956_ (.A1(_07118_),
    .A2(_07120_),
    .B(_04329_),
    .Y(_07121_));
 OAI21x1_ASAP7_75t_R _29957_ (.A1(_07116_),
    .A2(_07121_),
    .B(net667),
    .Y(_07122_));
 INVx1_ASAP7_75t_R _29958_ (.A(_07122_),
    .Y(_07123_));
 INVx2_ASAP7_75t_R _29959_ (.A(_01113_),
    .Y(_07124_));
 OAI21x1_ASAP7_75t_R _29960_ (.A1(_07123_),
    .A2(_07111_),
    .B(_07124_),
    .Y(_07125_));
 INVx3_ASAP7_75t_R _29961_ (.A(_07111_),
    .Y(_07126_));
 NAND3x2_ASAP7_75t_R _29962_ (.B(_01113_),
    .C(_07126_),
    .Y(_07127_),
    .A(_07122_));
 NAND2x2_ASAP7_75t_R _29963_ (.A(_07127_),
    .B(_07125_),
    .Y(_07128_));
 BUFx10_ASAP7_75t_R _29964_ (.A(_07128_),
    .Y(_07129_));
 BUFx10_ASAP7_75t_R _29965_ (.A(_07129_),
    .Y(_16077_));
 BUFx12_ASAP7_75t_R _29966_ (.A(_07110_),
    .Y(_16064_));
 NAND3x2_ASAP7_75t_R _29967_ (.B(_07124_),
    .C(_07126_),
    .Y(_07130_),
    .A(_07122_));
 AO21x1_ASAP7_75t_R _29968_ (.A1(_07122_),
    .A2(_07126_),
    .B(_07124_),
    .Y(_07131_));
 BUFx4f_ASAP7_75t_R _29969_ (.A(_07131_),
    .Y(_07132_));
 NAND2x2_ASAP7_75t_R _29970_ (.A(_07130_),
    .B(_07132_),
    .Y(_07133_));
 BUFx10_ASAP7_75t_R _29971_ (.A(_07133_),
    .Y(_16074_));
 BUFx5_ASAP7_75t_R _29972_ (.A(_00415_),
    .Y(_07134_));
 AO21x2_ASAP7_75t_R _29973_ (.A1(_07132_),
    .A2(_07130_),
    .B(_07134_),
    .Y(_07135_));
 INVx1_ASAP7_75t_R _29974_ (.A(_00414_),
    .Y(_07136_));
 AO21x2_ASAP7_75t_R _29975_ (.A1(_07127_),
    .A2(net948),
    .B(_07136_),
    .Y(_07137_));
 XOR2x1_ASAP7_75t_R _29976_ (.A(_12911_),
    .Y(_07138_),
    .B(_12913_));
 OAI21x1_ASAP7_75t_R _29977_ (.A1(_07138_),
    .A2(_04356_),
    .B(_12921_),
    .Y(_07139_));
 XNOR2x1_ASAP7_75t_R _29978_ (.B(_12911_),
    .Y(_07140_),
    .A(_12913_));
 INVx1_ASAP7_75t_R _29979_ (.A(_04356_),
    .Y(_07141_));
 NOR2x1_ASAP7_75t_R _29980_ (.A(_07140_),
    .B(_07141_),
    .Y(_07142_));
 NAND2x1_ASAP7_75t_R _29981_ (.A(_00685_),
    .B(net849),
    .Y(_07143_));
 OAI21x1_ASAP7_75t_R _29982_ (.A1(_07139_),
    .A2(_07142_),
    .B(_07143_),
    .Y(_07144_));
 XNOR2x2_ASAP7_75t_R _29983_ (.A(_01116_),
    .B(_07144_),
    .Y(_07145_));
 BUFx10_ASAP7_75t_R _29984_ (.A(_07145_),
    .Y(_07146_));
 BUFx6f_ASAP7_75t_R _29985_ (.A(_07146_),
    .Y(_07147_));
 AO21x1_ASAP7_75t_R _29986_ (.A1(_07135_),
    .A2(_07137_),
    .B(_07147_),
    .Y(_07148_));
 INVx2_ASAP7_75t_R _29987_ (.A(_00412_),
    .Y(_07149_));
 AO21x2_ASAP7_75t_R _29988_ (.A1(_07127_),
    .A2(net948),
    .B(_07149_),
    .Y(_07150_));
 AOI21x1_ASAP7_75t_R _29989_ (.A1(_07130_),
    .A2(_07132_),
    .B(_07136_),
    .Y(_07151_));
 INVx4_ASAP7_75t_R _29990_ (.A(_07151_),
    .Y(_07152_));
 XOR2x2_ASAP7_75t_R _29991_ (.A(_07144_),
    .B(_01116_),
    .Y(_07153_));
 BUFx12_ASAP7_75t_R _29992_ (.A(_07153_),
    .Y(_07154_));
 BUFx6f_ASAP7_75t_R _29993_ (.A(_07154_),
    .Y(_07155_));
 AO21x1_ASAP7_75t_R _29994_ (.A1(_07150_),
    .A2(_07152_),
    .B(_07155_),
    .Y(_07156_));
 XNOR2x1_ASAP7_75t_R _29995_ (.B(_12928_),
    .Y(_07157_),
    .A(_00824_));
 XOR2x1_ASAP7_75t_R _29996_ (.A(_12953_),
    .Y(_07158_),
    .B(_04369_));
 NOR2x1_ASAP7_75t_R _29997_ (.A(_07157_),
    .B(_07158_),
    .Y(_07159_));
 AO21x1_ASAP7_75t_R _29998_ (.A1(_07158_),
    .A2(_07157_),
    .B(_11370_),
    .Y(_07160_));
 NAND2x2_ASAP7_75t_R _29999_ (.A(_00679_),
    .B(_12092_),
    .Y(_07161_));
 OAI21x1_ASAP7_75t_R _30000_ (.A1(_07159_),
    .A2(_07160_),
    .B(_07161_),
    .Y(_07162_));
 XOR2x2_ASAP7_75t_R _30001_ (.A(_07162_),
    .B(_01117_),
    .Y(_07163_));
 BUFx6f_ASAP7_75t_R _30002_ (.A(_07163_),
    .Y(_07164_));
 AO21x1_ASAP7_75t_R _30003_ (.A1(_07148_),
    .A2(_07156_),
    .B(_07164_),
    .Y(_07165_));
 NAND2x2_ASAP7_75t_R _30004_ (.A(_07128_),
    .B(net938),
    .Y(_07166_));
 BUFx6f_ASAP7_75t_R _30005_ (.A(_07154_),
    .Y(_07167_));
 AO21x1_ASAP7_75t_R _30006_ (.A1(_07166_),
    .A2(_07135_),
    .B(_07167_),
    .Y(_07168_));
 INVx4_ASAP7_75t_R _30007_ (.A(_07134_),
    .Y(_07169_));
 AOI21x1_ASAP7_75t_R _30008_ (.A1(net950),
    .A2(_07127_),
    .B(_07169_),
    .Y(_07170_));
 NAND2x2_ASAP7_75t_R _30009_ (.A(_07154_),
    .B(net561),
    .Y(_07171_));
 XOR2x2_ASAP7_75t_R _30010_ (.A(_07162_),
    .B(_09507_),
    .Y(_07172_));
 BUFx6f_ASAP7_75t_R _30011_ (.A(_07172_),
    .Y(_07173_));
 BUFx6f_ASAP7_75t_R _30012_ (.A(_07173_),
    .Y(_07174_));
 AO21x1_ASAP7_75t_R _30013_ (.A1(_07168_),
    .A2(_07171_),
    .B(_07174_),
    .Y(_07175_));
 XOR2x1_ASAP7_75t_R _30014_ (.A(_12952_),
    .Y(_07176_),
    .B(_12902_));
 XOR2x1_ASAP7_75t_R _30015_ (.A(_07176_),
    .Y(_07177_),
    .B(_00856_));
 XOR2x1_ASAP7_75t_R _30016_ (.A(_07177_),
    .Y(_07178_),
    .B(_12954_));
 NOR2x2_ASAP7_75t_R _30017_ (.A(_11374_),
    .B(_07178_),
    .Y(_07179_));
 NOR2x2_ASAP7_75t_R _30018_ (.A(net585),
    .B(_00672_),
    .Y(_07180_));
 NOR3x2_ASAP7_75t_R _30019_ (.B(_01118_),
    .C(_07180_),
    .Y(_07181_),
    .A(_07179_));
 OA21x2_ASAP7_75t_R _30020_ (.A1(_07179_),
    .A2(_07180_),
    .B(_01118_),
    .Y(_07182_));
 NOR2x2_ASAP7_75t_R _30021_ (.A(_07181_),
    .B(_07182_),
    .Y(_07183_));
 CKINVDCx6p67_ASAP7_75t_R _30022_ (.A(_07183_),
    .Y(_07184_));
 BUFx10_ASAP7_75t_R _30023_ (.A(_07184_),
    .Y(_07185_));
 AOI21x1_ASAP7_75t_R _30024_ (.A1(_07165_),
    .A2(_07175_),
    .B(_07185_),
    .Y(_07186_));
 OAI21x1_ASAP7_75t_R _30025_ (.A1(_07129_),
    .A2(net74),
    .B(_07145_),
    .Y(_07187_));
 BUFx12_ASAP7_75t_R _30026_ (.A(net933),
    .Y(_07188_));
 AND2x4_ASAP7_75t_R _30027_ (.A(_07091_),
    .B(_07085_),
    .Y(_07189_));
 BUFx16f_ASAP7_75t_R _30028_ (.A(_07189_),
    .Y(_16065_));
 NAND2x2_ASAP7_75t_R _30029_ (.A(_07188_),
    .B(net943),
    .Y(_07190_));
 INVx2_ASAP7_75t_R _30030_ (.A(_07190_),
    .Y(_07191_));
 NOR2x2_ASAP7_75t_R _30031_ (.A(_07187_),
    .B(_07191_),
    .Y(_07192_));
 NOR2x2_ASAP7_75t_R _30032_ (.A(_07133_),
    .B(_07188_),
    .Y(_07193_));
 BUFx6f_ASAP7_75t_R _30033_ (.A(_07145_),
    .Y(_07194_));
 AO21x1_ASAP7_75t_R _30034_ (.A1(_16067_),
    .A2(_16064_),
    .B(_07194_),
    .Y(_07195_));
 BUFx10_ASAP7_75t_R _30035_ (.A(_07163_),
    .Y(_07196_));
 OAI21x1_ASAP7_75t_R _30036_ (.A1(_07193_),
    .A2(_07195_),
    .B(_07196_),
    .Y(_07197_));
 OAI21x1_ASAP7_75t_R _30037_ (.A1(_07192_),
    .A2(_07197_),
    .B(_07185_),
    .Y(_07198_));
 NOR2x2_ASAP7_75t_R _30038_ (.A(_16064_),
    .B(_07166_),
    .Y(_07199_));
 INVx1_ASAP7_75t_R _30039_ (.A(_07199_),
    .Y(_07200_));
 NOR2x2_ASAP7_75t_R _30040_ (.A(_07169_),
    .B(_07128_),
    .Y(_07201_));
 NOR2x2_ASAP7_75t_R _30041_ (.A(_07167_),
    .B(_07201_),
    .Y(_07202_));
 INVx1_ASAP7_75t_R _30042_ (.A(_07137_),
    .Y(_07203_));
 NOR2x2_ASAP7_75t_R _30043_ (.A(_07149_),
    .B(_07129_),
    .Y(_07204_));
 BUFx6f_ASAP7_75t_R _30044_ (.A(_07154_),
    .Y(_07205_));
 OA21x2_ASAP7_75t_R _30045_ (.A1(_07203_),
    .A2(_07204_),
    .B(_07205_),
    .Y(_07206_));
 BUFx6f_ASAP7_75t_R _30046_ (.A(_07163_),
    .Y(_07207_));
 BUFx6f_ASAP7_75t_R _30047_ (.A(_07207_),
    .Y(_07208_));
 AOI211x1_ASAP7_75t_R _30048_ (.A1(_07200_),
    .A2(_07202_),
    .B(_07206_),
    .C(_07208_),
    .Y(_07209_));
 XOR2x1_ASAP7_75t_R _30049_ (.A(_12902_),
    .Y(_07210_),
    .B(_00762_));
 XOR2x1_ASAP7_75t_R _30050_ (.A(_07210_),
    .Y(_07211_),
    .B(_12956_));
 XOR2x1_ASAP7_75t_R _30051_ (.A(_07211_),
    .Y(_07212_),
    .B(_12900_));
 NOR2x2_ASAP7_75t_R _30052_ (.A(_11450_),
    .B(_00664_),
    .Y(_07213_));
 AO21x1_ASAP7_75t_R _30053_ (.A1(_07212_),
    .A2(_10829_),
    .B(_07213_),
    .Y(_07214_));
 XOR2x2_ASAP7_75t_R _30054_ (.A(_07214_),
    .B(_01119_),
    .Y(_07215_));
 BUFx10_ASAP7_75t_R _30055_ (.A(_07215_),
    .Y(_07216_));
 OAI21x1_ASAP7_75t_R _30056_ (.A1(_07198_),
    .A2(_07209_),
    .B(_07216_),
    .Y(_07217_));
 NOR2x1_ASAP7_75t_R _30057_ (.A(_07186_),
    .B(_07217_),
    .Y(_07218_));
 BUFx6f_ASAP7_75t_R _30058_ (.A(_07172_),
    .Y(_07219_));
 BUFx6f_ASAP7_75t_R _30059_ (.A(_07219_),
    .Y(_07220_));
 BUFx6f_ASAP7_75t_R _30060_ (.A(_07194_),
    .Y(_07221_));
 AO21x2_ASAP7_75t_R _30061_ (.A1(_07132_),
    .A2(_07130_),
    .B(net940),
    .Y(_07222_));
 OAI21x1_ASAP7_75t_R _30062_ (.A1(_16067_),
    .A2(_16074_),
    .B(_07222_),
    .Y(_07223_));
 NAND2x2_ASAP7_75t_R _30063_ (.A(_07133_),
    .B(_07093_),
    .Y(_07224_));
 BUFx12_ASAP7_75t_R _30064_ (.A(_07128_),
    .Y(_07225_));
 BUFx6f_ASAP7_75t_R _30065_ (.A(_07145_),
    .Y(_07226_));
 AOI21x1_ASAP7_75t_R _30066_ (.A1(_07225_),
    .A2(_07188_),
    .B(_07226_),
    .Y(_07227_));
 OA21x2_ASAP7_75t_R _30067_ (.A1(_16064_),
    .A2(_07224_),
    .B(_07227_),
    .Y(_07228_));
 AOI21x1_ASAP7_75t_R _30068_ (.A1(_07221_),
    .A2(_07223_),
    .B(_07228_),
    .Y(_07229_));
 INVx2_ASAP7_75t_R _30069_ (.A(_01274_),
    .Y(_07230_));
 AO21x1_ASAP7_75t_R _30070_ (.A1(_07132_),
    .A2(_07130_),
    .B(_07230_),
    .Y(_07231_));
 BUFx4f_ASAP7_75t_R _30071_ (.A(_07231_),
    .Y(_07232_));
 BUFx6f_ASAP7_75t_R _30072_ (.A(_07172_),
    .Y(_07233_));
 AO21x1_ASAP7_75t_R _30073_ (.A1(_07227_),
    .A2(_07232_),
    .B(_07233_),
    .Y(_07234_));
 NAND2x2_ASAP7_75t_R _30074_ (.A(_07129_),
    .B(_07188_),
    .Y(_07235_));
 NOR2x2_ASAP7_75t_R _30075_ (.A(net943),
    .B(_07235_),
    .Y(_07236_));
 BUFx10_ASAP7_75t_R _30076_ (.A(_07133_),
    .Y(_07237_));
 BUFx6f_ASAP7_75t_R _30077_ (.A(_07153_),
    .Y(_07238_));
 AO21x2_ASAP7_75t_R _30078_ (.A1(net943),
    .A2(_07237_),
    .B(_07238_),
    .Y(_07239_));
 NOR2x1_ASAP7_75t_R _30079_ (.A(_07236_),
    .B(_07239_),
    .Y(_07240_));
 BUFx10_ASAP7_75t_R _30080_ (.A(_07183_),
    .Y(_07241_));
 OAI21x1_ASAP7_75t_R _30081_ (.A1(_07234_),
    .A2(_07240_),
    .B(_07241_),
    .Y(_07242_));
 AOI21x1_ASAP7_75t_R _30082_ (.A1(_07220_),
    .A2(_07229_),
    .B(_07242_),
    .Y(_07243_));
 NOR2x2_ASAP7_75t_R _30083_ (.A(_07230_),
    .B(_07133_),
    .Y(_07244_));
 AO21x1_ASAP7_75t_R _30084_ (.A1(_07132_),
    .A2(_07130_),
    .B(_07169_),
    .Y(_07245_));
 BUFx6f_ASAP7_75t_R _30085_ (.A(_07245_),
    .Y(_07246_));
 NAND2x2_ASAP7_75t_R _30086_ (.A(_07246_),
    .B(_07154_),
    .Y(_07247_));
 OAI21x1_ASAP7_75t_R _30087_ (.A1(_07244_),
    .A2(_07247_),
    .B(_07164_),
    .Y(_07248_));
 NOR2x2_ASAP7_75t_R _30088_ (.A(_07128_),
    .B(net933),
    .Y(_07249_));
 AOI21x1_ASAP7_75t_R _30089_ (.A1(net74),
    .A2(_07093_),
    .B(_07133_),
    .Y(_07250_));
 BUFx6f_ASAP7_75t_R _30090_ (.A(_07226_),
    .Y(_07251_));
 OAI21x1_ASAP7_75t_R _30091_ (.A1(_07249_),
    .A2(_07250_),
    .B(_07251_),
    .Y(_07252_));
 INVx1_ASAP7_75t_R _30092_ (.A(_07252_),
    .Y(_07253_));
 OAI21x1_ASAP7_75t_R _30093_ (.A1(_07248_),
    .A2(_07253_),
    .B(_07185_),
    .Y(_07254_));
 BUFx6f_ASAP7_75t_R _30094_ (.A(_01272_),
    .Y(_07255_));
 INVx1_ASAP7_75t_R _30095_ (.A(_07255_),
    .Y(_07256_));
 OAI21x1_ASAP7_75t_R _30096_ (.A1(_07256_),
    .A2(_07129_),
    .B(_07153_),
    .Y(_07257_));
 AOI21x1_ASAP7_75t_R _30097_ (.A1(_07128_),
    .A2(net74),
    .B(_07153_),
    .Y(_07258_));
 INVx2_ASAP7_75t_R _30098_ (.A(_07258_),
    .Y(_07259_));
 BUFx6f_ASAP7_75t_R _30099_ (.A(_07173_),
    .Y(_07260_));
 OA211x2_ASAP7_75t_R _30100_ (.A1(_07236_),
    .A2(_07257_),
    .B(_07259_),
    .C(_07260_),
    .Y(_07261_));
 INVx3_ASAP7_75t_R _30101_ (.A(_07215_),
    .Y(_07262_));
 BUFx10_ASAP7_75t_R _30102_ (.A(_07262_),
    .Y(_07263_));
 OAI21x1_ASAP7_75t_R _30103_ (.A1(_07254_),
    .A2(_07261_),
    .B(_07263_),
    .Y(_07264_));
 XOR2x1_ASAP7_75t_R _30104_ (.A(_13012_),
    .Y(_07265_),
    .B(_00858_));
 XNOR2x1_ASAP7_75t_R _30105_ (.B(net647),
    .Y(_07266_),
    .A(_00762_));
 XOR2x1_ASAP7_75t_R _30106_ (.A(_07265_),
    .Y(_07267_),
    .B(_07266_));
 NOR2x1_ASAP7_75t_R _30107_ (.A(_10830_),
    .B(_00656_),
    .Y(_07268_));
 AO21x1_ASAP7_75t_R _30108_ (.A1(_07267_),
    .A2(_10830_),
    .B(_07268_),
    .Y(_07269_));
 XOR2x2_ASAP7_75t_R _30109_ (.A(_07269_),
    .B(_01120_),
    .Y(_07270_));
 BUFx10_ASAP7_75t_R _30110_ (.A(_07270_),
    .Y(_07271_));
 OAI21x1_ASAP7_75t_R _30111_ (.A1(_07243_),
    .A2(_07264_),
    .B(_07271_),
    .Y(_07272_));
 AOI21x1_ASAP7_75t_R _30112_ (.A1(_07130_),
    .A2(_07132_),
    .B(_01273_),
    .Y(_07273_));
 AOI21x1_ASAP7_75t_R _30113_ (.A1(_07147_),
    .A2(_07273_),
    .B(_07219_),
    .Y(_07274_));
 NAND2x1_ASAP7_75t_R _30114_ (.A(_07247_),
    .B(_07274_),
    .Y(_07275_));
 NAND2x2_ASAP7_75t_R _30115_ (.A(net947),
    .B(_07249_),
    .Y(_07276_));
 BUFx6f_ASAP7_75t_R _30116_ (.A(_07163_),
    .Y(_07277_));
 AO21x1_ASAP7_75t_R _30117_ (.A1(_07276_),
    .A2(_07227_),
    .B(_07277_),
    .Y(_07278_));
 AOI21x1_ASAP7_75t_R _30118_ (.A1(net948),
    .A2(_07127_),
    .B(_07255_),
    .Y(_07279_));
 AO21x1_ASAP7_75t_R _30119_ (.A1(_07251_),
    .A2(_07279_),
    .B(_07184_),
    .Y(_07280_));
 AOI21x1_ASAP7_75t_R _30120_ (.A1(_07275_),
    .A2(_07278_),
    .B(_07280_),
    .Y(_07281_));
 BUFx6f_ASAP7_75t_R _30121_ (.A(_07153_),
    .Y(_07282_));
 AO21x1_ASAP7_75t_R _30122_ (.A1(_07222_),
    .A2(_07137_),
    .B(_07282_),
    .Y(_07283_));
 AND2x2_ASAP7_75t_R _30123_ (.A(_07257_),
    .B(_07163_),
    .Y(_07284_));
 NAND2x1_ASAP7_75t_R _30124_ (.A(_07283_),
    .B(_07284_),
    .Y(_07285_));
 NOR2x2_ASAP7_75t_R _30125_ (.A(_07134_),
    .B(_07237_),
    .Y(_07286_));
 AOI21x1_ASAP7_75t_R _30126_ (.A1(_07237_),
    .A2(_07093_),
    .B(_07154_),
    .Y(_07287_));
 INVx1_ASAP7_75t_R _30127_ (.A(_07287_),
    .Y(_07288_));
 AO21x1_ASAP7_75t_R _30128_ (.A1(_07127_),
    .A2(net949),
    .B(_00412_),
    .Y(_07289_));
 AOI21x1_ASAP7_75t_R _30129_ (.A1(_16074_),
    .A2(_16064_),
    .B(_07194_),
    .Y(_07290_));
 AOI21x1_ASAP7_75t_R _30130_ (.A1(_07289_),
    .A2(_07290_),
    .B(_07277_),
    .Y(_07291_));
 OAI21x1_ASAP7_75t_R _30131_ (.A1(_07286_),
    .A2(_07288_),
    .B(_07291_),
    .Y(_07292_));
 BUFx10_ASAP7_75t_R _30132_ (.A(_07183_),
    .Y(_07293_));
 AOI21x1_ASAP7_75t_R _30133_ (.A1(_07285_),
    .A2(_07292_),
    .B(_07293_),
    .Y(_07294_));
 OAI21x1_ASAP7_75t_R _30134_ (.A1(_07281_),
    .A2(_07294_),
    .B(_07263_),
    .Y(_07295_));
 NAND2x2_ASAP7_75t_R _30135_ (.A(net934),
    .B(net937),
    .Y(_07296_));
 INVx1_ASAP7_75t_R _30136_ (.A(_01273_),
    .Y(_07297_));
 AOI21x1_ASAP7_75t_R _30137_ (.A1(net950),
    .A2(_07127_),
    .B(_07297_),
    .Y(_07298_));
 NOR2x2_ASAP7_75t_R _30138_ (.A(_07146_),
    .B(_07298_),
    .Y(_07299_));
 OAI21x1_ASAP7_75t_R _30139_ (.A1(_16077_),
    .A2(_07296_),
    .B(_07299_),
    .Y(_07300_));
 OA21x2_ASAP7_75t_R _30140_ (.A1(_07222_),
    .A2(_07282_),
    .B(_07173_),
    .Y(_07301_));
 BUFx6f_ASAP7_75t_R _30141_ (.A(_07183_),
    .Y(_07302_));
 AOI21x1_ASAP7_75t_R _30142_ (.A1(_07300_),
    .A2(_07301_),
    .B(_07302_),
    .Y(_07303_));
 OA21x2_ASAP7_75t_R _30143_ (.A1(_07237_),
    .A2(_00412_),
    .B(_07145_),
    .Y(_07304_));
 INVx1_ASAP7_75t_R _30144_ (.A(_07304_),
    .Y(_07305_));
 NOR2x2_ASAP7_75t_R _30145_ (.A(_07225_),
    .B(_07296_),
    .Y(_07306_));
 NOR2x2_ASAP7_75t_R _30146_ (.A(_07146_),
    .B(_07222_),
    .Y(_07307_));
 NOR2x2_ASAP7_75t_R _30147_ (.A(_07173_),
    .B(_07307_),
    .Y(_07308_));
 OAI21x1_ASAP7_75t_R _30148_ (.A1(_07305_),
    .A2(_07306_),
    .B(_07308_),
    .Y(_07309_));
 BUFx10_ASAP7_75t_R _30149_ (.A(_07262_),
    .Y(_07310_));
 AOI21x1_ASAP7_75t_R _30150_ (.A1(_07303_),
    .A2(_07309_),
    .B(_07310_),
    .Y(_07311_));
 NOR2x2_ASAP7_75t_R _30151_ (.A(net941),
    .B(_07237_),
    .Y(_07312_));
 NAND2x1_ASAP7_75t_R _30152_ (.A(_07194_),
    .B(_07312_),
    .Y(_07313_));
 AOI21x1_ASAP7_75t_R _30153_ (.A1(_07188_),
    .A2(_07093_),
    .B(_07129_),
    .Y(_07314_));
 OAI21x1_ASAP7_75t_R _30154_ (.A1(_07279_),
    .A2(_07314_),
    .B(_07194_),
    .Y(_07315_));
 NAND2x1_ASAP7_75t_R _30155_ (.A(_07313_),
    .B(_07315_),
    .Y(_07316_));
 NOR2x1_ASAP7_75t_R _30156_ (.A(_07188_),
    .B(_07226_),
    .Y(_07317_));
 OAI21x1_ASAP7_75t_R _30157_ (.A1(_07226_),
    .A2(_07152_),
    .B(_07173_),
    .Y(_07318_));
 AOI21x1_ASAP7_75t_R _30158_ (.A1(_16077_),
    .A2(_07317_),
    .B(_07318_),
    .Y(_07319_));
 INVx1_ASAP7_75t_R _30159_ (.A(_07319_),
    .Y(_07320_));
 INVx1_ASAP7_75t_R _30160_ (.A(_01276_),
    .Y(_07321_));
 AO21x2_ASAP7_75t_R _30161_ (.A1(_07127_),
    .A2(net950),
    .B(_07134_),
    .Y(_07322_));
 NAND2x2_ASAP7_75t_R _30162_ (.A(_07146_),
    .B(_07322_),
    .Y(_07323_));
 OAI21x1_ASAP7_75t_R _30163_ (.A1(_07321_),
    .A2(_07251_),
    .B(_07323_),
    .Y(_07324_));
 BUFx10_ASAP7_75t_R _30164_ (.A(_07184_),
    .Y(_07325_));
 AOI21x1_ASAP7_75t_R _30165_ (.A1(_07164_),
    .A2(_07324_),
    .B(_07325_),
    .Y(_07326_));
 OAI21x1_ASAP7_75t_R _30166_ (.A1(_07316_),
    .A2(_07320_),
    .B(_07326_),
    .Y(_07327_));
 AOI21x1_ASAP7_75t_R _30167_ (.A1(_07311_),
    .A2(_07327_),
    .B(_07271_),
    .Y(_07328_));
 NAND2x1_ASAP7_75t_R _30168_ (.A(_07328_),
    .B(_07295_),
    .Y(_07329_));
 OAI21x1_ASAP7_75t_R _30169_ (.A1(_07218_),
    .A2(_07272_),
    .B(_07329_),
    .Y(_00152_));
 OAI21x1_ASAP7_75t_R _30170_ (.A1(_16064_),
    .A2(_07166_),
    .B(_07167_),
    .Y(_07330_));
 NOR2x2_ASAP7_75t_R _30171_ (.A(_07134_),
    .B(_07225_),
    .Y(_07331_));
 AO21x2_ASAP7_75t_R _30172_ (.A1(_07132_),
    .A2(_07130_),
    .B(_07255_),
    .Y(_07332_));
 OA21x2_ASAP7_75t_R _30173_ (.A1(_07332_),
    .A2(_07155_),
    .B(_07219_),
    .Y(_07333_));
 OA21x2_ASAP7_75t_R _30174_ (.A1(_07330_),
    .A2(_07331_),
    .B(_07333_),
    .Y(_07334_));
 NAND2x2_ASAP7_75t_R _30175_ (.A(_07237_),
    .B(_16065_),
    .Y(_07335_));
 NOR2x2_ASAP7_75t_R _30176_ (.A(_07146_),
    .B(_07244_),
    .Y(_07336_));
 AOI21x1_ASAP7_75t_R _30177_ (.A1(_07335_),
    .A2(_07336_),
    .B(_07219_),
    .Y(_07337_));
 BUFx6f_ASAP7_75t_R _30178_ (.A(_07146_),
    .Y(_07338_));
 AOI21x1_ASAP7_75t_R _30179_ (.A1(net947),
    .A2(_16069_),
    .B(_07225_),
    .Y(_07339_));
 NAND2x1_ASAP7_75t_R _30180_ (.A(_07338_),
    .B(_07339_),
    .Y(_07340_));
 AO21x1_ASAP7_75t_R _30181_ (.A1(_07337_),
    .A2(_07340_),
    .B(_07302_),
    .Y(_07341_));
 OAI21x1_ASAP7_75t_R _30182_ (.A1(_07334_),
    .A2(_07341_),
    .B(_07310_),
    .Y(_07342_));
 OAI21x1_ASAP7_75t_R _30183_ (.A1(net946),
    .A2(_16074_),
    .B(_07238_),
    .Y(_07343_));
 OAI21x1_ASAP7_75t_R _30184_ (.A1(_07237_),
    .A2(_07188_),
    .B(_07226_),
    .Y(_07344_));
 OA22x2_ASAP7_75t_R _30185_ (.A1(_07201_),
    .A2(_07343_),
    .B1(_07344_),
    .B2(_07151_),
    .Y(_07345_));
 NAND2x2_ASAP7_75t_R _30186_ (.A(net947),
    .B(_16069_),
    .Y(_07346_));
 NAND2x2_ASAP7_75t_R _30187_ (.A(_07133_),
    .B(net74),
    .Y(_07347_));
 AO21x1_ASAP7_75t_R _30188_ (.A1(_07346_),
    .A2(_07347_),
    .B(_07147_),
    .Y(_07348_));
 INVx2_ASAP7_75t_R _30189_ (.A(_07347_),
    .Y(_07349_));
 OA21x2_ASAP7_75t_R _30190_ (.A1(_07323_),
    .A2(_07349_),
    .B(_07219_),
    .Y(_07350_));
 AOI21x1_ASAP7_75t_R _30191_ (.A1(_07348_),
    .A2(_07350_),
    .B(_07325_),
    .Y(_07351_));
 OA21x2_ASAP7_75t_R _30192_ (.A1(_07220_),
    .A2(_07345_),
    .B(_07351_),
    .Y(_07352_));
 NOR2x2_ASAP7_75t_R _30193_ (.A(_07170_),
    .B(_07145_),
    .Y(_07353_));
 AOI21x1_ASAP7_75t_R _30194_ (.A1(_07232_),
    .A2(_07353_),
    .B(_07207_),
    .Y(_07354_));
 NAND2x1_ASAP7_75t_R _30195_ (.A(_07354_),
    .B(_07315_),
    .Y(_07355_));
 AOI21x1_ASAP7_75t_R _30196_ (.A1(_07155_),
    .A2(_07166_),
    .B(_07219_),
    .Y(_07356_));
 NOR2x2_ASAP7_75t_R _30197_ (.A(net946),
    .B(_07154_),
    .Y(_07357_));
 NOR2x2_ASAP7_75t_R _30198_ (.A(_07225_),
    .B(net947),
    .Y(_07358_));
 AOI21x1_ASAP7_75t_R _30199_ (.A1(_16077_),
    .A2(_07357_),
    .B(_07358_),
    .Y(_07359_));
 BUFx6f_ASAP7_75t_R _30200_ (.A(_07184_),
    .Y(_07360_));
 AOI21x1_ASAP7_75t_R _30201_ (.A1(_07356_),
    .A2(_07359_),
    .B(_07360_),
    .Y(_07361_));
 AOI21x1_ASAP7_75t_R _30202_ (.A1(_07355_),
    .A2(_07361_),
    .B(_07310_),
    .Y(_07362_));
 NOR2x2_ASAP7_75t_R _30203_ (.A(_07237_),
    .B(_07145_),
    .Y(_07363_));
 NAND2x1_ASAP7_75t_R _30204_ (.A(_07363_),
    .B(_07296_),
    .Y(_07364_));
 NAND2x2_ASAP7_75t_R _30205_ (.A(_07190_),
    .B(_07287_),
    .Y(_07365_));
 NAND2x1_ASAP7_75t_R _30206_ (.A(_07364_),
    .B(_07365_),
    .Y(_07366_));
 AOI21x1_ASAP7_75t_R _30207_ (.A1(_07246_),
    .A2(_07227_),
    .B(_07233_),
    .Y(_07367_));
 AO21x1_ASAP7_75t_R _30208_ (.A1(_07235_),
    .A2(_07332_),
    .B(_07155_),
    .Y(_07368_));
 AOI21x1_ASAP7_75t_R _30209_ (.A1(_07367_),
    .A2(_07368_),
    .B(_07302_),
    .Y(_07369_));
 OAI21x1_ASAP7_75t_R _30210_ (.A1(_07208_),
    .A2(_07366_),
    .B(_07369_),
    .Y(_07370_));
 AOI21x1_ASAP7_75t_R _30211_ (.A1(_07362_),
    .A2(_07370_),
    .B(_07271_),
    .Y(_07371_));
 OAI21x1_ASAP7_75t_R _30212_ (.A1(_07342_),
    .A2(_07352_),
    .B(_07371_),
    .Y(_07372_));
 AO21x1_ASAP7_75t_R _30213_ (.A1(_07136_),
    .A2(_07129_),
    .B(_07154_),
    .Y(_07373_));
 OA21x2_ASAP7_75t_R _30214_ (.A1(_07373_),
    .A2(_07349_),
    .B(_07184_),
    .Y(_07374_));
 INVx1_ASAP7_75t_R _30215_ (.A(_07250_),
    .Y(_07375_));
 OAI21x1_ASAP7_75t_R _30216_ (.A1(_07188_),
    .A2(net943),
    .B(_07237_),
    .Y(_07376_));
 AO21x1_ASAP7_75t_R _30217_ (.A1(_07375_),
    .A2(_07376_),
    .B(_07194_),
    .Y(_07377_));
 AND2x2_ASAP7_75t_R _30218_ (.A(_07374_),
    .B(_07377_),
    .Y(_07378_));
 NOR2x2_ASAP7_75t_R _30219_ (.A(_07133_),
    .B(net938),
    .Y(_07379_));
 NOR2x2_ASAP7_75t_R _30220_ (.A(_07379_),
    .B(_07257_),
    .Y(_07380_));
 INVx2_ASAP7_75t_R _30221_ (.A(_07166_),
    .Y(_07381_));
 NOR2x2_ASAP7_75t_R _30222_ (.A(_07187_),
    .B(_07381_),
    .Y(_07382_));
 NOR2x1_ASAP7_75t_R _30223_ (.A(_07380_),
    .B(_07382_),
    .Y(_07383_));
 AO21x1_ASAP7_75t_R _30224_ (.A1(_07383_),
    .A2(_07302_),
    .B(_07174_),
    .Y(_07384_));
 NAND2x1_ASAP7_75t_R _30225_ (.A(_00417_),
    .B(_07155_),
    .Y(_07385_));
 NAND2x2_ASAP7_75t_R _30226_ (.A(_07304_),
    .B(_07276_),
    .Y(_07386_));
 OAI21x1_ASAP7_75t_R _30227_ (.A1(_07360_),
    .A2(_07385_),
    .B(_07386_),
    .Y(_07387_));
 AOI21x1_ASAP7_75t_R _30228_ (.A1(_07220_),
    .A2(_07387_),
    .B(_07310_),
    .Y(_07388_));
 OAI21x1_ASAP7_75t_R _30229_ (.A1(_07378_),
    .A2(_07384_),
    .B(_07388_),
    .Y(_07389_));
 INVx2_ASAP7_75t_R _30230_ (.A(_07222_),
    .Y(_07390_));
 OAI21x1_ASAP7_75t_R _30231_ (.A1(_07193_),
    .A2(_07390_),
    .B(_07338_),
    .Y(_07391_));
 AO21x1_ASAP7_75t_R _30232_ (.A1(_07322_),
    .A2(_07152_),
    .B(_07194_),
    .Y(_07392_));
 AOI21x1_ASAP7_75t_R _30233_ (.A1(_07391_),
    .A2(_07392_),
    .B(_07260_),
    .Y(_07393_));
 INVx1_ASAP7_75t_R _30234_ (.A(_07380_),
    .Y(_07394_));
 AO21x1_ASAP7_75t_R _30235_ (.A1(_07347_),
    .A2(_07137_),
    .B(_07282_),
    .Y(_07395_));
 AOI21x1_ASAP7_75t_R _30236_ (.A1(_07394_),
    .A2(_07395_),
    .B(_07196_),
    .Y(_07396_));
 OAI21x1_ASAP7_75t_R _30237_ (.A1(_07393_),
    .A2(_07396_),
    .B(_07325_),
    .Y(_07397_));
 NAND2x2_ASAP7_75t_R _30238_ (.A(net940),
    .B(_07225_),
    .Y(_07398_));
 OA21x2_ASAP7_75t_R _30239_ (.A1(_07129_),
    .A2(_07230_),
    .B(_07146_),
    .Y(_07399_));
 AOI21x1_ASAP7_75t_R _30240_ (.A1(_07398_),
    .A2(_07399_),
    .B(_07219_),
    .Y(_07400_));
 OAI21x1_ASAP7_75t_R _30241_ (.A1(_07331_),
    .A2(_07330_),
    .B(_07400_),
    .Y(_07401_));
 NOR2x2_ASAP7_75t_R _30242_ (.A(_07146_),
    .B(_07201_),
    .Y(_07402_));
 NOR2x1_ASAP7_75t_R _30243_ (.A(_07207_),
    .B(_07402_),
    .Y(_07403_));
 NAND2x1_ASAP7_75t_R _30244_ (.A(_07258_),
    .B(_07276_),
    .Y(_07404_));
 AOI21x1_ASAP7_75t_R _30245_ (.A1(_07403_),
    .A2(_07404_),
    .B(_07360_),
    .Y(_07405_));
 AOI21x1_ASAP7_75t_R _30246_ (.A1(_07401_),
    .A2(_07405_),
    .B(_07215_),
    .Y(_07406_));
 INVx5_ASAP7_75t_R _30247_ (.A(_07270_),
    .Y(_07407_));
 AOI21x1_ASAP7_75t_R _30248_ (.A1(_07397_),
    .A2(_07406_),
    .B(_07407_),
    .Y(_07408_));
 NAND2x1_ASAP7_75t_R _30249_ (.A(_07389_),
    .B(_07408_),
    .Y(_07409_));
 NAND2x1_ASAP7_75t_R _30250_ (.A(_07372_),
    .B(_07409_),
    .Y(_00153_));
 OAI21x1_ASAP7_75t_R _30251_ (.A1(_07343_),
    .A2(_07314_),
    .B(_07233_),
    .Y(_07410_));
 AO21x1_ASAP7_75t_R _30252_ (.A1(_07322_),
    .A2(_07287_),
    .B(_07410_),
    .Y(_07411_));
 OAI21x1_ASAP7_75t_R _30253_ (.A1(_16074_),
    .A2(_07188_),
    .B(_16067_),
    .Y(_07412_));
 NAND2x1_ASAP7_75t_R _30254_ (.A(_07155_),
    .B(_07412_),
    .Y(_07413_));
 AOI21x1_ASAP7_75t_R _30255_ (.A1(net950),
    .A2(_07127_),
    .B(_01274_),
    .Y(_07414_));
 NOR2x1_ASAP7_75t_R _30256_ (.A(net946),
    .B(_07225_),
    .Y(_07415_));
 OAI21x1_ASAP7_75t_R _30257_ (.A1(net932),
    .A2(_07415_),
    .B(_07147_),
    .Y(_07416_));
 AO21x1_ASAP7_75t_R _30258_ (.A1(_07416_),
    .A2(_07413_),
    .B(_07174_),
    .Y(_07417_));
 NAND3x1_ASAP7_75t_R _30259_ (.A(_07411_),
    .B(_07241_),
    .C(_07417_),
    .Y(_07418_));
 OAI21x1_ASAP7_75t_R _30260_ (.A1(net943),
    .A2(_07235_),
    .B(_07338_),
    .Y(_07419_));
 NAND2x1_ASAP7_75t_R _30261_ (.A(_07174_),
    .B(_07419_),
    .Y(_07420_));
 AO21x1_ASAP7_75t_R _30262_ (.A1(_07132_),
    .A2(_07130_),
    .B(_01274_),
    .Y(_07421_));
 AO21x2_ASAP7_75t_R _30263_ (.A1(_16069_),
    .A2(_16067_),
    .B(_16074_),
    .Y(_07422_));
 AOI21x1_ASAP7_75t_R _30264_ (.A1(_07421_),
    .A2(_07422_),
    .B(_07221_),
    .Y(_07423_));
 OAI21x1_ASAP7_75t_R _30265_ (.A1(_07134_),
    .A2(_07129_),
    .B(_07145_),
    .Y(_07424_));
 NOR2x1_ASAP7_75t_R _30266_ (.A(_07379_),
    .B(_07424_),
    .Y(_07425_));
 OAI21x1_ASAP7_75t_R _30267_ (.A1(_16077_),
    .A2(_16064_),
    .B(_07282_),
    .Y(_07426_));
 NOR2x1_ASAP7_75t_R _30268_ (.A(_07312_),
    .B(_07426_),
    .Y(_07427_));
 OAI21x1_ASAP7_75t_R _30269_ (.A1(_07425_),
    .A2(_07427_),
    .B(_07164_),
    .Y(_07428_));
 OAI21x1_ASAP7_75t_R _30270_ (.A1(_07420_),
    .A2(_07423_),
    .B(_07428_),
    .Y(_07429_));
 AOI21x1_ASAP7_75t_R _30271_ (.A1(_07185_),
    .A2(_07429_),
    .B(_07263_),
    .Y(_07430_));
 OAI21x1_ASAP7_75t_R _30272_ (.A1(_07279_),
    .A2(_07273_),
    .B(_07147_),
    .Y(_07431_));
 AOI21x1_ASAP7_75t_R _30273_ (.A1(net946),
    .A2(_07225_),
    .B(_07226_),
    .Y(_07432_));
 AOI21x1_ASAP7_75t_R _30274_ (.A1(_07432_),
    .A2(_07335_),
    .B(_07207_),
    .Y(_07433_));
 NAND2x1_ASAP7_75t_R _30275_ (.A(_07431_),
    .B(_07433_),
    .Y(_07434_));
 OAI21x1_ASAP7_75t_R _30276_ (.A1(net936),
    .A2(_16074_),
    .B(_07194_),
    .Y(_07435_));
 OAI21x1_ASAP7_75t_R _30277_ (.A1(_07249_),
    .A2(_07343_),
    .B(_07435_),
    .Y(_07436_));
 AOI21x1_ASAP7_75t_R _30278_ (.A1(_07274_),
    .A2(_07436_),
    .B(_07360_),
    .Y(_07437_));
 NAND2x1_ASAP7_75t_R _30279_ (.A(_07434_),
    .B(_07437_),
    .Y(_07438_));
 NOR2x2_ASAP7_75t_R _30280_ (.A(_07153_),
    .B(_07298_),
    .Y(_07439_));
 NAND2x2_ASAP7_75t_R _30281_ (.A(_07347_),
    .B(_07439_),
    .Y(_07440_));
 OAI21x1_ASAP7_75t_R _30282_ (.A1(net561),
    .A2(_07331_),
    .B(_07205_),
    .Y(_07441_));
 AOI21x1_ASAP7_75t_R _30283_ (.A1(_07440_),
    .A2(_07441_),
    .B(_07196_),
    .Y(_07442_));
 OAI21x1_ASAP7_75t_R _30284_ (.A1(_07133_),
    .A2(net947),
    .B(_07154_),
    .Y(_07443_));
 NOR2x1_ASAP7_75t_R _30285_ (.A(_07273_),
    .B(_07443_),
    .Y(_07444_));
 OAI21x1_ASAP7_75t_R _30286_ (.A1(net932),
    .A2(_07187_),
    .B(_07207_),
    .Y(_07445_));
 NOR2x1_ASAP7_75t_R _30287_ (.A(_07444_),
    .B(_07445_),
    .Y(_07446_));
 OAI21x1_ASAP7_75t_R _30288_ (.A1(_07442_),
    .A2(_07446_),
    .B(_07185_),
    .Y(_07447_));
 AOI21x1_ASAP7_75t_R _30289_ (.A1(_07438_),
    .A2(_07447_),
    .B(_07216_),
    .Y(_07448_));
 AOI21x1_ASAP7_75t_R _30290_ (.A1(_07418_),
    .A2(_07430_),
    .B(_07448_),
    .Y(_07449_));
 INVx2_ASAP7_75t_R _30291_ (.A(_07224_),
    .Y(_07450_));
 OAI21x1_ASAP7_75t_R _30292_ (.A1(_16067_),
    .A2(_16069_),
    .B(_07155_),
    .Y(_07451_));
 OAI21x1_ASAP7_75t_R _30293_ (.A1(_07450_),
    .A2(_07451_),
    .B(_07260_),
    .Y(_07452_));
 AOI21x1_ASAP7_75t_R _30294_ (.A1(_00417_),
    .A2(_07221_),
    .B(_07452_),
    .Y(_07453_));
 NOR2x1_ASAP7_75t_R _30295_ (.A(_07147_),
    .B(_07204_),
    .Y(_07454_));
 AOI22x1_ASAP7_75t_R _30296_ (.A1(_07454_),
    .A2(_07322_),
    .B1(_07137_),
    .B2(_07287_),
    .Y(_07455_));
 OAI21x1_ASAP7_75t_R _30297_ (.A1(_07220_),
    .A2(_07455_),
    .B(_07310_),
    .Y(_07456_));
 NOR2x1_ASAP7_75t_R _30298_ (.A(_07453_),
    .B(_07456_),
    .Y(_07457_));
 NAND2x1_ASAP7_75t_R _30299_ (.A(_00418_),
    .B(_07167_),
    .Y(_07458_));
 AOI21x1_ASAP7_75t_R _30300_ (.A1(_07458_),
    .A2(_07419_),
    .B(_07196_),
    .Y(_07459_));
 OR2x2_ASAP7_75t_R _30301_ (.A(_01278_),
    .B(_07238_),
    .Y(_07460_));
 AOI21x1_ASAP7_75t_R _30302_ (.A1(_07460_),
    .A2(_07413_),
    .B(_07174_),
    .Y(_07461_));
 OAI21x1_ASAP7_75t_R _30303_ (.A1(_07459_),
    .A2(_07461_),
    .B(_07216_),
    .Y(_07462_));
 NAND2x1_ASAP7_75t_R _30304_ (.A(_07241_),
    .B(_07462_),
    .Y(_07463_));
 OA21x2_ASAP7_75t_R _30305_ (.A1(_01276_),
    .A2(_07282_),
    .B(_07173_),
    .Y(_07464_));
 OAI21x1_ASAP7_75t_R _30306_ (.A1(_16077_),
    .A2(_07296_),
    .B(_07353_),
    .Y(_07465_));
 AOI21x1_ASAP7_75t_R _30307_ (.A1(_07464_),
    .A2(_07465_),
    .B(_07215_),
    .Y(_07466_));
 AOI21x1_ASAP7_75t_R _30308_ (.A1(_07322_),
    .A2(_07287_),
    .B(_07233_),
    .Y(_07467_));
 OAI21x1_ASAP7_75t_R _30309_ (.A1(_07249_),
    .A2(_07381_),
    .B(_07205_),
    .Y(_07468_));
 NAND2x1_ASAP7_75t_R _30310_ (.A(_07467_),
    .B(_07468_),
    .Y(_07469_));
 AOI21x1_ASAP7_75t_R _30311_ (.A1(_07466_),
    .A2(_07469_),
    .B(_07241_),
    .Y(_07470_));
 NAND2x2_ASAP7_75t_R _30312_ (.A(_07255_),
    .B(net940),
    .Y(_07471_));
 NAND2x2_ASAP7_75t_R _30313_ (.A(_07471_),
    .B(_07133_),
    .Y(_07472_));
 AOI21x1_ASAP7_75t_R _30314_ (.A1(_07472_),
    .A2(_07422_),
    .B(_07221_),
    .Y(_07473_));
 AO21x1_ASAP7_75t_R _30315_ (.A1(_07276_),
    .A2(_07304_),
    .B(_07260_),
    .Y(_07474_));
 INVx2_ASAP7_75t_R _30316_ (.A(_07279_),
    .Y(_07475_));
 AO21x1_ASAP7_75t_R _30317_ (.A1(_07135_),
    .A2(_07475_),
    .B(_07147_),
    .Y(_07476_));
 NAND2x1_ASAP7_75t_R _30318_ (.A(_07146_),
    .B(_07151_),
    .Y(_07477_));
 AND2x2_ASAP7_75t_R _30319_ (.A(_07477_),
    .B(_07173_),
    .Y(_07478_));
 AOI21x1_ASAP7_75t_R _30320_ (.A1(_07476_),
    .A2(_07478_),
    .B(_07262_),
    .Y(_07479_));
 OAI21x1_ASAP7_75t_R _30321_ (.A1(_07473_),
    .A2(_07474_),
    .B(_07479_),
    .Y(_07480_));
 AOI21x1_ASAP7_75t_R _30322_ (.A1(_07470_),
    .A2(_07480_),
    .B(_07271_),
    .Y(_07481_));
 OAI21x1_ASAP7_75t_R _30323_ (.A1(_07457_),
    .A2(_07463_),
    .B(_07481_),
    .Y(_07482_));
 OAI21x1_ASAP7_75t_R _30324_ (.A1(_07407_),
    .A2(_07449_),
    .B(_07482_),
    .Y(_00154_));
 INVx1_ASAP7_75t_R _30325_ (.A(_07171_),
    .Y(_07483_));
 OAI21x1_ASAP7_75t_R _30326_ (.A1(_07483_),
    .A2(_07382_),
    .B(_07277_),
    .Y(_07484_));
 AO21x1_ASAP7_75t_R _30327_ (.A1(_16067_),
    .A2(_16064_),
    .B(_07187_),
    .Y(_07485_));
 OA21x2_ASAP7_75t_R _30328_ (.A1(_07443_),
    .A2(_07201_),
    .B(_07173_),
    .Y(_07486_));
 AOI21x1_ASAP7_75t_R _30329_ (.A1(_07485_),
    .A2(_07486_),
    .B(_07360_),
    .Y(_07487_));
 NAND2x1_ASAP7_75t_R _30330_ (.A(_07484_),
    .B(_07487_),
    .Y(_07488_));
 NOR2x1_ASAP7_75t_R _30331_ (.A(_07204_),
    .B(_07344_),
    .Y(_07489_));
 AND2x2_ASAP7_75t_R _30332_ (.A(_07152_),
    .B(_07353_),
    .Y(_07490_));
 OAI21x1_ASAP7_75t_R _30333_ (.A1(_07489_),
    .A2(_07490_),
    .B(_07277_),
    .Y(_07491_));
 NAND2x1_ASAP7_75t_R _30334_ (.A(_07232_),
    .B(_07432_),
    .Y(_07492_));
 OA21x2_ASAP7_75t_R _30335_ (.A1(_07424_),
    .A2(_07379_),
    .B(_07173_),
    .Y(_07493_));
 AOI21x1_ASAP7_75t_R _30336_ (.A1(_07492_),
    .A2(_07493_),
    .B(_07302_),
    .Y(_07494_));
 AOI21x1_ASAP7_75t_R _30337_ (.A1(_07494_),
    .A2(_07491_),
    .B(_07262_),
    .Y(_07495_));
 NAND2x1_ASAP7_75t_R _30338_ (.A(_07495_),
    .B(_07488_),
    .Y(_07496_));
 AO21x1_ASAP7_75t_R _30339_ (.A1(_07237_),
    .A2(_00412_),
    .B(_07146_),
    .Y(_07497_));
 NOR2x1_ASAP7_75t_R _30340_ (.A(_07250_),
    .B(_07497_),
    .Y(_07498_));
 OAI21x1_ASAP7_75t_R _30341_ (.A1(_07323_),
    .A2(_07339_),
    .B(_07219_),
    .Y(_07499_));
 NOR2x1_ASAP7_75t_R _30342_ (.A(_07498_),
    .B(_07499_),
    .Y(_07500_));
 AO21x1_ASAP7_75t_R _30343_ (.A1(_07246_),
    .A2(_07150_),
    .B(_07282_),
    .Y(_07501_));
 INVx1_ASAP7_75t_R _30344_ (.A(_07296_),
    .Y(_07502_));
 OAI21x1_ASAP7_75t_R _30345_ (.A1(_07193_),
    .A2(_07502_),
    .B(_07167_),
    .Y(_07503_));
 AOI21x1_ASAP7_75t_R _30346_ (.A1(_07501_),
    .A2(_07503_),
    .B(_07260_),
    .Y(_07504_));
 OAI21x1_ASAP7_75t_R _30347_ (.A1(_07500_),
    .A2(_07504_),
    .B(_07325_),
    .Y(_07505_));
 NOR2x1_ASAP7_75t_R _30348_ (.A(_07225_),
    .B(_07226_),
    .Y(_07506_));
 NOR2x1_ASAP7_75t_R _30349_ (.A(_07207_),
    .B(_07506_),
    .Y(_07507_));
 INVx2_ASAP7_75t_R _30350_ (.A(_07249_),
    .Y(_07508_));
 NAND2x1_ASAP7_75t_R _30351_ (.A(_07296_),
    .B(_07508_),
    .Y(_07509_));
 AOI21x1_ASAP7_75t_R _30352_ (.A1(_07507_),
    .A2(_07509_),
    .B(_07360_),
    .Y(_07510_));
 AO21x1_ASAP7_75t_R _30353_ (.A1(_07127_),
    .A2(net950),
    .B(_01273_),
    .Y(_07511_));
 AO21x1_ASAP7_75t_R _30354_ (.A1(_07246_),
    .A2(_07511_),
    .B(_07238_),
    .Y(_07512_));
 NAND2x1_ASAP7_75t_R _30355_ (.A(_07512_),
    .B(_07337_),
    .Y(_07513_));
 AOI21x1_ASAP7_75t_R _30356_ (.A1(_07510_),
    .A2(_07513_),
    .B(_07215_),
    .Y(_07514_));
 AOI21x1_ASAP7_75t_R _30357_ (.A1(_07505_),
    .A2(_07514_),
    .B(_07271_),
    .Y(_07515_));
 NAND2x1_ASAP7_75t_R _30358_ (.A(_07515_),
    .B(_07496_),
    .Y(_07516_));
 INVx3_ASAP7_75t_R _30359_ (.A(_07414_),
    .Y(_07517_));
 AO21x1_ASAP7_75t_R _30360_ (.A1(_07472_),
    .A2(_07517_),
    .B(_07226_),
    .Y(_07518_));
 AOI21x1_ASAP7_75t_R _30361_ (.A1(_07246_),
    .A2(_07258_),
    .B(_07184_),
    .Y(_07519_));
 NAND2x1_ASAP7_75t_R _30362_ (.A(_07518_),
    .B(_07519_),
    .Y(_07520_));
 NAND2x2_ASAP7_75t_R _30363_ (.A(_07238_),
    .B(_07273_),
    .Y(_07521_));
 NAND3x1_ASAP7_75t_R _30364_ (.A(_07440_),
    .B(_07184_),
    .C(_07521_),
    .Y(_07522_));
 AOI21x1_ASAP7_75t_R _30365_ (.A1(_07520_),
    .A2(_07522_),
    .B(_07164_),
    .Y(_07523_));
 NOR2x2_ASAP7_75t_R _30366_ (.A(_07154_),
    .B(_07246_),
    .Y(_07524_));
 NAND2x1_ASAP7_75t_R _30367_ (.A(_07184_),
    .B(_07524_),
    .Y(_07525_));
 NAND2x1_ASAP7_75t_R _30368_ (.A(_07308_),
    .B(_07525_),
    .Y(_07526_));
 NAND2x1_ASAP7_75t_R _30369_ (.A(_07224_),
    .B(_07304_),
    .Y(_07527_));
 AOI21x1_ASAP7_75t_R _30370_ (.A1(_07171_),
    .A2(_07527_),
    .B(_07360_),
    .Y(_07528_));
 OAI21x1_ASAP7_75t_R _30371_ (.A1(_07526_),
    .A2(_07528_),
    .B(_07215_),
    .Y(_07529_));
 NOR2x1_ASAP7_75t_R _30372_ (.A(_07523_),
    .B(_07529_),
    .Y(_07530_));
 NAND2x1_ASAP7_75t_R _30373_ (.A(_07302_),
    .B(_07445_),
    .Y(_07531_));
 AO21x2_ASAP7_75t_R _30374_ (.A1(_07472_),
    .A2(_07511_),
    .B(_07226_),
    .Y(_07532_));
 AOI21x1_ASAP7_75t_R _30375_ (.A1(_07532_),
    .A2(_07386_),
    .B(_07196_),
    .Y(_07533_));
 OAI21x1_ASAP7_75t_R _30376_ (.A1(_07531_),
    .A2(_07533_),
    .B(_07310_),
    .Y(_07534_));
 AO21x1_ASAP7_75t_R _30377_ (.A1(_07135_),
    .A2(_07517_),
    .B(_07238_),
    .Y(_07535_));
 NAND2x2_ASAP7_75t_R _30378_ (.A(_16064_),
    .B(_07363_),
    .Y(_07536_));
 AOI21x1_ASAP7_75t_R _30379_ (.A1(_07238_),
    .A2(_07273_),
    .B(_07173_),
    .Y(_07537_));
 NAND3x1_ASAP7_75t_R _30380_ (.A(_07535_),
    .B(_07536_),
    .C(_07537_),
    .Y(_07538_));
 NAND2x1_ASAP7_75t_R _30381_ (.A(_07365_),
    .B(_07319_),
    .Y(_07539_));
 AOI21x1_ASAP7_75t_R _30382_ (.A1(_07538_),
    .A2(_07539_),
    .B(_07293_),
    .Y(_07540_));
 NOR2x1_ASAP7_75t_R _30383_ (.A(_07534_),
    .B(_07540_),
    .Y(_07541_));
 OAI21x1_ASAP7_75t_R _30384_ (.A1(_07530_),
    .A2(_07541_),
    .B(_07271_),
    .Y(_07542_));
 NAND2x1_ASAP7_75t_R _30385_ (.A(_07542_),
    .B(_07516_),
    .Y(_00155_));
 BUFx6f_ASAP7_75t_R _30386_ (.A(_07238_),
    .Y(_07543_));
 AOI21x1_ASAP7_75t_R _30387_ (.A1(_07346_),
    .A2(_07335_),
    .B(_07543_),
    .Y(_07544_));
 AND2x2_ASAP7_75t_R _30388_ (.A(_07508_),
    .B(_07299_),
    .Y(_07545_));
 OAI21x1_ASAP7_75t_R _30389_ (.A1(_07544_),
    .A2(_07545_),
    .B(_07208_),
    .Y(_07546_));
 NOR2x1_ASAP7_75t_R _30390_ (.A(_07193_),
    .B(_07195_),
    .Y(_07547_));
 OA21x2_ASAP7_75t_R _30391_ (.A1(_07390_),
    .A2(_07203_),
    .B(_07251_),
    .Y(_07548_));
 OAI21x1_ASAP7_75t_R _30392_ (.A1(_07547_),
    .A2(_07548_),
    .B(_07220_),
    .Y(_07549_));
 AOI21x1_ASAP7_75t_R _30393_ (.A1(_07546_),
    .A2(_07549_),
    .B(_07263_),
    .Y(_07550_));
 AO21x1_ASAP7_75t_R _30394_ (.A1(_16077_),
    .A2(_07205_),
    .B(_07277_),
    .Y(_07551_));
 NOR2x1_ASAP7_75t_R _30395_ (.A(_07244_),
    .B(_07187_),
    .Y(_07552_));
 OAI21x1_ASAP7_75t_R _30396_ (.A1(_07551_),
    .A2(_07552_),
    .B(_07310_),
    .Y(_07553_));
 OA21x2_ASAP7_75t_R _30397_ (.A1(_07084_),
    .A2(_07076_),
    .B(_07090_),
    .Y(_07554_));
 OA21x2_ASAP7_75t_R _30398_ (.A1(_07089_),
    .A2(_07086_),
    .B(_01102_),
    .Y(_07555_));
 OAI21x1_ASAP7_75t_R _30399_ (.A1(_07554_),
    .A2(_07555_),
    .B(_07129_),
    .Y(_07556_));
 NAND2x2_ASAP7_75t_R _30400_ (.A(_07152_),
    .B(_07556_),
    .Y(_07557_));
 AOI211x1_ASAP7_75t_R _30401_ (.A1(_07557_),
    .A2(_07221_),
    .B(_07380_),
    .C(_07220_),
    .Y(_07558_));
 OAI21x1_ASAP7_75t_R _30402_ (.A1(_07553_),
    .A2(_07558_),
    .B(_07241_),
    .Y(_07559_));
 OAI21x1_ASAP7_75t_R _30403_ (.A1(_07550_),
    .A2(_07559_),
    .B(_07271_),
    .Y(_07560_));
 NAND2x2_ASAP7_75t_R _30404_ (.A(_07238_),
    .B(_07286_),
    .Y(_07561_));
 OA21x2_ASAP7_75t_R _30405_ (.A1(_00419_),
    .A2(_07167_),
    .B(_07233_),
    .Y(_07562_));
 AOI21x1_ASAP7_75t_R _30406_ (.A1(_07561_),
    .A2(_07562_),
    .B(_07310_),
    .Y(_07563_));
 NAND2x1_ASAP7_75t_R _30407_ (.A(_07338_),
    .B(_07314_),
    .Y(_07564_));
 NAND2x2_ASAP7_75t_R _30408_ (.A(_07299_),
    .B(_07335_),
    .Y(_07565_));
 AO21x1_ASAP7_75t_R _30409_ (.A1(_07564_),
    .A2(_07565_),
    .B(_07174_),
    .Y(_07566_));
 NAND2x1_ASAP7_75t_R _30410_ (.A(_07563_),
    .B(_07566_),
    .Y(_07567_));
 AO21x1_ASAP7_75t_R _30411_ (.A1(_07398_),
    .A2(_07251_),
    .B(_07233_),
    .Y(_07568_));
 AOI21x1_ASAP7_75t_R _30412_ (.A1(_07543_),
    .A2(_07200_),
    .B(_07568_),
    .Y(_07569_));
 AO21x1_ASAP7_75t_R _30413_ (.A1(_16074_),
    .A2(net946),
    .B(_07238_),
    .Y(_07570_));
 OAI21x1_ASAP7_75t_R _30414_ (.A1(_07286_),
    .A2(_07570_),
    .B(_07260_),
    .Y(_07571_));
 NOR2x1_ASAP7_75t_R _30415_ (.A(_07571_),
    .B(_07228_),
    .Y(_07572_));
 OAI21x1_ASAP7_75t_R _30416_ (.A1(_07569_),
    .A2(_07572_),
    .B(_07263_),
    .Y(_07573_));
 AOI21x1_ASAP7_75t_R _30417_ (.A1(_07567_),
    .A2(_07573_),
    .B(_07241_),
    .Y(_07574_));
 OAI21x1_ASAP7_75t_R _30418_ (.A1(_07382_),
    .A2(_07452_),
    .B(_07293_),
    .Y(_07575_));
 OA21x2_ASAP7_75t_R _30419_ (.A1(_07450_),
    .A2(_07203_),
    .B(_07205_),
    .Y(_07576_));
 NOR2x2_ASAP7_75t_R _30420_ (.A(_07188_),
    .B(net943),
    .Y(_07577_));
 OAI21x1_ASAP7_75t_R _30421_ (.A1(_07577_),
    .A2(_07239_),
    .B(_07196_),
    .Y(_07578_));
 NOR2x1_ASAP7_75t_R _30422_ (.A(_07576_),
    .B(_07578_),
    .Y(_07579_));
 AO21x1_ASAP7_75t_R _30423_ (.A1(_16067_),
    .A2(_07225_),
    .B(_07226_),
    .Y(_07580_));
 AOI21x1_ASAP7_75t_R _30424_ (.A1(_07373_),
    .A2(_07580_),
    .B(_07349_),
    .Y(_07581_));
 NOR2x1_ASAP7_75t_R _30425_ (.A(_07390_),
    .B(_07299_),
    .Y(_07582_));
 AOI21x1_ASAP7_75t_R _30426_ (.A1(_07196_),
    .A2(_07582_),
    .B(_07302_),
    .Y(_07583_));
 OAI21x1_ASAP7_75t_R _30427_ (.A1(_07208_),
    .A2(_07581_),
    .B(_07583_),
    .Y(_07584_));
 OAI21x1_ASAP7_75t_R _30428_ (.A1(_07575_),
    .A2(_07579_),
    .B(_07584_),
    .Y(_07585_));
 NOR2x1_ASAP7_75t_R _30429_ (.A(_07216_),
    .B(_07585_),
    .Y(_07586_));
 NAND2x1_ASAP7_75t_R _30430_ (.A(_07282_),
    .B(_16067_),
    .Y(_07587_));
 AOI21x1_ASAP7_75t_R _30431_ (.A1(_07155_),
    .A2(_07151_),
    .B(_07207_),
    .Y(_07588_));
 OAI21x1_ASAP7_75t_R _30432_ (.A1(_16074_),
    .A2(_07587_),
    .B(_07588_),
    .Y(_07589_));
 INVx1_ASAP7_75t_R _30433_ (.A(_07315_),
    .Y(_07590_));
 OAI21x1_ASAP7_75t_R _30434_ (.A1(_07589_),
    .A2(_07590_),
    .B(_07293_),
    .Y(_07591_));
 OAI21x1_ASAP7_75t_R _30435_ (.A1(_07443_),
    .A2(_07306_),
    .B(_07416_),
    .Y(_07592_));
 NOR2x1_ASAP7_75t_R _30436_ (.A(_07220_),
    .B(_07592_),
    .Y(_07593_));
 NOR2x1_ASAP7_75t_R _30437_ (.A(_07591_),
    .B(_07593_),
    .Y(_07594_));
 INVx1_ASAP7_75t_R _30438_ (.A(_07300_),
    .Y(_07595_));
 NAND2x1_ASAP7_75t_R _30439_ (.A(_07147_),
    .B(_07232_),
    .Y(_07596_));
 OAI21x1_ASAP7_75t_R _30440_ (.A1(net562),
    .A2(_07596_),
    .B(_07174_),
    .Y(_07597_));
 NOR2x1_ASAP7_75t_R _30441_ (.A(_07595_),
    .B(_07597_),
    .Y(_07598_));
 AO31x2_ASAP7_75t_R _30442_ (.A1(_07561_),
    .A2(_07431_),
    .A3(_07537_),
    .B(_07302_),
    .Y(_07599_));
 OAI21x1_ASAP7_75t_R _30443_ (.A1(_07598_),
    .A2(_07599_),
    .B(_07216_),
    .Y(_07600_));
 OAI21x1_ASAP7_75t_R _30444_ (.A1(_07594_),
    .A2(_07600_),
    .B(_07407_),
    .Y(_07601_));
 OAI22x1_ASAP7_75t_R _30445_ (.A1(_07560_),
    .A2(_07574_),
    .B1(_07586_),
    .B2(_07601_),
    .Y(_00156_));
 AO21x1_ASAP7_75t_R _30446_ (.A1(net942),
    .A2(_16077_),
    .B(_07282_),
    .Y(_07602_));
 OAI21x1_ASAP7_75t_R _30447_ (.A1(_07450_),
    .A2(_07602_),
    .B(_07561_),
    .Y(_07603_));
 OAI21x1_ASAP7_75t_R _30448_ (.A1(_07155_),
    .A2(_07414_),
    .B(_07219_),
    .Y(_07604_));
 AOI21x1_ASAP7_75t_R _30449_ (.A1(_07137_),
    .A2(_07402_),
    .B(_07604_),
    .Y(_07605_));
 AOI21x1_ASAP7_75t_R _30450_ (.A1(_07208_),
    .A2(_07603_),
    .B(_07605_),
    .Y(_07606_));
 OAI21x1_ASAP7_75t_R _30451_ (.A1(_07185_),
    .A2(_07606_),
    .B(_07216_),
    .Y(_07607_));
 NAND2x1_ASAP7_75t_R _30452_ (.A(_07150_),
    .B(_07376_),
    .Y(_07608_));
 OAI22x1_ASAP7_75t_R _30453_ (.A1(_07608_),
    .A2(_07221_),
    .B1(_07577_),
    .B2(_07259_),
    .Y(_07609_));
 NAND2x1_ASAP7_75t_R _30454_ (.A(_07260_),
    .B(_07587_),
    .Y(_07610_));
 NOR2x1_ASAP7_75t_R _30455_ (.A(_07577_),
    .B(_07239_),
    .Y(_07611_));
 OAI21x1_ASAP7_75t_R _30456_ (.A1(_07610_),
    .A2(_07611_),
    .B(_07325_),
    .Y(_07612_));
 AOI21x1_ASAP7_75t_R _30457_ (.A1(_07208_),
    .A2(_07609_),
    .B(_07612_),
    .Y(_07613_));
 NOR2x1_ASAP7_75t_R _30458_ (.A(_07607_),
    .B(_07613_),
    .Y(_07614_));
 AOI21x1_ASAP7_75t_R _30459_ (.A1(_07282_),
    .A2(_07273_),
    .B(_07163_),
    .Y(_07615_));
 NAND2x1_ASAP7_75t_R _30460_ (.A(_07615_),
    .B(_07536_),
    .Y(_07616_));
 NOR2x1_ASAP7_75t_R _30461_ (.A(_07202_),
    .B(_07616_),
    .Y(_07617_));
 NAND2x1_ASAP7_75t_R _30462_ (.A(_07570_),
    .B(_07364_),
    .Y(_07618_));
 OAI21x1_ASAP7_75t_R _30463_ (.A1(_07220_),
    .A2(_07618_),
    .B(_07293_),
    .Y(_07619_));
 NOR2x1_ASAP7_75t_R _30464_ (.A(_07617_),
    .B(_07619_),
    .Y(_07620_));
 AOI21x1_ASAP7_75t_R _30465_ (.A1(_07517_),
    .A2(_07332_),
    .B(_07251_),
    .Y(_07621_));
 AOI211x1_ASAP7_75t_R _30466_ (.A1(_07223_),
    .A2(_07221_),
    .B(_07621_),
    .C(_07208_),
    .Y(_07622_));
 NOR2x1_ASAP7_75t_R _30467_ (.A(_07256_),
    .B(_16074_),
    .Y(_07623_));
 NAND2x1_ASAP7_75t_R _30468_ (.A(_07471_),
    .B(_07167_),
    .Y(_07624_));
 OAI21x1_ASAP7_75t_R _30469_ (.A1(_07623_),
    .A2(_07624_),
    .B(_07196_),
    .Y(_07625_));
 OA21x2_ASAP7_75t_R _30470_ (.A1(_07296_),
    .A2(_16077_),
    .B(_07439_),
    .Y(_07626_));
 OAI21x1_ASAP7_75t_R _30471_ (.A1(_07625_),
    .A2(_07626_),
    .B(_07185_),
    .Y(_07627_));
 OAI21x1_ASAP7_75t_R _30472_ (.A1(_07622_),
    .A2(_07627_),
    .B(_07263_),
    .Y(_07628_));
 OAI21x1_ASAP7_75t_R _30473_ (.A1(_07620_),
    .A2(_07628_),
    .B(_07407_),
    .Y(_07629_));
 AO21x1_ASAP7_75t_R _30474_ (.A1(_16069_),
    .A2(_07205_),
    .B(_07277_),
    .Y(_07630_));
 OAI21x1_ASAP7_75t_R _30475_ (.A1(_07630_),
    .A2(_07192_),
    .B(_07185_),
    .Y(_07631_));
 NOR2x1_ASAP7_75t_R _30476_ (.A(_07236_),
    .B(_07247_),
    .Y(_07632_));
 AO21x1_ASAP7_75t_R _30477_ (.A1(_07335_),
    .A2(_07439_),
    .B(_07233_),
    .Y(_07633_));
 NOR2x1_ASAP7_75t_R _30478_ (.A(_07633_),
    .B(_07632_),
    .Y(_07634_));
 OAI21x1_ASAP7_75t_R _30479_ (.A1(_07631_),
    .A2(_07634_),
    .B(_07263_),
    .Y(_07635_));
 INVx1_ASAP7_75t_R _30480_ (.A(_07150_),
    .Y(_07636_));
 AO21x1_ASAP7_75t_R _30481_ (.A1(_07636_),
    .A2(_07205_),
    .B(_07233_),
    .Y(_07637_));
 AOI21x1_ASAP7_75t_R _30482_ (.A1(_07517_),
    .A2(_07376_),
    .B(_07543_),
    .Y(_07638_));
 OAI21x1_ASAP7_75t_R _30483_ (.A1(_07637_),
    .A2(_07638_),
    .B(_07293_),
    .Y(_07639_));
 AOI21x1_ASAP7_75t_R _30484_ (.A1(_07475_),
    .A2(_07508_),
    .B(_07543_),
    .Y(_07640_));
 AOI211x1_ASAP7_75t_R _30485_ (.A1(_07227_),
    .A2(_07276_),
    .B(_07640_),
    .C(_07208_),
    .Y(_07641_));
 NOR2x1_ASAP7_75t_R _30486_ (.A(_07639_),
    .B(_07641_),
    .Y(_07642_));
 OAI21x1_ASAP7_75t_R _30487_ (.A1(_07642_),
    .A2(_07635_),
    .B(_07271_),
    .Y(_07643_));
 OAI21x1_ASAP7_75t_R _30488_ (.A1(_07244_),
    .A2(_07424_),
    .B(_07164_),
    .Y(_07644_));
 AO21x1_ASAP7_75t_R _30489_ (.A1(_07402_),
    .A2(_07289_),
    .B(_07644_),
    .Y(_07645_));
 OA21x2_ASAP7_75t_R _30490_ (.A1(_07149_),
    .A2(_07251_),
    .B(_07260_),
    .Y(_07646_));
 AO21x1_ASAP7_75t_R _30491_ (.A1(_07249_),
    .A2(_16067_),
    .B(_07543_),
    .Y(_07647_));
 AOI21x1_ASAP7_75t_R _30492_ (.A1(_07646_),
    .A2(_07647_),
    .B(_07185_),
    .Y(_07648_));
 OA21x2_ASAP7_75t_R _30493_ (.A1(_16077_),
    .A2(_07471_),
    .B(_07167_),
    .Y(_07649_));
 NOR2x1_ASAP7_75t_R _30494_ (.A(_07164_),
    .B(_07649_),
    .Y(_07650_));
 AO21x1_ASAP7_75t_R _30495_ (.A1(_07375_),
    .A2(_07376_),
    .B(_07543_),
    .Y(_07651_));
 AO21x1_ASAP7_75t_R _30496_ (.A1(_07338_),
    .A2(_07279_),
    .B(_07233_),
    .Y(_07652_));
 OAI21x1_ASAP7_75t_R _30497_ (.A1(_07336_),
    .A2(_07652_),
    .B(_07325_),
    .Y(_07653_));
 AOI21x1_ASAP7_75t_R _30498_ (.A1(_07650_),
    .A2(_07651_),
    .B(_07653_),
    .Y(_07654_));
 AOI211x1_ASAP7_75t_R _30499_ (.A1(_07645_),
    .A2(_07648_),
    .B(_07654_),
    .C(_07263_),
    .Y(_07655_));
 OAI22x1_ASAP7_75t_R _30500_ (.A1(_07614_),
    .A2(_07629_),
    .B1(_07643_),
    .B2(_07655_),
    .Y(_00157_));
 AOI21x1_ASAP7_75t_R _30501_ (.A1(_07147_),
    .A2(net562),
    .B(_07207_),
    .Y(_07656_));
 OAI21x1_ASAP7_75t_R _30502_ (.A1(_07543_),
    .A2(_07472_),
    .B(_07656_),
    .Y(_07657_));
 INVx1_ASAP7_75t_R _30503_ (.A(_07314_),
    .Y(_07658_));
 AOI21x1_ASAP7_75t_R _30504_ (.A1(_07235_),
    .A2(_07658_),
    .B(_07221_),
    .Y(_07659_));
 NOR2x1_ASAP7_75t_R _30505_ (.A(_07659_),
    .B(_07657_),
    .Y(_07660_));
 AO21x1_ASAP7_75t_R _30506_ (.A1(_07636_),
    .A2(_07251_),
    .B(_07260_),
    .Y(_07661_));
 OA21x2_ASAP7_75t_R _30507_ (.A1(_07249_),
    .A2(net943),
    .B(_07543_),
    .Y(_07662_));
 OAI21x1_ASAP7_75t_R _30508_ (.A1(_07661_),
    .A2(_07662_),
    .B(_07241_),
    .Y(_07663_));
 OAI21x1_ASAP7_75t_R _30509_ (.A1(_07660_),
    .A2(_07663_),
    .B(_07216_),
    .Y(_07664_));
 AO21x1_ASAP7_75t_R _30510_ (.A1(_07419_),
    .A2(_07458_),
    .B(_07524_),
    .Y(_07665_));
 OA21x2_ASAP7_75t_R _30511_ (.A1(_07450_),
    .A2(_07250_),
    .B(_07543_),
    .Y(_07666_));
 INVx1_ASAP7_75t_R _30512_ (.A(_07424_),
    .Y(_07667_));
 AO21x1_ASAP7_75t_R _30513_ (.A1(_07667_),
    .A2(_07398_),
    .B(_07277_),
    .Y(_07668_));
 OAI21x1_ASAP7_75t_R _30514_ (.A1(_07666_),
    .A2(_07668_),
    .B(_07185_),
    .Y(_07669_));
 AOI21x1_ASAP7_75t_R _30515_ (.A1(_07208_),
    .A2(_07665_),
    .B(_07669_),
    .Y(_07670_));
 OAI21x1_ASAP7_75t_R _30516_ (.A1(_07664_),
    .A2(_07670_),
    .B(_07407_),
    .Y(_07671_));
 AND2x2_ASAP7_75t_R _30517_ (.A(_07439_),
    .B(_07232_),
    .Y(_07672_));
 AO21x1_ASAP7_75t_R _30518_ (.A1(_07363_),
    .A2(_07346_),
    .B(_07307_),
    .Y(_07673_));
 OAI21x1_ASAP7_75t_R _30519_ (.A1(_07672_),
    .A2(_07673_),
    .B(_07293_),
    .Y(_07674_));
 AO21x1_ASAP7_75t_R _30520_ (.A1(_01277_),
    .A2(_01275_),
    .B(_07282_),
    .Y(_07675_));
 OAI21x1_ASAP7_75t_R _30521_ (.A1(_07358_),
    .A2(_07577_),
    .B(_07167_),
    .Y(_07676_));
 NAND2x1_ASAP7_75t_R _30522_ (.A(_07675_),
    .B(_07676_),
    .Y(_07677_));
 AOI21x1_ASAP7_75t_R _30523_ (.A1(_07325_),
    .A2(_07677_),
    .B(_07208_),
    .Y(_07678_));
 NAND2x1_ASAP7_75t_R _30524_ (.A(_07674_),
    .B(_07678_),
    .Y(_07679_));
 OA21x2_ASAP7_75t_R _30525_ (.A1(_07338_),
    .A2(_07475_),
    .B(_07521_),
    .Y(_07680_));
 OAI21x1_ASAP7_75t_R _30526_ (.A1(_07249_),
    .A2(_07323_),
    .B(_07680_),
    .Y(_07681_));
 NAND2x1_ASAP7_75t_R _30527_ (.A(_07477_),
    .B(_07521_),
    .Y(_07682_));
 AO21x1_ASAP7_75t_R _30528_ (.A1(_07312_),
    .A2(_07155_),
    .B(_07219_),
    .Y(_07683_));
 AO21x1_ASAP7_75t_R _30529_ (.A1(_07360_),
    .A2(_07682_),
    .B(_07683_),
    .Y(_07684_));
 AO21x1_ASAP7_75t_R _30530_ (.A1(_07241_),
    .A2(_07681_),
    .B(_07684_),
    .Y(_07685_));
 AOI21x1_ASAP7_75t_R _30531_ (.A1(_07679_),
    .A2(_07685_),
    .B(_07216_),
    .Y(_07686_));
 NAND2x1_ASAP7_75t_R _30532_ (.A(_07338_),
    .B(_07331_),
    .Y(_07687_));
 AND3x1_ASAP7_75t_R _30533_ (.A(_07536_),
    .B(_07615_),
    .C(_07687_),
    .Y(_07688_));
 AO21x1_ASAP7_75t_R _30534_ (.A1(_07252_),
    .A2(_07356_),
    .B(_07325_),
    .Y(_07689_));
 OAI21x1_ASAP7_75t_R _30535_ (.A1(_07688_),
    .A2(_07689_),
    .B(_07263_),
    .Y(_07690_));
 OAI21x1_ASAP7_75t_R _30536_ (.A1(_07193_),
    .A2(_07191_),
    .B(_07543_),
    .Y(_07691_));
 NAND2x1_ASAP7_75t_R _30537_ (.A(_07251_),
    .B(_07412_),
    .Y(_07692_));
 AO21x1_ASAP7_75t_R _30538_ (.A1(_07691_),
    .A2(_07692_),
    .B(_07164_),
    .Y(_07693_));
 AO21x1_ASAP7_75t_R _30539_ (.A1(_07508_),
    .A2(_07296_),
    .B(_07338_),
    .Y(_07694_));
 AO21x1_ASAP7_75t_R _30540_ (.A1(_07235_),
    .A2(_07421_),
    .B(_07205_),
    .Y(_07695_));
 AO21x1_ASAP7_75t_R _30541_ (.A1(_07694_),
    .A2(_07695_),
    .B(_07220_),
    .Y(_07696_));
 AOI21x1_ASAP7_75t_R _30542_ (.A1(_07693_),
    .A2(_07696_),
    .B(_07241_),
    .Y(_07697_));
 AOI21x1_ASAP7_75t_R _30543_ (.A1(_07338_),
    .A2(_07193_),
    .B(_07233_),
    .Y(_07698_));
 AO21x1_ASAP7_75t_R _30544_ (.A1(_07517_),
    .A2(_07246_),
    .B(_07147_),
    .Y(_07699_));
 NAND2x1_ASAP7_75t_R _30545_ (.A(_07698_),
    .B(_07699_),
    .Y(_07700_));
 AOI21x1_ASAP7_75t_R _30546_ (.A1(_00421_),
    .A2(_07205_),
    .B(_07277_),
    .Y(_07701_));
 NAND2x1_ASAP7_75t_R _30547_ (.A(_07439_),
    .B(_07335_),
    .Y(_07702_));
 AOI21x1_ASAP7_75t_R _30548_ (.A1(_07701_),
    .A2(_07702_),
    .B(_07302_),
    .Y(_07703_));
 AOI21x1_ASAP7_75t_R _30549_ (.A1(_07703_),
    .A2(_07700_),
    .B(_07310_),
    .Y(_07704_));
 INVx1_ASAP7_75t_R _30550_ (.A(_07410_),
    .Y(_07705_));
 AOI21x1_ASAP7_75t_R _30551_ (.A1(_07305_),
    .A2(_07565_),
    .B(_07174_),
    .Y(_07706_));
 OAI21x1_ASAP7_75t_R _30552_ (.A1(_07705_),
    .A2(_07706_),
    .B(_07241_),
    .Y(_07707_));
 AOI21x1_ASAP7_75t_R _30553_ (.A1(_07704_),
    .A2(_07707_),
    .B(_07407_),
    .Y(_07708_));
 OAI21x1_ASAP7_75t_R _30554_ (.A1(_07690_),
    .A2(_07697_),
    .B(_07708_),
    .Y(_07709_));
 OAI21x1_ASAP7_75t_R _30555_ (.A1(_07671_),
    .A2(_07686_),
    .B(_07709_),
    .Y(_00158_));
 AOI211x1_ASAP7_75t_R _30556_ (.A1(_07346_),
    .A2(_07506_),
    .B(_07524_),
    .C(_07164_),
    .Y(_07710_));
 NOR2x1_ASAP7_75t_R _30557_ (.A(_07424_),
    .B(_07199_),
    .Y(_07711_));
 OAI21x1_ASAP7_75t_R _30558_ (.A1(_07221_),
    .A2(_07306_),
    .B(_07196_),
    .Y(_07712_));
 OAI21x1_ASAP7_75t_R _30559_ (.A1(_07711_),
    .A2(_07712_),
    .B(_07293_),
    .Y(_07713_));
 OAI21x1_ASAP7_75t_R _30560_ (.A1(_07710_),
    .A2(_07713_),
    .B(_07216_),
    .Y(_07714_));
 NOR2x1_ASAP7_75t_R _30561_ (.A(_07199_),
    .B(_07239_),
    .Y(_07715_));
 NAND2x1_ASAP7_75t_R _30562_ (.A(_16064_),
    .B(_07194_),
    .Y(_07716_));
 OAI21x1_ASAP7_75t_R _30563_ (.A1(_07349_),
    .A2(_07580_),
    .B(_07716_),
    .Y(_07717_));
 AOI21x1_ASAP7_75t_R _30564_ (.A1(_07164_),
    .A2(_07717_),
    .B(_07293_),
    .Y(_07718_));
 OA21x2_ASAP7_75t_R _30565_ (.A1(_07452_),
    .A2(_07715_),
    .B(_07718_),
    .Y(_07719_));
 NOR2x1_ASAP7_75t_R _30566_ (.A(_07714_),
    .B(_07719_),
    .Y(_07720_));
 NAND2x1_ASAP7_75t_R _30567_ (.A(_07174_),
    .B(_07468_),
    .Y(_07721_));
 NAND2x1_ASAP7_75t_R _30568_ (.A(_07246_),
    .B(_07258_),
    .Y(_07722_));
 AOI21x1_ASAP7_75t_R _30569_ (.A1(_07232_),
    .A2(_07353_),
    .B(_07260_),
    .Y(_07723_));
 AOI21x1_ASAP7_75t_R _30570_ (.A1(_07722_),
    .A2(_07723_),
    .B(_07325_),
    .Y(_07724_));
 OA21x2_ASAP7_75t_R _30571_ (.A1(_07721_),
    .A2(_07672_),
    .B(_07724_),
    .Y(_07725_));
 OAI21x1_ASAP7_75t_R _30572_ (.A1(_07259_),
    .A2(_07306_),
    .B(_07196_),
    .Y(_07726_));
 AOI21x1_ASAP7_75t_R _30573_ (.A1(_07152_),
    .A2(_07422_),
    .B(_07221_),
    .Y(_07727_));
 NOR2x1_ASAP7_75t_R _30574_ (.A(_07726_),
    .B(_07727_),
    .Y(_07728_));
 NOR2x1_ASAP7_75t_R _30575_ (.A(_07277_),
    .B(_07399_),
    .Y(_07729_));
 AO21x1_ASAP7_75t_R _30576_ (.A1(_07729_),
    .A2(_07565_),
    .B(_07293_),
    .Y(_07730_));
 OAI21x1_ASAP7_75t_R _30577_ (.A1(_07728_),
    .A2(_07730_),
    .B(_07263_),
    .Y(_07731_));
 OAI21x1_ASAP7_75t_R _30578_ (.A1(_07725_),
    .A2(_07731_),
    .B(_07271_),
    .Y(_07732_));
 NOR2x1_ASAP7_75t_R _30579_ (.A(_07151_),
    .B(_07184_),
    .Y(_07733_));
 OAI21x1_ASAP7_75t_R _30580_ (.A1(_07167_),
    .A2(_07312_),
    .B(_07443_),
    .Y(_07734_));
 AOI21x1_ASAP7_75t_R _30581_ (.A1(_07733_),
    .A2(_07734_),
    .B(_07277_),
    .Y(_07735_));
 NOR2x1_ASAP7_75t_R _30582_ (.A(_07636_),
    .B(_07247_),
    .Y(_07736_));
 NOR2x1_ASAP7_75t_R _30583_ (.A(_07259_),
    .B(_07557_),
    .Y(_07737_));
 OAI21x1_ASAP7_75t_R _30584_ (.A1(_07737_),
    .A2(_07736_),
    .B(_07360_),
    .Y(_07738_));
 NAND2x1_ASAP7_75t_R _30585_ (.A(_07735_),
    .B(_07738_),
    .Y(_07739_));
 NOR2x1_ASAP7_75t_R _30586_ (.A(_07357_),
    .B(_07184_),
    .Y(_07740_));
 AOI21x1_ASAP7_75t_R _30587_ (.A1(_07740_),
    .A2(_07676_),
    .B(_07174_),
    .Y(_07741_));
 NAND2x1_ASAP7_75t_R _30588_ (.A(_07346_),
    .B(_07287_),
    .Y(_07742_));
 NAND3x1_ASAP7_75t_R _30589_ (.A(_07532_),
    .B(_07360_),
    .C(_07742_),
    .Y(_07743_));
 AOI21x1_ASAP7_75t_R _30590_ (.A1(_07741_),
    .A2(_07743_),
    .B(_07216_),
    .Y(_07744_));
 NAND2x1_ASAP7_75t_R _30591_ (.A(_07744_),
    .B(_07739_),
    .Y(_07745_));
 AO22x1_ASAP7_75t_R _30592_ (.A1(_07135_),
    .A2(_07353_),
    .B1(_07335_),
    .B2(_07258_),
    .Y(_07746_));
 NOR2x1_ASAP7_75t_R _30593_ (.A(_01277_),
    .B(_07194_),
    .Y(_07747_));
 AOI21x1_ASAP7_75t_R _30594_ (.A1(_07251_),
    .A2(_07273_),
    .B(_07747_),
    .Y(_07748_));
 AOI21x1_ASAP7_75t_R _30595_ (.A1(_07656_),
    .A2(_07748_),
    .B(_07325_),
    .Y(_07749_));
 OAI21x1_ASAP7_75t_R _30596_ (.A1(_07220_),
    .A2(_07746_),
    .B(_07749_),
    .Y(_07750_));
 AOI21x1_ASAP7_75t_R _30597_ (.A1(_00419_),
    .A2(_07205_),
    .B(_07207_),
    .Y(_07751_));
 AOI21x1_ASAP7_75t_R _30598_ (.A1(_07751_),
    .A2(_07313_),
    .B(_07302_),
    .Y(_07752_));
 OAI21x1_ASAP7_75t_R _30599_ (.A1(net943),
    .A2(_07249_),
    .B(_07338_),
    .Y(_07753_));
 OA21x2_ASAP7_75t_R _30600_ (.A1(_07257_),
    .A2(_07379_),
    .B(_07207_),
    .Y(_07754_));
 NAND2x1_ASAP7_75t_R _30601_ (.A(_07753_),
    .B(_07754_),
    .Y(_07755_));
 AOI21x1_ASAP7_75t_R _30602_ (.A1(_07752_),
    .A2(_07755_),
    .B(_07310_),
    .Y(_07756_));
 AOI21x1_ASAP7_75t_R _30603_ (.A1(_07750_),
    .A2(_07756_),
    .B(_07271_),
    .Y(_07757_));
 NAND2x1_ASAP7_75t_R _30604_ (.A(_07757_),
    .B(_07745_),
    .Y(_07758_));
 OAI21x1_ASAP7_75t_R _30605_ (.A1(_07720_),
    .A2(_07732_),
    .B(_07758_),
    .Y(_00159_));
 INVx1_ASAP7_75t_R _30606_ (.A(_00728_),
    .Y(_07759_));
 AND5x1_ASAP7_75t_R _30607_ (.A(_08080_),
    .B(_07759_),
    .C(_00726_),
    .D(_00727_),
    .E(_00729_),
    .Y(_00160_));
 XOR2x1_ASAP7_75t_R _30608_ (.A(net25),
    .Y(_00185_),
    .B(_01011_));
 XOR2x1_ASAP7_75t_R _30609_ (.A(net52),
    .Y(_00186_),
    .B(_08185_));
 XOR2x1_ASAP7_75t_R _30610_ (.A(_10711_),
    .Y(_00187_),
    .B(_01013_));
 XOR2x1_ASAP7_75t_R _30611_ (.A(_00735_),
    .Y(_00188_),
    .B(_01014_));
 XOR2x1_ASAP7_75t_R _30612_ (.A(_10756_),
    .Y(_00189_),
    .B(_01015_));
 XOR2x1_ASAP7_75t_R _30613_ (.A(_10783_),
    .Y(_00190_),
    .B(_01016_));
 XOR2x1_ASAP7_75t_R _30614_ (.A(_00738_),
    .Y(_00191_),
    .B(_01018_));
 XOR2x1_ASAP7_75t_R _30615_ (.A(net50),
    .Y(_00192_),
    .B(_01019_));
 XOR2x1_ASAP7_75t_R _30616_ (.A(net19),
    .Y(_00281_),
    .B(_01043_));
 XOR2x1_ASAP7_75t_R _30617_ (.A(_11404_),
    .Y(_00282_),
    .B(_08186_));
 XOR2x1_ASAP7_75t_R _30618_ (.A(_11433_),
    .Y(_00283_),
    .B(_01045_));
 XOR2x1_ASAP7_75t_R _30619_ (.A(_00743_),
    .Y(_00284_),
    .B(_01046_));
 XOR2x1_ASAP7_75t_R _30620_ (.A(_00744_),
    .Y(_00285_),
    .B(_08220_));
 XOR2x1_ASAP7_75t_R _30621_ (.A(_00745_),
    .Y(_00286_),
    .B(_01048_));
 XOR2x1_ASAP7_75t_R _30622_ (.A(_00746_),
    .Y(_00287_),
    .B(_01050_));
 XOR2x1_ASAP7_75t_R _30623_ (.A(_11363_),
    .Y(_00288_),
    .B(_01051_));
 XOR2x1_ASAP7_75t_R _30624_ (.A(net38),
    .Y(_00241_),
    .B(_08177_));
 XOR2x1_ASAP7_75t_R _30625_ (.A(net59),
    .Y(_00242_),
    .B(_08190_));
 XOR2x1_ASAP7_75t_R _30626_ (.A(_12169_),
    .Y(_00243_),
    .B(_08197_));
 XOR2x1_ASAP7_75t_R _30627_ (.A(_00751_),
    .Y(_00244_),
    .B(_08211_));
 XOR2x1_ASAP7_75t_R _30628_ (.A(_00752_),
    .Y(_00245_),
    .B(_01079_));
 XOR2x1_ASAP7_75t_R _30629_ (.A(_00753_),
    .Y(_00246_),
    .B(_01080_));
 XOR2x1_ASAP7_75t_R _30630_ (.A(_00754_),
    .Y(_00247_),
    .B(_01082_));
 XOR2x1_ASAP7_75t_R _30631_ (.A(_12085_),
    .Y(_00248_),
    .B(_01083_));
 XOR2x1_ASAP7_75t_R _30632_ (.A(net35),
    .Y(_00209_),
    .B(_01107_));
 XOR2x2_ASAP7_75t_R _30633_ (.A(_12870_),
    .B(_08191_),
    .Y(_00210_));
 XOR2x1_ASAP7_75t_R _30634_ (.A(_12910_),
    .Y(_00211_),
    .B(_08198_));
 XOR2x1_ASAP7_75t_R _30635_ (.A(_00759_),
    .Y(_00212_),
    .B(_01110_));
 XOR2x1_ASAP7_75t_R _30636_ (.A(_12952_),
    .Y(_00213_),
    .B(_01111_));
 XOR2x1_ASAP7_75t_R _30637_ (.A(_12902_),
    .Y(_00214_),
    .B(_01112_));
 XOR2x1_ASAP7_75t_R _30638_ (.A(_00762_),
    .Y(_00215_),
    .B(_01114_));
 XOR2x1_ASAP7_75t_R _30639_ (.A(net647),
    .Y(_00216_),
    .B(_01115_));
 XOR2x1_ASAP7_75t_R _30640_ (.A(net49),
    .Y(_00177_),
    .B(_07958_));
 XOR2x1_ASAP7_75t_R _30641_ (.A(_00765_),
    .Y(_00178_),
    .B(_07969_));
 XOR2x1_ASAP7_75t_R _30642_ (.A(_10674_),
    .Y(_00179_),
    .B(_08002_));
 XOR2x1_ASAP7_75t_R _30643_ (.A(_10710_),
    .Y(_00180_),
    .B(_07942_));
 XOR2x1_ASAP7_75t_R _30644_ (.A(_00768_),
    .Y(_00181_),
    .B(_01007_));
 XOR2x1_ASAP7_75t_R _30645_ (.A(_00769_),
    .Y(_00182_),
    .B(_01008_));
 XOR2x1_ASAP7_75t_R _30646_ (.A(_00770_),
    .Y(_00183_),
    .B(_01009_));
 XOR2x1_ASAP7_75t_R _30647_ (.A(_10825_),
    .Y(_00184_),
    .B(_01010_));
 XOR2x1_ASAP7_75t_R _30648_ (.A(net689),
    .Y(_00273_),
    .B(_07960_));
 XOR2x1_ASAP7_75t_R _30649_ (.A(_00773_),
    .Y(_00274_),
    .B(_07970_));
 XOR2x1_ASAP7_75t_R _30650_ (.A(_11402_),
    .Y(_00275_),
    .B(_08004_));
 XOR2x1_ASAP7_75t_R _30651_ (.A(_00775_),
    .Y(_00276_),
    .B(_01037_));
 XOR2x1_ASAP7_75t_R _30652_ (.A(_00776_),
    .Y(_00277_),
    .B(_01039_));
 XOR2x1_ASAP7_75t_R _30653_ (.A(_00777_),
    .Y(_00278_),
    .B(_01040_));
 XOR2x1_ASAP7_75t_R _30654_ (.A(_00778_),
    .Y(_00279_),
    .B(_01041_));
 XOR2x1_ASAP7_75t_R _30655_ (.A(_11383_),
    .Y(_00280_),
    .B(_01042_));
 XOR2x1_ASAP7_75t_R _30656_ (.A(net20),
    .Y(_00233_),
    .B(_07961_));
 XOR2x1_ASAP7_75t_R _30657_ (.A(_00781_),
    .Y(_00234_),
    .B(_07972_));
 XOR2x1_ASAP7_75t_R _30658_ (.A(_12125_),
    .Y(_00235_),
    .B(_08007_));
 XOR2x1_ASAP7_75t_R _30659_ (.A(_00783_),
    .Y(_00236_),
    .B(_01069_));
 XOR2x1_ASAP7_75t_R _30660_ (.A(_00784_),
    .Y(_00237_),
    .B(_07994_));
 XOR2x1_ASAP7_75t_R _30661_ (.A(_00785_),
    .Y(_00238_),
    .B(_07984_));
 XOR2x1_ASAP7_75t_R _30662_ (.A(_00786_),
    .Y(_00239_),
    .B(_01073_));
 XOR2x1_ASAP7_75t_R _30663_ (.A(_12108_),
    .Y(_00240_),
    .B(_01074_));
 XOR2x1_ASAP7_75t_R _30664_ (.A(_12834_),
    .Y(_00201_),
    .B(_01098_));
 XOR2x1_ASAP7_75t_R _30665_ (.A(net640),
    .Y(_00202_),
    .B(_07973_));
 XOR2x1_ASAP7_75t_R _30666_ (.A(_12868_),
    .Y(_00203_),
    .B(_08008_));
 XOR2x1_ASAP7_75t_R _30667_ (.A(_00791_),
    .Y(_00204_),
    .B(_07945_));
 XOR2x1_ASAP7_75t_R _30668_ (.A(_00792_),
    .Y(_00205_),
    .B(_07996_));
 XOR2x1_ASAP7_75t_R _30669_ (.A(_00793_),
    .Y(_00206_),
    .B(_01104_));
 XOR2x1_ASAP7_75t_R _30670_ (.A(_00794_),
    .Y(_00207_),
    .B(_01105_));
 XOR2x1_ASAP7_75t_R _30671_ (.A(net72),
    .Y(_00208_),
    .B(_01106_));
 XOR2x1_ASAP7_75t_R _30672_ (.A(_00796_),
    .Y(_00169_),
    .B(_01025_));
 XOR2x1_ASAP7_75t_R _30673_ (.A(_10628_),
    .Y(_00170_),
    .B(_08101_));
 XOR2x1_ASAP7_75t_R _30674_ (.A(_10681_),
    .Y(_00171_),
    .B(_08106_));
 XOR2x1_ASAP7_75t_R _30675_ (.A(_10714_),
    .Y(_00172_),
    .B(_00997_));
 XOR2x1_ASAP7_75t_R _30676_ (.A(_00800_),
    .Y(_00173_),
    .B(_00998_));
 XOR2x1_ASAP7_75t_R _30677_ (.A(_00801_),
    .Y(_00174_),
    .B(_00999_));
 XOR2x2_ASAP7_75t_R _30678_ (.A(_00802_),
    .B(_01000_),
    .Y(_00175_));
 XOR2x1_ASAP7_75t_R _30679_ (.A(net58),
    .Y(_00176_),
    .B(_01001_));
 XOR2x1_ASAP7_75t_R _30680_ (.A(_11388_),
    .Y(_00257_),
    .B(_01057_));
 XOR2x1_ASAP7_75t_R _30681_ (.A(_11365_),
    .Y(_00258_),
    .B(net930));
 XOR2x1_ASAP7_75t_R _30682_ (.A(_11409_),
    .Y(_00259_),
    .B(_08108_));
 XOR2x2_ASAP7_75t_R _30683_ (.A(_00807_),
    .B(_01029_),
    .Y(_00260_));
 XOR2x1_ASAP7_75t_R _30684_ (.A(_00808_),
    .Y(_00261_),
    .B(_01030_));
 XOR2x1_ASAP7_75t_R _30685_ (.A(_00809_),
    .Y(_00262_),
    .B(_01031_));
 XOR2x2_ASAP7_75t_R _30686_ (.A(_00810_),
    .B(_01032_),
    .Y(_00263_));
 XOR2x1_ASAP7_75t_R _30687_ (.A(net28),
    .Y(_00264_),
    .B(_01033_));
 XOR2x1_ASAP7_75t_R _30688_ (.A(net806),
    .Y(_00225_),
    .B(_01089_));
 XOR2x1_ASAP7_75t_R _30689_ (.A(_12087_),
    .Y(_00226_),
    .B(_08099_));
 XOR2x2_ASAP7_75t_R _30690_ (.A(_12132_),
    .B(_08110_),
    .Y(_00227_));
 XOR2x1_ASAP7_75t_R _30691_ (.A(_00815_),
    .Y(_00228_),
    .B(_01061_));
 XOR2x1_ASAP7_75t_R _30692_ (.A(_00816_),
    .Y(_00229_),
    .B(_01062_));
 XOR2x1_ASAP7_75t_R _30693_ (.A(_00817_),
    .Y(_00230_),
    .B(_01063_));
 XOR2x1_ASAP7_75t_R _30694_ (.A(_00818_),
    .Y(_00231_),
    .B(_01064_));
 XOR2x1_ASAP7_75t_R _30695_ (.A(net40),
    .Y(_00232_),
    .B(_01065_));
 XOR2x1_ASAP7_75t_R _30696_ (.A(net910),
    .Y(_00193_),
    .B(_01121_));
 XOR2x1_ASAP7_75t_R _30697_ (.A(_00642_),
    .Y(_00194_),
    .B(_12831_));
 XOR2x1_ASAP7_75t_R _30698_ (.A(_12879_),
    .Y(_00195_),
    .B(_08111_));
 XOR2x1_ASAP7_75t_R _30699_ (.A(_12913_),
    .Y(_00196_),
    .B(_08124_));
 XOR2x1_ASAP7_75t_R _30700_ (.A(_00824_),
    .Y(_00197_),
    .B(_08133_));
 XOR2x2_ASAP7_75t_R _30701_ (.A(_00825_),
    .B(_01095_),
    .Y(_00198_));
 XOR2x2_ASAP7_75t_R _30702_ (.A(_00826_),
    .B(_01096_),
    .Y(_00199_));
 XOR2x1_ASAP7_75t_R _30703_ (.A(net908),
    .Y(_00200_),
    .B(_01097_));
 XOR2x1_ASAP7_75t_R _30704_ (.A(_10651_),
    .Y(_00161_),
    .B(net617));
 XOR2x1_ASAP7_75t_R _30705_ (.A(_10624_),
    .Y(_00162_),
    .B(_08023_));
 XOR2x1_ASAP7_75t_R _30706_ (.A(_10682_),
    .Y(_00163_),
    .B(_08031_));
 XOR2x1_ASAP7_75t_R _30707_ (.A(_10715_),
    .Y(_00164_),
    .B(_01020_));
 XOR2x1_ASAP7_75t_R _30708_ (.A(_00832_),
    .Y(_00165_),
    .B(_01021_));
 XOR2x1_ASAP7_75t_R _30709_ (.A(_10758_),
    .Y(_00166_),
    .B(_01022_));
 XOR2x1_ASAP7_75t_R _30710_ (.A(_00834_),
    .Y(_00167_),
    .B(_01023_));
 XOR2x1_ASAP7_75t_R _30711_ (.A(_10822_),
    .Y(_00168_),
    .B(_01024_));
 XOR2x1_ASAP7_75t_R _30712_ (.A(_11381_),
    .Y(_00249_),
    .B(net859));
 XOR2x2_ASAP7_75t_R _30713_ (.A(_11360_),
    .B(_08024_),
    .Y(_00250_));
 XOR2x1_ASAP7_75t_R _30714_ (.A(_11410_),
    .Y(_00251_),
    .B(_08033_));
 XOR2x1_ASAP7_75t_R _30715_ (.A(_00839_),
    .Y(_00252_),
    .B(_01052_));
 XOR2x1_ASAP7_75t_R _30716_ (.A(_00840_),
    .Y(_00253_),
    .B(_01053_));
 XOR2x1_ASAP7_75t_R _30717_ (.A(_00841_),
    .Y(_00254_),
    .B(_01054_));
 XOR2x1_ASAP7_75t_R _30718_ (.A(_00842_),
    .Y(_00255_),
    .B(_01055_));
 XOR2x1_ASAP7_75t_R _30719_ (.A(_11536_),
    .Y(_00256_),
    .B(_01056_));
 XOR2x1_ASAP7_75t_R _30720_ (.A(_12104_),
    .Y(_00217_),
    .B(net856));
 XOR2x1_ASAP7_75t_R _30721_ (.A(net844),
    .Y(_00218_),
    .B(_08026_));
 XOR2x1_ASAP7_75t_R _30722_ (.A(_12133_),
    .Y(_00219_),
    .B(_08035_));
 XOR2x1_ASAP7_75t_R _30723_ (.A(_00847_),
    .Y(_00220_),
    .B(_08047_));
 XOR2x1_ASAP7_75t_R _30724_ (.A(_00848_),
    .Y(_00221_),
    .B(_01085_));
 XOR2x1_ASAP7_75t_R _30725_ (.A(_12259_),
    .Y(_00222_),
    .B(_01086_));
 XOR2x1_ASAP7_75t_R _30726_ (.A(_00850_),
    .Y(_00223_),
    .B(_01087_));
 XOR2x1_ASAP7_75t_R _30727_ (.A(_12275_),
    .Y(_00224_),
    .B(_01088_));
 XOR2x1_ASAP7_75t_R _30728_ (.A(net665),
    .Y(_00265_),
    .B(_01091_));
 XOR2x1_ASAP7_75t_R _30729_ (.A(_12836_),
    .Y(_00266_),
    .B(_01102_));
 XOR2x2_ASAP7_75t_R _30730_ (.A(_12880_),
    .B(_01113_),
    .Y(_00267_));
 XOR2x1_ASAP7_75t_R _30731_ (.A(_00855_),
    .Y(_00268_),
    .B(_01116_));
 XOR2x1_ASAP7_75t_R _30732_ (.A(_00856_),
    .Y(_00269_),
    .B(_01117_));
 XOR2x1_ASAP7_75t_R _30733_ (.A(_12955_),
    .Y(_00270_),
    .B(_01118_));
 XOR2x1_ASAP7_75t_R _30734_ (.A(_00858_),
    .Y(_00271_),
    .B(_01119_));
 XOR2x1_ASAP7_75t_R _30735_ (.A(_13013_),
    .Y(_00272_),
    .B(_01120_));
 INVx2_ASAP7_75t_R _30736_ (.A(_00644_),
    .Y(net453));
 INVx1_ASAP7_75t_R _30737_ (.A(_00730_),
    .Y(net325));
 INVx2_ASAP7_75t_R _30738_ (.A(_00859_),
    .Y(net326));
 INVx2_ASAP7_75t_R _30739_ (.A(_00860_),
    .Y(net327));
 INVx3_ASAP7_75t_R _30740_ (.A(_00861_),
    .Y(net328));
 INVx2_ASAP7_75t_R _30741_ (.A(_00862_),
    .Y(net329));
 INVx3_ASAP7_75t_R _30742_ (.A(_00863_),
    .Y(net330));
 INVx2_ASAP7_75t_R _30743_ (.A(_00864_),
    .Y(net331));
 INVx1_ASAP7_75t_R _30744_ (.A(_00865_),
    .Y(net332));
 INVx2_ASAP7_75t_R _30745_ (.A(_00866_),
    .Y(net333));
 INVx2_ASAP7_75t_R _30746_ (.A(_00867_),
    .Y(net334));
 INVx2_ASAP7_75t_R _30747_ (.A(_00868_),
    .Y(net335));
 INVx1_ASAP7_75t_R _30748_ (.A(_00869_),
    .Y(net336));
 INVx2_ASAP7_75t_R _30749_ (.A(_00870_),
    .Y(net337));
 INVx1_ASAP7_75t_R _30750_ (.A(_00871_),
    .Y(net338));
 INVx1_ASAP7_75t_R _30751_ (.A(_00872_),
    .Y(net339));
 INVx1_ASAP7_75t_R _30752_ (.A(_00873_),
    .Y(net340));
 INVx1_ASAP7_75t_R _30753_ (.A(_00874_),
    .Y(net341));
 INVx1_ASAP7_75t_R _30754_ (.A(_00875_),
    .Y(net342));
 INVx1_ASAP7_75t_R _30755_ (.A(_00876_),
    .Y(net343));
 INVx1_ASAP7_75t_R _30756_ (.A(_00877_),
    .Y(net344));
 INVx1_ASAP7_75t_R _30757_ (.A(_00878_),
    .Y(net345));
 INVx1_ASAP7_75t_R _30758_ (.A(_00879_),
    .Y(net346));
 INVx1_ASAP7_75t_R _30759_ (.A(_00880_),
    .Y(net347));
 INVx2_ASAP7_75t_R _30760_ (.A(_00881_),
    .Y(net348));
 INVx1_ASAP7_75t_R _30761_ (.A(_00882_),
    .Y(net349));
 INVx1_ASAP7_75t_R _30762_ (.A(_00883_),
    .Y(net350));
 INVx1_ASAP7_75t_R _30763_ (.A(_00884_),
    .Y(net351));
 INVx1_ASAP7_75t_R _30764_ (.A(_00885_),
    .Y(net352));
 INVx1_ASAP7_75t_R _30765_ (.A(_00886_),
    .Y(net353));
 INVx2_ASAP7_75t_R _30766_ (.A(_00887_),
    .Y(net354));
 INVx2_ASAP7_75t_R _30767_ (.A(_00888_),
    .Y(net355));
 INVx2_ASAP7_75t_R _30768_ (.A(_00889_),
    .Y(net356));
 INVx2_ASAP7_75t_R _30769_ (.A(_00890_),
    .Y(net357));
 INVx1_ASAP7_75t_R _30770_ (.A(_00891_),
    .Y(net358));
 INVx1_ASAP7_75t_R _30771_ (.A(_00892_),
    .Y(net359));
 INVx2_ASAP7_75t_R _30772_ (.A(_00893_),
    .Y(net360));
 INVx2_ASAP7_75t_R _30773_ (.A(_00894_),
    .Y(net361));
 INVx1_ASAP7_75t_R _30774_ (.A(_00895_),
    .Y(net362));
 INVx1_ASAP7_75t_R _30775_ (.A(_00896_),
    .Y(net363));
 INVx1_ASAP7_75t_R _30776_ (.A(_00897_),
    .Y(net364));
 INVx2_ASAP7_75t_R _30777_ (.A(_00898_),
    .Y(net365));
 INVx1_ASAP7_75t_R _30778_ (.A(_00899_),
    .Y(net366));
 INVx2_ASAP7_75t_R _30779_ (.A(_00900_),
    .Y(net367));
 INVx2_ASAP7_75t_R _30780_ (.A(_00901_),
    .Y(net368));
 INVx1_ASAP7_75t_R _30781_ (.A(_00902_),
    .Y(net369));
 INVx2_ASAP7_75t_R _30782_ (.A(_00903_),
    .Y(net370));
 INVx1_ASAP7_75t_R _30783_ (.A(_00904_),
    .Y(net371));
 INVx2_ASAP7_75t_R _30784_ (.A(_00905_),
    .Y(net372));
 INVx2_ASAP7_75t_R _30785_ (.A(_00906_),
    .Y(net373));
 INVx2_ASAP7_75t_R _30786_ (.A(_00907_),
    .Y(net374));
 INVx1_ASAP7_75t_R _30787_ (.A(_00908_),
    .Y(net375));
 INVx1_ASAP7_75t_R _30788_ (.A(_00909_),
    .Y(net376));
 INVx1_ASAP7_75t_R _30789_ (.A(_00910_),
    .Y(net377));
 INVx2_ASAP7_75t_R _30790_ (.A(_00911_),
    .Y(net378));
 INVx1_ASAP7_75t_R _30791_ (.A(_00912_),
    .Y(net379));
 INVx1_ASAP7_75t_R _30792_ (.A(_00913_),
    .Y(net380));
 INVx1_ASAP7_75t_R _30793_ (.A(_00914_),
    .Y(net381));
 INVx1_ASAP7_75t_R _30794_ (.A(_00915_),
    .Y(net382));
 INVx1_ASAP7_75t_R _30795_ (.A(_00916_),
    .Y(net383));
 INVx1_ASAP7_75t_R _30796_ (.A(_00917_),
    .Y(net384));
 INVx1_ASAP7_75t_R _30797_ (.A(_00918_),
    .Y(net385));
 INVx1_ASAP7_75t_R _30798_ (.A(_00919_),
    .Y(net386));
 INVx2_ASAP7_75t_R _30799_ (.A(_00920_),
    .Y(net387));
 INVx2_ASAP7_75t_R _30800_ (.A(_00921_),
    .Y(net388));
 INVx2_ASAP7_75t_R _30801_ (.A(_00922_),
    .Y(net389));
 INVx1_ASAP7_75t_R _30802_ (.A(_00923_),
    .Y(net390));
 INVx2_ASAP7_75t_R _30803_ (.A(_00924_),
    .Y(net391));
 INVx2_ASAP7_75t_R _30804_ (.A(_00925_),
    .Y(net392));
 INVx2_ASAP7_75t_R _30805_ (.A(_00926_),
    .Y(net393));
 INVx2_ASAP7_75t_R _30806_ (.A(_00927_),
    .Y(net394));
 INVx2_ASAP7_75t_R _30807_ (.A(_00928_),
    .Y(net395));
 INVx2_ASAP7_75t_R _30808_ (.A(_00929_),
    .Y(net396));
 INVx2_ASAP7_75t_R _30809_ (.A(_00930_),
    .Y(net397));
 INVx2_ASAP7_75t_R _30810_ (.A(_00931_),
    .Y(net398));
 INVx2_ASAP7_75t_R _30811_ (.A(_00932_),
    .Y(net399));
 INVx1_ASAP7_75t_R _30812_ (.A(_00933_),
    .Y(net400));
 INVx2_ASAP7_75t_R _30813_ (.A(_00934_),
    .Y(net401));
 INVx1_ASAP7_75t_R _30814_ (.A(_00935_),
    .Y(net402));
 INVx1_ASAP7_75t_R _30815_ (.A(_00936_),
    .Y(net403));
 INVx2_ASAP7_75t_R _30816_ (.A(_00937_),
    .Y(net404));
 INVx2_ASAP7_75t_R _30817_ (.A(_00938_),
    .Y(net405));
 INVx1_ASAP7_75t_R _30818_ (.A(_00939_),
    .Y(net406));
 INVx1_ASAP7_75t_R _30819_ (.A(_00940_),
    .Y(net407));
 INVx1_ASAP7_75t_R _30820_ (.A(_00941_),
    .Y(net408));
 INVx1_ASAP7_75t_R _30821_ (.A(_00942_),
    .Y(net409));
 INVx1_ASAP7_75t_R _30822_ (.A(_00943_),
    .Y(net410));
 INVx1_ASAP7_75t_R _30823_ (.A(_00944_),
    .Y(net411));
 INVx1_ASAP7_75t_R _30824_ (.A(_00945_),
    .Y(net412));
 INVx2_ASAP7_75t_R _30825_ (.A(_00946_),
    .Y(net413));
 INVx2_ASAP7_75t_R _30826_ (.A(_00947_),
    .Y(net414));
 INVx1_ASAP7_75t_R _30827_ (.A(_00948_),
    .Y(net415));
 INVx2_ASAP7_75t_R _30828_ (.A(_00949_),
    .Y(net416));
 INVx2_ASAP7_75t_R _30829_ (.A(_00950_),
    .Y(net417));
 INVx1_ASAP7_75t_R _30830_ (.A(_00951_),
    .Y(net418));
 INVx2_ASAP7_75t_R _30831_ (.A(_00952_),
    .Y(net419));
 INVx2_ASAP7_75t_R _30832_ (.A(_00953_),
    .Y(net420));
 INVx1_ASAP7_75t_R _30833_ (.A(_00954_),
    .Y(net421));
 INVx1_ASAP7_75t_R _30834_ (.A(_00955_),
    .Y(net422));
 INVx2_ASAP7_75t_R _30835_ (.A(_00956_),
    .Y(net423));
 INVx2_ASAP7_75t_R _30836_ (.A(_00957_),
    .Y(net424));
 INVx2_ASAP7_75t_R _30837_ (.A(_00958_),
    .Y(net425));
 INVx1_ASAP7_75t_R _30838_ (.A(_00959_),
    .Y(net426));
 INVx2_ASAP7_75t_R _30839_ (.A(_00960_),
    .Y(net427));
 INVx2_ASAP7_75t_R _30840_ (.A(_00961_),
    .Y(net428));
 INVx1_ASAP7_75t_R _30841_ (.A(_00962_),
    .Y(net429));
 INVx2_ASAP7_75t_R _30842_ (.A(_00963_),
    .Y(net430));
 INVx2_ASAP7_75t_R _30843_ (.A(_00964_),
    .Y(net431));
 INVx2_ASAP7_75t_R _30844_ (.A(_00965_),
    .Y(net432));
 INVx2_ASAP7_75t_R _30845_ (.A(_00966_),
    .Y(net433));
 INVx2_ASAP7_75t_R _30846_ (.A(_00967_),
    .Y(net434));
 INVx1_ASAP7_75t_R _30847_ (.A(_00968_),
    .Y(net435));
 INVx1_ASAP7_75t_R _30848_ (.A(_00969_),
    .Y(net436));
 INVx2_ASAP7_75t_R _30849_ (.A(_00970_),
    .Y(net437));
 INVx2_ASAP7_75t_R _30850_ (.A(_00971_),
    .Y(net438));
 INVx2_ASAP7_75t_R _30851_ (.A(_00972_),
    .Y(net439));
 INVx2_ASAP7_75t_R _30852_ (.A(_00973_),
    .Y(net440));
 INVx2_ASAP7_75t_R _30853_ (.A(_00974_),
    .Y(net441));
 INVx2_ASAP7_75t_R _30854_ (.A(_00975_),
    .Y(net442));
 INVx2_ASAP7_75t_R _30855_ (.A(_00976_),
    .Y(net443));
 INVx1_ASAP7_75t_R _30856_ (.A(_00977_),
    .Y(net444));
 INVx2_ASAP7_75t_R _30857_ (.A(_00978_),
    .Y(net445));
 INVx2_ASAP7_75t_R _30858_ (.A(_00979_),
    .Y(net446));
 INVx1_ASAP7_75t_R _30859_ (.A(_00980_),
    .Y(net447));
 INVx2_ASAP7_75t_R _30860_ (.A(_00981_),
    .Y(net448));
 INVx2_ASAP7_75t_R _30861_ (.A(_00982_),
    .Y(net449));
 INVx2_ASAP7_75t_R _30862_ (.A(_00983_),
    .Y(net450));
 INVx1_ASAP7_75t_R _30863_ (.A(_00984_),
    .Y(net451));
 INVx2_ASAP7_75t_R _30864_ (.A(_00985_),
    .Y(net452));
 NOR2x1_ASAP7_75t_R _30865_ (.A(_08409_),
    .B(_00411_),
    .Y(_07760_));
 AO21x1_ASAP7_75t_R _30866_ (.A1(_08398_),
    .A2(net197),
    .B(_07760_),
    .Y(_01287_));
 NOR2x1_ASAP7_75t_R _30867_ (.A(_08409_),
    .B(_00724_),
    .Y(_07761_));
 AO21x1_ASAP7_75t_R _30868_ (.A1(_08398_),
    .A2(net198),
    .B(_07761_),
    .Y(_01288_));
 BUFx6f_ASAP7_75t_R _30869_ (.A(_08379_),
    .Y(_07762_));
 NOR2x1_ASAP7_75t_R _30870_ (.A(_08409_),
    .B(_00723_),
    .Y(_07763_));
 AO21x1_ASAP7_75t_R _30871_ (.A1(_07762_),
    .A2(net199),
    .B(_07763_),
    .Y(_01289_));
 NOR2x1_ASAP7_75t_R _30872_ (.A(_08409_),
    .B(_00722_),
    .Y(_07764_));
 AO21x1_ASAP7_75t_R _30873_ (.A1(_07762_),
    .A2(net200),
    .B(_07764_),
    .Y(_01290_));
 NOR2x1_ASAP7_75t_R _30874_ (.A(_08409_),
    .B(_00721_),
    .Y(_07765_));
 AO21x1_ASAP7_75t_R _30875_ (.A1(_07762_),
    .A2(net201),
    .B(_07765_),
    .Y(_01291_));
 NOR2x1_ASAP7_75t_R _30876_ (.A(_08409_),
    .B(_00570_),
    .Y(_07766_));
 AO21x1_ASAP7_75t_R _30877_ (.A1(_07762_),
    .A2(net202),
    .B(_07766_),
    .Y(_01292_));
 BUFx12f_ASAP7_75t_R _30878_ (.A(_07967_),
    .Y(_07767_));
 BUFx10_ASAP7_75t_R _30879_ (.A(_07767_),
    .Y(_07768_));
 NOR2x1_ASAP7_75t_R _30880_ (.A(_07768_),
    .B(_00569_),
    .Y(_07769_));
 AO21x1_ASAP7_75t_R _30881_ (.A1(_07762_),
    .A2(net203),
    .B(_07769_),
    .Y(_01293_));
 NOR2x1_ASAP7_75t_R _30882_ (.A(_07768_),
    .B(_00572_),
    .Y(_07770_));
 AO21x1_ASAP7_75t_R _30883_ (.A1(_07762_),
    .A2(net204),
    .B(_07770_),
    .Y(_01294_));
 NOR2x1_ASAP7_75t_R _30884_ (.A(_07768_),
    .B(_00720_),
    .Y(_07771_));
 AO21x1_ASAP7_75t_R _30885_ (.A1(_07762_),
    .A2(net205),
    .B(_07771_),
    .Y(_01295_));
 NOR2x1_ASAP7_75t_R _30886_ (.A(_07768_),
    .B(_00719_),
    .Y(_07772_));
 AO21x1_ASAP7_75t_R _30887_ (.A1(_07762_),
    .A2(net206),
    .B(_07772_),
    .Y(_01296_));
 NOR2x1_ASAP7_75t_R _30888_ (.A(_07768_),
    .B(_00718_),
    .Y(_07773_));
 AO21x1_ASAP7_75t_R _30889_ (.A1(_07762_),
    .A2(net207),
    .B(_07773_),
    .Y(_01297_));
 NOR2x1_ASAP7_75t_R _30890_ (.A(_07768_),
    .B(_00608_),
    .Y(_07774_));
 AO21x1_ASAP7_75t_R _30891_ (.A1(_07762_),
    .A2(net208),
    .B(_07774_),
    .Y(_01298_));
 BUFx6f_ASAP7_75t_R _30892_ (.A(_08379_),
    .Y(_07775_));
 NOR2x1_ASAP7_75t_R _30893_ (.A(_07768_),
    .B(_00717_),
    .Y(_07776_));
 AO21x1_ASAP7_75t_R _30894_ (.A1(_07775_),
    .A2(net209),
    .B(_07776_),
    .Y(_01299_));
 NOR2x1_ASAP7_75t_R _30895_ (.A(_07768_),
    .B(_00716_),
    .Y(_07777_));
 AO21x1_ASAP7_75t_R _30896_ (.A1(_07775_),
    .A2(net210),
    .B(_07777_),
    .Y(_01300_));
 NOR2x1_ASAP7_75t_R _30897_ (.A(_07768_),
    .B(_00530_),
    .Y(_07778_));
 AO21x1_ASAP7_75t_R _30898_ (.A1(_07775_),
    .A2(net211),
    .B(_07778_),
    .Y(_01301_));
 NOR2x1_ASAP7_75t_R _30899_ (.A(_07768_),
    .B(_00529_),
    .Y(_07779_));
 AO21x1_ASAP7_75t_R _30900_ (.A1(_07775_),
    .A2(net212),
    .B(_07779_),
    .Y(_01302_));
 BUFx10_ASAP7_75t_R _30901_ (.A(_07767_),
    .Y(_07780_));
 NOR2x1_ASAP7_75t_R _30902_ (.A(_07780_),
    .B(_00532_),
    .Y(_07781_));
 AO21x1_ASAP7_75t_R _30903_ (.A1(_07775_),
    .A2(net213),
    .B(_07781_),
    .Y(_01303_));
 NOR2x1_ASAP7_75t_R _30904_ (.A(_07780_),
    .B(_00715_),
    .Y(_07782_));
 AO21x1_ASAP7_75t_R _30905_ (.A1(_07775_),
    .A2(net214),
    .B(_07782_),
    .Y(_01304_));
 NOR2x1_ASAP7_75t_R _30906_ (.A(_07780_),
    .B(_00714_),
    .Y(_07783_));
 AO21x1_ASAP7_75t_R _30907_ (.A1(_07775_),
    .A2(net215),
    .B(_07783_),
    .Y(_01305_));
 NOR2x1_ASAP7_75t_R _30908_ (.A(_07780_),
    .B(_00713_),
    .Y(_07784_));
 AO21x1_ASAP7_75t_R _30909_ (.A1(_07775_),
    .A2(net216),
    .B(_07784_),
    .Y(_01306_));
 NOR2x1_ASAP7_75t_R _30910_ (.A(_07780_),
    .B(_00712_),
    .Y(_07785_));
 AO21x1_ASAP7_75t_R _30911_ (.A1(_07775_),
    .A2(net217),
    .B(_07785_),
    .Y(_01307_));
 NOR2x1_ASAP7_75t_R _30912_ (.A(_07780_),
    .B(_00711_),
    .Y(_07786_));
 AO21x1_ASAP7_75t_R _30913_ (.A1(_07775_),
    .A2(net218),
    .B(_07786_),
    .Y(_01308_));
 BUFx6f_ASAP7_75t_R _30914_ (.A(_08379_),
    .Y(_07787_));
 NOR2x1_ASAP7_75t_R _30915_ (.A(_07780_),
    .B(_00710_),
    .Y(_07788_));
 AO21x1_ASAP7_75t_R _30916_ (.A1(_07787_),
    .A2(net219),
    .B(_07788_),
    .Y(_01309_));
 NOR2x1_ASAP7_75t_R _30917_ (.A(_07780_),
    .B(_00490_),
    .Y(_07789_));
 AO21x1_ASAP7_75t_R _30918_ (.A1(_07787_),
    .A2(net220),
    .B(_07789_),
    .Y(_01310_));
 NOR2x1_ASAP7_75t_R _30919_ (.A(_07780_),
    .B(_00489_),
    .Y(_07790_));
 AO21x1_ASAP7_75t_R _30920_ (.A1(_07787_),
    .A2(net221),
    .B(_07790_),
    .Y(_01311_));
 NOR2x1_ASAP7_75t_R _30921_ (.A(_07780_),
    .B(_00492_),
    .Y(_07791_));
 AO21x1_ASAP7_75t_R _30922_ (.A1(_07787_),
    .A2(net222),
    .B(_07791_),
    .Y(_01312_));
 BUFx10_ASAP7_75t_R _30923_ (.A(_07767_),
    .Y(_07792_));
 NOR2x1_ASAP7_75t_R _30924_ (.A(_07792_),
    .B(_00709_),
    .Y(_07793_));
 AO21x1_ASAP7_75t_R _30925_ (.A1(_07787_),
    .A2(net223),
    .B(_07793_),
    .Y(_01313_));
 NOR2x1_ASAP7_75t_R _30926_ (.A(_07792_),
    .B(_00708_),
    .Y(_07794_));
 AO21x1_ASAP7_75t_R _30927_ (.A1(_07787_),
    .A2(net224),
    .B(_07794_),
    .Y(_01314_));
 NOR2x1_ASAP7_75t_R _30928_ (.A(_07792_),
    .B(_00707_),
    .Y(_07795_));
 AO21x1_ASAP7_75t_R _30929_ (.A1(_07787_),
    .A2(net225),
    .B(_07795_),
    .Y(_01315_));
 NOR2x1_ASAP7_75t_R _30930_ (.A(_07792_),
    .B(_00706_),
    .Y(_07796_));
 AO21x1_ASAP7_75t_R _30931_ (.A1(_07787_),
    .A2(net226),
    .B(_07796_),
    .Y(_01316_));
 NOR2x1_ASAP7_75t_R _30932_ (.A(_07792_),
    .B(_00705_),
    .Y(_07797_));
 AO21x1_ASAP7_75t_R _30933_ (.A1(_07787_),
    .A2(net227),
    .B(_07797_),
    .Y(_01317_));
 NOR2x1_ASAP7_75t_R _30934_ (.A(_07792_),
    .B(_00704_),
    .Y(_07798_));
 AO21x1_ASAP7_75t_R _30935_ (.A1(_07787_),
    .A2(net228),
    .B(_07798_),
    .Y(_01318_));
 BUFx6f_ASAP7_75t_R _30936_ (.A(_08379_),
    .Y(_07799_));
 NOR2x1_ASAP7_75t_R _30937_ (.A(_07792_),
    .B(_00703_),
    .Y(_07800_));
 AO21x1_ASAP7_75t_R _30938_ (.A1(_07799_),
    .A2(net229),
    .B(_07800_),
    .Y(_01319_));
 NOR2x1_ASAP7_75t_R _30939_ (.A(_07792_),
    .B(_00702_),
    .Y(_07801_));
 AO21x1_ASAP7_75t_R _30940_ (.A1(_07799_),
    .A2(net230),
    .B(_07801_),
    .Y(_01320_));
 NOR2x1_ASAP7_75t_R _30941_ (.A(_07792_),
    .B(_00701_),
    .Y(_07802_));
 AO21x1_ASAP7_75t_R _30942_ (.A1(_07799_),
    .A2(net231),
    .B(_07802_),
    .Y(_01321_));
 NOR2x1_ASAP7_75t_R _30943_ (.A(_07792_),
    .B(_00560_),
    .Y(_07803_));
 AO21x1_ASAP7_75t_R _30944_ (.A1(_07799_),
    .A2(net232),
    .B(_07803_),
    .Y(_01322_));
 BUFx6f_ASAP7_75t_R _30945_ (.A(_07767_),
    .Y(_07804_));
 NOR2x1_ASAP7_75t_R _30946_ (.A(_07804_),
    .B(_00559_),
    .Y(_07805_));
 AO21x1_ASAP7_75t_R _30947_ (.A1(_07799_),
    .A2(net233),
    .B(_07805_),
    .Y(_01323_));
 NOR2x1_ASAP7_75t_R _30948_ (.A(_07804_),
    .B(_00562_),
    .Y(_07806_));
 AO21x1_ASAP7_75t_R _30949_ (.A1(_07799_),
    .A2(net234),
    .B(_07806_),
    .Y(_01324_));
 NOR2x1_ASAP7_75t_R _30950_ (.A(_07804_),
    .B(_00700_),
    .Y(_07807_));
 AO21x1_ASAP7_75t_R _30951_ (.A1(_07799_),
    .A2(net235),
    .B(_07807_),
    .Y(_01325_));
 NOR2x1_ASAP7_75t_R _30952_ (.A(_07804_),
    .B(_00410_),
    .Y(_07808_));
 AO21x1_ASAP7_75t_R _30953_ (.A1(_07799_),
    .A2(net236),
    .B(_07808_),
    .Y(_01326_));
 NOR2x1_ASAP7_75t_R _30954_ (.A(_07804_),
    .B(_00699_),
    .Y(_07809_));
 AO21x1_ASAP7_75t_R _30955_ (.A1(_07799_),
    .A2(net237),
    .B(_07809_),
    .Y(_01327_));
 NOR2x1_ASAP7_75t_R _30956_ (.A(_07804_),
    .B(_00698_),
    .Y(_07810_));
 AO21x1_ASAP7_75t_R _30957_ (.A1(_07799_),
    .A2(net238),
    .B(_07810_),
    .Y(_01328_));
 BUFx6f_ASAP7_75t_R _30958_ (.A(_08379_),
    .Y(_07811_));
 NOR2x1_ASAP7_75t_R _30959_ (.A(_07804_),
    .B(_00697_),
    .Y(_07812_));
 AO21x1_ASAP7_75t_R _30960_ (.A1(_07811_),
    .A2(net239),
    .B(_07812_),
    .Y(_01329_));
 NOR2x1_ASAP7_75t_R _30961_ (.A(_07804_),
    .B(_00696_),
    .Y(_07813_));
 AO21x1_ASAP7_75t_R _30962_ (.A1(_07811_),
    .A2(net240),
    .B(_07813_),
    .Y(_01330_));
 NOR2x1_ASAP7_75t_R _30963_ (.A(_07804_),
    .B(_00520_),
    .Y(_07814_));
 AO21x1_ASAP7_75t_R _30964_ (.A1(_07811_),
    .A2(net241),
    .B(_07814_),
    .Y(_01331_));
 NOR2x1_ASAP7_75t_R _30965_ (.A(_07804_),
    .B(_00519_),
    .Y(_07815_));
 AO21x1_ASAP7_75t_R _30966_ (.A1(_07811_),
    .A2(net242),
    .B(_07815_),
    .Y(_01332_));
 BUFx6f_ASAP7_75t_R _30967_ (.A(_07767_),
    .Y(_07816_));
 NOR2x1_ASAP7_75t_R _30968_ (.A(_07816_),
    .B(_00522_),
    .Y(_07817_));
 AO21x1_ASAP7_75t_R _30969_ (.A1(_07811_),
    .A2(net243),
    .B(_07817_),
    .Y(_01333_));
 NOR2x1_ASAP7_75t_R _30970_ (.A(_07816_),
    .B(_00695_),
    .Y(_07818_));
 AO21x1_ASAP7_75t_R _30971_ (.A1(_07811_),
    .A2(net244),
    .B(_07818_),
    .Y(_01334_));
 NOR2x1_ASAP7_75t_R _30972_ (.A(_07816_),
    .B(_00694_),
    .Y(_07819_));
 AO21x1_ASAP7_75t_R _30973_ (.A1(_07811_),
    .A2(net245),
    .B(_07819_),
    .Y(_01335_));
 NOR2x1_ASAP7_75t_R _30974_ (.A(_07816_),
    .B(_00693_),
    .Y(_07820_));
 AO21x1_ASAP7_75t_R _30975_ (.A1(_07811_),
    .A2(net246),
    .B(_07820_),
    .Y(_01336_));
 NOR2x1_ASAP7_75t_R _30976_ (.A(_07816_),
    .B(_00413_),
    .Y(_07821_));
 AO21x1_ASAP7_75t_R _30977_ (.A1(_07811_),
    .A2(net247),
    .B(_07821_),
    .Y(_01337_));
 NOR2x1_ASAP7_75t_R _30978_ (.A(_07816_),
    .B(_00692_),
    .Y(_07822_));
 AO21x1_ASAP7_75t_R _30979_ (.A1(_07811_),
    .A2(net248),
    .B(_07822_),
    .Y(_01338_));
 BUFx4f_ASAP7_75t_R _30980_ (.A(_08379_),
    .Y(_07823_));
 NOR2x1_ASAP7_75t_R _30981_ (.A(_07816_),
    .B(_00691_),
    .Y(_07824_));
 AO21x1_ASAP7_75t_R _30982_ (.A1(_07823_),
    .A2(net249),
    .B(_07824_),
    .Y(_01339_));
 NOR2x1_ASAP7_75t_R _30983_ (.A(_07816_),
    .B(_00638_),
    .Y(_07825_));
 AO21x1_ASAP7_75t_R _30984_ (.A1(_07823_),
    .A2(net250),
    .B(_07825_),
    .Y(_01340_));
 NOR2x1_ASAP7_75t_R _30985_ (.A(_07816_),
    .B(_00637_),
    .Y(_07826_));
 AO21x1_ASAP7_75t_R _30986_ (.A1(_07823_),
    .A2(net251),
    .B(_07826_),
    .Y(_01341_));
 NOR2x1_ASAP7_75t_R _30987_ (.A(_07816_),
    .B(_00639_),
    .Y(_07827_));
 AO21x1_ASAP7_75t_R _30988_ (.A1(_07823_),
    .A2(net252),
    .B(_07827_),
    .Y(_01342_));
 BUFx6f_ASAP7_75t_R _30989_ (.A(_07767_),
    .Y(_07828_));
 NOR2x1_ASAP7_75t_R _30990_ (.A(_07828_),
    .B(_00690_),
    .Y(_07829_));
 AO21x1_ASAP7_75t_R _30991_ (.A1(_07823_),
    .A2(net253),
    .B(_07829_),
    .Y(_01343_));
 NOR2x1_ASAP7_75t_R _30992_ (.A(_07828_),
    .B(_00689_),
    .Y(_07830_));
 AO21x1_ASAP7_75t_R _30993_ (.A1(_07823_),
    .A2(net254),
    .B(_07830_),
    .Y(_01344_));
 NOR2x1_ASAP7_75t_R _30994_ (.A(_07828_),
    .B(_00688_),
    .Y(_07831_));
 AO21x1_ASAP7_75t_R _30995_ (.A1(_07823_),
    .A2(net255),
    .B(_07831_),
    .Y(_01345_));
 NOR2x1_ASAP7_75t_R _30996_ (.A(_07828_),
    .B(_00687_),
    .Y(_07832_));
 AO21x1_ASAP7_75t_R _30997_ (.A1(_07823_),
    .A2(net256),
    .B(_07832_),
    .Y(_01346_));
 NOR2x1_ASAP7_75t_R _30998_ (.A(_07828_),
    .B(_00686_),
    .Y(_07833_));
 AO21x1_ASAP7_75t_R _30999_ (.A1(_07823_),
    .A2(net257),
    .B(_07833_),
    .Y(_01347_));
 NOR2x1_ASAP7_75t_R _31000_ (.A(_07828_),
    .B(_00685_),
    .Y(_07834_));
 AO21x1_ASAP7_75t_R _31001_ (.A1(_07823_),
    .A2(net258),
    .B(_07834_),
    .Y(_01348_));
 BUFx4f_ASAP7_75t_R _31002_ (.A(_08379_),
    .Y(_07835_));
 NOR2x1_ASAP7_75t_R _31003_ (.A(_07828_),
    .B(_00594_),
    .Y(_07836_));
 AO21x1_ASAP7_75t_R _31004_ (.A1(_07835_),
    .A2(net259),
    .B(_07836_),
    .Y(_01349_));
 NOR2x1_ASAP7_75t_R _31005_ (.A(_07828_),
    .B(_00593_),
    .Y(_07837_));
 AO21x1_ASAP7_75t_R _31006_ (.A1(_07835_),
    .A2(net260),
    .B(_07837_),
    .Y(_01350_));
 NOR2x1_ASAP7_75t_R _31007_ (.A(_07828_),
    .B(_00596_),
    .Y(_07838_));
 AO21x1_ASAP7_75t_R _31008_ (.A1(_07835_),
    .A2(net261),
    .B(_07838_),
    .Y(_01351_));
 NOR2x1_ASAP7_75t_R _31009_ (.A(_07828_),
    .B(_00684_),
    .Y(_07839_));
 AO21x1_ASAP7_75t_R _31010_ (.A1(_07835_),
    .A2(net262),
    .B(_07839_),
    .Y(_01352_));
 BUFx6f_ASAP7_75t_R _31011_ (.A(_07767_),
    .Y(_07840_));
 NOR2x1_ASAP7_75t_R _31012_ (.A(_07840_),
    .B(_00683_),
    .Y(_07841_));
 AO21x1_ASAP7_75t_R _31013_ (.A1(_07835_),
    .A2(net263),
    .B(_07841_),
    .Y(_01353_));
 NOR2x1_ASAP7_75t_R _31014_ (.A(_07840_),
    .B(_00682_),
    .Y(_07842_));
 AO21x1_ASAP7_75t_R _31015_ (.A1(_07835_),
    .A2(net264),
    .B(_07842_),
    .Y(_01354_));
 NOR2x1_ASAP7_75t_R _31016_ (.A(_07840_),
    .B(_00681_),
    .Y(_07843_));
 AO21x1_ASAP7_75t_R _31017_ (.A1(_07835_),
    .A2(net265),
    .B(_07843_),
    .Y(_01355_));
 NOR2x1_ASAP7_75t_R _31018_ (.A(_07840_),
    .B(_00680_),
    .Y(_07844_));
 AO21x1_ASAP7_75t_R _31019_ (.A1(_07835_),
    .A2(net266),
    .B(_07844_),
    .Y(_01356_));
 NOR2x1_ASAP7_75t_R _31020_ (.A(_07840_),
    .B(_00550_),
    .Y(_07845_));
 AO21x1_ASAP7_75t_R _31021_ (.A1(_07835_),
    .A2(net267),
    .B(_07845_),
    .Y(_01357_));
 NOR2x1_ASAP7_75t_R _31022_ (.A(_07840_),
    .B(_00549_),
    .Y(_07846_));
 AO21x1_ASAP7_75t_R _31023_ (.A1(_07835_),
    .A2(net268),
    .B(_07846_),
    .Y(_01358_));
 BUFx6f_ASAP7_75t_R _31024_ (.A(_08379_),
    .Y(_07847_));
 NOR2x1_ASAP7_75t_R _31025_ (.A(_07840_),
    .B(_00679_),
    .Y(_07848_));
 AO21x1_ASAP7_75t_R _31026_ (.A1(_07847_),
    .A2(net269),
    .B(_07848_),
    .Y(_01359_));
 NOR2x1_ASAP7_75t_R _31027_ (.A(_07840_),
    .B(_00552_),
    .Y(_07849_));
 AO21x1_ASAP7_75t_R _31028_ (.A1(_07847_),
    .A2(net270),
    .B(_07849_),
    .Y(_01360_));
 NOR2x1_ASAP7_75t_R _31029_ (.A(_07840_),
    .B(_00678_),
    .Y(_07850_));
 AO21x1_ASAP7_75t_R _31030_ (.A1(_07847_),
    .A2(net271),
    .B(_07850_),
    .Y(_01361_));
 NOR2x1_ASAP7_75t_R _31031_ (.A(_07840_),
    .B(_00677_),
    .Y(_07851_));
 AO21x1_ASAP7_75t_R _31032_ (.A1(_07847_),
    .A2(net272),
    .B(_07851_),
    .Y(_01362_));
 BUFx6f_ASAP7_75t_R _31033_ (.A(_07767_),
    .Y(_07852_));
 NOR2x1_ASAP7_75t_R _31034_ (.A(_07852_),
    .B(_00676_),
    .Y(_07853_));
 AO21x1_ASAP7_75t_R _31035_ (.A1(_07847_),
    .A2(net273),
    .B(_07853_),
    .Y(_01363_));
 NOR2x1_ASAP7_75t_R _31036_ (.A(_07852_),
    .B(_00675_),
    .Y(_07854_));
 AO21x1_ASAP7_75t_R _31037_ (.A1(_07847_),
    .A2(net274),
    .B(_07854_),
    .Y(_01364_));
 NOR2x1_ASAP7_75t_R _31038_ (.A(_07852_),
    .B(_00674_),
    .Y(_07855_));
 AO21x1_ASAP7_75t_R _31039_ (.A1(_07847_),
    .A2(net275),
    .B(_07855_),
    .Y(_01365_));
 NOR2x1_ASAP7_75t_R _31040_ (.A(_07852_),
    .B(_00510_),
    .Y(_07856_));
 AO21x1_ASAP7_75t_R _31041_ (.A1(_07847_),
    .A2(net276),
    .B(_07856_),
    .Y(_01366_));
 NOR2x1_ASAP7_75t_R _31042_ (.A(_07852_),
    .B(_00509_),
    .Y(_07857_));
 AO21x1_ASAP7_75t_R _31043_ (.A1(_07847_),
    .A2(net277),
    .B(_07857_),
    .Y(_01367_));
 NOR2x1_ASAP7_75t_R _31044_ (.A(_07852_),
    .B(_00512_),
    .Y(_07858_));
 AO21x1_ASAP7_75t_R _31045_ (.A1(_07847_),
    .A2(net278),
    .B(_07858_),
    .Y(_01368_));
 BUFx6f_ASAP7_75t_R _31046_ (.A(_08319_),
    .Y(_07859_));
 NOR2x1_ASAP7_75t_R _31047_ (.A(_07852_),
    .B(_00673_),
    .Y(_07860_));
 AO21x1_ASAP7_75t_R _31048_ (.A1(_07859_),
    .A2(net279),
    .B(_07860_),
    .Y(_01369_));
 NOR2x1_ASAP7_75t_R _31049_ (.A(_07852_),
    .B(_00672_),
    .Y(_07861_));
 AO21x1_ASAP7_75t_R _31050_ (.A1(_07859_),
    .A2(net280),
    .B(_07861_),
    .Y(_01370_));
 NOR2x1_ASAP7_75t_R _31051_ (.A(_07852_),
    .B(_00671_),
    .Y(_07862_));
 AO21x1_ASAP7_75t_R _31052_ (.A1(_07859_),
    .A2(net281),
    .B(_07862_),
    .Y(_01371_));
 NOR2x1_ASAP7_75t_R _31053_ (.A(_07852_),
    .B(_00670_),
    .Y(_07863_));
 AO21x1_ASAP7_75t_R _31054_ (.A1(_07859_),
    .A2(net282),
    .B(_07863_),
    .Y(_01372_));
 BUFx6f_ASAP7_75t_R _31055_ (.A(_07767_),
    .Y(_07864_));
 NOR2x1_ASAP7_75t_R _31056_ (.A(_07864_),
    .B(_00669_),
    .Y(_07865_));
 AO21x1_ASAP7_75t_R _31057_ (.A1(_07859_),
    .A2(net283),
    .B(_07865_),
    .Y(_01373_));
 NOR2x1_ASAP7_75t_R _31058_ (.A(_07864_),
    .B(_00668_),
    .Y(_07866_));
 AO21x1_ASAP7_75t_R _31059_ (.A1(_07859_),
    .A2(net284),
    .B(_07866_),
    .Y(_01374_));
 NOR2x1_ASAP7_75t_R _31060_ (.A(_07864_),
    .B(_00628_),
    .Y(_07867_));
 AO21x1_ASAP7_75t_R _31061_ (.A1(_07859_),
    .A2(net285),
    .B(_07867_),
    .Y(_01375_));
 NOR2x1_ASAP7_75t_R _31062_ (.A(_07864_),
    .B(_00627_),
    .Y(_07868_));
 AO21x1_ASAP7_75t_R _31063_ (.A1(_07859_),
    .A2(net286),
    .B(_07868_),
    .Y(_01376_));
 NOR2x1_ASAP7_75t_R _31064_ (.A(_07864_),
    .B(_00630_),
    .Y(_07869_));
 AO21x1_ASAP7_75t_R _31065_ (.A1(_07859_),
    .A2(net287),
    .B(_07869_),
    .Y(_01377_));
 NOR2x1_ASAP7_75t_R _31066_ (.A(_07864_),
    .B(_00667_),
    .Y(_07870_));
 AO21x1_ASAP7_75t_R _31067_ (.A1(_07859_),
    .A2(net288),
    .B(_07870_),
    .Y(_01378_));
 BUFx6f_ASAP7_75t_R _31068_ (.A(_08319_),
    .Y(_07871_));
 NOR2x1_ASAP7_75t_R _31069_ (.A(_07864_),
    .B(_00666_),
    .Y(_07872_));
 AO21x1_ASAP7_75t_R _31070_ (.A1(_07871_),
    .A2(net289),
    .B(_07872_),
    .Y(_01379_));
 NOR2x1_ASAP7_75t_R _31071_ (.A(_07864_),
    .B(_00665_),
    .Y(_07873_));
 AO21x1_ASAP7_75t_R _31072_ (.A1(_07871_),
    .A2(net290),
    .B(_07873_),
    .Y(_01380_));
 NOR2x1_ASAP7_75t_R _31073_ (.A(_07864_),
    .B(_00664_),
    .Y(_07874_));
 AO21x1_ASAP7_75t_R _31074_ (.A1(_07871_),
    .A2(net291),
    .B(_07874_),
    .Y(_01381_));
 NOR2x1_ASAP7_75t_R _31075_ (.A(_07864_),
    .B(_00663_),
    .Y(_07875_));
 AO21x1_ASAP7_75t_R _31076_ (.A1(_07871_),
    .A2(net292),
    .B(_07875_),
    .Y(_01382_));
 BUFx6f_ASAP7_75t_R _31077_ (.A(_07767_),
    .Y(_07876_));
 NOR2x1_ASAP7_75t_R _31078_ (.A(_07876_),
    .B(_00662_),
    .Y(_07877_));
 AO21x1_ASAP7_75t_R _31079_ (.A1(_07871_),
    .A2(net293),
    .B(_07877_),
    .Y(_01383_));
 NOR2x1_ASAP7_75t_R _31080_ (.A(_07876_),
    .B(_00582_),
    .Y(_07878_));
 AO21x1_ASAP7_75t_R _31081_ (.A1(_07871_),
    .A2(net294),
    .B(_07878_),
    .Y(_01384_));
 NOR2x1_ASAP7_75t_R _31082_ (.A(_07876_),
    .B(_00581_),
    .Y(_07879_));
 AO21x1_ASAP7_75t_R _31083_ (.A1(_07871_),
    .A2(net295),
    .B(_07879_),
    .Y(_01385_));
 NOR2x1_ASAP7_75t_R _31084_ (.A(_07876_),
    .B(_00584_),
    .Y(_07880_));
 AO21x1_ASAP7_75t_R _31085_ (.A1(_07871_),
    .A2(net296),
    .B(_07880_),
    .Y(_01386_));
 NOR2x1_ASAP7_75t_R _31086_ (.A(_07876_),
    .B(_00661_),
    .Y(_07881_));
 AO21x1_ASAP7_75t_R _31087_ (.A1(_07871_),
    .A2(net297),
    .B(_07881_),
    .Y(_01387_));
 NOR2x1_ASAP7_75t_R _31088_ (.A(_07876_),
    .B(_00660_),
    .Y(_07882_));
 AO21x1_ASAP7_75t_R _31089_ (.A1(_07871_),
    .A2(net298),
    .B(_07882_),
    .Y(_01388_));
 BUFx6f_ASAP7_75t_R _31090_ (.A(_08319_),
    .Y(_07883_));
 NOR2x1_ASAP7_75t_R _31091_ (.A(_07876_),
    .B(_00659_),
    .Y(_07884_));
 AO21x1_ASAP7_75t_R _31092_ (.A1(_07883_),
    .A2(net299),
    .B(_07884_),
    .Y(_01389_));
 NOR2x1_ASAP7_75t_R _31093_ (.A(_07876_),
    .B(_00658_),
    .Y(_07885_));
 AO21x1_ASAP7_75t_R _31094_ (.A1(_07883_),
    .A2(net300),
    .B(_07885_),
    .Y(_01390_));
 NOR2x1_ASAP7_75t_R _31095_ (.A(_07876_),
    .B(_00657_),
    .Y(_07886_));
 AO21x1_ASAP7_75t_R _31096_ (.A1(_07883_),
    .A2(net301),
    .B(_07886_),
    .Y(_01391_));
 NOR2x1_ASAP7_75t_R _31097_ (.A(_07876_),
    .B(_00656_),
    .Y(_07887_));
 AO21x1_ASAP7_75t_R _31098_ (.A1(_07883_),
    .A2(net302),
    .B(_07887_),
    .Y(_01392_));
 BUFx6f_ASAP7_75t_R _31099_ (.A(_08252_),
    .Y(_07888_));
 NOR2x1_ASAP7_75t_R _31100_ (.A(_07888_),
    .B(_00540_),
    .Y(_07889_));
 AO21x1_ASAP7_75t_R _31101_ (.A1(_07883_),
    .A2(net303),
    .B(_07889_),
    .Y(_01393_));
 NOR2x1_ASAP7_75t_R _31102_ (.A(_07888_),
    .B(_00539_),
    .Y(_07890_));
 AO21x1_ASAP7_75t_R _31103_ (.A1(_07883_),
    .A2(net304),
    .B(_07890_),
    .Y(_01394_));
 NOR2x1_ASAP7_75t_R _31104_ (.A(_07888_),
    .B(_00542_),
    .Y(_07891_));
 AO21x1_ASAP7_75t_R _31105_ (.A1(_07883_),
    .A2(net305),
    .B(_07891_),
    .Y(_01395_));
 NOR2x1_ASAP7_75t_R _31106_ (.A(_07888_),
    .B(_00655_),
    .Y(_07892_));
 AO21x1_ASAP7_75t_R _31107_ (.A1(_07883_),
    .A2(net306),
    .B(_07892_),
    .Y(_01396_));
 NOR2x1_ASAP7_75t_R _31108_ (.A(_07888_),
    .B(_00654_),
    .Y(_07893_));
 AO21x1_ASAP7_75t_R _31109_ (.A1(_07883_),
    .A2(net307),
    .B(_07893_),
    .Y(_01397_));
 NOR2x1_ASAP7_75t_R _31110_ (.A(_07888_),
    .B(_00653_),
    .Y(_07894_));
 AO21x1_ASAP7_75t_R _31111_ (.A1(_07883_),
    .A2(net308),
    .B(_07894_),
    .Y(_01398_));
 BUFx4f_ASAP7_75t_R _31112_ (.A(_08319_),
    .Y(_07895_));
 NOR2x1_ASAP7_75t_R _31113_ (.A(_07888_),
    .B(_00652_),
    .Y(_07896_));
 AO21x1_ASAP7_75t_R _31114_ (.A1(_07895_),
    .A2(net309),
    .B(_07896_),
    .Y(_01399_));
 NOR2x1_ASAP7_75t_R _31115_ (.A(_07888_),
    .B(_00651_),
    .Y(_07897_));
 AO21x1_ASAP7_75t_R _31116_ (.A1(_07895_),
    .A2(net310),
    .B(_07897_),
    .Y(_01400_));
 NOR2x1_ASAP7_75t_R _31117_ (.A(_07888_),
    .B(_00500_),
    .Y(_07898_));
 AO21x1_ASAP7_75t_R _31118_ (.A1(_07895_),
    .A2(net311),
    .B(_07898_),
    .Y(_01401_));
 NOR2x1_ASAP7_75t_R _31119_ (.A(_07888_),
    .B(_00499_),
    .Y(_07899_));
 AO21x1_ASAP7_75t_R _31120_ (.A1(_07895_),
    .A2(net312),
    .B(_07899_),
    .Y(_01402_));
 BUFx6f_ASAP7_75t_R _31121_ (.A(_08252_),
    .Y(_07900_));
 NOR2x1_ASAP7_75t_R _31122_ (.A(_07900_),
    .B(_00606_),
    .Y(_07901_));
 AO21x1_ASAP7_75t_R _31123_ (.A1(_07895_),
    .A2(net313),
    .B(_07901_),
    .Y(_01403_));
 NOR2x1_ASAP7_75t_R _31124_ (.A(_07900_),
    .B(_00502_),
    .Y(_07902_));
 AO21x1_ASAP7_75t_R _31125_ (.A1(_07895_),
    .A2(net314),
    .B(_07902_),
    .Y(_01404_));
 NOR2x1_ASAP7_75t_R _31126_ (.A(_07900_),
    .B(_00650_),
    .Y(_07903_));
 AO21x1_ASAP7_75t_R _31127_ (.A1(_07895_),
    .A2(net315),
    .B(_07903_),
    .Y(_01405_));
 NOR2x1_ASAP7_75t_R _31128_ (.A(_07900_),
    .B(_00649_),
    .Y(_07904_));
 AO21x1_ASAP7_75t_R _31129_ (.A1(_07895_),
    .A2(net316),
    .B(_07904_),
    .Y(_01406_));
 NOR2x1_ASAP7_75t_R _31130_ (.A(_07900_),
    .B(_00648_),
    .Y(_07905_));
 AO21x1_ASAP7_75t_R _31131_ (.A1(_07895_),
    .A2(net317),
    .B(_07905_),
    .Y(_01407_));
 NOR2x1_ASAP7_75t_R _31132_ (.A(_07900_),
    .B(_00647_),
    .Y(_07906_));
 AO21x1_ASAP7_75t_R _31133_ (.A1(_07895_),
    .A2(net318),
    .B(_07906_),
    .Y(_01408_));
 NOR2x1_ASAP7_75t_R _31134_ (.A(_07900_),
    .B(_00646_),
    .Y(_07907_));
 AO21x1_ASAP7_75t_R _31135_ (.A1(_08321_),
    .A2(net319),
    .B(_07907_),
    .Y(_01409_));
 NOR2x1_ASAP7_75t_R _31136_ (.A(_07900_),
    .B(_00618_),
    .Y(_07908_));
 AO21x1_ASAP7_75t_R _31137_ (.A1(_08321_),
    .A2(net320),
    .B(_07908_),
    .Y(_01410_));
 NOR2x1_ASAP7_75t_R _31138_ (.A(_07900_),
    .B(_00617_),
    .Y(_07909_));
 AO21x1_ASAP7_75t_R _31139_ (.A1(_08321_),
    .A2(net321),
    .B(_07909_),
    .Y(_01411_));
 NOR2x1_ASAP7_75t_R _31140_ (.A(_07900_),
    .B(_00620_),
    .Y(_07910_));
 AO21x1_ASAP7_75t_R _31141_ (.A1(_08321_),
    .A2(net322),
    .B(_07910_),
    .Y(_01412_));
 NOR2x1_ASAP7_75t_R _31142_ (.A(_08253_),
    .B(_00645_),
    .Y(_07911_));
 AO21x1_ASAP7_75t_R _31143_ (.A1(_08321_),
    .A2(net323),
    .B(_07911_),
    .Y(_01413_));
 NOR2x1_ASAP7_75t_R _31144_ (.A(_08253_),
    .B(_00605_),
    .Y(_07912_));
 AO21x1_ASAP7_75t_R _31145_ (.A1(_08321_),
    .A2(net324),
    .B(_07912_),
    .Y(_01414_));
 AND3x1_ASAP7_75t_R _31146_ (.A(_00726_),
    .B(_00727_),
    .C(_00728_),
    .Y(_07913_));
 AOI21x1_ASAP7_75t_R _31147_ (.A1(_00727_),
    .A2(_00728_),
    .B(_00726_),
    .Y(_07914_));
 INVx1_ASAP7_75t_R _31148_ (.A(_07913_),
    .Y(_07915_));
 INVx1_ASAP7_75t_R _31149_ (.A(_00729_),
    .Y(_07916_));
 OA21x2_ASAP7_75t_R _31150_ (.A1(_07915_),
    .A2(_07916_),
    .B(net196),
    .Y(_07917_));
 OA211x2_ASAP7_75t_R _31151_ (.A1(_07913_),
    .A2(_07914_),
    .B(_07917_),
    .C(_08080_),
    .Y(_01285_));
 XNOR2x2_ASAP7_75t_R _31152_ (.A(_00643_),
    .B(_01282_),
    .Y(_07918_));
 INVx2_ASAP7_75t_R _31153_ (.A(_07918_),
    .Y(_07919_));
 OAI21x1_ASAP7_75t_R _31154_ (.A1(_00420_),
    .A2(_07919_),
    .B(_08251_),
    .Y(_01415_));
 OR3x1_ASAP7_75t_R _31155_ (.A(_00643_),
    .B(_16081_),
    .C(\u0.r0.rcnt_next[0] ),
    .Y(_07920_));
 XNOR2x2_ASAP7_75t_R _31156_ (.A(_00986_),
    .B(_07920_),
    .Y(_07921_));
 INVx1_ASAP7_75t_R _31157_ (.A(_01279_),
    .Y(_07922_));
 OR3x2_ASAP7_75t_R _31158_ (.A(_07921_),
    .B(_07922_),
    .C(_07919_),
    .Y(_07923_));
 INVx2_ASAP7_75t_R _31159_ (.A(_07921_),
    .Y(_07924_));
 OR3x1_ASAP7_75t_R _31160_ (.A(_07924_),
    .B(_00422_),
    .C(_07919_),
    .Y(_07925_));
 AOI21x1_ASAP7_75t_R _31161_ (.A1(_07923_),
    .A2(_07925_),
    .B(_08360_),
    .Y(_01416_));
 OR3x2_ASAP7_75t_R _31162_ (.A(_07921_),
    .B(_00422_),
    .C(_07919_),
    .Y(_07926_));
 OR3x1_ASAP7_75t_R _31163_ (.A(_07924_),
    .B(_01281_),
    .C(_07919_),
    .Y(_07927_));
 AOI21x1_ASAP7_75t_R _31164_ (.A1(_07926_),
    .A2(_07927_),
    .B(_08360_),
    .Y(_01417_));
 OR3x1_ASAP7_75t_R _31165_ (.A(_07921_),
    .B(_00420_),
    .C(_07919_),
    .Y(_07928_));
 OR3x1_ASAP7_75t_R _31166_ (.A(_07924_),
    .B(_01280_),
    .C(_07919_),
    .Y(_07929_));
 AOI21x1_ASAP7_75t_R _31167_ (.A1(_07928_),
    .A2(_07929_),
    .B(_08360_),
    .Y(_01418_));
 OR3x1_ASAP7_75t_R _31168_ (.A(_07924_),
    .B(_00420_),
    .C(_07918_),
    .Y(_07930_));
 AOI21x1_ASAP7_75t_R _31169_ (.A1(_07923_),
    .A2(_07930_),
    .B(_08360_),
    .Y(_01419_));
 OR3x1_ASAP7_75t_R _31170_ (.A(_07924_),
    .B(_00422_),
    .C(_07918_),
    .Y(_07931_));
 AOI21x1_ASAP7_75t_R _31171_ (.A1(_07926_),
    .A2(_07931_),
    .B(_08360_),
    .Y(_01420_));
 NOR2x1_ASAP7_75t_R _31172_ (.A(_07918_),
    .B(_07924_),
    .Y(_07932_));
 INVx1_ASAP7_75t_R _31173_ (.A(_01281_),
    .Y(_07933_));
 AND3x1_ASAP7_75t_R _31174_ (.A(_07932_),
    .B(_08367_),
    .C(_07933_),
    .Y(_01421_));
 INVx1_ASAP7_75t_R _31175_ (.A(_01280_),
    .Y(_07934_));
 AND3x1_ASAP7_75t_R _31176_ (.A(_07932_),
    .B(_08080_),
    .C(_07934_),
    .Y(_01422_));
 NOR2x1_ASAP7_75t_R _31177_ (.A(_08360_),
    .B(\u0.r0.rcnt[0] ),
    .Y(_01423_));
 NOR2x1_ASAP7_75t_R _31178_ (.A(_08360_),
    .B(_01279_),
    .Y(_01424_));
 NOR2x1_ASAP7_75t_R _31179_ (.A(_08360_),
    .B(_07918_),
    .Y(_01425_));
 NOR2x1_ASAP7_75t_R _31180_ (.A(_08360_),
    .B(_07921_),
    .Y(_01426_));
 AO22x1_ASAP7_75t_R _31181_ (.A1(_08321_),
    .A2(net196),
    .B1(_07917_),
    .B2(_00728_),
    .Y(_01283_));
 NAND2x1_ASAP7_75t_R _31182_ (.A(_00727_),
    .B(_00728_),
    .Y(_07935_));
 AO21x1_ASAP7_75t_R _31183_ (.A1(_00726_),
    .A2(_00729_),
    .B(_07935_),
    .Y(_07936_));
 OAI21x1_ASAP7_75t_R _31184_ (.A1(_00727_),
    .A2(_00728_),
    .B(_07936_),
    .Y(_07937_));
 OA21x2_ASAP7_75t_R _31185_ (.A1(_07937_),
    .A2(_08320_),
    .B(net196),
    .Y(_01284_));
 AO21x1_ASAP7_75t_R _31186_ (.A1(_07915_),
    .A2(_07916_),
    .B(_08253_),
    .Y(_07938_));
 AND2x2_ASAP7_75t_R _31187_ (.A(_07938_),
    .B(net196),
    .Y(_01286_));
 HAxp5_ASAP7_75t_R _31188_ (.A(_15729_),
    .B(_15730_),
    .CON(_00457_),
    .SN(_00456_));
 HAxp5_ASAP7_75t_R _31189_ (.A(_15729_),
    .B(_15730_),
    .CON(_01122_),
    .SN(_15731_));
 HAxp5_ASAP7_75t_R _31190_ (.A(_15729_),
    .B(_15732_),
    .CON(_00458_),
    .SN(_15733_));
 HAxp5_ASAP7_75t_R _31191_ (.A(_15729_),
    .B(_15732_),
    .CON(_01123_),
    .SN(_15734_));
 HAxp5_ASAP7_75t_R _31192_ (.A(_15735_),
    .B(_15730_),
    .CON(_00454_),
    .SN(_15736_));
 HAxp5_ASAP7_75t_R _31193_ (.A(_15735_),
    .B(_15730_),
    .CON(_01124_),
    .SN(_15737_));
 HAxp5_ASAP7_75t_R _31194_ (.A(_15735_),
    .B(_15732_),
    .CON(_00455_),
    .SN(_15738_));
 HAxp5_ASAP7_75t_R _31195_ (.A(_15735_),
    .B(_15732_),
    .CON(_01125_),
    .SN(_15739_));
 HAxp5_ASAP7_75t_R _31196_ (.A(_15729_),
    .B(_15740_),
    .CON(_00460_),
    .SN(_00462_));
 HAxp5_ASAP7_75t_R _31197_ (.A(_15729_),
    .B(_15740_),
    .CON(_01126_),
    .SN(_15741_));
 HAxp5_ASAP7_75t_R _31198_ (.A(_15729_),
    .B(_15742_),
    .CON(_00461_),
    .SN(_15743_));
 HAxp5_ASAP7_75t_R _31199_ (.A(_15729_),
    .B(_15742_),
    .CON(_01127_),
    .SN(_15744_));
 HAxp5_ASAP7_75t_R _31200_ (.A(_15735_),
    .B(_15740_),
    .CON(_00459_),
    .SN(_15745_));
 HAxp5_ASAP7_75t_R _31201_ (.A(_15735_),
    .B(_15740_),
    .CON(_01128_),
    .SN(_15746_));
 HAxp5_ASAP7_75t_R _31202_ (.A(_15747_),
    .B(_15748_),
    .CON(_00466_),
    .SN(_00465_));
 HAxp5_ASAP7_75t_R _31203_ (.A(_15747_),
    .B(_15748_),
    .CON(_01129_),
    .SN(_15749_));
 HAxp5_ASAP7_75t_R _31204_ (.A(_15750_),
    .B(_15747_),
    .CON(_00467_),
    .SN(_15751_));
 HAxp5_ASAP7_75t_R _31205_ (.A(_15747_),
    .B(_15750_),
    .CON(_01130_),
    .SN(_15752_));
 HAxp5_ASAP7_75t_R _31206_ (.A(_15753_),
    .B(_15748_),
    .CON(_00463_),
    .SN(_15754_));
 HAxp5_ASAP7_75t_R _31207_ (.A(_15753_),
    .B(_15748_),
    .CON(_01131_),
    .SN(_15755_));
 HAxp5_ASAP7_75t_R _31208_ (.A(_15753_),
    .B(_15750_),
    .CON(_00464_),
    .SN(_15756_));
 HAxp5_ASAP7_75t_R _31209_ (.A(_15753_),
    .B(_15750_),
    .CON(_01132_),
    .SN(_15757_));
 HAxp5_ASAP7_75t_R _31210_ (.A(_15747_),
    .B(_15758_),
    .CON(_00469_),
    .SN(_00471_));
 HAxp5_ASAP7_75t_R _31211_ (.A(_15747_),
    .B(_15758_),
    .CON(_01133_),
    .SN(_15759_));
 HAxp5_ASAP7_75t_R _31212_ (.A(_15747_),
    .B(_15760_),
    .CON(_00470_),
    .SN(_15761_));
 HAxp5_ASAP7_75t_R _31213_ (.A(_15747_),
    .B(_15760_),
    .CON(_01134_),
    .SN(_15762_));
 HAxp5_ASAP7_75t_R _31214_ (.A(net927),
    .B(_15758_),
    .CON(_00468_),
    .SN(_15763_));
 HAxp5_ASAP7_75t_R _31215_ (.A(net927),
    .B(_15758_),
    .CON(_01135_),
    .SN(_15764_));
 HAxp5_ASAP7_75t_R _31216_ (.A(_15766_),
    .B(_15765_),
    .CON(_00475_),
    .SN(_00474_));
 HAxp5_ASAP7_75t_R _31217_ (.A(_15765_),
    .B(_15766_),
    .CON(_01136_),
    .SN(_15767_));
 HAxp5_ASAP7_75t_R _31218_ (.A(_15765_),
    .B(_15768_),
    .CON(_00476_),
    .SN(_15769_));
 HAxp5_ASAP7_75t_R _31219_ (.A(_15765_),
    .B(_15768_),
    .CON(_01137_),
    .SN(_15770_));
 HAxp5_ASAP7_75t_R _31220_ (.A(_15771_),
    .B(_15766_),
    .CON(_00472_),
    .SN(_15772_));
 HAxp5_ASAP7_75t_R _31221_ (.A(_15771_),
    .B(_15766_),
    .CON(_01138_),
    .SN(_15773_));
 HAxp5_ASAP7_75t_R _31222_ (.A(_15771_),
    .B(_15768_),
    .CON(_00473_),
    .SN(_15774_));
 HAxp5_ASAP7_75t_R _31223_ (.A(_15771_),
    .B(_15768_),
    .CON(_01139_),
    .SN(_15775_));
 HAxp5_ASAP7_75t_R _31224_ (.A(net2),
    .B(_15776_),
    .CON(_00478_),
    .SN(_00480_));
 HAxp5_ASAP7_75t_R _31225_ (.A(net17),
    .B(_15776_),
    .CON(_01140_),
    .SN(_15777_));
 HAxp5_ASAP7_75t_R _31226_ (.A(net2),
    .B(_15778_),
    .CON(_00479_),
    .SN(_15779_));
 HAxp5_ASAP7_75t_R _31227_ (.A(net17),
    .B(_15778_),
    .CON(_01141_),
    .SN(_15780_));
 HAxp5_ASAP7_75t_R _31228_ (.A(_15771_),
    .B(_15776_),
    .CON(_00477_),
    .SN(_15781_));
 HAxp5_ASAP7_75t_R _31229_ (.A(_15771_),
    .B(_15776_),
    .CON(_01142_),
    .SN(_15782_));
 HAxp5_ASAP7_75t_R _31230_ (.A(net822),
    .B(_15783_),
    .CON(_00484_),
    .SN(_00483_));
 HAxp5_ASAP7_75t_R _31231_ (.A(_15783_),
    .B(net822),
    .CON(_01143_),
    .SN(_15785_));
 HAxp5_ASAP7_75t_R _31232_ (.A(_15786_),
    .B(_15783_),
    .CON(_00485_),
    .SN(_15787_));
 HAxp5_ASAP7_75t_R _31233_ (.A(_15783_),
    .B(_15786_),
    .CON(_01144_),
    .SN(_15788_));
 HAxp5_ASAP7_75t_R _31234_ (.A(net493),
    .B(net822),
    .CON(_00481_),
    .SN(_15790_));
 HAxp5_ASAP7_75t_R _31235_ (.A(net493),
    .B(net822),
    .CON(_01145_),
    .SN(_15791_));
 HAxp5_ASAP7_75t_R _31236_ (.A(_15789_),
    .B(_15786_),
    .CON(_00482_),
    .SN(_15792_));
 HAxp5_ASAP7_75t_R _31237_ (.A(net494),
    .B(_15786_),
    .CON(_01146_),
    .SN(_15793_));
 HAxp5_ASAP7_75t_R _31238_ (.A(_15794_),
    .B(net18),
    .CON(_00488_),
    .SN(_01147_));
 HAxp5_ASAP7_75t_R _31239_ (.A(_15794_),
    .B(_15783_),
    .CON(_01148_),
    .SN(_15795_));
 HAxp5_ASAP7_75t_R _31240_ (.A(_15796_),
    .B(_15783_),
    .CON(_00487_),
    .SN(_15797_));
 HAxp5_ASAP7_75t_R _31241_ (.A(_15796_),
    .B(net18),
    .CON(_01149_),
    .SN(_15798_));
 HAxp5_ASAP7_75t_R _31242_ (.A(_15796_),
    .B(net11),
    .CON(_00486_),
    .SN(_15799_));
 HAxp5_ASAP7_75t_R _31243_ (.A(_15796_),
    .B(net11),
    .CON(_01150_),
    .SN(_15800_));
 HAxp5_ASAP7_75t_R _31244_ (.A(_15801_),
    .B(_15802_),
    .CON(_00493_),
    .SN(_00494_));
 HAxp5_ASAP7_75t_R _31245_ (.A(_15801_),
    .B(_15802_),
    .CON(_01151_),
    .SN(_15803_));
 HAxp5_ASAP7_75t_R _31246_ (.A(_15801_),
    .B(_15804_),
    .CON(_01152_),
    .SN(_15805_));
 HAxp5_ASAP7_75t_R _31247_ (.A(_15806_),
    .B(_15802_),
    .CON(_00491_),
    .SN(_15807_));
 HAxp5_ASAP7_75t_R _31248_ (.A(_15806_),
    .B(_15802_),
    .CON(_01153_),
    .SN(_15808_));
 HAxp5_ASAP7_75t_R _31249_ (.A(_15806_),
    .B(_15804_),
    .CON(_00497_),
    .SN(_15809_));
 HAxp5_ASAP7_75t_R _31250_ (.A(_15806_),
    .B(_15804_),
    .CON(_01154_),
    .SN(_15810_));
 HAxp5_ASAP7_75t_R _31251_ (.A(_15811_),
    .B(_15802_),
    .CON(_01155_),
    .SN(_00498_));
 HAxp5_ASAP7_75t_R _31252_ (.A(_15811_),
    .B(_15804_),
    .CON(_00496_),
    .SN(_15812_));
 HAxp5_ASAP7_75t_R _31253_ (.A(_15811_),
    .B(_15804_),
    .CON(_01156_),
    .SN(_15813_));
 HAxp5_ASAP7_75t_R _31254_ (.A(_15814_),
    .B(_15802_),
    .CON(_00495_),
    .SN(_15815_));
 HAxp5_ASAP7_75t_R _31255_ (.A(_15814_),
    .B(_15802_),
    .CON(_01157_),
    .SN(_15816_));
 HAxp5_ASAP7_75t_R _31256_ (.A(_15814_),
    .B(_15804_),
    .CON(_01158_),
    .SN(_15817_));
 HAxp5_ASAP7_75t_R _31257_ (.A(_15818_),
    .B(_15819_),
    .CON(_00503_),
    .SN(_00504_));
 HAxp5_ASAP7_75t_R _31258_ (.A(_15818_),
    .B(_15819_),
    .CON(_01159_),
    .SN(_15820_));
 HAxp5_ASAP7_75t_R _31259_ (.A(_15821_),
    .B(_15818_),
    .CON(_01160_),
    .SN(_15822_));
 HAxp5_ASAP7_75t_R _31260_ (.A(_15823_),
    .B(_15819_),
    .CON(_00501_),
    .SN(_15824_));
 HAxp5_ASAP7_75t_R _31261_ (.A(_15823_),
    .B(_15819_),
    .CON(_01161_),
    .SN(_15825_));
 HAxp5_ASAP7_75t_R _31262_ (.A(_15823_),
    .B(_15821_),
    .CON(_00507_),
    .SN(_15826_));
 HAxp5_ASAP7_75t_R _31263_ (.A(_15823_),
    .B(_15821_),
    .CON(_01162_),
    .SN(_15827_));
 HAxp5_ASAP7_75t_R _31264_ (.A(_15828_),
    .B(net603),
    .CON(_01163_),
    .SN(_00508_));
 HAxp5_ASAP7_75t_R _31265_ (.A(_15828_),
    .B(_15821_),
    .CON(_00506_),
    .SN(_15829_));
 HAxp5_ASAP7_75t_R _31266_ (.A(_15828_),
    .B(_15821_),
    .CON(_01164_),
    .SN(_15830_));
 HAxp5_ASAP7_75t_R _31267_ (.A(_15831_),
    .B(_15819_),
    .CON(_00505_),
    .SN(_15832_));
 HAxp5_ASAP7_75t_R _31268_ (.A(_15831_),
    .B(net603),
    .CON(_01165_),
    .SN(_15833_));
 HAxp5_ASAP7_75t_R _31269_ (.A(_15831_),
    .B(_15821_),
    .CON(_01166_),
    .SN(_15834_));
 HAxp5_ASAP7_75t_R _31270_ (.A(_15835_),
    .B(_15836_),
    .CON(_00513_),
    .SN(_00514_));
 HAxp5_ASAP7_75t_R _31271_ (.A(_15835_),
    .B(_15836_),
    .CON(_01167_),
    .SN(_15837_));
 HAxp5_ASAP7_75t_R _31272_ (.A(_15835_),
    .B(_15838_),
    .CON(_01168_),
    .SN(_15839_));
 HAxp5_ASAP7_75t_R _31273_ (.A(_15840_),
    .B(_15836_),
    .CON(_00511_),
    .SN(_15841_));
 HAxp5_ASAP7_75t_R _31274_ (.A(_15840_),
    .B(_15836_),
    .CON(_01169_),
    .SN(_15842_));
 HAxp5_ASAP7_75t_R _31275_ (.A(_15840_),
    .B(_15838_),
    .CON(_00517_),
    .SN(_15843_));
 HAxp5_ASAP7_75t_R _31276_ (.A(_15840_),
    .B(_15838_),
    .CON(_01170_),
    .SN(_15844_));
 HAxp5_ASAP7_75t_R _31277_ (.A(_15845_),
    .B(_15836_),
    .CON(_01171_),
    .SN(_00518_));
 HAxp5_ASAP7_75t_R _31278_ (.A(_15845_),
    .B(_15838_),
    .CON(_00516_),
    .SN(_15846_));
 HAxp5_ASAP7_75t_R _31279_ (.A(_15845_),
    .B(_15838_),
    .CON(_01172_),
    .SN(_15847_));
 HAxp5_ASAP7_75t_R _31280_ (.A(_15848_),
    .B(_15836_),
    .CON(_00515_),
    .SN(_15849_));
 HAxp5_ASAP7_75t_R _31281_ (.A(_15848_),
    .B(_15836_),
    .CON(_01173_),
    .SN(_15850_));
 HAxp5_ASAP7_75t_R _31282_ (.A(_15848_),
    .B(_15838_),
    .CON(_01174_),
    .SN(_15851_));
 HAxp5_ASAP7_75t_R _31283_ (.A(_15852_),
    .B(_15853_),
    .CON(_00523_),
    .SN(_00524_));
 HAxp5_ASAP7_75t_R _31284_ (.A(_15853_),
    .B(_15852_),
    .CON(_01175_),
    .SN(_15854_));
 HAxp5_ASAP7_75t_R _31285_ (.A(_15855_),
    .B(_15852_),
    .CON(_01176_),
    .SN(_15856_));
 HAxp5_ASAP7_75t_R _31286_ (.A(_15857_),
    .B(_15853_),
    .CON(_00521_),
    .SN(_15858_));
 HAxp5_ASAP7_75t_R _31287_ (.A(_15857_),
    .B(_15853_),
    .CON(_01177_),
    .SN(_15859_));
 HAxp5_ASAP7_75t_R _31288_ (.A(_15857_),
    .B(_15855_),
    .CON(_00527_),
    .SN(_15860_));
 HAxp5_ASAP7_75t_R _31289_ (.A(_15855_),
    .B(_15857_),
    .CON(_01178_),
    .SN(_15861_));
 HAxp5_ASAP7_75t_R _31290_ (.A(_15862_),
    .B(_15853_),
    .CON(_01179_),
    .SN(_00528_));
 HAxp5_ASAP7_75t_R _31291_ (.A(_15862_),
    .B(_15855_),
    .CON(_00526_),
    .SN(_15863_));
 HAxp5_ASAP7_75t_R _31292_ (.A(_15862_),
    .B(_15855_),
    .CON(_01180_),
    .SN(_15864_));
 HAxp5_ASAP7_75t_R _31293_ (.A(_15865_),
    .B(_15853_),
    .CON(_00525_),
    .SN(_15866_));
 HAxp5_ASAP7_75t_R _31294_ (.A(_15865_),
    .B(_15853_),
    .CON(_01181_),
    .SN(_15867_));
 HAxp5_ASAP7_75t_R _31295_ (.A(_15865_),
    .B(_15855_),
    .CON(_01182_),
    .SN(_15868_));
 HAxp5_ASAP7_75t_R _31296_ (.A(_15870_),
    .B(_15869_),
    .CON(_00533_),
    .SN(_00534_));
 HAxp5_ASAP7_75t_R _31297_ (.A(_15869_),
    .B(_15870_),
    .CON(_01183_),
    .SN(_15871_));
 HAxp5_ASAP7_75t_R _31298_ (.A(_15872_),
    .B(_15869_),
    .CON(_01184_),
    .SN(_15873_));
 HAxp5_ASAP7_75t_R _31299_ (.A(_15874_),
    .B(_15870_),
    .CON(_00531_),
    .SN(_15875_));
 HAxp5_ASAP7_75t_R _31300_ (.A(_15874_),
    .B(_15870_),
    .CON(_01185_),
    .SN(_15876_));
 HAxp5_ASAP7_75t_R _31301_ (.A(_15874_),
    .B(net541),
    .CON(_00537_),
    .SN(_15877_));
 HAxp5_ASAP7_75t_R _31302_ (.A(_15874_),
    .B(_15872_),
    .CON(_01186_),
    .SN(_15878_));
 HAxp5_ASAP7_75t_R _31303_ (.A(_15879_),
    .B(_15870_),
    .CON(_01187_),
    .SN(_00538_));
 HAxp5_ASAP7_75t_R _31304_ (.A(_15879_),
    .B(net69),
    .CON(_00536_),
    .SN(_15880_));
 HAxp5_ASAP7_75t_R _31305_ (.A(_15879_),
    .B(net69),
    .CON(_01188_),
    .SN(_15881_));
 HAxp5_ASAP7_75t_R _31306_ (.A(_15882_),
    .B(_15870_),
    .CON(_00535_),
    .SN(_15883_));
 HAxp5_ASAP7_75t_R _31307_ (.A(_15882_),
    .B(_15870_),
    .CON(_01189_),
    .SN(_15884_));
 HAxp5_ASAP7_75t_R _31308_ (.A(_15882_),
    .B(net69),
    .CON(_01190_),
    .SN(_15885_));
 HAxp5_ASAP7_75t_R _31309_ (.A(_15886_),
    .B(_15887_),
    .CON(_00543_),
    .SN(_00544_));
 HAxp5_ASAP7_75t_R _31310_ (.A(_15886_),
    .B(_15887_),
    .CON(_01191_),
    .SN(_15888_));
 HAxp5_ASAP7_75t_R _31311_ (.A(_15889_),
    .B(_15886_),
    .CON(_01192_),
    .SN(_15890_));
 HAxp5_ASAP7_75t_R _31312_ (.A(_15887_),
    .B(_15891_),
    .CON(_00541_),
    .SN(_15892_));
 HAxp5_ASAP7_75t_R _31313_ (.A(_15887_),
    .B(_15891_),
    .CON(_01193_),
    .SN(_15893_));
 HAxp5_ASAP7_75t_R _31314_ (.A(_15891_),
    .B(net720),
    .CON(_00547_),
    .SN(_15894_));
 HAxp5_ASAP7_75t_R _31315_ (.A(_15891_),
    .B(_15889_),
    .CON(_01194_),
    .SN(_15895_));
 HAxp5_ASAP7_75t_R _31316_ (.A(_15896_),
    .B(net56),
    .CON(_01195_),
    .SN(_00548_));
 HAxp5_ASAP7_75t_R _31317_ (.A(_15896_),
    .B(net722),
    .CON(_00546_),
    .SN(_15897_));
 HAxp5_ASAP7_75t_R _31318_ (.A(_15896_),
    .B(net720),
    .CON(_01196_),
    .SN(_15898_));
 HAxp5_ASAP7_75t_R _31319_ (.A(_15899_),
    .B(_15887_),
    .CON(_00545_),
    .SN(_15900_));
 HAxp5_ASAP7_75t_R _31320_ (.A(_15899_),
    .B(net56),
    .CON(_01197_),
    .SN(_15901_));
 HAxp5_ASAP7_75t_R _31321_ (.A(_15899_),
    .B(net722),
    .CON(_01198_),
    .SN(_15902_));
 HAxp5_ASAP7_75t_R _31322_ (.A(_15903_),
    .B(_15904_),
    .CON(_00553_),
    .SN(_00554_));
 HAxp5_ASAP7_75t_R _31323_ (.A(_15904_),
    .B(_15903_),
    .CON(_01199_),
    .SN(_15905_));
 HAxp5_ASAP7_75t_R _31324_ (.A(_15903_),
    .B(_15906_),
    .CON(_01200_),
    .SN(_15907_));
 HAxp5_ASAP7_75t_R _31325_ (.A(_15908_),
    .B(_15904_),
    .CON(_00551_),
    .SN(_15909_));
 HAxp5_ASAP7_75t_R _31326_ (.A(_15908_),
    .B(_15904_),
    .CON(_01201_),
    .SN(_15910_));
 HAxp5_ASAP7_75t_R _31327_ (.A(_15908_),
    .B(_15906_),
    .CON(_00557_),
    .SN(_15911_));
 HAxp5_ASAP7_75t_R _31328_ (.A(_15908_),
    .B(_15906_),
    .CON(_01202_),
    .SN(_15912_));
 HAxp5_ASAP7_75t_R _31329_ (.A(_15913_),
    .B(_15904_),
    .CON(_01203_),
    .SN(_00558_));
 HAxp5_ASAP7_75t_R _31330_ (.A(_15913_),
    .B(_15906_),
    .CON(_00556_),
    .SN(_15914_));
 HAxp5_ASAP7_75t_R _31331_ (.A(_15913_),
    .B(_15906_),
    .CON(_01204_),
    .SN(_15915_));
 HAxp5_ASAP7_75t_R _31332_ (.A(_15916_),
    .B(_15904_),
    .CON(_00555_),
    .SN(_15917_));
 HAxp5_ASAP7_75t_R _31333_ (.A(_15916_),
    .B(_15904_),
    .CON(_01205_),
    .SN(_15918_));
 HAxp5_ASAP7_75t_R _31334_ (.A(_15916_),
    .B(_15906_),
    .CON(_01206_),
    .SN(_15919_));
 HAxp5_ASAP7_75t_R _31335_ (.A(_15920_),
    .B(_15921_),
    .CON(_00563_),
    .SN(_00564_));
 HAxp5_ASAP7_75t_R _31336_ (.A(_15920_),
    .B(_15921_),
    .CON(_01207_),
    .SN(_15922_));
 HAxp5_ASAP7_75t_R _31337_ (.A(_15923_),
    .B(_15920_),
    .CON(_01208_),
    .SN(_15924_));
 HAxp5_ASAP7_75t_R _31338_ (.A(_15925_),
    .B(_15921_),
    .CON(_00561_),
    .SN(_15926_));
 HAxp5_ASAP7_75t_R _31339_ (.A(_15925_),
    .B(_15921_),
    .CON(_01209_),
    .SN(_15927_));
 HAxp5_ASAP7_75t_R _31340_ (.A(_15925_),
    .B(_15923_),
    .CON(_00567_),
    .SN(_15928_));
 HAxp5_ASAP7_75t_R _31341_ (.A(_15925_),
    .B(_15923_),
    .CON(_01210_),
    .SN(_15929_));
 HAxp5_ASAP7_75t_R _31342_ (.A(_15930_),
    .B(_15921_),
    .CON(_01211_),
    .SN(_00568_));
 HAxp5_ASAP7_75t_R _31343_ (.A(_15930_),
    .B(_15923_),
    .CON(_00566_),
    .SN(_15931_));
 HAxp5_ASAP7_75t_R _31344_ (.A(_15930_),
    .B(_15923_),
    .CON(_01212_),
    .SN(_15932_));
 HAxp5_ASAP7_75t_R _31345_ (.A(_15933_),
    .B(_15921_),
    .CON(_00565_),
    .SN(_15934_));
 HAxp5_ASAP7_75t_R _31346_ (.A(_15933_),
    .B(_15921_),
    .CON(_01213_),
    .SN(_15935_));
 HAxp5_ASAP7_75t_R _31347_ (.A(_15933_),
    .B(_15923_),
    .CON(_01214_),
    .SN(_15936_));
 HAxp5_ASAP7_75t_R _31348_ (.A(_15937_),
    .B(_15938_),
    .CON(_00573_),
    .SN(_00574_));
 HAxp5_ASAP7_75t_R _31349_ (.A(_15937_),
    .B(_15938_),
    .CON(_01215_),
    .SN(_15939_));
 HAxp5_ASAP7_75t_R _31350_ (.A(_15937_),
    .B(_15940_),
    .CON(_00576_),
    .SN(_15941_));
 HAxp5_ASAP7_75t_R _31351_ (.A(_15937_),
    .B(_15940_),
    .CON(_01216_),
    .SN(_15942_));
 HAxp5_ASAP7_75t_R _31352_ (.A(_15943_),
    .B(_15938_),
    .CON(_00571_),
    .SN(_15944_));
 HAxp5_ASAP7_75t_R _31353_ (.A(_15943_),
    .B(_15938_),
    .CON(_01217_),
    .SN(_15945_));
 HAxp5_ASAP7_75t_R _31354_ (.A(_15940_),
    .B(_15943_),
    .CON(_00575_),
    .SN(_15946_));
 HAxp5_ASAP7_75t_R _31355_ (.A(_15943_),
    .B(_15940_),
    .CON(_01218_),
    .SN(_15947_));
 HAxp5_ASAP7_75t_R _31356_ (.A(_15948_),
    .B(_15938_),
    .CON(_01219_),
    .SN(_00580_));
 HAxp5_ASAP7_75t_R _31357_ (.A(_15948_),
    .B(_15940_),
    .CON(_00579_),
    .SN(_15949_));
 HAxp5_ASAP7_75t_R _31358_ (.A(_15948_),
    .B(_15940_),
    .CON(_01220_),
    .SN(_15950_));
 HAxp5_ASAP7_75t_R _31359_ (.A(_15951_),
    .B(_15938_),
    .CON(_00577_),
    .SN(_15952_));
 HAxp5_ASAP7_75t_R _31360_ (.A(_15951_),
    .B(net57),
    .CON(_01221_),
    .SN(_15953_));
 HAxp5_ASAP7_75t_R _31361_ (.A(_15951_),
    .B(_15940_),
    .CON(_00578_),
    .SN(_15954_));
 HAxp5_ASAP7_75t_R _31362_ (.A(_15951_),
    .B(_15940_),
    .CON(_01222_),
    .SN(_15955_));
 HAxp5_ASAP7_75t_R _31363_ (.A(_15956_),
    .B(_15957_),
    .CON(_00585_),
    .SN(_00586_));
 HAxp5_ASAP7_75t_R _31364_ (.A(_15956_),
    .B(_15957_),
    .CON(_01223_),
    .SN(_15958_));
 HAxp5_ASAP7_75t_R _31365_ (.A(_15956_),
    .B(net638),
    .CON(_00588_),
    .SN(_15960_));
 HAxp5_ASAP7_75t_R _31366_ (.A(_15956_),
    .B(_15959_),
    .CON(_01224_),
    .SN(_15961_));
 HAxp5_ASAP7_75t_R _31367_ (.A(_15962_),
    .B(net827),
    .CON(_00583_),
    .SN(_15963_));
 HAxp5_ASAP7_75t_R _31368_ (.A(_15962_),
    .B(net827),
    .CON(_01225_),
    .SN(_15964_));
 HAxp5_ASAP7_75t_R _31369_ (.A(_15959_),
    .B(_15962_),
    .CON(_00587_),
    .SN(_15965_));
 HAxp5_ASAP7_75t_R _31370_ (.A(_15962_),
    .B(_15959_),
    .CON(_01226_),
    .SN(_15966_));
 HAxp5_ASAP7_75t_R _31371_ (.A(_15967_),
    .B(_15957_),
    .CON(_01227_),
    .SN(_00592_));
 HAxp5_ASAP7_75t_R _31372_ (.A(_15967_),
    .B(net637),
    .CON(_00591_),
    .SN(_15968_));
 HAxp5_ASAP7_75t_R _31373_ (.A(_15967_),
    .B(_15959_),
    .CON(_01228_),
    .SN(_15969_));
 HAxp5_ASAP7_75t_R _31374_ (.A(_15970_),
    .B(net7),
    .CON(_00589_),
    .SN(_15971_));
 HAxp5_ASAP7_75t_R _31375_ (.A(_15970_),
    .B(_15957_),
    .CON(_01229_),
    .SN(_15972_));
 HAxp5_ASAP7_75t_R _31376_ (.A(_15970_),
    .B(net637),
    .CON(_00590_),
    .SN(_15973_));
 HAxp5_ASAP7_75t_R _31377_ (.A(_15970_),
    .B(net636),
    .CON(_01230_),
    .SN(_15974_));
 HAxp5_ASAP7_75t_R _31378_ (.A(_15975_),
    .B(_15976_),
    .CON(_00597_),
    .SN(_00598_));
 HAxp5_ASAP7_75t_R _31379_ (.A(_15975_),
    .B(_15976_),
    .CON(_01231_),
    .SN(_15977_));
 HAxp5_ASAP7_75t_R _31380_ (.A(_15975_),
    .B(_15978_),
    .CON(_00600_),
    .SN(_15979_));
 HAxp5_ASAP7_75t_R _31381_ (.A(_15975_),
    .B(_15978_),
    .CON(_01232_),
    .SN(_15980_));
 HAxp5_ASAP7_75t_R _31382_ (.A(_15981_),
    .B(_15976_),
    .CON(_00595_),
    .SN(_15982_));
 HAxp5_ASAP7_75t_R _31383_ (.A(_15976_),
    .B(_15981_),
    .CON(_01233_),
    .SN(_15983_));
 HAxp5_ASAP7_75t_R _31384_ (.A(_15978_),
    .B(_15981_),
    .CON(_00599_),
    .SN(_15984_));
 HAxp5_ASAP7_75t_R _31385_ (.A(_15978_),
    .B(_15981_),
    .CON(_01234_),
    .SN(_15985_));
 HAxp5_ASAP7_75t_R _31386_ (.A(_15986_),
    .B(_15976_),
    .CON(_01235_),
    .SN(_00604_));
 HAxp5_ASAP7_75t_R _31387_ (.A(_15986_),
    .B(net587),
    .CON(_00603_),
    .SN(_15987_));
 HAxp5_ASAP7_75t_R _31388_ (.A(_15986_),
    .B(net587),
    .CON(_01236_),
    .SN(_15988_));
 HAxp5_ASAP7_75t_R _31389_ (.A(_15989_),
    .B(net46),
    .CON(_00601_),
    .SN(_15990_));
 HAxp5_ASAP7_75t_R _31390_ (.A(_15989_),
    .B(_15976_),
    .CON(_01237_),
    .SN(_15991_));
 HAxp5_ASAP7_75t_R _31391_ (.A(_15989_),
    .B(net587),
    .CON(_00602_),
    .SN(_15992_));
 HAxp5_ASAP7_75t_R _31392_ (.A(_15989_),
    .B(net589),
    .CON(_01238_),
    .SN(_15993_));
 HAxp5_ASAP7_75t_R _31393_ (.A(_15994_),
    .B(_15995_),
    .CON(_00609_),
    .SN(_00610_));
 HAxp5_ASAP7_75t_R _31394_ (.A(_15994_),
    .B(_15995_),
    .CON(_01239_),
    .SN(_15996_));
 HAxp5_ASAP7_75t_R _31395_ (.A(_15994_),
    .B(_15997_),
    .CON(_00612_),
    .SN(_15998_));
 HAxp5_ASAP7_75t_R _31396_ (.A(_15994_),
    .B(_15997_),
    .CON(_01240_),
    .SN(_15999_));
 HAxp5_ASAP7_75t_R _31397_ (.A(_16000_),
    .B(_15995_),
    .CON(_00607_),
    .SN(_16001_));
 HAxp5_ASAP7_75t_R _31398_ (.A(_16000_),
    .B(_15995_),
    .CON(_01241_),
    .SN(_16002_));
 HAxp5_ASAP7_75t_R _31399_ (.A(_16000_),
    .B(_15997_),
    .CON(_00611_),
    .SN(_16003_));
 HAxp5_ASAP7_75t_R _31400_ (.A(_16000_),
    .B(_15997_),
    .CON(_01242_),
    .SN(_16004_));
 HAxp5_ASAP7_75t_R _31401_ (.A(_16005_),
    .B(net36),
    .CON(_01243_),
    .SN(_00616_));
 HAxp5_ASAP7_75t_R _31402_ (.A(_16005_),
    .B(_15997_),
    .CON(_00615_),
    .SN(_16006_));
 HAxp5_ASAP7_75t_R _31403_ (.A(_16005_),
    .B(_15997_),
    .CON(_01244_),
    .SN(_16007_));
 HAxp5_ASAP7_75t_R _31404_ (.A(_16008_),
    .B(_15995_),
    .CON(_00613_),
    .SN(_16009_));
 HAxp5_ASAP7_75t_R _31405_ (.A(_16008_),
    .B(_15995_),
    .CON(_01245_),
    .SN(_16010_));
 HAxp5_ASAP7_75t_R _31406_ (.A(_16008_),
    .B(_15997_),
    .CON(_00614_),
    .SN(_16011_));
 HAxp5_ASAP7_75t_R _31407_ (.A(_16008_),
    .B(_15997_),
    .CON(_01246_),
    .SN(_16012_));
 HAxp5_ASAP7_75t_R _31408_ (.A(_05057_),
    .B(_16014_),
    .CON(_00621_),
    .SN(_00622_));
 HAxp5_ASAP7_75t_R _31409_ (.A(net765),
    .B(_16014_),
    .CON(_01247_),
    .SN(_16015_));
 HAxp5_ASAP7_75t_R _31410_ (.A(net765),
    .B(_16016_),
    .CON(_01248_),
    .SN(_16017_));
 HAxp5_ASAP7_75t_R _31411_ (.A(_16018_),
    .B(_16014_),
    .CON(_00619_),
    .SN(_16019_));
 HAxp5_ASAP7_75t_R _31412_ (.A(_16014_),
    .B(_16018_),
    .CON(_01249_),
    .SN(_16020_));
 HAxp5_ASAP7_75t_R _31413_ (.A(_16018_),
    .B(_16016_),
    .CON(_00625_),
    .SN(_16021_));
 HAxp5_ASAP7_75t_R _31414_ (.A(_16018_),
    .B(_16016_),
    .CON(_01250_),
    .SN(_16022_));
 HAxp5_ASAP7_75t_R _31415_ (.A(_16023_),
    .B(_16014_),
    .CON(_01251_),
    .SN(_00626_));
 HAxp5_ASAP7_75t_R _31416_ (.A(_16023_),
    .B(_16016_),
    .CON(_00624_),
    .SN(_16024_));
 HAxp5_ASAP7_75t_R _31417_ (.A(_16023_),
    .B(_16016_),
    .CON(_01252_),
    .SN(_16025_));
 HAxp5_ASAP7_75t_R _31418_ (.A(_16026_),
    .B(net43),
    .CON(_00623_),
    .SN(_16027_));
 HAxp5_ASAP7_75t_R _31419_ (.A(_16026_),
    .B(net43),
    .CON(_01253_),
    .SN(_16028_));
 HAxp5_ASAP7_75t_R _31420_ (.A(_16026_),
    .B(_16016_),
    .CON(_01254_),
    .SN(_16029_));
 HAxp5_ASAP7_75t_R _31421_ (.A(_16030_),
    .B(_16031_),
    .CON(_00631_),
    .SN(_00632_));
 HAxp5_ASAP7_75t_R _31422_ (.A(_16030_),
    .B(_16031_),
    .CON(_01255_),
    .SN(_16032_));
 HAxp5_ASAP7_75t_R _31423_ (.A(_16030_),
    .B(_16033_),
    .CON(_01256_),
    .SN(_16034_));
 HAxp5_ASAP7_75t_R _31424_ (.A(_16035_),
    .B(_16031_),
    .CON(_00629_),
    .SN(_16036_));
 HAxp5_ASAP7_75t_R _31425_ (.A(_16035_),
    .B(_16031_),
    .CON(_01257_),
    .SN(_16037_));
 HAxp5_ASAP7_75t_R _31426_ (.A(_16035_),
    .B(_16033_),
    .CON(_00635_),
    .SN(_16038_));
 HAxp5_ASAP7_75t_R _31427_ (.A(_16035_),
    .B(_16033_),
    .CON(_01258_),
    .SN(_16039_));
 HAxp5_ASAP7_75t_R _31428_ (.A(_16040_),
    .B(_16031_),
    .CON(_01259_),
    .SN(_00636_));
 HAxp5_ASAP7_75t_R _31429_ (.A(_16040_),
    .B(_16033_),
    .CON(_00634_),
    .SN(_16041_));
 HAxp5_ASAP7_75t_R _31430_ (.A(_16040_),
    .B(_16033_),
    .CON(_01260_),
    .SN(_16042_));
 HAxp5_ASAP7_75t_R _31431_ (.A(_16043_),
    .B(_16031_),
    .CON(_00633_),
    .SN(_16044_));
 HAxp5_ASAP7_75t_R _31432_ (.A(_16043_),
    .B(_16031_),
    .CON(_01261_),
    .SN(_16045_));
 HAxp5_ASAP7_75t_R _31433_ (.A(_16043_),
    .B(_16033_),
    .CON(_01262_),
    .SN(_16046_));
 HAxp5_ASAP7_75t_R _31434_ (.A(_16048_),
    .B(_16047_),
    .CON(_00640_),
    .SN(_00641_));
 HAxp5_ASAP7_75t_R _31435_ (.A(_16047_),
    .B(_16048_),
    .CON(_01263_),
    .SN(_16049_));
 HAxp5_ASAP7_75t_R _31436_ (.A(_16047_),
    .B(_16050_),
    .CON(_01264_),
    .SN(_16051_));
 HAxp5_ASAP7_75t_R _31437_ (.A(_16052_),
    .B(_16048_),
    .CON(_00408_),
    .SN(_16053_));
 HAxp5_ASAP7_75t_R _31438_ (.A(_16052_),
    .B(_16048_),
    .CON(_01265_),
    .SN(_16054_));
 HAxp5_ASAP7_75t_R _31439_ (.A(_16052_),
    .B(_16050_),
    .CON(_00407_),
    .SN(_16055_));
 HAxp5_ASAP7_75t_R _31440_ (.A(_16052_),
    .B(_16050_),
    .CON(_01266_),
    .SN(_16056_));
 HAxp5_ASAP7_75t_R _31441_ (.A(_16057_),
    .B(net26),
    .CON(_01267_),
    .SN(_00409_));
 HAxp5_ASAP7_75t_R _31442_ (.A(_16057_),
    .B(_16050_),
    .CON(_00406_),
    .SN(_16058_));
 HAxp5_ASAP7_75t_R _31443_ (.A(_16057_),
    .B(_16050_),
    .CON(_01268_),
    .SN(_16059_));
 HAxp5_ASAP7_75t_R _31444_ (.A(_16060_),
    .B(_16048_),
    .CON(_00405_),
    .SN(_16061_));
 HAxp5_ASAP7_75t_R _31445_ (.A(_16060_),
    .B(_16048_),
    .CON(_01269_),
    .SN(_16062_));
 HAxp5_ASAP7_75t_R _31446_ (.A(_16060_),
    .B(_16050_),
    .CON(_01270_),
    .SN(_16063_));
 HAxp5_ASAP7_75t_R _31447_ (.A(_16065_),
    .B(_16064_),
    .CON(_00414_),
    .SN(_00415_));
 HAxp5_ASAP7_75t_R _31448_ (.A(_16065_),
    .B(_16064_),
    .CON(_01271_),
    .SN(_16066_));
 HAxp5_ASAP7_75t_R _31449_ (.A(_16064_),
    .B(_16067_),
    .CON(_01272_),
    .SN(_16068_));
 HAxp5_ASAP7_75t_R _31450_ (.A(_16069_),
    .B(_16065_),
    .CON(_00412_),
    .SN(_16070_));
 HAxp5_ASAP7_75t_R _31451_ (.A(_16069_),
    .B(_16065_),
    .CON(_01273_),
    .SN(_16071_));
 HAxp5_ASAP7_75t_R _31452_ (.A(_16069_),
    .B(_16067_),
    .CON(_00419_),
    .SN(_16072_));
 HAxp5_ASAP7_75t_R _31453_ (.A(_16069_),
    .B(_16067_),
    .CON(_01274_),
    .SN(_16073_));
 HAxp5_ASAP7_75t_R _31454_ (.A(_16074_),
    .B(_16065_),
    .CON(_01275_),
    .SN(_00421_));
 HAxp5_ASAP7_75t_R _31455_ (.A(_16074_),
    .B(_16067_),
    .CON(_00418_),
    .SN(_16075_));
 HAxp5_ASAP7_75t_R _31456_ (.A(_16074_),
    .B(_16067_),
    .CON(_01276_),
    .SN(_16076_));
 HAxp5_ASAP7_75t_R _31457_ (.A(_16077_),
    .B(_16065_),
    .CON(_00417_),
    .SN(_16078_));
 HAxp5_ASAP7_75t_R _31458_ (.A(_16077_),
    .B(_16065_),
    .CON(_01277_),
    .SN(_16079_));
 HAxp5_ASAP7_75t_R _31459_ (.A(_16077_),
    .B(_16067_),
    .CON(_01278_),
    .SN(_16080_));
 HAxp5_ASAP7_75t_R _31460_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_16081_),
    .CON(_00422_),
    .SN(_01279_));
 HAxp5_ASAP7_75t_R _31461_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_01280_),
    .SN(_16082_));
 HAxp5_ASAP7_75t_R _31462_ (.A(\u0.r0.rcnt[0] ),
    .B(_16081_),
    .CON(_01281_),
    .SN(_16083_));
 HAxp5_ASAP7_75t_R _31463_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00420_),
    .SN(_16084_));
 HAxp5_ASAP7_75t_R _31464_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_01282_),
    .SN(_16085_));
 DFFHQNx2_ASAP7_75t_R \dcnt[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_01283_),
    .QN(_00728_));
 DFFHQNx2_ASAP7_75t_R \dcnt[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_01284_),
    .QN(_00727_));
 DFFHQNx2_ASAP7_75t_R \dcnt[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .D(_01285_),
    .QN(_00726_));
 DFFHQNx2_ASAP7_75t_R \dcnt[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_01286_),
    .QN(_00729_));
 DFFHQNx3_ASAP7_75t_R \done$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00160_),
    .QN(_00730_));
 DFFHQNx1_ASAP7_75t_R \ld_r$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net195),
    .QN(_00731_));
 DFFHQNx2_ASAP7_75t_R \sa00_sr[0]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00032_),
    .QN(_00732_));
 DFFHQNx2_ASAP7_75t_R \sa00_sr[1]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00033_),
    .QN(_00733_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[2]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00034_),
    .QN(_00734_));
 DFFHQNx2_ASAP7_75t_R \sa00_sr[3]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00035_),
    .QN(_00735_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[4]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00036_),
    .QN(_00736_));
 DFFHQNx2_ASAP7_75t_R \sa00_sr[5]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00037_),
    .QN(_00737_));
 DFFHQNx2_ASAP7_75t_R \sa00_sr[6]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00038_),
    .QN(_00738_));
 DFFHQNx2_ASAP7_75t_R \sa00_sr[7]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00039_),
    .QN(_00739_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[0]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00040_),
    .QN(_00740_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[1]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00041_),
    .QN(_00741_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[2]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00042_),
    .QN(_00742_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[3]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00043_),
    .QN(_00743_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[4]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00044_),
    .QN(_00744_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[5]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00045_),
    .QN(_00745_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[6]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00046_),
    .QN(_00746_));
 DFFHQNx2_ASAP7_75t_R \sa01_sr[7]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00047_),
    .QN(_00747_));
 DFFHQNx2_ASAP7_75t_R \sa02_sr[0]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00048_),
    .QN(_00748_));
 DFFHQNx2_ASAP7_75t_R \sa02_sr[1]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00049_),
    .QN(_00749_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[2]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00050_),
    .QN(_00750_));
 DFFHQNx2_ASAP7_75t_R \sa02_sr[3]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00051_),
    .QN(_00751_));
 DFFHQNx2_ASAP7_75t_R \sa02_sr[4]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00052_),
    .QN(_00752_));
 DFFHQNx2_ASAP7_75t_R \sa02_sr[5]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00053_),
    .QN(_00753_));
 DFFHQNx2_ASAP7_75t_R \sa02_sr[6]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00054_),
    .QN(_00754_));
 DFFHQNx2_ASAP7_75t_R \sa02_sr[7]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00055_),
    .QN(_00755_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[0]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00056_),
    .QN(_00756_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[1]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00057_),
    .QN(_00757_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[2]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00058_),
    .QN(_00758_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[3]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00059_),
    .QN(_00759_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[4]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00060_),
    .QN(_00760_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[5]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00061_),
    .QN(_00761_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[6]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00062_),
    .QN(_00762_));
 DFFHQNx2_ASAP7_75t_R \sa03_sr[7]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00063_),
    .QN(_00763_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[0]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00072_),
    .QN(_00764_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[1]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00073_),
    .QN(_00765_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[2]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00074_),
    .QN(_00766_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[3]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00075_),
    .QN(_00767_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[4]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00076_),
    .QN(_00768_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[5]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00077_),
    .QN(_00769_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[6]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00078_),
    .QN(_00770_));
 DFFHQNx2_ASAP7_75t_R \sa10_sr[7]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00079_),
    .QN(_00771_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[0]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00080_),
    .QN(_00772_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[1]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00081_),
    .QN(_00773_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[2]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00082_),
    .QN(_00774_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[3]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00083_),
    .QN(_00775_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[4]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00084_),
    .QN(_00776_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[5]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00085_),
    .QN(_00777_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[6]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00086_),
    .QN(_00778_));
 DFFHQNx2_ASAP7_75t_R \sa11_sr[7]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00087_),
    .QN(_00779_));
 DFFHQNx2_ASAP7_75t_R \sa12_sr[0]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00088_),
    .QN(_00780_));
 DFFHQNx2_ASAP7_75t_R \sa12_sr[1]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00089_),
    .QN(_00781_));
 DFFHQNx2_ASAP7_75t_R \sa12_sr[2]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00090_),
    .QN(_00782_));
 DFFHQNx2_ASAP7_75t_R \sa12_sr[3]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00091_),
    .QN(_00783_));
 DFFHQNx2_ASAP7_75t_R \sa12_sr[4]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00092_),
    .QN(_00784_));
 DFFHQNx2_ASAP7_75t_R \sa12_sr[5]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00093_),
    .QN(_00785_));
 DFFHQNx2_ASAP7_75t_R \sa12_sr[6]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00094_),
    .QN(_00786_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[7]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00095_),
    .QN(_00787_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[0]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00064_),
    .QN(_00788_));
 DFFHQNx2_ASAP7_75t_R \sa13_sr[1]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00065_),
    .QN(_00789_));
 DFFHQNx2_ASAP7_75t_R \sa13_sr[2]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00066_),
    .QN(_00790_));
 DFFHQNx2_ASAP7_75t_R \sa13_sr[3]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00067_),
    .QN(_00791_));
 DFFHQNx2_ASAP7_75t_R \sa13_sr[4]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00068_),
    .QN(_00792_));
 DFFHQNx2_ASAP7_75t_R \sa13_sr[5]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00069_),
    .QN(_00793_));
 DFFHQNx2_ASAP7_75t_R \sa13_sr[6]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00070_),
    .QN(_00794_));
 DFFHQNx2_ASAP7_75t_R \sa13_sr[7]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00071_),
    .QN(_00795_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[0]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00112_),
    .QN(_00796_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[1]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00113_),
    .QN(_00797_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[2]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00114_),
    .QN(_00798_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[3]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00115_),
    .QN(_00799_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[4]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00116_),
    .QN(_00800_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[5]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00117_),
    .QN(_00801_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[6]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00118_),
    .QN(_00802_));
 DFFHQNx2_ASAP7_75t_R \sa20_sr[7]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00119_),
    .QN(_00803_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[0]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00120_),
    .QN(_00804_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[1]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00121_),
    .QN(_00805_));
 DFFHQNx2_ASAP7_75t_R \sa21_sr[2]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00122_),
    .QN(_00806_));
 DFFHQNx2_ASAP7_75t_R \sa21_sr[3]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00123_),
    .QN(_00807_));
 DFFHQNx2_ASAP7_75t_R \sa21_sr[4]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00124_),
    .QN(_00808_));
 DFFHQNx2_ASAP7_75t_R \sa21_sr[5]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00125_),
    .QN(_00809_));
 DFFHQNx2_ASAP7_75t_R \sa21_sr[6]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00126_),
    .QN(_00810_));
 DFFHQNx2_ASAP7_75t_R \sa21_sr[7]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00127_),
    .QN(_00811_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[0]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00096_),
    .QN(_00812_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[1]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00097_),
    .QN(_00813_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[2]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00098_),
    .QN(_00814_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[3]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00099_),
    .QN(_00815_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[4]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00100_),
    .QN(_00816_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[5]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00101_),
    .QN(_00817_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[6]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00102_),
    .QN(_00818_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[7]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00103_),
    .QN(_00819_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[0]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00104_),
    .QN(_00820_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[1]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00105_),
    .QN(_00821_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00106_),
    .QN(_00822_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[3]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00107_),
    .QN(_00823_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[4]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00108_),
    .QN(_00824_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[5]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00109_),
    .QN(_00825_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[6]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00110_),
    .QN(_00826_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[7]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00111_),
    .QN(_00827_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[0]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00152_),
    .QN(_00828_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[1]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00153_),
    .QN(_00829_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[2]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00154_),
    .QN(_00830_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[3]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00155_),
    .QN(_00831_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[4]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00156_),
    .QN(_00832_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[5]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00157_),
    .QN(_00833_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[6]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00158_),
    .QN(_00834_));
 DFFHQNx2_ASAP7_75t_R \sa30_sr[7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00159_),
    .QN(_00835_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[0]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00128_),
    .QN(_00836_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[1]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00129_),
    .QN(_00837_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[2]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00130_),
    .QN(_00838_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[3]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00131_),
    .QN(_00839_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[4]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00132_),
    .QN(_00840_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[5]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00133_),
    .QN(_00841_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[6]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00134_),
    .QN(_00842_));
 DFFHQNx2_ASAP7_75t_R \sa31_sr[7]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00135_),
    .QN(_00843_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[0]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00136_),
    .QN(_00844_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[1]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00137_),
    .QN(_00845_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[2]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00138_),
    .QN(_00846_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[3]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00139_),
    .QN(_00847_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[4]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00140_),
    .QN(_00848_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[5]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00141_),
    .QN(_00849_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[6]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00142_),
    .QN(_00850_));
 DFFHQNx2_ASAP7_75t_R \sa32_sr[7]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00143_),
    .QN(_00851_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[0]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00144_),
    .QN(_00852_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[1]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00145_),
    .QN(_00853_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[2]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00146_),
    .QN(_00854_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[3]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00147_),
    .QN(_00855_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[4]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00148_),
    .QN(_00856_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[5]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00149_),
    .QN(_00857_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[6]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00150_),
    .QN(_00858_));
 DFFHQNx2_ASAP7_75t_R \sa33_sr[7]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00151_),
    .QN(_00725_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[0]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01287_),
    .QN(_00411_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[100]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01288_),
    .QN(_00724_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[101]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01289_),
    .QN(_00723_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[102]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01290_),
    .QN(_00722_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[103]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01291_),
    .QN(_00721_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[104]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01292_),
    .QN(_00570_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[105]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01293_),
    .QN(_00569_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[106]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01294_),
    .QN(_00572_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[107]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01295_),
    .QN(_00720_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[108]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01296_),
    .QN(_00719_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[109]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01297_),
    .QN(_00718_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[10]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01298_),
    .QN(_00608_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[110]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01299_),
    .QN(_00717_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[111]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01300_),
    .QN(_00716_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[112]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01301_),
    .QN(_00530_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[113]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01302_),
    .QN(_00529_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[114]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01303_),
    .QN(_00532_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[115]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01304_),
    .QN(_00715_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[116]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01305_),
    .QN(_00714_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[117]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01306_),
    .QN(_00713_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[118]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01307_),
    .QN(_00712_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[119]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01308_),
    .QN(_00711_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[11]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01309_),
    .QN(_00710_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[120]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01310_),
    .QN(_00490_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[121]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01311_),
    .QN(_00489_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[122]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01312_),
    .QN(_00492_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[123]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01313_),
    .QN(_00709_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[124]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01314_),
    .QN(_00708_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[125]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01315_),
    .QN(_00707_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[126]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01316_),
    .QN(_00706_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[127]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01317_),
    .QN(_00705_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[12]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01318_),
    .QN(_00704_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[13]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01319_),
    .QN(_00703_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[14]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01320_),
    .QN(_00702_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[15]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01321_),
    .QN(_00701_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[16]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01322_),
    .QN(_00560_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01323_),
    .QN(_00559_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[18]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01324_),
    .QN(_00562_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[19]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01325_),
    .QN(_00700_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01326_),
    .QN(_00410_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[20]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01327_),
    .QN(_00699_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[21]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01328_),
    .QN(_00698_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[22]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01329_),
    .QN(_00697_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[23]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01330_),
    .QN(_00696_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[24]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01331_),
    .QN(_00520_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[25]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01332_),
    .QN(_00519_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[26]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01333_),
    .QN(_00522_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[27]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01334_),
    .QN(_00695_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[28]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01335_),
    .QN(_00694_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[29]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01336_),
    .QN(_00693_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01337_),
    .QN(_00413_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[30]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01338_),
    .QN(_00692_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[31]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01339_),
    .QN(_00691_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[32]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01340_),
    .QN(_00638_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[33]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .D(_01341_),
    .QN(_00637_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[34]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01342_),
    .QN(_00639_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[35]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01343_),
    .QN(_00690_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[36]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01344_),
    .QN(_00689_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[37]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .D(_01345_),
    .QN(_00688_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[38]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01346_),
    .QN(_00687_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[39]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .D(_01347_),
    .QN(_00686_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .D(_01348_),
    .QN(_00685_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[40]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01349_),
    .QN(_00594_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[41]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01350_),
    .QN(_00593_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[42]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01351_),
    .QN(_00596_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[43]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01352_),
    .QN(_00684_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[44]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01353_),
    .QN(_00683_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[45]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01354_),
    .QN(_00682_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[46]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01355_),
    .QN(_00681_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[47]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01356_),
    .QN(_00680_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[48]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01357_),
    .QN(_00550_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[49]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01358_),
    .QN(_00549_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[4]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01359_),
    .QN(_00679_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[50]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01360_),
    .QN(_00552_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[51]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01361_),
    .QN(_00678_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[52]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01362_),
    .QN(_00677_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[53]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01363_),
    .QN(_00676_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[54]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01364_),
    .QN(_00675_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[55]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01365_),
    .QN(_00674_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[56]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01366_),
    .QN(_00510_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[57]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01367_),
    .QN(_00509_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[58]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .D(_01368_),
    .QN(_00512_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[59]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01369_),
    .QN(_00673_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[5]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .D(_01370_),
    .QN(_00672_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[60]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01371_),
    .QN(_00671_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[61]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .D(_01372_),
    .QN(_00670_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[62]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01373_),
    .QN(_00669_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[63]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01374_),
    .QN(_00668_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[64]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01375_),
    .QN(_00628_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[65]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01376_),
    .QN(_00627_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[66]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01377_),
    .QN(_00630_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[67]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01378_),
    .QN(_00667_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[68]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01379_),
    .QN(_00666_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[69]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01380_),
    .QN(_00665_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[6]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01381_),
    .QN(_00664_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[70]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01382_),
    .QN(_00663_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[71]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01383_),
    .QN(_00662_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[72]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01384_),
    .QN(_00582_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[73]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01385_),
    .QN(_00581_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[74]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01386_),
    .QN(_00584_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[75]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01387_),
    .QN(_00661_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[76]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01388_),
    .QN(_00660_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[77]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01389_),
    .QN(_00659_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[78]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01390_),
    .QN(_00658_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[79]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01391_),
    .QN(_00657_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01392_),
    .QN(_00656_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[80]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01393_),
    .QN(_00540_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[81]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01394_),
    .QN(_00539_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[82]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01395_),
    .QN(_00542_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[83]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01396_),
    .QN(_00655_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[84]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01397_),
    .QN(_00654_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[85]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01398_),
    .QN(_00653_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[86]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01399_),
    .QN(_00652_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[87]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01400_),
    .QN(_00651_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[88]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01401_),
    .QN(_00500_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[89]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01402_),
    .QN(_00499_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[8]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01403_),
    .QN(_00606_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[90]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01404_),
    .QN(_00502_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[91]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01405_),
    .QN(_00650_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[92]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01406_),
    .QN(_00649_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[93]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01407_),
    .QN(_00648_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[94]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01408_),
    .QN(_00647_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[95]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01409_),
    .QN(_00646_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[96]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01410_),
    .QN(_00618_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[97]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01411_),
    .QN(_00617_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[98]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01412_),
    .QN(_00620_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[99]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01413_),
    .QN(_00645_));
 DFFHQNx2_ASAP7_75t_R \text_in_r[9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01414_),
    .QN(_00605_));
 DFFHQNx2_ASAP7_75t_R \text_out[0]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00265_),
    .QN(_00859_));
 DFFHQNx2_ASAP7_75t_R \text_out[100]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00165_),
    .QN(_00860_));
 DFFHQNx2_ASAP7_75t_R \text_out[101]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00166_),
    .QN(_00861_));
 DFFHQNx2_ASAP7_75t_R \text_out[102]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00167_),
    .QN(_00862_));
 DFFHQNx2_ASAP7_75t_R \text_out[103]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00168_),
    .QN(_00863_));
 DFFHQNx2_ASAP7_75t_R \text_out[104]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00169_),
    .QN(_00864_));
 DFFHQNx3_ASAP7_75t_R \text_out[105]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00170_),
    .QN(_00865_));
 DFFHQNx2_ASAP7_75t_R \text_out[106]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00171_),
    .QN(_00866_));
 DFFHQNx2_ASAP7_75t_R \text_out[107]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00172_),
    .QN(_00867_));
 DFFHQNx2_ASAP7_75t_R \text_out[108]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00173_),
    .QN(_00868_));
 DFFHQNx3_ASAP7_75t_R \text_out[109]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00174_),
    .QN(_00869_));
 DFFHQNx2_ASAP7_75t_R \text_out[10]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00195_),
    .QN(_00870_));
 DFFHQNx3_ASAP7_75t_R \text_out[110]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00175_),
    .QN(_00871_));
 DFFHQNx3_ASAP7_75t_R \text_out[111]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00176_),
    .QN(_00872_));
 DFFHQNx3_ASAP7_75t_R \text_out[112]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00177_),
    .QN(_00873_));
 DFFHQNx3_ASAP7_75t_R \text_out[113]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00178_),
    .QN(_00874_));
 DFFHQNx3_ASAP7_75t_R \text_out[114]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00179_),
    .QN(_00875_));
 DFFHQNx3_ASAP7_75t_R \text_out[115]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00180_),
    .QN(_00876_));
 DFFHQNx3_ASAP7_75t_R \text_out[116]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00181_),
    .QN(_00877_));
 DFFHQNx3_ASAP7_75t_R \text_out[117]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00182_),
    .QN(_00878_));
 DFFHQNx3_ASAP7_75t_R \text_out[118]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00183_),
    .QN(_00879_));
 DFFHQNx3_ASAP7_75t_R \text_out[119]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00184_),
    .QN(_00880_));
 DFFHQNx2_ASAP7_75t_R \text_out[11]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00196_),
    .QN(_00881_));
 DFFHQNx3_ASAP7_75t_R \text_out[120]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00185_),
    .QN(_00882_));
 DFFHQNx3_ASAP7_75t_R \text_out[121]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00186_),
    .QN(_00883_));
 DFFHQNx3_ASAP7_75t_R \text_out[122]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00187_),
    .QN(_00884_));
 DFFHQNx3_ASAP7_75t_R \text_out[123]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00188_),
    .QN(_00885_));
 DFFHQNx3_ASAP7_75t_R \text_out[124]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00189_),
    .QN(_00886_));
 DFFHQNx2_ASAP7_75t_R \text_out[125]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00190_),
    .QN(_00887_));
 DFFHQNx2_ASAP7_75t_R \text_out[126]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00191_),
    .QN(_00888_));
 DFFHQNx2_ASAP7_75t_R \text_out[127]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00192_),
    .QN(_00889_));
 DFFHQNx2_ASAP7_75t_R \text_out[12]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00197_),
    .QN(_00890_));
 DFFHQNx3_ASAP7_75t_R \text_out[13]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00198_),
    .QN(_00891_));
 DFFHQNx3_ASAP7_75t_R \text_out[14]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00199_),
    .QN(_00892_));
 DFFHQNx2_ASAP7_75t_R \text_out[15]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00200_),
    .QN(_00893_));
 DFFHQNx2_ASAP7_75t_R \text_out[16]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00201_),
    .QN(_00894_));
 DFFHQNx3_ASAP7_75t_R \text_out[17]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00202_),
    .QN(_00895_));
 DFFHQNx3_ASAP7_75t_R \text_out[18]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00203_),
    .QN(_00896_));
 DFFHQNx3_ASAP7_75t_R \text_out[19]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00204_),
    .QN(_00897_));
 DFFHQNx2_ASAP7_75t_R \text_out[1]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00266_),
    .QN(_00898_));
 DFFHQNx3_ASAP7_75t_R \text_out[20]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00205_),
    .QN(_00899_));
 DFFHQNx2_ASAP7_75t_R \text_out[21]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00206_),
    .QN(_00900_));
 DFFHQNx2_ASAP7_75t_R \text_out[22]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00207_),
    .QN(_00901_));
 DFFHQNx3_ASAP7_75t_R \text_out[23]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00208_),
    .QN(_00902_));
 DFFHQNx2_ASAP7_75t_R \text_out[24]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00209_),
    .QN(_00903_));
 DFFHQNx3_ASAP7_75t_R \text_out[25]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00210_),
    .QN(_00904_));
 DFFHQNx2_ASAP7_75t_R \text_out[26]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00211_),
    .QN(_00905_));
 DFFHQNx2_ASAP7_75t_R \text_out[27]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00212_),
    .QN(_00906_));
 DFFHQNx2_ASAP7_75t_R \text_out[28]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00213_),
    .QN(_00907_));
 DFFHQNx3_ASAP7_75t_R \text_out[29]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00214_),
    .QN(_00908_));
 DFFHQNx3_ASAP7_75t_R \text_out[2]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00267_),
    .QN(_00909_));
 DFFHQNx3_ASAP7_75t_R \text_out[30]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00215_),
    .QN(_00910_));
 DFFHQNx2_ASAP7_75t_R \text_out[31]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00216_),
    .QN(_00911_));
 DFFHQNx3_ASAP7_75t_R \text_out[32]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00217_),
    .QN(_00912_));
 DFFHQNx3_ASAP7_75t_R \text_out[33]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00218_),
    .QN(_00913_));
 DFFHQNx3_ASAP7_75t_R \text_out[34]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00219_),
    .QN(_00914_));
 DFFHQNx3_ASAP7_75t_R \text_out[35]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00220_),
    .QN(_00915_));
 DFFHQNx3_ASAP7_75t_R \text_out[36]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00221_),
    .QN(_00916_));
 DFFHQNx3_ASAP7_75t_R \text_out[37]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00222_),
    .QN(_00917_));
 DFFHQNx3_ASAP7_75t_R \text_out[38]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00223_),
    .QN(_00918_));
 DFFHQNx3_ASAP7_75t_R \text_out[39]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00224_),
    .QN(_00919_));
 DFFHQNx2_ASAP7_75t_R \text_out[3]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00268_),
    .QN(_00920_));
 DFFHQNx2_ASAP7_75t_R \text_out[40]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00225_),
    .QN(_00921_));
 DFFHQNx2_ASAP7_75t_R \text_out[41]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00226_),
    .QN(_00922_));
 DFFHQNx3_ASAP7_75t_R \text_out[42]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00227_),
    .QN(_00923_));
 DFFHQNx2_ASAP7_75t_R \text_out[43]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00228_),
    .QN(_00924_));
 DFFHQNx2_ASAP7_75t_R \text_out[44]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00229_),
    .QN(_00925_));
 DFFHQNx2_ASAP7_75t_R \text_out[45]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00230_),
    .QN(_00926_));
 DFFHQNx2_ASAP7_75t_R \text_out[46]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00231_),
    .QN(_00927_));
 DFFHQNx2_ASAP7_75t_R \text_out[47]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00232_),
    .QN(_00928_));
 DFFHQNx2_ASAP7_75t_R \text_out[48]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00233_),
    .QN(_00929_));
 DFFHQNx2_ASAP7_75t_R \text_out[49]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00234_),
    .QN(_00930_));
 DFFHQNx2_ASAP7_75t_R \text_out[4]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00269_),
    .QN(_00931_));
 DFFHQNx2_ASAP7_75t_R \text_out[50]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00235_),
    .QN(_00932_));
 DFFHQNx3_ASAP7_75t_R \text_out[51]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00236_),
    .QN(_00933_));
 DFFHQNx2_ASAP7_75t_R \text_out[52]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00237_),
    .QN(_00934_));
 DFFHQNx3_ASAP7_75t_R \text_out[53]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00238_),
    .QN(_00935_));
 DFFHQNx3_ASAP7_75t_R \text_out[54]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00239_),
    .QN(_00936_));
 DFFHQNx2_ASAP7_75t_R \text_out[55]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00240_),
    .QN(_00937_));
 DFFHQNx2_ASAP7_75t_R \text_out[56]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00241_),
    .QN(_00938_));
 DFFHQNx3_ASAP7_75t_R \text_out[57]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00242_),
    .QN(_00939_));
 DFFHQNx3_ASAP7_75t_R \text_out[58]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00243_),
    .QN(_00940_));
 DFFHQNx3_ASAP7_75t_R \text_out[59]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00244_),
    .QN(_00941_));
 DFFHQNx3_ASAP7_75t_R \text_out[5]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00270_),
    .QN(_00942_));
 DFFHQNx3_ASAP7_75t_R \text_out[60]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00245_),
    .QN(_00943_));
 DFFHQNx3_ASAP7_75t_R \text_out[61]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00246_),
    .QN(_00944_));
 DFFHQNx3_ASAP7_75t_R \text_out[62]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00247_),
    .QN(_00945_));
 DFFHQNx2_ASAP7_75t_R \text_out[63]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00248_),
    .QN(_00946_));
 DFFHQNx2_ASAP7_75t_R \text_out[64]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00249_),
    .QN(_00947_));
 DFFHQNx3_ASAP7_75t_R \text_out[65]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00250_),
    .QN(_00948_));
 DFFHQNx2_ASAP7_75t_R \text_out[66]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00251_),
    .QN(_00949_));
 DFFHQNx2_ASAP7_75t_R \text_out[67]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00252_),
    .QN(_00950_));
 DFFHQNx3_ASAP7_75t_R \text_out[68]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00253_),
    .QN(_00951_));
 DFFHQNx2_ASAP7_75t_R \text_out[69]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00254_),
    .QN(_00952_));
 DFFHQNx2_ASAP7_75t_R \text_out[6]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00271_),
    .QN(_00953_));
 DFFHQNx3_ASAP7_75t_R \text_out[70]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00255_),
    .QN(_00954_));
 DFFHQNx3_ASAP7_75t_R \text_out[71]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00256_),
    .QN(_00955_));
 DFFHQNx2_ASAP7_75t_R \text_out[72]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00257_),
    .QN(_00956_));
 DFFHQNx2_ASAP7_75t_R \text_out[73]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00258_),
    .QN(_00957_));
 DFFHQNx2_ASAP7_75t_R \text_out[74]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00259_),
    .QN(_00958_));
 DFFHQNx3_ASAP7_75t_R \text_out[75]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00260_),
    .QN(_00959_));
 DFFHQNx2_ASAP7_75t_R \text_out[76]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00261_),
    .QN(_00960_));
 DFFHQNx2_ASAP7_75t_R \text_out[77]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00262_),
    .QN(_00961_));
 DFFHQNx3_ASAP7_75t_R \text_out[78]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00263_),
    .QN(_00962_));
 DFFHQNx2_ASAP7_75t_R \text_out[79]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00264_),
    .QN(_00963_));
 DFFHQNx2_ASAP7_75t_R \text_out[7]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00272_),
    .QN(_00964_));
 DFFHQNx2_ASAP7_75t_R \text_out[80]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00273_),
    .QN(_00965_));
 DFFHQNx2_ASAP7_75t_R \text_out[81]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00274_),
    .QN(_00966_));
 DFFHQNx2_ASAP7_75t_R \text_out[82]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00275_),
    .QN(_00967_));
 DFFHQNx3_ASAP7_75t_R \text_out[83]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00276_),
    .QN(_00968_));
 DFFHQNx3_ASAP7_75t_R \text_out[84]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00277_),
    .QN(_00969_));
 DFFHQNx2_ASAP7_75t_R \text_out[85]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00278_),
    .QN(_00970_));
 DFFHQNx2_ASAP7_75t_R \text_out[86]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00279_),
    .QN(_00971_));
 DFFHQNx2_ASAP7_75t_R \text_out[87]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00280_),
    .QN(_00972_));
 DFFHQNx2_ASAP7_75t_R \text_out[88]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00281_),
    .QN(_00973_));
 DFFHQNx2_ASAP7_75t_R \text_out[89]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00282_),
    .QN(_00974_));
 DFFHQNx2_ASAP7_75t_R \text_out[8]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00193_),
    .QN(_00975_));
 DFFHQNx2_ASAP7_75t_R \text_out[90]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00283_),
    .QN(_00976_));
 DFFHQNx3_ASAP7_75t_R \text_out[91]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00284_),
    .QN(_00977_));
 DFFHQNx2_ASAP7_75t_R \text_out[92]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00285_),
    .QN(_00978_));
 DFFHQNx2_ASAP7_75t_R \text_out[93]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00286_),
    .QN(_00979_));
 DFFHQNx3_ASAP7_75t_R \text_out[94]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00287_),
    .QN(_00980_));
 DFFHQNx2_ASAP7_75t_R \text_out[95]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00288_),
    .QN(_00981_));
 DFFHQNx2_ASAP7_75t_R \text_out[96]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00161_),
    .QN(_00982_));
 DFFHQNx2_ASAP7_75t_R \text_out[97]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00162_),
    .QN(_00983_));
 DFFHQNx3_ASAP7_75t_R \text_out[98]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00163_),
    .QN(_00984_));
 DFFHQNx2_ASAP7_75t_R \text_out[99]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00164_),
    .QN(_00985_));
 DFFHQNx2_ASAP7_75t_R \text_out[9]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00194_),
    .QN(_00644_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[24]$_SDFF_PP1_  (.CLK(clknet_leaf_31_clk),
    .D(_01415_),
    .QN(_00446_));
 DFFHQNx2_ASAP7_75t_R \u0.r0.out[25]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_01416_),
    .QN(_00447_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[26]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01417_),
    .QN(_00448_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[27]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01418_),
    .QN(_00449_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[28]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .D(_01419_),
    .QN(_00450_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[29]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01420_),
    .QN(_00451_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[30]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_01421_),
    .QN(_00452_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[31]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_01422_),
    .QN(_00453_));
 DFFHQNx2_ASAP7_75t_R \u0.r0.rcnt[0]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_01423_),
    .QN(\u0.r0.rcnt_next[0] ));
 DFFHQNx2_ASAP7_75t_R \u0.r0.rcnt[1]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_01424_),
    .QN(_16081_));
 DFFHQNx2_ASAP7_75t_R \u0.r0.rcnt[2]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_01425_),
    .QN(_00643_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.rcnt[3]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_01426_),
    .QN(_00986_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[0]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00000_),
    .QN(_00987_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[1]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00001_),
    .QN(_00988_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[2]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00002_),
    .QN(_00989_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[3]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00003_),
    .QN(_00990_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[4]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00004_),
    .QN(_00991_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[5]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00005_),
    .QN(_00992_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[6]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00006_),
    .QN(_00993_));
 DFFHQNx2_ASAP7_75t_R \u0.u0.d[7]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00007_),
    .QN(_00994_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[0]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00008_),
    .QN(_00439_));
 DFFHQNx2_ASAP7_75t_R \u0.u1.d[1]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00009_),
    .QN(_00440_));
 DFFHQNx2_ASAP7_75t_R \u0.u1.d[2]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00010_),
    .QN(_00416_));
 DFFHQNx2_ASAP7_75t_R \u0.u1.d[3]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00011_),
    .QN(_00441_));
 DFFHQNx2_ASAP7_75t_R \u0.u1.d[4]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00012_),
    .QN(_00442_));
 DFFHQNx2_ASAP7_75t_R \u0.u1.d[5]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00013_),
    .QN(_00443_));
 DFFHQNx2_ASAP7_75t_R \u0.u1.d[6]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00014_),
    .QN(_00444_));
 DFFHQNx2_ASAP7_75t_R \u0.u1.d[7]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00015_),
    .QN(_00445_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[0]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00016_),
    .QN(_00432_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[1]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00017_),
    .QN(_00433_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00018_),
    .QN(_00424_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00019_),
    .QN(_00434_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[4]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00020_),
    .QN(_00435_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[5]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00021_),
    .QN(_00436_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[6]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00022_),
    .QN(_00437_));
 DFFHQNx2_ASAP7_75t_R \u0.u2.d[7]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00023_),
    .QN(_00438_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[0]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00024_),
    .QN(_00425_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[1]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00025_),
    .QN(_00426_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[2]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00026_),
    .QN(_00423_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[3]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00027_),
    .QN(_00427_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[4]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00028_),
    .QN(_00428_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[5]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00029_),
    .QN(_00429_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[6]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00030_),
    .QN(_00430_));
 DFFHQNx2_ASAP7_75t_R \u0.u3.d[7]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00031_),
    .QN(_00431_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][0]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00289_),
    .QN(_00995_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][10]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00290_),
    .QN(_00996_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][11]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00291_),
    .QN(_00997_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][12]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00292_),
    .QN(_00998_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][13]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00293_),
    .QN(_00999_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][14]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00294_),
    .QN(_01000_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][15]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00295_),
    .QN(_01001_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][16]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00296_),
    .QN(_01002_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][17]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00297_),
    .QN(_01003_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][18]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00298_),
    .QN(_01004_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][19]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00299_),
    .QN(_01005_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][1]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00300_),
    .QN(_01006_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][20]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00301_),
    .QN(_01007_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][21]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00302_),
    .QN(_01008_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][22]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00303_),
    .QN(_01009_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][23]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00304_),
    .QN(_01010_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][24]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00305_),
    .QN(_01011_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][25]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00306_),
    .QN(_01012_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][26]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00307_),
    .QN(_01013_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][27]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00308_),
    .QN(_01014_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][28]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00309_),
    .QN(_01015_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][29]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00310_),
    .QN(_01016_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][2]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00311_),
    .QN(_01017_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][30]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00312_),
    .QN(_01018_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][31]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00313_),
    .QN(_01019_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][3]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00314_),
    .QN(_01020_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][4]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00315_),
    .QN(_01021_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][5]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00316_),
    .QN(_01022_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][6]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00317_),
    .QN(_01023_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00318_),
    .QN(_01024_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][8]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00319_),
    .QN(_01025_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][9]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00320_),
    .QN(_01026_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][0]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00321_),
    .QN(_01027_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][10]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00322_),
    .QN(_01028_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][11]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00323_),
    .QN(_01029_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][12]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00324_),
    .QN(_01030_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][13]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00325_),
    .QN(_01031_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][14]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00326_),
    .QN(_01032_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][15]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00327_),
    .QN(_01033_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][16]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00328_),
    .QN(_01034_));
 DFFHQNx3_ASAP7_75t_R \u0.w[1][17]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00329_),
    .QN(_01035_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][18]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00330_),
    .QN(_01036_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][19]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00331_),
    .QN(_01037_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][1]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00332_),
    .QN(_01038_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][20]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00333_),
    .QN(_01039_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][21]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00334_),
    .QN(_01040_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][22]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00335_),
    .QN(_01041_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][23]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00336_),
    .QN(_01042_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][24]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00337_),
    .QN(_01043_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][25]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00338_),
    .QN(_01044_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][26]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00339_),
    .QN(_01045_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][27]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00340_),
    .QN(_01046_));
 DFFHQNx3_ASAP7_75t_R \u0.w[1][28]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00341_),
    .QN(_01047_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][29]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00342_),
    .QN(_01048_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00343_),
    .QN(_01049_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][30]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00344_),
    .QN(_01050_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][31]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00345_),
    .QN(_01051_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][3]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00346_),
    .QN(_01052_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][4]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00347_),
    .QN(_01053_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][5]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00348_),
    .QN(_01054_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][6]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00349_),
    .QN(_01055_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00350_),
    .QN(_01056_));
 DFFHQNx2_ASAP7_75t_R \u0.w[1][8]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00351_),
    .QN(_01057_));
 DFFHQNx3_ASAP7_75t_R \u0.w[1][9]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00352_),
    .QN(_01058_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][0]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00353_),
    .QN(_01059_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][10]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00354_),
    .QN(_01060_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][11]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00355_),
    .QN(_01061_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][12]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00356_),
    .QN(_01062_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][13]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00357_),
    .QN(_01063_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][14]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00358_),
    .QN(_01064_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][15]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00359_),
    .QN(_01065_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][16]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00360_),
    .QN(_01066_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][17]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00361_),
    .QN(_01067_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][18]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00362_),
    .QN(_01068_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][19]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00363_),
    .QN(_01069_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][1]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00364_),
    .QN(_01070_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][20]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00365_),
    .QN(_01071_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][21]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00366_),
    .QN(_01072_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][22]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00367_),
    .QN(_01073_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][23]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00368_),
    .QN(_01074_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][24]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00369_),
    .QN(_01075_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][25]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00370_),
    .QN(_01076_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][26]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00371_),
    .QN(_01077_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][27]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00372_),
    .QN(_01078_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][28]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00373_),
    .QN(_01079_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][29]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00374_),
    .QN(_01080_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][2]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00375_),
    .QN(_01081_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][30]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00376_),
    .QN(_01082_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][31]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00377_),
    .QN(_01083_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][3]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00378_),
    .QN(_01084_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][4]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00379_),
    .QN(_01085_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][5]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00380_),
    .QN(_01086_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][6]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00381_),
    .QN(_01087_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][7]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00382_),
    .QN(_01088_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][8]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00383_),
    .QN(_01089_));
 DFFHQNx2_ASAP7_75t_R \u0.w[2][9]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00384_),
    .QN(_01090_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][0]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(net16),
    .QN(_01091_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][10]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_15760_),
    .QN(_01092_));
 DFFHQNx3_ASAP7_75t_R \u0.w[3][11]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00385_),
    .QN(_01093_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][12]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00386_),
    .QN(_01094_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][13]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00387_),
    .QN(_01095_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][14]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00388_),
    .QN(_01096_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][15]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00389_),
    .QN(_01097_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][16]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_15730_),
    .QN(_01098_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][17]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_15729_),
    .QN(_01099_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][18]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_15742_),
    .QN(_01100_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][19]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00390_),
    .QN(_01101_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][1]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(net2),
    .QN(_01102_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][20]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00391_),
    .QN(_01103_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][21]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00392_),
    .QN(_01104_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][22]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00393_),
    .QN(_01105_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][23]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00394_),
    .QN(_01106_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][24]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_15784_),
    .QN(_01107_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][25]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(net18),
    .QN(_01108_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][26]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_15794_),
    .QN(_01109_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][27]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00395_),
    .QN(_01110_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][28]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00396_),
    .QN(_01111_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][29]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00397_),
    .QN(_01112_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][2]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_15778_),
    .QN(_01113_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][30]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00398_),
    .QN(_01114_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][31]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00399_),
    .QN(_01115_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][3]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00400_),
    .QN(_01116_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][4]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00401_),
    .QN(_01117_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][5]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00402_),
    .QN(_01118_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][6]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00403_),
    .QN(_01119_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][7]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00404_),
    .QN(_01120_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][8]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_15748_),
    .QN(_01121_));
 DFFHQNx2_ASAP7_75t_R \u0.w[3][9]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_15747_),
    .QN(_00642_));
 NOR2x2_ASAP7_75t_R clone1 (.A(net486),
    .B(_10727_),
    .Y(net1));
 NOR2x2_ASAP7_75t_R clone2 (.A(_08030_),
    .B(_08022_),
    .Y(net2));
 NAND2x2_ASAP7_75t_R clone3 (.A(net728),
    .B(net782),
    .Y(net3));
 NAND2x2_ASAP7_75t_R clone4 (.A(net686),
    .B(net896),
    .Y(net4));
 OAI21x1_ASAP7_75t_R clone5 (.A1(_15090_),
    .A2(_15091_),
    .B(_15189_),
    .Y(net5));
 OAI21x1_ASAP7_75t_R clone6 (.A1(_13641_),
    .A2(_13642_),
    .B(_13706_),
    .Y(net6));
 NAND2x2_ASAP7_75t_R clone7 (.A(net775),
    .B(net773),
    .Y(net7));
 AOI21x1_ASAP7_75t_R clone8 (.A1(_04385_),
    .A2(_04384_),
    .B(_04488_),
    .Y(net8));
 BUFx6f_ASAP7_75t_R clone9 (.A(net568),
    .Y(net9));
 BUFx4f_ASAP7_75t_R clone10 (.A(_12338_),
    .Y(net10));
 NAND2x2_ASAP7_75t_R clone11 (.A(net825),
    .B(_08183_),
    .Y(net11));
 BUFx6f_ASAP7_75t_R clone13 (.A(_08021_),
    .Y(net13));
 BUFx6f_ASAP7_75t_R clone14 (.A(_07939_),
    .Y(net14));
 BUFx2_ASAP7_75t_R clone15 (.A(_09516_),
    .Y(net15));
 INVx4_ASAP7_75t_R clone16 (.A(_15768_),
    .Y(net16));
 NOR2x2_ASAP7_75t_R clone17 (.A(_08030_),
    .B(_08022_),
    .Y(net17));
 INVx4_ASAP7_75t_R clone18 (.A(net492),
    .Y(net18));
 BUFx2_ASAP7_75t_R clone19 (.A(_00740_),
    .Y(net19));
 BUFx6f_ASAP7_75t_R clone20 (.A(net618),
    .Y(net20));
 BUFx4f_ASAP7_75t_R clone21 (.A(_06441_),
    .Y(net21));
 BUFx6f_ASAP7_75t_R clone22 (.A(_06570_),
    .Y(net22));
 BUFx4_ASAP7_75t_R clone23 (.A(net808),
    .Y(net23));
 BUFx4f_ASAP7_75t_R clone24 (.A(_10838_),
    .Y(net24));
 BUFx3_ASAP7_75t_R clone25 (.A(net602),
    .Y(net25));
 BUFx6f_ASAP7_75t_R clone26 (.A(_06475_),
    .Y(net26));
 BUFx6f_ASAP7_75t_R clone27 (.A(_02942_),
    .Y(net27));
 BUFx4f_ASAP7_75t_R clone28 (.A(net697),
    .Y(net28));
 BUFx6f_ASAP7_75t_R clone29 (.A(_05823_),
    .Y(net29));
 BUFx3_ASAP7_75t_R clone30 (.A(net522),
    .Y(net30));
 OAI21x1_ASAP7_75t_R clone32 (.A1(_02968_),
    .A2(_02969_),
    .B(_03005_),
    .Y(net32));
 OAI21x1_ASAP7_75t_R clone33 (.A1(_02972_),
    .A2(_02963_),
    .B(_03005_),
    .Y(net33));
 BUFx6f_ASAP7_75t_R clone34 (.A(_12944_),
    .Y(net34));
 BUFx3_ASAP7_75t_R clone35 (.A(_00756_),
    .Y(net35));
 INVx5_ASAP7_75t_R clone36 (.A(net605),
    .Y(net36));
 BUFx2_ASAP7_75t_R clone37 (.A(_04496_),
    .Y(net37));
 BUFx3_ASAP7_75t_R clone38 (.A(_00748_),
    .Y(net38));
 XOR2x2_ASAP7_75t_R clone39 (.A(_15139_),
    .B(_15038_),
    .Y(net39));
 BUFx4f_ASAP7_75t_R clone40 (.A(net778),
    .Y(net40));
 BUFx4f_ASAP7_75t_R clone41 (.A(net564),
    .Y(net41));
 BUFx6f_ASAP7_75t_R clone43 (.A(_05081_),
    .Y(net43));
 BUFx4f_ASAP7_75t_R clone44 (.A(_05057_),
    .Y(net44));
 BUFx6f_ASAP7_75t_R clone46 (.A(net832),
    .Y(net46));
 NAND2x2_ASAP7_75t_R clone48 (.A(_04426_),
    .B(_04425_),
    .Y(net48));
 BUFx3_ASAP7_75t_R clone49 (.A(_00764_),
    .Y(net49));
 BUFx3_ASAP7_75t_R clone50 (.A(_00739_),
    .Y(net50));
 BUFx3_ASAP7_75t_R clone52 (.A(_00733_),
    .Y(net52));
 BUFx4f_ASAP7_75t_R clone53 (.A(_12148_),
    .Y(net53));
 OAI21x1_ASAP7_75t_R clone54 (.A1(_14356_),
    .A2(_14365_),
    .B(net465),
    .Y(net54));
 OAI21x1_ASAP7_75t_R clone55 (.A1(_14356_),
    .A2(_14365_),
    .B(_14499_),
    .Y(net55));
 BUFx6f_ASAP7_75t_R clone56 (.A(net693),
    .Y(net56));
 BUFx4f_ASAP7_75t_R clone57 (.A(net549),
    .Y(net57));
 BUFx3_ASAP7_75t_R clone58 (.A(_00803_),
    .Y(net58));
 BUFx3_ASAP7_75t_R clone59 (.A(_00749_),
    .Y(net59));
 BUFx3_ASAP7_75t_R clone60 (.A(net62),
    .Y(net60));
 BUFx6f_ASAP7_75t_R clone61 (.A(_13704_),
    .Y(net61));
 NAND2x2_ASAP7_75t_R clone62 (.A(_13638_),
    .B(net818),
    .Y(net62));
 XOR2x2_ASAP7_75t_R clone63 (.A(_13703_),
    .B(net817),
    .Y(net63));
 BUFx4f_ASAP7_75t_R clone65 (.A(net783),
    .Y(net65));
 AOI21x1_ASAP7_75t_R clone66 (.A1(_12886_),
    .A2(_12888_),
    .B(net455),
    .Y(net66));
 BUFx3_ASAP7_75t_R clone67 (.A(_13707_),
    .Y(net67));
 XOR2x2_ASAP7_75t_R clone69 (.A(net816),
    .B(_07969_),
    .Y(net69));
 BUFx6f_ASAP7_75t_R clone70 (.A(net875),
    .Y(net70));
 BUFx4f_ASAP7_75t_R clone71 (.A(net533),
    .Y(net71));
 BUFx3_ASAP7_75t_R clone72 (.A(_00795_),
    .Y(net72));
 BUFx2_ASAP7_75t_R clone73 (.A(_02306_),
    .Y(net73));
 NAND2x2_ASAP7_75t_R clone74 (.A(_07109_),
    .B(_07102_),
    .Y(net74));
 BUFx2_ASAP7_75t_R input1 (.A(key[0]),
    .Y(net12));
 BUFx2_ASAP7_75t_R input2 (.A(key[100]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input3 (.A(key[101]),
    .Y(net42));
 BUFx2_ASAP7_75t_R input4 (.A(key[102]),
    .Y(net45));
 BUFx2_ASAP7_75t_R input5 (.A(key[103]),
    .Y(net47));
 BUFx2_ASAP7_75t_R input6 (.A(key[104]),
    .Y(net51));
 BUFx2_ASAP7_75t_R input7 (.A(key[105]),
    .Y(net64));
 BUFx2_ASAP7_75t_R input8 (.A(key[106]),
    .Y(net68));
 BUFx2_ASAP7_75t_R input9 (.A(key[107]),
    .Y(net75));
 BUFx2_ASAP7_75t_R input10 (.A(key[108]),
    .Y(net76));
 BUFx2_ASAP7_75t_R input11 (.A(key[109]),
    .Y(net77));
 BUFx2_ASAP7_75t_R input12 (.A(key[10]),
    .Y(net78));
 BUFx2_ASAP7_75t_R input13 (.A(key[110]),
    .Y(net79));
 BUFx2_ASAP7_75t_R input14 (.A(key[111]),
    .Y(net80));
 BUFx2_ASAP7_75t_R input15 (.A(key[112]),
    .Y(net81));
 BUFx2_ASAP7_75t_R input16 (.A(key[113]),
    .Y(net82));
 BUFx2_ASAP7_75t_R input17 (.A(key[114]),
    .Y(net83));
 BUFx2_ASAP7_75t_R input18 (.A(key[115]),
    .Y(net84));
 BUFx2_ASAP7_75t_R input19 (.A(key[116]),
    .Y(net85));
 BUFx2_ASAP7_75t_R input20 (.A(key[117]),
    .Y(net86));
 BUFx2_ASAP7_75t_R input21 (.A(key[118]),
    .Y(net87));
 BUFx2_ASAP7_75t_R input22 (.A(key[119]),
    .Y(net88));
 BUFx2_ASAP7_75t_R input23 (.A(key[11]),
    .Y(net89));
 BUFx2_ASAP7_75t_R input24 (.A(key[120]),
    .Y(net90));
 BUFx2_ASAP7_75t_R input25 (.A(key[121]),
    .Y(net91));
 BUFx2_ASAP7_75t_R input26 (.A(key[122]),
    .Y(net92));
 BUFx2_ASAP7_75t_R input27 (.A(key[123]),
    .Y(net93));
 BUFx2_ASAP7_75t_R input28 (.A(key[124]),
    .Y(net94));
 BUFx2_ASAP7_75t_R input29 (.A(key[125]),
    .Y(net95));
 BUFx2_ASAP7_75t_R input30 (.A(key[126]),
    .Y(net96));
 BUFx2_ASAP7_75t_R input31 (.A(key[127]),
    .Y(net97));
 BUFx2_ASAP7_75t_R input32 (.A(key[12]),
    .Y(net98));
 BUFx2_ASAP7_75t_R input33 (.A(key[13]),
    .Y(net99));
 BUFx2_ASAP7_75t_R input34 (.A(key[14]),
    .Y(net100));
 BUFx2_ASAP7_75t_R input35 (.A(key[15]),
    .Y(net101));
 BUFx2_ASAP7_75t_R input36 (.A(key[16]),
    .Y(net102));
 BUFx2_ASAP7_75t_R input37 (.A(key[17]),
    .Y(net103));
 BUFx2_ASAP7_75t_R input38 (.A(key[18]),
    .Y(net104));
 BUFx2_ASAP7_75t_R input39 (.A(key[19]),
    .Y(net105));
 BUFx2_ASAP7_75t_R input40 (.A(key[1]),
    .Y(net106));
 BUFx2_ASAP7_75t_R input41 (.A(key[20]),
    .Y(net107));
 BUFx2_ASAP7_75t_R input42 (.A(key[21]),
    .Y(net108));
 BUFx2_ASAP7_75t_R input43 (.A(key[22]),
    .Y(net109));
 BUFx2_ASAP7_75t_R input44 (.A(key[23]),
    .Y(net110));
 BUFx3_ASAP7_75t_R input45 (.A(key[24]),
    .Y(net111));
 BUFx2_ASAP7_75t_R input46 (.A(key[25]),
    .Y(net112));
 BUFx2_ASAP7_75t_R input47 (.A(key[26]),
    .Y(net113));
 BUFx2_ASAP7_75t_R input48 (.A(key[27]),
    .Y(net114));
 BUFx2_ASAP7_75t_R input49 (.A(key[28]),
    .Y(net115));
 BUFx2_ASAP7_75t_R input50 (.A(key[29]),
    .Y(net116));
 BUFx2_ASAP7_75t_R input51 (.A(key[2]),
    .Y(net117));
 BUFx2_ASAP7_75t_R input52 (.A(key[30]),
    .Y(net118));
 BUFx2_ASAP7_75t_R input53 (.A(key[31]),
    .Y(net119));
 BUFx2_ASAP7_75t_R input54 (.A(key[32]),
    .Y(net120));
 BUFx2_ASAP7_75t_R input55 (.A(key[33]),
    .Y(net121));
 BUFx2_ASAP7_75t_R input56 (.A(key[34]),
    .Y(net122));
 BUFx2_ASAP7_75t_R input57 (.A(key[35]),
    .Y(net123));
 BUFx2_ASAP7_75t_R input58 (.A(key[36]),
    .Y(net124));
 BUFx2_ASAP7_75t_R input59 (.A(key[37]),
    .Y(net125));
 BUFx2_ASAP7_75t_R input60 (.A(key[38]),
    .Y(net126));
 BUFx2_ASAP7_75t_R input61 (.A(key[39]),
    .Y(net127));
 BUFx2_ASAP7_75t_R input62 (.A(key[3]),
    .Y(net128));
 BUFx2_ASAP7_75t_R input63 (.A(key[40]),
    .Y(net129));
 BUFx2_ASAP7_75t_R input64 (.A(key[41]),
    .Y(net130));
 BUFx2_ASAP7_75t_R input65 (.A(key[42]),
    .Y(net131));
 BUFx2_ASAP7_75t_R input66 (.A(key[43]),
    .Y(net132));
 BUFx2_ASAP7_75t_R input67 (.A(key[44]),
    .Y(net133));
 BUFx2_ASAP7_75t_R input68 (.A(key[45]),
    .Y(net134));
 BUFx2_ASAP7_75t_R input69 (.A(key[46]),
    .Y(net135));
 BUFx2_ASAP7_75t_R input70 (.A(key[47]),
    .Y(net136));
 BUFx2_ASAP7_75t_R input71 (.A(key[48]),
    .Y(net137));
 BUFx2_ASAP7_75t_R input72 (.A(key[49]),
    .Y(net138));
 BUFx2_ASAP7_75t_R input73 (.A(key[4]),
    .Y(net139));
 BUFx2_ASAP7_75t_R input74 (.A(key[50]),
    .Y(net140));
 BUFx2_ASAP7_75t_R input75 (.A(key[51]),
    .Y(net141));
 BUFx3_ASAP7_75t_R input76 (.A(key[52]),
    .Y(net142));
 BUFx3_ASAP7_75t_R input77 (.A(key[53]),
    .Y(net143));
 BUFx2_ASAP7_75t_R input78 (.A(key[54]),
    .Y(net144));
 BUFx2_ASAP7_75t_R input79 (.A(key[55]),
    .Y(net145));
 BUFx2_ASAP7_75t_R input80 (.A(key[56]),
    .Y(net146));
 BUFx2_ASAP7_75t_R input81 (.A(key[57]),
    .Y(net147));
 BUFx2_ASAP7_75t_R input82 (.A(key[58]),
    .Y(net148));
 BUFx2_ASAP7_75t_R input83 (.A(key[59]),
    .Y(net149));
 BUFx2_ASAP7_75t_R input84 (.A(key[5]),
    .Y(net150));
 BUFx2_ASAP7_75t_R input85 (.A(key[60]),
    .Y(net151));
 BUFx2_ASAP7_75t_R input86 (.A(key[61]),
    .Y(net152));
 BUFx2_ASAP7_75t_R input87 (.A(key[62]),
    .Y(net153));
 BUFx2_ASAP7_75t_R input88 (.A(key[63]),
    .Y(net154));
 BUFx2_ASAP7_75t_R input89 (.A(key[64]),
    .Y(net155));
 BUFx2_ASAP7_75t_R input90 (.A(key[65]),
    .Y(net156));
 BUFx2_ASAP7_75t_R input91 (.A(key[66]),
    .Y(net157));
 BUFx2_ASAP7_75t_R input92 (.A(key[67]),
    .Y(net158));
 BUFx2_ASAP7_75t_R input93 (.A(key[68]),
    .Y(net159));
 BUFx2_ASAP7_75t_R input94 (.A(key[69]),
    .Y(net160));
 BUFx2_ASAP7_75t_R input95 (.A(key[6]),
    .Y(net161));
 BUFx3_ASAP7_75t_R input96 (.A(key[70]),
    .Y(net162));
 BUFx2_ASAP7_75t_R input97 (.A(key[71]),
    .Y(net163));
 BUFx2_ASAP7_75t_R input98 (.A(key[72]),
    .Y(net164));
 BUFx2_ASAP7_75t_R input99 (.A(key[73]),
    .Y(net165));
 BUFx2_ASAP7_75t_R input100 (.A(key[74]),
    .Y(net166));
 BUFx2_ASAP7_75t_R input101 (.A(key[75]),
    .Y(net167));
 BUFx2_ASAP7_75t_R input102 (.A(key[76]),
    .Y(net168));
 BUFx2_ASAP7_75t_R input103 (.A(key[77]),
    .Y(net169));
 BUFx2_ASAP7_75t_R input104 (.A(key[78]),
    .Y(net170));
 BUFx2_ASAP7_75t_R input105 (.A(key[79]),
    .Y(net171));
 BUFx2_ASAP7_75t_R input106 (.A(key[7]),
    .Y(net172));
 BUFx2_ASAP7_75t_R input107 (.A(key[80]),
    .Y(net173));
 BUFx2_ASAP7_75t_R input108 (.A(key[81]),
    .Y(net174));
 BUFx2_ASAP7_75t_R input109 (.A(key[82]),
    .Y(net175));
 BUFx2_ASAP7_75t_R input110 (.A(key[83]),
    .Y(net176));
 BUFx2_ASAP7_75t_R input111 (.A(key[84]),
    .Y(net177));
 BUFx2_ASAP7_75t_R input112 (.A(key[85]),
    .Y(net178));
 BUFx2_ASAP7_75t_R input113 (.A(key[86]),
    .Y(net179));
 BUFx2_ASAP7_75t_R input114 (.A(key[87]),
    .Y(net180));
 BUFx2_ASAP7_75t_R input115 (.A(key[88]),
    .Y(net181));
 BUFx2_ASAP7_75t_R input116 (.A(key[89]),
    .Y(net182));
 BUFx2_ASAP7_75t_R input117 (.A(key[8]),
    .Y(net183));
 BUFx2_ASAP7_75t_R input118 (.A(key[90]),
    .Y(net184));
 BUFx2_ASAP7_75t_R input119 (.A(key[91]),
    .Y(net185));
 BUFx2_ASAP7_75t_R input120 (.A(key[92]),
    .Y(net186));
 BUFx2_ASAP7_75t_R input121 (.A(key[93]),
    .Y(net187));
 BUFx2_ASAP7_75t_R input122 (.A(key[94]),
    .Y(net188));
 BUFx2_ASAP7_75t_R input123 (.A(key[95]),
    .Y(net189));
 BUFx2_ASAP7_75t_R input124 (.A(key[96]),
    .Y(net190));
 BUFx2_ASAP7_75t_R input125 (.A(key[97]),
    .Y(net191));
 BUFx2_ASAP7_75t_R input126 (.A(key[98]),
    .Y(net192));
 BUFx2_ASAP7_75t_R input127 (.A(key[99]),
    .Y(net193));
 BUFx2_ASAP7_75t_R input128 (.A(key[9]),
    .Y(net194));
 BUFx4f_ASAP7_75t_R input129 (.A(ld),
    .Y(net195));
 BUFx2_ASAP7_75t_R input130 (.A(rst),
    .Y(net196));
 BUFx2_ASAP7_75t_R input131 (.A(text_in[0]),
    .Y(net197));
 BUFx2_ASAP7_75t_R input132 (.A(text_in[100]),
    .Y(net198));
 BUFx2_ASAP7_75t_R input133 (.A(text_in[101]),
    .Y(net199));
 BUFx2_ASAP7_75t_R input134 (.A(text_in[102]),
    .Y(net200));
 BUFx2_ASAP7_75t_R input135 (.A(text_in[103]),
    .Y(net201));
 BUFx2_ASAP7_75t_R input136 (.A(text_in[104]),
    .Y(net202));
 BUFx2_ASAP7_75t_R input137 (.A(text_in[105]),
    .Y(net203));
 BUFx2_ASAP7_75t_R input138 (.A(text_in[106]),
    .Y(net204));
 BUFx2_ASAP7_75t_R input139 (.A(text_in[107]),
    .Y(net205));
 BUFx2_ASAP7_75t_R input140 (.A(text_in[108]),
    .Y(net206));
 BUFx2_ASAP7_75t_R input141 (.A(text_in[109]),
    .Y(net207));
 BUFx2_ASAP7_75t_R input142 (.A(text_in[10]),
    .Y(net208));
 BUFx2_ASAP7_75t_R input143 (.A(text_in[110]),
    .Y(net209));
 BUFx2_ASAP7_75t_R input144 (.A(text_in[111]),
    .Y(net210));
 BUFx2_ASAP7_75t_R input145 (.A(text_in[112]),
    .Y(net211));
 BUFx2_ASAP7_75t_R input146 (.A(text_in[113]),
    .Y(net212));
 BUFx2_ASAP7_75t_R input147 (.A(text_in[114]),
    .Y(net213));
 BUFx2_ASAP7_75t_R input148 (.A(text_in[115]),
    .Y(net214));
 BUFx2_ASAP7_75t_R input149 (.A(text_in[116]),
    .Y(net215));
 BUFx2_ASAP7_75t_R input150 (.A(text_in[117]),
    .Y(net216));
 BUFx2_ASAP7_75t_R input151 (.A(text_in[118]),
    .Y(net217));
 BUFx2_ASAP7_75t_R input152 (.A(text_in[119]),
    .Y(net218));
 BUFx2_ASAP7_75t_R input153 (.A(text_in[11]),
    .Y(net219));
 BUFx2_ASAP7_75t_R input154 (.A(text_in[120]),
    .Y(net220));
 BUFx2_ASAP7_75t_R input155 (.A(text_in[121]),
    .Y(net221));
 BUFx2_ASAP7_75t_R input156 (.A(text_in[122]),
    .Y(net222));
 BUFx2_ASAP7_75t_R input157 (.A(text_in[123]),
    .Y(net223));
 BUFx2_ASAP7_75t_R input158 (.A(text_in[124]),
    .Y(net224));
 BUFx2_ASAP7_75t_R input159 (.A(text_in[125]),
    .Y(net225));
 BUFx2_ASAP7_75t_R input160 (.A(text_in[126]),
    .Y(net226));
 BUFx2_ASAP7_75t_R input161 (.A(text_in[127]),
    .Y(net227));
 BUFx2_ASAP7_75t_R input162 (.A(text_in[12]),
    .Y(net228));
 BUFx2_ASAP7_75t_R input163 (.A(text_in[13]),
    .Y(net229));
 BUFx2_ASAP7_75t_R input164 (.A(text_in[14]),
    .Y(net230));
 BUFx2_ASAP7_75t_R input165 (.A(text_in[15]),
    .Y(net231));
 BUFx2_ASAP7_75t_R input166 (.A(text_in[16]),
    .Y(net232));
 BUFx2_ASAP7_75t_R input167 (.A(text_in[17]),
    .Y(net233));
 BUFx2_ASAP7_75t_R input168 (.A(text_in[18]),
    .Y(net234));
 BUFx2_ASAP7_75t_R input169 (.A(text_in[19]),
    .Y(net235));
 BUFx2_ASAP7_75t_R input170 (.A(text_in[1]),
    .Y(net236));
 BUFx2_ASAP7_75t_R input171 (.A(text_in[20]),
    .Y(net237));
 BUFx2_ASAP7_75t_R input172 (.A(text_in[21]),
    .Y(net238));
 BUFx2_ASAP7_75t_R input173 (.A(text_in[22]),
    .Y(net239));
 BUFx2_ASAP7_75t_R input174 (.A(text_in[23]),
    .Y(net240));
 BUFx2_ASAP7_75t_R input175 (.A(text_in[24]),
    .Y(net241));
 BUFx2_ASAP7_75t_R input176 (.A(text_in[25]),
    .Y(net242));
 BUFx2_ASAP7_75t_R input177 (.A(text_in[26]),
    .Y(net243));
 BUFx2_ASAP7_75t_R input178 (.A(text_in[27]),
    .Y(net244));
 BUFx2_ASAP7_75t_R input179 (.A(text_in[28]),
    .Y(net245));
 BUFx2_ASAP7_75t_R input180 (.A(text_in[29]),
    .Y(net246));
 BUFx2_ASAP7_75t_R input181 (.A(text_in[2]),
    .Y(net247));
 BUFx2_ASAP7_75t_R input182 (.A(text_in[30]),
    .Y(net248));
 BUFx2_ASAP7_75t_R input183 (.A(text_in[31]),
    .Y(net249));
 BUFx2_ASAP7_75t_R input184 (.A(text_in[32]),
    .Y(net250));
 BUFx2_ASAP7_75t_R input185 (.A(text_in[33]),
    .Y(net251));
 BUFx2_ASAP7_75t_R input186 (.A(text_in[34]),
    .Y(net252));
 BUFx2_ASAP7_75t_R input187 (.A(text_in[35]),
    .Y(net253));
 BUFx2_ASAP7_75t_R input188 (.A(text_in[36]),
    .Y(net254));
 BUFx2_ASAP7_75t_R input189 (.A(text_in[37]),
    .Y(net255));
 BUFx2_ASAP7_75t_R input190 (.A(text_in[38]),
    .Y(net256));
 BUFx2_ASAP7_75t_R input191 (.A(text_in[39]),
    .Y(net257));
 BUFx2_ASAP7_75t_R input192 (.A(text_in[3]),
    .Y(net258));
 BUFx2_ASAP7_75t_R input193 (.A(text_in[40]),
    .Y(net259));
 BUFx2_ASAP7_75t_R input194 (.A(text_in[41]),
    .Y(net260));
 BUFx2_ASAP7_75t_R input195 (.A(text_in[42]),
    .Y(net261));
 BUFx2_ASAP7_75t_R input196 (.A(text_in[43]),
    .Y(net262));
 BUFx2_ASAP7_75t_R input197 (.A(text_in[44]),
    .Y(net263));
 BUFx2_ASAP7_75t_R input198 (.A(text_in[45]),
    .Y(net264));
 BUFx2_ASAP7_75t_R input199 (.A(text_in[46]),
    .Y(net265));
 BUFx2_ASAP7_75t_R input200 (.A(text_in[47]),
    .Y(net266));
 BUFx2_ASAP7_75t_R input201 (.A(text_in[48]),
    .Y(net267));
 BUFx2_ASAP7_75t_R input202 (.A(text_in[49]),
    .Y(net268));
 BUFx2_ASAP7_75t_R input203 (.A(text_in[4]),
    .Y(net269));
 BUFx2_ASAP7_75t_R input204 (.A(text_in[50]),
    .Y(net270));
 BUFx3_ASAP7_75t_R input205 (.A(text_in[51]),
    .Y(net271));
 BUFx2_ASAP7_75t_R input206 (.A(text_in[52]),
    .Y(net272));
 BUFx2_ASAP7_75t_R input207 (.A(text_in[53]),
    .Y(net273));
 BUFx2_ASAP7_75t_R input208 (.A(text_in[54]),
    .Y(net274));
 BUFx2_ASAP7_75t_R input209 (.A(text_in[55]),
    .Y(net275));
 BUFx2_ASAP7_75t_R input210 (.A(text_in[56]),
    .Y(net276));
 BUFx2_ASAP7_75t_R input211 (.A(text_in[57]),
    .Y(net277));
 BUFx2_ASAP7_75t_R input212 (.A(text_in[58]),
    .Y(net278));
 BUFx2_ASAP7_75t_R input213 (.A(text_in[59]),
    .Y(net279));
 BUFx2_ASAP7_75t_R input214 (.A(text_in[5]),
    .Y(net280));
 BUFx2_ASAP7_75t_R input215 (.A(text_in[60]),
    .Y(net281));
 BUFx2_ASAP7_75t_R input216 (.A(text_in[61]),
    .Y(net282));
 BUFx2_ASAP7_75t_R input217 (.A(text_in[62]),
    .Y(net283));
 BUFx2_ASAP7_75t_R input218 (.A(text_in[63]),
    .Y(net284));
 BUFx2_ASAP7_75t_R input219 (.A(text_in[64]),
    .Y(net285));
 BUFx2_ASAP7_75t_R input220 (.A(text_in[65]),
    .Y(net286));
 BUFx2_ASAP7_75t_R input221 (.A(text_in[66]),
    .Y(net287));
 BUFx2_ASAP7_75t_R input222 (.A(text_in[67]),
    .Y(net288));
 BUFx2_ASAP7_75t_R input223 (.A(text_in[68]),
    .Y(net289));
 BUFx2_ASAP7_75t_R input224 (.A(text_in[69]),
    .Y(net290));
 BUFx2_ASAP7_75t_R input225 (.A(text_in[6]),
    .Y(net291));
 BUFx2_ASAP7_75t_R input226 (.A(text_in[70]),
    .Y(net292));
 BUFx2_ASAP7_75t_R input227 (.A(text_in[71]),
    .Y(net293));
 BUFx2_ASAP7_75t_R input228 (.A(text_in[72]),
    .Y(net294));
 BUFx2_ASAP7_75t_R input229 (.A(text_in[73]),
    .Y(net295));
 BUFx2_ASAP7_75t_R input230 (.A(text_in[74]),
    .Y(net296));
 BUFx2_ASAP7_75t_R input231 (.A(text_in[75]),
    .Y(net297));
 BUFx2_ASAP7_75t_R input232 (.A(text_in[76]),
    .Y(net298));
 BUFx2_ASAP7_75t_R input233 (.A(text_in[77]),
    .Y(net299));
 BUFx2_ASAP7_75t_R input234 (.A(text_in[78]),
    .Y(net300));
 BUFx2_ASAP7_75t_R input235 (.A(text_in[79]),
    .Y(net301));
 BUFx2_ASAP7_75t_R input236 (.A(text_in[7]),
    .Y(net302));
 BUFx2_ASAP7_75t_R input237 (.A(text_in[80]),
    .Y(net303));
 BUFx2_ASAP7_75t_R input238 (.A(text_in[81]),
    .Y(net304));
 BUFx2_ASAP7_75t_R input239 (.A(text_in[82]),
    .Y(net305));
 BUFx2_ASAP7_75t_R input240 (.A(text_in[83]),
    .Y(net306));
 BUFx2_ASAP7_75t_R input241 (.A(text_in[84]),
    .Y(net307));
 BUFx2_ASAP7_75t_R input242 (.A(text_in[85]),
    .Y(net308));
 BUFx2_ASAP7_75t_R input243 (.A(text_in[86]),
    .Y(net309));
 BUFx2_ASAP7_75t_R input244 (.A(text_in[87]),
    .Y(net310));
 BUFx2_ASAP7_75t_R input245 (.A(text_in[88]),
    .Y(net311));
 BUFx2_ASAP7_75t_R input246 (.A(text_in[89]),
    .Y(net312));
 BUFx2_ASAP7_75t_R input247 (.A(text_in[8]),
    .Y(net313));
 BUFx2_ASAP7_75t_R input248 (.A(text_in[90]),
    .Y(net314));
 BUFx2_ASAP7_75t_R input249 (.A(text_in[91]),
    .Y(net315));
 BUFx2_ASAP7_75t_R input250 (.A(text_in[92]),
    .Y(net316));
 BUFx2_ASAP7_75t_R input251 (.A(text_in[93]),
    .Y(net317));
 BUFx2_ASAP7_75t_R input252 (.A(text_in[94]),
    .Y(net318));
 BUFx2_ASAP7_75t_R input253 (.A(text_in[95]),
    .Y(net319));
 BUFx2_ASAP7_75t_R input254 (.A(text_in[96]),
    .Y(net320));
 BUFx2_ASAP7_75t_R input255 (.A(text_in[97]),
    .Y(net321));
 BUFx2_ASAP7_75t_R input256 (.A(text_in[98]),
    .Y(net322));
 BUFx2_ASAP7_75t_R input257 (.A(text_in[99]),
    .Y(net323));
 BUFx2_ASAP7_75t_R input258 (.A(text_in[9]),
    .Y(net324));
 BUFx2_ASAP7_75t_R output259 (.A(net325),
    .Y(done));
 BUFx2_ASAP7_75t_R output260 (.A(net326),
    .Y(text_out[0]));
 BUFx2_ASAP7_75t_R output261 (.A(net327),
    .Y(text_out[100]));
 BUFx2_ASAP7_75t_R output262 (.A(net328),
    .Y(text_out[101]));
 BUFx2_ASAP7_75t_R output263 (.A(net329),
    .Y(text_out[102]));
 BUFx2_ASAP7_75t_R output264 (.A(net330),
    .Y(text_out[103]));
 BUFx2_ASAP7_75t_R output265 (.A(net331),
    .Y(text_out[104]));
 BUFx2_ASAP7_75t_R output266 (.A(net332),
    .Y(text_out[105]));
 BUFx2_ASAP7_75t_R output267 (.A(net333),
    .Y(text_out[106]));
 BUFx2_ASAP7_75t_R output268 (.A(net334),
    .Y(text_out[107]));
 BUFx2_ASAP7_75t_R output269 (.A(net335),
    .Y(text_out[108]));
 BUFx2_ASAP7_75t_R output270 (.A(net336),
    .Y(text_out[109]));
 BUFx2_ASAP7_75t_R output271 (.A(net337),
    .Y(text_out[10]));
 BUFx2_ASAP7_75t_R output272 (.A(net338),
    .Y(text_out[110]));
 BUFx2_ASAP7_75t_R output273 (.A(net339),
    .Y(text_out[111]));
 BUFx2_ASAP7_75t_R output274 (.A(net340),
    .Y(text_out[112]));
 BUFx2_ASAP7_75t_R output275 (.A(net341),
    .Y(text_out[113]));
 BUFx2_ASAP7_75t_R output276 (.A(net342),
    .Y(text_out[114]));
 BUFx2_ASAP7_75t_R output277 (.A(net343),
    .Y(text_out[115]));
 BUFx2_ASAP7_75t_R output278 (.A(net344),
    .Y(text_out[116]));
 BUFx2_ASAP7_75t_R output279 (.A(net345),
    .Y(text_out[117]));
 BUFx2_ASAP7_75t_R output280 (.A(net346),
    .Y(text_out[118]));
 BUFx2_ASAP7_75t_R output281 (.A(net347),
    .Y(text_out[119]));
 BUFx2_ASAP7_75t_R output282 (.A(net348),
    .Y(text_out[11]));
 BUFx2_ASAP7_75t_R output283 (.A(net349),
    .Y(text_out[120]));
 BUFx2_ASAP7_75t_R output284 (.A(net350),
    .Y(text_out[121]));
 BUFx2_ASAP7_75t_R output285 (.A(net351),
    .Y(text_out[122]));
 BUFx2_ASAP7_75t_R output286 (.A(net352),
    .Y(text_out[123]));
 BUFx2_ASAP7_75t_R output287 (.A(net353),
    .Y(text_out[124]));
 BUFx2_ASAP7_75t_R output288 (.A(net354),
    .Y(text_out[125]));
 BUFx2_ASAP7_75t_R output289 (.A(net355),
    .Y(text_out[126]));
 BUFx2_ASAP7_75t_R output290 (.A(net356),
    .Y(text_out[127]));
 BUFx2_ASAP7_75t_R output291 (.A(net357),
    .Y(text_out[12]));
 BUFx2_ASAP7_75t_R output292 (.A(net358),
    .Y(text_out[13]));
 BUFx2_ASAP7_75t_R output293 (.A(net359),
    .Y(text_out[14]));
 BUFx2_ASAP7_75t_R output294 (.A(net360),
    .Y(text_out[15]));
 BUFx2_ASAP7_75t_R output295 (.A(net361),
    .Y(text_out[16]));
 BUFx2_ASAP7_75t_R output296 (.A(net362),
    .Y(text_out[17]));
 BUFx2_ASAP7_75t_R output297 (.A(net363),
    .Y(text_out[18]));
 BUFx2_ASAP7_75t_R output298 (.A(net364),
    .Y(text_out[19]));
 BUFx2_ASAP7_75t_R output299 (.A(net365),
    .Y(text_out[1]));
 BUFx2_ASAP7_75t_R output300 (.A(net366),
    .Y(text_out[20]));
 BUFx2_ASAP7_75t_R output301 (.A(net367),
    .Y(text_out[21]));
 BUFx2_ASAP7_75t_R output302 (.A(net368),
    .Y(text_out[22]));
 BUFx2_ASAP7_75t_R output303 (.A(net369),
    .Y(text_out[23]));
 BUFx2_ASAP7_75t_R output304 (.A(net370),
    .Y(text_out[24]));
 BUFx2_ASAP7_75t_R output305 (.A(net371),
    .Y(text_out[25]));
 BUFx2_ASAP7_75t_R output306 (.A(net372),
    .Y(text_out[26]));
 BUFx2_ASAP7_75t_R output307 (.A(net373),
    .Y(text_out[27]));
 BUFx2_ASAP7_75t_R output308 (.A(net374),
    .Y(text_out[28]));
 BUFx2_ASAP7_75t_R output309 (.A(net375),
    .Y(text_out[29]));
 BUFx2_ASAP7_75t_R output310 (.A(net376),
    .Y(text_out[2]));
 BUFx2_ASAP7_75t_R output311 (.A(net377),
    .Y(text_out[30]));
 BUFx2_ASAP7_75t_R output312 (.A(net378),
    .Y(text_out[31]));
 BUFx2_ASAP7_75t_R output313 (.A(net379),
    .Y(text_out[32]));
 BUFx2_ASAP7_75t_R output314 (.A(net380),
    .Y(text_out[33]));
 BUFx2_ASAP7_75t_R output315 (.A(net381),
    .Y(text_out[34]));
 BUFx2_ASAP7_75t_R output316 (.A(net382),
    .Y(text_out[35]));
 BUFx2_ASAP7_75t_R output317 (.A(net383),
    .Y(text_out[36]));
 BUFx2_ASAP7_75t_R output318 (.A(net384),
    .Y(text_out[37]));
 BUFx2_ASAP7_75t_R output319 (.A(net385),
    .Y(text_out[38]));
 BUFx2_ASAP7_75t_R output320 (.A(net386),
    .Y(text_out[39]));
 BUFx2_ASAP7_75t_R output321 (.A(net387),
    .Y(text_out[3]));
 BUFx2_ASAP7_75t_R output322 (.A(net388),
    .Y(text_out[40]));
 BUFx2_ASAP7_75t_R output323 (.A(net389),
    .Y(text_out[41]));
 BUFx2_ASAP7_75t_R output324 (.A(net390),
    .Y(text_out[42]));
 BUFx2_ASAP7_75t_R output325 (.A(net391),
    .Y(text_out[43]));
 BUFx2_ASAP7_75t_R output326 (.A(net392),
    .Y(text_out[44]));
 BUFx2_ASAP7_75t_R output327 (.A(net393),
    .Y(text_out[45]));
 BUFx2_ASAP7_75t_R output328 (.A(net394),
    .Y(text_out[46]));
 BUFx2_ASAP7_75t_R output329 (.A(net395),
    .Y(text_out[47]));
 BUFx2_ASAP7_75t_R output330 (.A(net396),
    .Y(text_out[48]));
 BUFx2_ASAP7_75t_R output331 (.A(net397),
    .Y(text_out[49]));
 BUFx2_ASAP7_75t_R output332 (.A(net398),
    .Y(text_out[4]));
 BUFx2_ASAP7_75t_R output333 (.A(net399),
    .Y(text_out[50]));
 BUFx2_ASAP7_75t_R output334 (.A(net400),
    .Y(text_out[51]));
 BUFx2_ASAP7_75t_R output335 (.A(net401),
    .Y(text_out[52]));
 BUFx2_ASAP7_75t_R output336 (.A(net402),
    .Y(text_out[53]));
 BUFx2_ASAP7_75t_R output337 (.A(net403),
    .Y(text_out[54]));
 BUFx2_ASAP7_75t_R output338 (.A(net404),
    .Y(text_out[55]));
 BUFx2_ASAP7_75t_R output339 (.A(net405),
    .Y(text_out[56]));
 BUFx2_ASAP7_75t_R output340 (.A(net406),
    .Y(text_out[57]));
 BUFx2_ASAP7_75t_R output341 (.A(net407),
    .Y(text_out[58]));
 BUFx2_ASAP7_75t_R output342 (.A(net408),
    .Y(text_out[59]));
 BUFx2_ASAP7_75t_R output343 (.A(net409),
    .Y(text_out[5]));
 BUFx2_ASAP7_75t_R output344 (.A(net410),
    .Y(text_out[60]));
 BUFx2_ASAP7_75t_R output345 (.A(net411),
    .Y(text_out[61]));
 BUFx2_ASAP7_75t_R output346 (.A(net412),
    .Y(text_out[62]));
 BUFx2_ASAP7_75t_R output347 (.A(net413),
    .Y(text_out[63]));
 BUFx2_ASAP7_75t_R output348 (.A(net414),
    .Y(text_out[64]));
 BUFx2_ASAP7_75t_R output349 (.A(net415),
    .Y(text_out[65]));
 BUFx2_ASAP7_75t_R output350 (.A(net416),
    .Y(text_out[66]));
 BUFx2_ASAP7_75t_R output351 (.A(net417),
    .Y(text_out[67]));
 BUFx2_ASAP7_75t_R output352 (.A(net418),
    .Y(text_out[68]));
 BUFx2_ASAP7_75t_R output353 (.A(net419),
    .Y(text_out[69]));
 BUFx2_ASAP7_75t_R output354 (.A(net420),
    .Y(text_out[6]));
 BUFx2_ASAP7_75t_R output355 (.A(net421),
    .Y(text_out[70]));
 BUFx2_ASAP7_75t_R output356 (.A(net422),
    .Y(text_out[71]));
 BUFx2_ASAP7_75t_R output357 (.A(net423),
    .Y(text_out[72]));
 BUFx2_ASAP7_75t_R output358 (.A(net424),
    .Y(text_out[73]));
 BUFx2_ASAP7_75t_R output359 (.A(net425),
    .Y(text_out[74]));
 BUFx2_ASAP7_75t_R output360 (.A(net426),
    .Y(text_out[75]));
 BUFx2_ASAP7_75t_R output361 (.A(net427),
    .Y(text_out[76]));
 BUFx2_ASAP7_75t_R output362 (.A(net428),
    .Y(text_out[77]));
 BUFx2_ASAP7_75t_R output363 (.A(net429),
    .Y(text_out[78]));
 BUFx2_ASAP7_75t_R output364 (.A(net430),
    .Y(text_out[79]));
 BUFx2_ASAP7_75t_R output365 (.A(net431),
    .Y(text_out[7]));
 BUFx2_ASAP7_75t_R output366 (.A(net432),
    .Y(text_out[80]));
 BUFx2_ASAP7_75t_R output367 (.A(net433),
    .Y(text_out[81]));
 BUFx2_ASAP7_75t_R output368 (.A(net434),
    .Y(text_out[82]));
 BUFx2_ASAP7_75t_R output369 (.A(net435),
    .Y(text_out[83]));
 BUFx2_ASAP7_75t_R output370 (.A(net436),
    .Y(text_out[84]));
 BUFx2_ASAP7_75t_R output371 (.A(net437),
    .Y(text_out[85]));
 BUFx2_ASAP7_75t_R output372 (.A(net438),
    .Y(text_out[86]));
 BUFx2_ASAP7_75t_R output373 (.A(net439),
    .Y(text_out[87]));
 BUFx2_ASAP7_75t_R output374 (.A(net440),
    .Y(text_out[88]));
 BUFx2_ASAP7_75t_R output375 (.A(net441),
    .Y(text_out[89]));
 BUFx2_ASAP7_75t_R output376 (.A(net442),
    .Y(text_out[8]));
 BUFx2_ASAP7_75t_R output377 (.A(net443),
    .Y(text_out[90]));
 BUFx2_ASAP7_75t_R output378 (.A(net444),
    .Y(text_out[91]));
 BUFx2_ASAP7_75t_R output379 (.A(net445),
    .Y(text_out[92]));
 BUFx2_ASAP7_75t_R output380 (.A(net446),
    .Y(text_out[93]));
 BUFx2_ASAP7_75t_R output381 (.A(net447),
    .Y(text_out[94]));
 BUFx2_ASAP7_75t_R output382 (.A(net448),
    .Y(text_out[95]));
 BUFx2_ASAP7_75t_R output383 (.A(net449),
    .Y(text_out[96]));
 BUFx2_ASAP7_75t_R output384 (.A(net450),
    .Y(text_out[97]));
 BUFx2_ASAP7_75t_R output385 (.A(net451),
    .Y(text_out[98]));
 BUFx2_ASAP7_75t_R output386 (.A(net452),
    .Y(text_out[99]));
 BUFx2_ASAP7_75t_R output387 (.A(net453),
    .Y(text_out[9]));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_1_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_2_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_3_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_4_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_5_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_6_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_7_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_8_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_9_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_11_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_14_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_15_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_18_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_19_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_21_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_23_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_24_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_25_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_26_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_27_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_28_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_28_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_29_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_29_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_30_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_30_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_31_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_31_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_32_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_32_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_33_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_33_clk));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_0_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_1_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_2_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_3_0_clk));
 BUFx24_ASAP7_75t_R clkload0 (.A(clknet_2_0_0_clk));
 INVx8_ASAP7_75t_R clkload1 (.A(clknet_2_1_0_clk));
 CKINVDCx12_ASAP7_75t_R clkload2 (.A(clknet_2_3_0_clk));
 INVx5_ASAP7_75t_R clkload3 (.A(clknet_leaf_0_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload4 (.A(clknet_leaf_1_clk));
 INVxp67_ASAP7_75t_R clkload5 (.A(clknet_leaf_3_clk));
 INVxp33_ASAP7_75t_R clkload6 (.A(clknet_leaf_29_clk));
 INVx3_ASAP7_75t_R clkload7 (.A(clknet_leaf_30_clk));
 INVx5_ASAP7_75t_R clkload8 (.A(clknet_leaf_31_clk));
 INVx8_ASAP7_75t_R clkload9 (.A(clknet_leaf_32_clk));
 CKINVDCx9p33_ASAP7_75t_R clkload10 (.A(clknet_leaf_33_clk));
 INVx3_ASAP7_75t_R clkload11 (.A(clknet_leaf_4_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload12 (.A(clknet_leaf_6_clk));
 CKINVDCx14_ASAP7_75t_R clkload13 (.A(clknet_leaf_7_clk));
 CKINVDCx9p33_ASAP7_75t_R clkload14 (.A(clknet_leaf_8_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload15 (.A(clknet_leaf_9_clk));
 CKINVDCx10_ASAP7_75t_R clkload16 (.A(clknet_leaf_10_clk));
 INVxp67_ASAP7_75t_R clkload17 (.A(clknet_leaf_11_clk));
 BUFx4f_ASAP7_75t_R clkload18 (.A(clknet_leaf_19_clk));
 INVx3_ASAP7_75t_R clkload19 (.A(clknet_leaf_20_clk));
 INVx3_ASAP7_75t_R clkload20 (.A(clknet_leaf_21_clk));
 CKINVDCx11_ASAP7_75t_R clkload21 (.A(clknet_leaf_22_clk));
 INVx8_ASAP7_75t_R clkload22 (.A(clknet_leaf_23_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload23 (.A(clknet_leaf_24_clk));
 INVx5_ASAP7_75t_R clkload24 (.A(clknet_leaf_25_clk));
 INVx6_ASAP7_75t_R clkload25 (.A(clknet_leaf_26_clk));
 INVxp33_ASAP7_75t_R clkload26 (.A(clknet_leaf_27_clk));
 INVx3_ASAP7_75t_R clkload27 (.A(clknet_leaf_13_clk));
 INVx6_ASAP7_75t_R clkload28 (.A(clknet_leaf_14_clk));
 INVx6_ASAP7_75t_R clkload29 (.A(clknet_leaf_15_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload30 (.A(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkload31 (.A(clknet_leaf_17_clk));
 INVxp33_ASAP7_75t_R clkload32 (.A(clknet_leaf_18_clk));
 BUFx3_ASAP7_75t_R rebuffer1 (.A(_00524_),
    .Y(net454));
 BUFx6f_ASAP7_75t_R rebuffer2 (.A(net454),
    .Y(net455));
 BUFx3_ASAP7_75t_R rebuffer3 (.A(_00574_),
    .Y(net456));
 BUFx6f_ASAP7_75t_R rebuffer4 (.A(net456),
    .Y(net457));
 BUFx6f_ASAP7_75t_R rebuffer5 (.A(_04413_),
    .Y(net458));
 BUFx6f_ASAP7_75t_R rebuffer6 (.A(_05785_),
    .Y(net459));
 BUFx2_ASAP7_75t_R rebuffer7 (.A(_00504_),
    .Y(net460));
 BUFx2_ASAP7_75t_R rebuffer8 (.A(net460),
    .Y(net461));
 BUFx2_ASAP7_75t_R rebuffer9 (.A(net461),
    .Y(net462));
 BUFx6f_ASAP7_75t_R rebuffer10 (.A(_02445_),
    .Y(net463));
 BUFx3_ASAP7_75t_R rebuffer11 (.A(_00544_),
    .Y(net464));
 BUFx6f_ASAP7_75t_R rebuffer12 (.A(net464),
    .Y(net465));
 BUFx3_ASAP7_75t_R rebuffer13 (.A(_00494_),
    .Y(net466));
 BUFx6f_ASAP7_75t_R rebuffer14 (.A(_00609_),
    .Y(net467));
 BUFx3_ASAP7_75t_R rebuffer15 (.A(net467),
    .Y(net468));
 BUFx3_ASAP7_75t_R rebuffer16 (.A(_00534_),
    .Y(net469));
 BUFx3_ASAP7_75t_R rebuffer17 (.A(net469),
    .Y(net470));
 BUFx3_ASAP7_75t_R rebuffer18 (.A(net469),
    .Y(net471));
 BUFx2_ASAP7_75t_R rebuffer19 (.A(_00622_),
    .Y(net472));
 BUFx3_ASAP7_75t_R rebuffer20 (.A(_00622_),
    .Y(net473));
 BUFx2_ASAP7_75t_R rebuffer21 (.A(_00586_),
    .Y(net474));
 BUFx2_ASAP7_75t_R rebuffer22 (.A(net474),
    .Y(net475));
 BUFx3_ASAP7_75t_R rebuffer23 (.A(_00586_),
    .Y(net476));
 BUFx3_ASAP7_75t_R rebuffer24 (.A(_00554_),
    .Y(net477));
 BUFx2_ASAP7_75t_R rebuffer25 (.A(net477),
    .Y(net478));
 BUFx3_ASAP7_75t_R rebuffer26 (.A(net477),
    .Y(net479));
 BUFx3_ASAP7_75t_R rebuffer27 (.A(_00456_),
    .Y(net480));
 BUFx2_ASAP7_75t_R rebuffer28 (.A(net480),
    .Y(net481));
 BUFx3_ASAP7_75t_R rebuffer29 (.A(_06516_),
    .Y(net482));
 BUFx2_ASAP7_75t_R rebuffer30 (.A(net482),
    .Y(net483));
 BUFx3_ASAP7_75t_R rebuffer31 (.A(_00641_),
    .Y(net484));
 BUFx2_ASAP7_75t_R rebuffer32 (.A(net484),
    .Y(net485));
 BUFx6f_ASAP7_75t_R rebuffer33 (.A(_10814_),
    .Y(net486));
 BUFx3_ASAP7_75t_R rebuffer34 (.A(net486),
    .Y(net487));
 BUFx2_ASAP7_75t_R rebuffer35 (.A(net486),
    .Y(net488));
 BUFx2_ASAP7_75t_R rebuffer36 (.A(_00573_),
    .Y(net489));
 BUFx3_ASAP7_75t_R rebuffer37 (.A(_00610_),
    .Y(net490));
 BUFx2_ASAP7_75t_R rebuffer38 (.A(net490),
    .Y(net491));
 BUFx2_ASAP7_75t_R rebuffer39 (.A(_15789_),
    .Y(net492));
 BUFx2_ASAP7_75t_R rebuffer40 (.A(_15789_),
    .Y(net493));
 BUFx2_ASAP7_75t_R rebuffer41 (.A(net493),
    .Y(net494));
 BUFx3_ASAP7_75t_R rebuffer42 (.A(_00598_),
    .Y(net495));
 BUFx2_ASAP7_75t_R rebuffer43 (.A(_00632_),
    .Y(net496));
 BUFx2_ASAP7_75t_R rebuffer44 (.A(_00514_),
    .Y(net497));
 BUFx3_ASAP7_75t_R rebuffer45 (.A(_00514_),
    .Y(net498));
 BUFx2_ASAP7_75t_R rebuffer46 (.A(_00474_),
    .Y(net499));
 BUFx2_ASAP7_75t_R rebuffer47 (.A(_00484_),
    .Y(net500));
 BUFx2_ASAP7_75t_R rebuffer48 (.A(net500),
    .Y(net501));
 BUFx2_ASAP7_75t_R rebuffer49 (.A(_00484_),
    .Y(net502));
 BUFx2_ASAP7_75t_R rebuffer50 (.A(_00564_),
    .Y(net503));
 BUFx2_ASAP7_75t_R rebuffer51 (.A(net503),
    .Y(net504));
 BUFx3_ASAP7_75t_R rebuffer52 (.A(_01160_),
    .Y(net505));
 BUFx2_ASAP7_75t_R rebuffer53 (.A(net505),
    .Y(net506));
 BUFx2_ASAP7_75t_R rebuffer54 (.A(net505),
    .Y(net507));
 BUFx3_ASAP7_75t_R rebuffer55 (.A(_11461_),
    .Y(net508));
 BUFx6f_ASAP7_75t_R rebuffer56 (.A(net508),
    .Y(net509));
 BUFx2_ASAP7_75t_R rebuffer57 (.A(_11461_),
    .Y(net510));
 BUFx2_ASAP7_75t_R rebuffer58 (.A(_00640_),
    .Y(net511));
 BUFx3_ASAP7_75t_R rebuffer59 (.A(_00597_),
    .Y(net512));
 BUFx2_ASAP7_75t_R rebuffer60 (.A(_00597_),
    .Y(net513));
 BUFx2_ASAP7_75t_R rebuffer61 (.A(_05823_),
    .Y(net514));
 BUFx2_ASAP7_75t_R rebuffer62 (.A(_05823_),
    .Y(net515));
 BUFx2_ASAP7_75t_R rebuffer63 (.A(net515),
    .Y(net516));
 BUFx2_ASAP7_75t_R rebuffer64 (.A(_12893_),
    .Y(net517));
 BUFx2_ASAP7_75t_R rebuffer65 (.A(net517),
    .Y(net518));
 BUFx2_ASAP7_75t_R rebuffer66 (.A(net517),
    .Y(net519));
 BUFx2_ASAP7_75t_R rebuffer67 (.A(_12893_),
    .Y(net520));
 BUFx2_ASAP7_75t_R rebuffer68 (.A(net520),
    .Y(net521));
 BUFx4_ASAP7_75t_R rebuffer69 (.A(_05755_),
    .Y(net522));
 BUFx4f_ASAP7_75t_R rebuffer70 (.A(net522),
    .Y(net523));
 BUFx2_ASAP7_75t_R rebuffer71 (.A(net522),
    .Y(net524));
 BUFx2_ASAP7_75t_R rebuffer72 (.A(_13704_),
    .Y(net525));
 BUFx6f_ASAP7_75t_R rebuffer73 (.A(net525),
    .Y(net526));
 BUFx2_ASAP7_75t_R rebuffer74 (.A(_00475_),
    .Y(net527));
 BUFx2_ASAP7_75t_R rebuffer75 (.A(net527),
    .Y(net528));
 BUFx2_ASAP7_75t_R rebuffer76 (.A(_12148_),
    .Y(net529));
 BUFx2_ASAP7_75t_R rebuffer77 (.A(_02273_),
    .Y(net530));
 BUFx6f_ASAP7_75t_R rebuffer78 (.A(net530),
    .Y(net531));
 BUFx2_ASAP7_75t_R rebuffer79 (.A(_00483_),
    .Y(net532));
 BUFx2_ASAP7_75t_R rebuffer80 (.A(_01518_),
    .Y(net533));
 BUFx3_ASAP7_75t_R rebuffer81 (.A(net533),
    .Y(net534));
 BUFx2_ASAP7_75t_R rebuffer82 (.A(_01518_),
    .Y(net535));
 BUFx6f_ASAP7_75t_R rebuffer83 (.A(net535),
    .Y(net536));
 BUFx3_ASAP7_75t_R rebuffer84 (.A(_10911_),
    .Y(net537));
 BUFx6f_ASAP7_75t_R rebuffer85 (.A(_10911_),
    .Y(net538));
 BUFx2_ASAP7_75t_R rebuffer86 (.A(_00533_),
    .Y(net539));
 BUFx2_ASAP7_75t_R rebuffer87 (.A(_15872_),
    .Y(net540));
 BUFx2_ASAP7_75t_R rebuffer88 (.A(_15872_),
    .Y(net541));
 BUFx2_ASAP7_75t_R rebuffer89 (.A(_15872_),
    .Y(net542));
 BUFx2_ASAP7_75t_R rebuffer90 (.A(_00585_),
    .Y(net543));
 BUFx6f_ASAP7_75t_R rebuffer91 (.A(_10667_),
    .Y(net544));
 BUFx2_ASAP7_75t_R rebuffer92 (.A(net544),
    .Y(net545));
 BUFx2_ASAP7_75t_R rebuffer93 (.A(_02226_),
    .Y(net546));
 BUFx3_ASAP7_75t_R rebuffer94 (.A(_02226_),
    .Y(net547));
 BUFx2_ASAP7_75t_R rebuffer95 (.A(net547),
    .Y(net548));
 BUFx2_ASAP7_75t_R rebuffer96 (.A(net547),
    .Y(net549));
 BUFx2_ASAP7_75t_R rebuffer97 (.A(_10650_),
    .Y(net550));
 BUFx2_ASAP7_75t_R rebuffer98 (.A(_05057_),
    .Y(net551));
 BUFx2_ASAP7_75t_R rebuffer99 (.A(_05057_),
    .Y(net552));
 BUFx2_ASAP7_75t_R rebuffer100 (.A(_00465_),
    .Y(net553));
 BUFx2_ASAP7_75t_R rebuffer101 (.A(_00465_),
    .Y(net554));
 BUFx2_ASAP7_75t_R rebuffer102 (.A(_06441_),
    .Y(net555));
 BUFx2_ASAP7_75t_R rebuffer103 (.A(_06441_),
    .Y(net556));
 BUFx2_ASAP7_75t_R rebuffer104 (.A(_00599_),
    .Y(net557));
 BUFx2_ASAP7_75t_R rebuffer105 (.A(_15284_),
    .Y(net558));
 BUFx2_ASAP7_75t_R rebuffer106 (.A(_10650_),
    .Y(net559));
 BUFx2_ASAP7_75t_R rebuffer107 (.A(_12327_),
    .Y(net560));
 BUFx4f_ASAP7_75t_R rebuffer108 (.A(_07170_),
    .Y(net561));
 BUFx3_ASAP7_75t_R rebuffer109 (.A(_07170_),
    .Y(net562));
 BUFx2_ASAP7_75t_R rebuffer110 (.A(_01256_),
    .Y(net563));
 BUFx2_ASAP7_75t_R rebuffer111 (.A(_11380_),
    .Y(net564));
 BUFx2_ASAP7_75t_R rebuffer112 (.A(net564),
    .Y(net565));
 BUFx2_ASAP7_75t_R rebuffer113 (.A(net564),
    .Y(net566));
 BUFx2_ASAP7_75t_R rebuffer114 (.A(_15140_),
    .Y(net567));
 BUFx3_ASAP7_75t_R rebuffer115 (.A(net567),
    .Y(net568));
 BUFx2_ASAP7_75t_R rebuffer116 (.A(_15140_),
    .Y(net569));
 BUFx3_ASAP7_75t_R rebuffer117 (.A(_13089_),
    .Y(net570));
 BUFx2_ASAP7_75t_R rebuffer118 (.A(_01474_),
    .Y(net571));
 BUFx2_ASAP7_75t_R rebuffer119 (.A(net571),
    .Y(net572));
 BUFx2_ASAP7_75t_R rebuffer120 (.A(_01474_),
    .Y(net573));
 BUFx2_ASAP7_75t_R rebuffer121 (.A(net573),
    .Y(net574));
 BUFx2_ASAP7_75t_R rebuffer122 (.A(_00543_),
    .Y(net575));
 BUFx6f_ASAP7_75t_R rebuffer123 (.A(net774),
    .Y(net576));
 BUFx2_ASAP7_75t_R rebuffer124 (.A(_12234_),
    .Y(net577));
 BUFx2_ASAP7_75t_R rebuffer125 (.A(_13639_),
    .Y(net578));
 BUFx2_ASAP7_75t_R rebuffer126 (.A(_13639_),
    .Y(net579));
 BUFx3_ASAP7_75t_R rebuffer127 (.A(_01178_),
    .Y(net580));
 BUFx2_ASAP7_75t_R rebuffer128 (.A(net580),
    .Y(net581));
 BUFx2_ASAP7_75t_R rebuffer129 (.A(_00504_),
    .Y(net582));
 BUFx2_ASAP7_75t_R rebuffer130 (.A(net708),
    .Y(net583));
 BUFx2_ASAP7_75t_R rebuffer131 (.A(net583),
    .Y(net584));
 BUFx4_ASAP7_75t_R clone132 (.A(net650),
    .Y(net585));
 BUFx2_ASAP7_75t_R rebuffer133 (.A(_15978_),
    .Y(net586));
 BUFx2_ASAP7_75t_R rebuffer134 (.A(_15978_),
    .Y(net587));
 BUFx2_ASAP7_75t_R rebuffer135 (.A(net587),
    .Y(net588));
 BUFx2_ASAP7_75t_R rebuffer136 (.A(net587),
    .Y(net589));
 BUFx2_ASAP7_75t_R rebuffer137 (.A(net587),
    .Y(net590));
 BUFx2_ASAP7_75t_R rebuffer138 (.A(net597),
    .Y(net591));
 BUFx2_ASAP7_75t_R rebuffer139 (.A(_12148_),
    .Y(net592));
 BUFx6f_ASAP7_75t_R rebuffer140 (.A(_06558_),
    .Y(net593));
 BUFx3_ASAP7_75t_R rebuffer141 (.A(_03126_),
    .Y(net594));
 BUFx6f_ASAP7_75t_R rebuffer142 (.A(_05932_),
    .Y(net595));
 BUFx2_ASAP7_75t_R rebuffer143 (.A(_06569_),
    .Y(net596));
 BUFx6f_ASAP7_75t_R rebuffer144 (.A(_12086_),
    .Y(net597));
 BUFx2_ASAP7_75t_R rebuffer145 (.A(_04337_),
    .Y(net598));
 BUFx2_ASAP7_75t_R rebuffer146 (.A(net598),
    .Y(net599));
 BUFx3_ASAP7_75t_R rebuffer147 (.A(_03808_),
    .Y(net600));
 BUFx2_ASAP7_75t_R rebuffer148 (.A(net781),
    .Y(net601));
 BUFx2_ASAP7_75t_R rebuffer149 (.A(_00732_),
    .Y(net602));
 BUFx2_ASAP7_75t_R rebuffer150 (.A(_15819_),
    .Y(net603));
 BUFx2_ASAP7_75t_R rebuffer151 (.A(_10838_),
    .Y(net604));
 BUFx2_ASAP7_75t_R rebuffer152 (.A(_04308_),
    .Y(net605));
 BUFx2_ASAP7_75t_R rebuffer153 (.A(_00563_),
    .Y(net606));
 BUFx2_ASAP7_75t_R rebuffer154 (.A(net606),
    .Y(net607));
 BUFx2_ASAP7_75t_R rebuffer155 (.A(_12088_),
    .Y(net608));
 BUFx2_ASAP7_75t_R rebuffer156 (.A(net608),
    .Y(net609));
 BUFx2_ASAP7_75t_R rebuffer157 (.A(net608),
    .Y(net610));
 BUFx2_ASAP7_75t_R rebuffer158 (.A(_12118_),
    .Y(net611));
 BUFx2_ASAP7_75t_R rebuffer159 (.A(_13572_),
    .Y(net612));
 BUFx3_ASAP7_75t_R rebuffer160 (.A(net612),
    .Y(net613));
 BUFx2_ASAP7_75t_R rebuffer161 (.A(_13643_),
    .Y(net614));
 BUFx2_ASAP7_75t_R rebuffer162 (.A(_11536_),
    .Y(net615));
 BUFx2_ASAP7_75t_R rebuffer163 (.A(_11536_),
    .Y(net616));
 BUFx4_ASAP7_75t_R rebuffer164 (.A(_00995_),
    .Y(net617));
 BUFx3_ASAP7_75t_R rebuffer165 (.A(_00780_),
    .Y(net618));
 BUFx3_ASAP7_75t_R rebuffer166 (.A(_12830_),
    .Y(net619));
 BUFx2_ASAP7_75t_R rebuffer167 (.A(_00553_),
    .Y(net620));
 BUFx8_ASAP7_75t_R clone168 (.A(_10665_),
    .Y(net621));
 BUFx2_ASAP7_75t_R rebuffer169 (.A(_00598_),
    .Y(net622));
 BUFx8_ASAP7_75t_R clone170 (.A(net624),
    .Y(net623));
 BUFx2_ASAP7_75t_R rebuffer171 (.A(_02273_),
    .Y(net624));
 BUFx3_ASAP7_75t_R rebuffer172 (.A(_11364_),
    .Y(net625));
 BUFx3_ASAP7_75t_R rebuffer173 (.A(net625),
    .Y(net626));
 BUFx2_ASAP7_75t_R rebuffer174 (.A(_06475_),
    .Y(net627));
 BUFx2_ASAP7_75t_R rebuffer175 (.A(_06475_),
    .Y(net628));
 BUFx2_ASAP7_75t_R rebuffer176 (.A(_11407_),
    .Y(net629));
 BUFx2_ASAP7_75t_R rebuffer177 (.A(_01192_),
    .Y(net630));
 BUFx2_ASAP7_75t_R rebuffer178 (.A(_10679_),
    .Y(net631));
 BUFx2_ASAP7_75t_R rebuffer179 (.A(_14339_),
    .Y(net632));
 BUFx2_ASAP7_75t_R rebuffer180 (.A(_06404_),
    .Y(net633));
 BUFx2_ASAP7_75t_R rebuffer181 (.A(_06404_),
    .Y(net634));
 BUFx2_ASAP7_75t_R rebuffer182 (.A(_12116_),
    .Y(net635));
 BUFx2_ASAP7_75t_R rebuffer183 (.A(_15959_),
    .Y(net636));
 BUFx2_ASAP7_75t_R rebuffer184 (.A(_15959_),
    .Y(net637));
 BUFx3_ASAP7_75t_R rebuffer185 (.A(_15959_),
    .Y(net638));
 BUFx3_ASAP7_75t_R rebuffer186 (.A(_13090_),
    .Y(net639));
 BUFx2_ASAP7_75t_R rebuffer187 (.A(_00789_),
    .Y(net640));
 BUFx8_ASAP7_75t_R clone188 (.A(_10762_),
    .Y(net641));
 BUFx2_ASAP7_75t_R rebuffer189 (.A(_12832_),
    .Y(net642));
 BUFx2_ASAP7_75t_R rebuffer190 (.A(net642),
    .Y(net643));
 BUFx2_ASAP7_75t_R rebuffer191 (.A(net642),
    .Y(net644));
 BUFx2_ASAP7_75t_R rebuffer192 (.A(_12835_),
    .Y(net645));
 BUFx2_ASAP7_75t_R rebuffer193 (.A(_12835_),
    .Y(net646));
 BUFx2_ASAP7_75t_R clone194 (.A(net649),
    .Y(net647));
 BUFx4_ASAP7_75t_R clone195 (.A(_12893_),
    .Y(net648));
 BUFx2_ASAP7_75t_R rebuffer196 (.A(_00763_),
    .Y(net649));
 BUFx8_ASAP7_75t_R clone197 (.A(_10741_),
    .Y(net650));
 BUFx4f_ASAP7_75t_R clone198 (.A(_10665_),
    .Y(net651));
 BUFx2_ASAP7_75t_R rebuffer205 (.A(_00756_),
    .Y(net658));
 BUFx2_ASAP7_75t_R rebuffer206 (.A(_12867_),
    .Y(net659));
 BUFx6f_ASAP7_75t_R rebuffer207 (.A(_12867_),
    .Y(net660));
 BUFx2_ASAP7_75t_R rebuffer208 (.A(net660),
    .Y(net661));
 BUFx2_ASAP7_75t_R rebuffer209 (.A(_12847_),
    .Y(net662));
 BUFx2_ASAP7_75t_R rebuffer210 (.A(_13013_),
    .Y(net663));
 BUFx3_ASAP7_75t_R rebuffer211 (.A(_12848_),
    .Y(net664));
 BUFx2_ASAP7_75t_R rebuffer212 (.A(net664),
    .Y(net665));
 BUFx2_ASAP7_75t_R rebuffer213 (.A(net664),
    .Y(net666));
 BUFx2_ASAP7_75t_R rebuffer214 (.A(_10741_),
    .Y(net667));
 BUFx8_ASAP7_75t_R clone215 (.A(net669),
    .Y(net668));
 BUFx2_ASAP7_75t_R rebuffer216 (.A(_10618_),
    .Y(net669));
 BUFx4f_ASAP7_75t_R rebuffer217 (.A(_10651_),
    .Y(net670));
 BUFx2_ASAP7_75t_R rebuffer218 (.A(net670),
    .Y(net671));
 BUFx2_ASAP7_75t_R rebuffer225 (.A(_13584_),
    .Y(net678));
 BUFx3_ASAP7_75t_R clone226 (.A(_02337_),
    .Y(net679));
 BUFx8_ASAP7_75t_R clone227 (.A(_10619_),
    .Y(net680));
 BUFx2_ASAP7_75t_R rebuffer228 (.A(_13584_),
    .Y(net681));
 BUFx2_ASAP7_75t_R rebuffer229 (.A(_10822_),
    .Y(net682));
 BUFx6f_ASAP7_75t_R rebuffer230 (.A(net682),
    .Y(net683));
 BUFx2_ASAP7_75t_R rebuffer231 (.A(_10677_),
    .Y(net684));
 BUFx2_ASAP7_75t_R rebuffer232 (.A(_00576_),
    .Y(net685));
 BUFx2_ASAP7_75t_R rebuffer233 (.A(_11512_),
    .Y(net686));
 BUFx4f_ASAP7_75t_R rebuffer234 (.A(_11395_),
    .Y(net687));
 BUFx3_ASAP7_75t_R rebuffer235 (.A(_00772_),
    .Y(net688));
 BUFx2_ASAP7_75t_R rebuffer236 (.A(net688),
    .Y(net689));
 BUFx3_ASAP7_75t_R rebuffer237 (.A(_11395_),
    .Y(net690));
 BUFx6f_ASAP7_75t_R rebuffer238 (.A(_13041_),
    .Y(net691));
 BUFx2_ASAP7_75t_R rebuffer239 (.A(_14390_),
    .Y(net692));
 BUFx2_ASAP7_75t_R rebuffer240 (.A(_14390_),
    .Y(net693));
 BUFx2_ASAP7_75t_R rebuffer241 (.A(_14318_),
    .Y(net694));
 BUFx2_ASAP7_75t_R rebuffer242 (.A(_14390_),
    .Y(net695));
 BUFx2_ASAP7_75t_R rebuffer243 (.A(_14322_),
    .Y(net696));
 BUFx2_ASAP7_75t_R rebuffer244 (.A(_00811_),
    .Y(net697));
 BUFx2_ASAP7_75t_R rebuffer245 (.A(net697),
    .Y(net698));
 BUFx6f_ASAP7_75t_R rebuffer246 (.A(_14369_),
    .Y(net699));
 BUFx3_ASAP7_75t_R rebuffer247 (.A(_11360_),
    .Y(net700));
 BUFx2_ASAP7_75t_R rebuffer248 (.A(net700),
    .Y(net701));
 BUFx2_ASAP7_75t_R rebuffer249 (.A(_11360_),
    .Y(net702));
 BUFx4_ASAP7_75t_R clone250 (.A(_14369_),
    .Y(net703));
 BUFx2_ASAP7_75t_R rebuffer251 (.A(_11539_),
    .Y(net704));
 BUFx2_ASAP7_75t_R rebuffer253 (.A(_14366_),
    .Y(net706));
 BUFx2_ASAP7_75t_R rebuffer254 (.A(_01193_),
    .Y(net707));
 BUFx2_ASAP7_75t_R rebuffer255 (.A(_10629_),
    .Y(net708));
 BUFx2_ASAP7_75t_R rebuffer265 (.A(_15889_),
    .Y(net718));
 BUFx2_ASAP7_75t_R rebuffer266 (.A(_15889_),
    .Y(net719));
 BUFx2_ASAP7_75t_R rebuffer267 (.A(_15889_),
    .Y(net720));
 BUFx2_ASAP7_75t_R rebuffer268 (.A(net720),
    .Y(net721));
 BUFx2_ASAP7_75t_R rebuffer269 (.A(net720),
    .Y(net722));
 BUFx2_ASAP7_75t_R rebuffer270 (.A(_13639_),
    .Y(net723));
 BUFx2_ASAP7_75t_R rebuffer271 (.A(_13571_),
    .Y(net724));
 BUFx2_ASAP7_75t_R rebuffer272 (.A(_13573_),
    .Y(net725));
 BUFx2_ASAP7_75t_R clone273 (.A(_00771_),
    .Y(net726));
 BUFx2_ASAP7_75t_R clone274 (.A(_13841_),
    .Y(net727));
 BUFx2_ASAP7_75t_R rebuffer275 (.A(_10649_),
    .Y(net728));
 BUFx2_ASAP7_75t_R rebuffer285 (.A(_00575_),
    .Y(net738));
 BUFx6f_ASAP7_75t_R rebuffer286 (.A(_02436_),
    .Y(net739));
 BUFx3_ASAP7_75t_R rebuffer287 (.A(_04493_),
    .Y(net740));
 BUFx3_ASAP7_75t_R rebuffer288 (.A(_00612_),
    .Y(net741));
 BUFx2_ASAP7_75t_R rebuffer289 (.A(net741),
    .Y(net742));
 BUFx2_ASAP7_75t_R rebuffer304 (.A(_11579_),
    .Y(net757));
 BUFx2_ASAP7_75t_R rebuffer305 (.A(_00541_),
    .Y(net758));
 BUFx3_ASAP7_75t_R rebuffer306 (.A(_00541_),
    .Y(net759));
 BUFx3_ASAP7_75t_R rebuffer307 (.A(_14345_),
    .Y(net760));
 BUFx3_ASAP7_75t_R rebuffer308 (.A(_10826_),
    .Y(net761));
 BUFx3_ASAP7_75t_R rebuffer309 (.A(_05081_),
    .Y(net762));
 BUFx2_ASAP7_75t_R rebuffer310 (.A(_10733_),
    .Y(net763));
 BUFx3_ASAP7_75t_R rebuffer311 (.A(_05084_),
    .Y(net764));
 BUFx2_ASAP7_75t_R rebuffer313 (.A(_01248_),
    .Y(net766));
 BUFx8_ASAP7_75t_R clone314 (.A(_10619_),
    .Y(net767));
 BUFx2_ASAP7_75t_R rebuffer316 (.A(_01175_),
    .Y(net769));
 BUFx2_ASAP7_75t_R rebuffer317 (.A(net769),
    .Y(net770));
 BUFx2_ASAP7_75t_R rebuffer318 (.A(_01175_),
    .Y(net771));
 BUFx4_ASAP7_75t_R clone319 (.A(_12847_),
    .Y(net772));
 BUFx2_ASAP7_75t_R rebuffer320 (.A(_02966_),
    .Y(net773));
 BUFx6f_ASAP7_75t_R rebuffer321 (.A(_02909_),
    .Y(net774));
 BUFx2_ASAP7_75t_R rebuffer322 (.A(_02967_),
    .Y(net775));
 BUFx3_ASAP7_75t_R rebuffer323 (.A(_11381_),
    .Y(net776));
 BUFx2_ASAP7_75t_R rebuffer324 (.A(net776),
    .Y(net777));
 BUFx2_ASAP7_75t_R rebuffer325 (.A(_00819_),
    .Y(net778));
 BUFx2_ASAP7_75t_R rebuffer326 (.A(net899),
    .Y(net779));
 BUFx8_ASAP7_75t_R clone327 (.A(_10619_),
    .Y(net780));
 BUFx6f_ASAP7_75t_R rebuffer328 (.A(_10627_),
    .Y(net781));
 BUFx2_ASAP7_75t_R rebuffer329 (.A(_10642_),
    .Y(net782));
 BUFx2_ASAP7_75t_R rebuffer330 (.A(_10704_),
    .Y(net783));
 BUFx2_ASAP7_75t_R rebuffer331 (.A(_10704_),
    .Y(net784));
 BUFx2_ASAP7_75t_R rebuffer332 (.A(_10635_),
    .Y(net785));
 BUFx2_ASAP7_75t_R rebuffer333 (.A(_10619_),
    .Y(net786));
 BUFx2_ASAP7_75t_R rebuffer334 (.A(_11407_),
    .Y(net787));
 BUFx2_ASAP7_75t_R rebuffer335 (.A(_11405_),
    .Y(net788));
 BUFx2_ASAP7_75t_R rebuffer336 (.A(_11404_),
    .Y(net789));
 BUFx2_ASAP7_75t_R rebuffer349 (.A(net804),
    .Y(net802));
 BUFx4_ASAP7_75t_R clone350 (.A(net804),
    .Y(net803));
 BUFx2_ASAP7_75t_R rebuffer351 (.A(net839),
    .Y(net804));
 BUFx2_ASAP7_75t_R rebuffer352 (.A(_07978_),
    .Y(net805));
 BUFx2_ASAP7_75t_R rebuffer353 (.A(_00812_),
    .Y(net806));
 BUFx2_ASAP7_75t_R rebuffer355 (.A(net807),
    .Y(net808));
 BUFx2_ASAP7_75t_R rebuffer356 (.A(net807),
    .Y(net809));
 BUFx2_ASAP7_75t_R rebuffer357 (.A(_04457_),
    .Y(net810));
 BUFx6f_ASAP7_75t_R rebuffer358 (.A(_04457_),
    .Y(net811));
 BUFx2_ASAP7_75t_R rebuffer359 (.A(_15872_),
    .Y(net812));
 OAI21x1_ASAP7_75t_R clone360 (.A1(_13641_),
    .A2(_13642_),
    .B(_13793_),
    .Y(net813));
 BUFx2_ASAP7_75t_R rebuffer361 (.A(_01186_),
    .Y(net814));
 BUFx2_ASAP7_75t_R rebuffer362 (.A(_01186_),
    .Y(net815));
 BUFx3_ASAP7_75t_R rebuffer363 (.A(_13588_),
    .Y(net816));
 BUFx2_ASAP7_75t_R rebuffer364 (.A(net816),
    .Y(net817));
 BUFx2_ASAP7_75t_R rebuffer365 (.A(_13637_),
    .Y(net818));
 BUFx3_ASAP7_75t_R rebuffer366 (.A(_13608_),
    .Y(net819));
 BUFx2_ASAP7_75t_R rebuffer367 (.A(_13612_),
    .Y(net820));
 BUFx3_ASAP7_75t_R rebuffer368 (.A(_06569_),
    .Y(net821));
 BUFx12f_ASAP7_75t_R rebuffer369 (.A(_15784_),
    .Y(net822));
 BUFx2_ASAP7_75t_R rebuffer370 (.A(net822),
    .Y(net823));
 BUFx2_ASAP7_75t_R rebuffer371 (.A(net823),
    .Y(net824));
 BUFx2_ASAP7_75t_R rebuffer372 (.A(_08196_),
    .Y(net825));
 BUFx2_ASAP7_75t_R rebuffer373 (.A(net825),
    .Y(net826));
 BUFx2_ASAP7_75t_R rebuffer374 (.A(_15957_),
    .Y(net827));
 BUFx2_ASAP7_75t_R rebuffer375 (.A(_06614_),
    .Y(net828));
 BUFx6f_ASAP7_75t_R rebuffer376 (.A(_03597_),
    .Y(net829));
 BUFx2_ASAP7_75t_R rebuffer377 (.A(_00819_),
    .Y(net830));
 BUFx2_ASAP7_75t_R rebuffer378 (.A(_03732_),
    .Y(net831));
 BUFx2_ASAP7_75t_R rebuffer379 (.A(_03651_),
    .Y(net832));
 BUFx4_ASAP7_75t_R clone380 (.A(_03732_),
    .Y(net833));
 BUFx6f_ASAP7_75t_R rebuffer382 (.A(_03597_),
    .Y(net835));
 BUFx3_ASAP7_75t_R rebuffer383 (.A(_03808_),
    .Y(net836));
 BUFx2_ASAP7_75t_R rebuffer384 (.A(_00458_),
    .Y(net837));
 BUFx6f_ASAP7_75t_R rebuffer385 (.A(_07966_),
    .Y(net838));
 BUFx6f_ASAP7_75t_R rebuffer386 (.A(_07966_),
    .Y(net839));
 BUFx2_ASAP7_75t_R rebuffer387 (.A(_15088_),
    .Y(net840));
 BUFx2_ASAP7_75t_R rebuffer388 (.A(net840),
    .Y(net841));
 BUFx2_ASAP7_75t_R rebuffer389 (.A(_15084_),
    .Y(net842));
 BUFx2_ASAP7_75t_R rebuffer390 (.A(_15084_),
    .Y(net843));
 BUFx4_ASAP7_75t_R clone391 (.A(net845),
    .Y(net844));
 BUFx2_ASAP7_75t_R rebuffer392 (.A(_00845_),
    .Y(net845));
 BUFx2_ASAP7_75t_R rebuffer393 (.A(_06565_),
    .Y(net846));
 BUFx2_ASAP7_75t_R rebuffer394 (.A(_12338_),
    .Y(net847));
 BUFx2_ASAP7_75t_R rebuffer395 (.A(_12099_),
    .Y(net848));
 BUFx4_ASAP7_75t_R clone396 (.A(net866),
    .Y(net849));
 BUFx2_ASAP7_75t_R rebuffer397 (.A(_12087_),
    .Y(net850));
 BUFx6f_ASAP7_75t_R rebuffer400 (.A(_11367_),
    .Y(net853));
 BUFx2_ASAP7_75t_R rebuffer401 (.A(_01059_),
    .Y(net854));
 BUFx3_ASAP7_75t_R rebuffer402 (.A(net854),
    .Y(net855));
 BUFx2_ASAP7_75t_R rebuffer403 (.A(net854),
    .Y(net856));
 BUFx2_ASAP7_75t_R rebuffer404 (.A(_09503_),
    .Y(net857));
 BUFx2_ASAP7_75t_R rebuffer405 (.A(_08016_),
    .Y(net858));
 BUFx2_ASAP7_75t_R rebuffer406 (.A(net858),
    .Y(net859));
 BUFx3_ASAP7_75t_R rebuffer407 (.A(net858),
    .Y(net860));
 BUFx2_ASAP7_75t_R rebuffer408 (.A(_08015_),
    .Y(net861));
 BUFx2_ASAP7_75t_R rebuffer409 (.A(_08015_),
    .Y(net862));
 BUFx2_ASAP7_75t_R rebuffer410 (.A(_03126_),
    .Y(net863));
 BUFx2_ASAP7_75t_R rebuffer411 (.A(_00485_),
    .Y(net864));
 BUFx2_ASAP7_75t_R rebuffer412 (.A(_12103_),
    .Y(net865));
 BUFx8_ASAP7_75t_R clone413 (.A(_10638_),
    .Y(net866));
 BUFx8_ASAP7_75t_R clone414 (.A(_10620_),
    .Y(net867));
 BUFx2_ASAP7_75t_R rebuffer415 (.A(_01199_),
    .Y(net868));
 BUFx2_ASAP7_75t_R rebuffer416 (.A(_01199_),
    .Y(net869));
 BUFx2_ASAP7_75t_R rebuffer417 (.A(_15023_),
    .Y(net870));
 BUFx2_ASAP7_75t_R rebuffer418 (.A(_05802_),
    .Y(net871));
 BUFx2_ASAP7_75t_R rebuffer419 (.A(_03652_),
    .Y(net872));
 BUFx2_ASAP7_75t_R rebuffer420 (.A(net872),
    .Y(net873));
 BUFx2_ASAP7_75t_R rebuffer421 (.A(net872),
    .Y(net874));
 BUFx2_ASAP7_75t_R rebuffer422 (.A(_01631_),
    .Y(net875));
 BUFx2_ASAP7_75t_R rebuffer423 (.A(_01631_),
    .Y(net876));
 BUFx2_ASAP7_75t_R rebuffer424 (.A(net876),
    .Y(net877));
 BUFx6f_ASAP7_75t_R rebuffer425 (.A(_01459_),
    .Y(net878));
 BUFx2_ASAP7_75t_R rebuffer431 (.A(_01233_),
    .Y(net884));
 BUFx3_ASAP7_75t_R rebuffer432 (.A(_01521_),
    .Y(net885));
 BUFx2_ASAP7_75t_R rebuffer433 (.A(net885),
    .Y(net886));
 BUFx2_ASAP7_75t_R rebuffer434 (.A(_01506_),
    .Y(net887));
 BUFx2_ASAP7_75t_R rebuffer435 (.A(net887),
    .Y(net888));
 BUFx2_ASAP7_75t_R rebuffer436 (.A(_01210_),
    .Y(net889));
 BUFx2_ASAP7_75t_R rebuffer437 (.A(_01210_),
    .Y(net890));
 BUFx2_ASAP7_75t_R rebuffer438 (.A(_06421_),
    .Y(net891));
 BUFx2_ASAP7_75t_R rebuffer439 (.A(net891),
    .Y(net892));
 BUFx2_ASAP7_75t_R rebuffer440 (.A(_11615_),
    .Y(net893));
 BUFx3_ASAP7_75t_R rebuffer441 (.A(_11615_),
    .Y(net894));
 BUFx3_ASAP7_75t_R rebuffer442 (.A(net894),
    .Y(net895));
 BUFx2_ASAP7_75t_R rebuffer443 (.A(_11511_),
    .Y(net896));
 BUFx2_ASAP7_75t_R rebuffer444 (.A(_11594_),
    .Y(net897));
 BUFx3_ASAP7_75t_R rebuffer445 (.A(_11631_),
    .Y(net898));
 BUFx2_ASAP7_75t_R rebuffer446 (.A(_15022_),
    .Y(net899));
 BUFx2_ASAP7_75t_R clone447 (.A(_15211_),
    .Y(net900));
 BUFx3_ASAP7_75t_R rebuffer448 (.A(_03795_),
    .Y(net901));
 BUFx2_ASAP7_75t_R rebuffer449 (.A(_03943_),
    .Y(net902));
 BUFx6f_ASAP7_75t_R rebuffer450 (.A(_15034_),
    .Y(net903));
 BUFx4_ASAP7_75t_R clone451 (.A(_15088_),
    .Y(net904));
 BUFx4f_ASAP7_75t_R rebuffer452 (.A(_12082_),
    .Y(net905));
 BUFx2_ASAP7_75t_R rebuffer453 (.A(_05139_),
    .Y(net906));
 BUFx2_ASAP7_75t_R rebuffer454 (.A(_01463_),
    .Y(net907));
 BUFx2_ASAP7_75t_R clone455 (.A(net909),
    .Y(net908));
 BUFx2_ASAP7_75t_R rebuffer456 (.A(_00827_),
    .Y(net909));
 BUFx2_ASAP7_75t_R rebuffer457 (.A(_00820_),
    .Y(net910));
 BUFx6f_ASAP7_75t_R rebuffer458 (.A(_00820_),
    .Y(net911));
 BUFx6f_ASAP7_75t_R rebuffer462 (.A(net916),
    .Y(net915));
 BUFx6f_ASAP7_75t_R rebuffer463 (.A(_03769_),
    .Y(net916));
 BUFx2_ASAP7_75t_R rebuffer464 (.A(_01264_),
    .Y(net917));
 BUFx2_ASAP7_75t_R rebuffer465 (.A(_01249_),
    .Y(net918));
 BUFx2_ASAP7_75t_R rebuffer466 (.A(_01249_),
    .Y(net919));
 BUFx2_ASAP7_75t_R rebuffer467 (.A(_01249_),
    .Y(net920));
 BUFx4f_ASAP7_75t_R rebuffer468 (.A(_12084_),
    .Y(net921));
 BUFx2_ASAP7_75t_R rebuffer469 (.A(_12289_),
    .Y(net922));
 BUFx2_ASAP7_75t_R rebuffer470 (.A(_03648_),
    .Y(net923));
 BUFx3_ASAP7_75t_R rebuffer471 (.A(_03648_),
    .Y(net924));
 BUFx2_ASAP7_75t_R rebuffer472 (.A(net924),
    .Y(net925));
 BUFx8_ASAP7_75t_R clone474 (.A(net931),
    .Y(net927));
 BUFx2_ASAP7_75t_R rebuffer476 (.A(net928),
    .Y(net929));
 BUFx2_ASAP7_75t_R rebuffer477 (.A(net928),
    .Y(net930));
 BUFx2_ASAP7_75t_R rebuffer478 (.A(_08105_),
    .Y(net931));
 BUFx3_ASAP7_75t_R rebuffer479 (.A(_07414_),
    .Y(net932));
 BUFx2_ASAP7_75t_R rebuffer480 (.A(_07110_),
    .Y(net933));
 BUFx2_ASAP7_75t_R rebuffer481 (.A(net933),
    .Y(net934));
 BUFx2_ASAP7_75t_R rebuffer482 (.A(_07110_),
    .Y(net935));
 BUFx2_ASAP7_75t_R rebuffer483 (.A(_01274_),
    .Y(net936));
 BUFx2_ASAP7_75t_R rebuffer484 (.A(_07092_),
    .Y(net937));
 BUFx2_ASAP7_75t_R rebuffer485 (.A(_07092_),
    .Y(net938));
 BUFx6f_ASAP7_75t_R rebuffer486 (.A(_04293_),
    .Y(net939));
 BUFx6f_ASAP7_75t_R rebuffer487 (.A(_01271_),
    .Y(net940));
 BUFx2_ASAP7_75t_R rebuffer488 (.A(net940),
    .Y(net941));
 BUFx2_ASAP7_75t_R rebuffer489 (.A(net941),
    .Y(net942));
 BUFx8_ASAP7_75t_R clone490 (.A(_07189_),
    .Y(net943));
 BUFx6f_ASAP7_75t_R rebuffer491 (.A(_00467_),
    .Y(net944));
 BUFx2_ASAP7_75t_R rebuffer492 (.A(net944),
    .Y(net945));
 BUFx2_ASAP7_75t_R rebuffer493 (.A(_07255_),
    .Y(net946));
 BUFx4_ASAP7_75t_R clone494 (.A(_07092_),
    .Y(net947));
 BUFx2_ASAP7_75t_R rebuffer495 (.A(_07125_),
    .Y(net948));
 BUFx2_ASAP7_75t_R rebuffer496 (.A(net948),
    .Y(net949));
 BUFx2_ASAP7_75t_R rebuffer497 (.A(_07125_),
    .Y(net950));
endmodule
