module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire net3;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire net2013;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire net2008;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire net2;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire net8;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire net7;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire net6;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire net5;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire clk_i_regs;
 wire net305;
 wire \alu_adder_result_ex[0] ;
 wire \alu_adder_result_ex[10] ;
 wire \alu_adder_result_ex[11] ;
 wire \alu_adder_result_ex[12] ;
 wire \alu_adder_result_ex[13] ;
 wire \alu_adder_result_ex[14] ;
 wire \alu_adder_result_ex[15] ;
 wire \alu_adder_result_ex[16] ;
 wire \alu_adder_result_ex[17] ;
 wire \alu_adder_result_ex[18] ;
 wire \alu_adder_result_ex[19] ;
 wire \alu_adder_result_ex[1] ;
 wire \alu_adder_result_ex[20] ;
 wire \alu_adder_result_ex[21] ;
 wire \alu_adder_result_ex[22] ;
 wire \alu_adder_result_ex[23] ;
 wire \alu_adder_result_ex[24] ;
 wire \alu_adder_result_ex[25] ;
 wire \alu_adder_result_ex[26] ;
 wire \alu_adder_result_ex[27] ;
 wire \alu_adder_result_ex[28] ;
 wire \alu_adder_result_ex[29] ;
 wire \alu_adder_result_ex[2] ;
 wire \alu_adder_result_ex[30] ;
 wire \alu_adder_result_ex[31] ;
 wire \alu_adder_result_ex[3] ;
 wire \alu_adder_result_ex[4] ;
 wire \alu_adder_result_ex[5] ;
 wire \alu_adder_result_ex[6] ;
 wire \alu_adder_result_ex[7] ;
 wire \alu_adder_result_ex[8] ;
 wire \alu_adder_result_ex[9] ;
 wire clk;
 wire core_busy_d;
 wire \core_clock_gate_i.en_latch ;
 wire net199;
 wire \cs_registers_i.mcycle_counter_i.counter[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter[1] ;
 wire \cs_registers_i.mhpmcounter[2][0] ;
 wire \cs_registers_i.mhpmcounter[2][1] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.priv_lvl_q[0] ;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.load_err_d ;
 wire \id_stage_i.controller_i.store_err_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net1;
 wire net4;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net95;
 wire net145;
 wire net151;
 wire net152;
 wire net153;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_leaf_0_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_6_clk_i_regs;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_13_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_18_clk_i_regs;
 wire clknet_leaf_19_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_23_clk_i_regs;
 wire clknet_leaf_24_clk_i_regs;
 wire clknet_leaf_25_clk_i_regs;
 wire clknet_leaf_26_clk_i_regs;
 wire clknet_leaf_27_clk_i_regs;
 wire clknet_leaf_28_clk_i_regs;
 wire clknet_leaf_29_clk_i_regs;
 wire clknet_leaf_30_clk_i_regs;
 wire clknet_leaf_31_clk_i_regs;
 wire clknet_leaf_32_clk_i_regs;
 wire clknet_leaf_33_clk_i_regs;
 wire clknet_leaf_34_clk_i_regs;
 wire clknet_leaf_35_clk_i_regs;
 wire clknet_leaf_36_clk_i_regs;
 wire clknet_leaf_37_clk_i_regs;
 wire clknet_leaf_38_clk_i_regs;
 wire clknet_leaf_39_clk_i_regs;
 wire clknet_leaf_40_clk_i_regs;
 wire clknet_leaf_41_clk_i_regs;
 wire clknet_leaf_42_clk_i_regs;
 wire clknet_leaf_43_clk_i_regs;
 wire clknet_leaf_44_clk_i_regs;
 wire clknet_0_clk_i_regs;
 wire clknet_2_0__leaf_clk_i_regs;
 wire clknet_2_1__leaf_clk_i_regs;
 wire clknet_2_2__leaf_clk_i_regs;
 wire clknet_2_3__leaf_clk_i_regs;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire delaynet_0_core_clock;
 wire delaynet_1_core_clock;
 wire delaynet_2_core_clock;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;

 BUFx4f_ASAP7_75t_R _19086_ (.A(_01510_),
    .Y(_13357_));
 INVx2_ASAP7_75t_R _19087_ (.A(_13357_),
    .Y(_13358_));
 BUFx4f_ASAP7_75t_R _19088_ (.A(_01509_),
    .Y(_13359_));
 INVx1_ASAP7_75t_R _19089_ (.A(_00399_),
    .Y(_13360_));
 AO211x2_ASAP7_75t_R _19090_ (.A1(_18763_),
    .A2(_13358_),
    .B(_13359_),
    .C(_13360_),
    .Y(_13361_));
 NAND2x2_ASAP7_75t_R _19091_ (.A(_13359_),
    .B(_01510_),
    .Y(_13362_));
 OR2x2_ASAP7_75t_R _19092_ (.A(_00399_),
    .B(_13362_),
    .Y(_13363_));
 AND2x2_ASAP7_75t_R _19093_ (.A(_13361_),
    .B(_13363_),
    .Y(_13364_));
 BUFx4f_ASAP7_75t_R _19094_ (.A(_13364_),
    .Y(_13365_));
 BUFx4f_ASAP7_75t_R _19095_ (.A(_13365_),
    .Y(_13366_));
 BUFx4f_ASAP7_75t_R _19096_ (.A(_13366_),
    .Y(_13367_));
 INVx2_ASAP7_75t_R _19097_ (.A(_01776_),
    .Y(_13368_));
 BUFx6f_ASAP7_75t_R _19098_ (.A(_00400_),
    .Y(_13369_));
 BUFx6f_ASAP7_75t_R _19099_ (.A(_00024_),
    .Y(_13370_));
 NOR2x2_ASAP7_75t_R _19100_ (.A(_13369_),
    .B(_13370_),
    .Y(_13371_));
 OA211x2_ASAP7_75t_R _19101_ (.A1(_13368_),
    .A2(net2018),
    .B(_00021_),
    .C(_13371_),
    .Y(_13372_));
 BUFx6f_ASAP7_75t_R _19102_ (.A(_13372_),
    .Y(_13373_));
 BUFx12f_ASAP7_75t_R _19103_ (.A(_13370_),
    .Y(_13374_));
 INVx3_ASAP7_75t_R _19104_ (.A(_13369_),
    .Y(_13375_));
 BUFx6f_ASAP7_75t_R _19105_ (.A(_00021_),
    .Y(_13376_));
 INVx3_ASAP7_75t_R _19106_ (.A(_13376_),
    .Y(_13377_));
 AND3x1_ASAP7_75t_R _19107_ (.A(_13369_),
    .B(net2001),
    .C(_13376_),
    .Y(_13378_));
 AO21x1_ASAP7_75t_R _19108_ (.A1(_13375_),
    .A2(_13377_),
    .B(_13378_),
    .Y(_13379_));
 BUFx4f_ASAP7_75t_R _19109_ (.A(_01553_),
    .Y(_13380_));
 NOR2x2_ASAP7_75t_R _19110_ (.A(_00013_),
    .B(_13380_),
    .Y(_13381_));
 BUFx6f_ASAP7_75t_R _19111_ (.A(_00015_),
    .Y(_13382_));
 BUFx6f_ASAP7_75t_R _19112_ (.A(_00018_),
    .Y(_13383_));
 AND2x4_ASAP7_75t_R _19113_ (.A(_13382_),
    .B(_13383_),
    .Y(_13384_));
 NAND2x1_ASAP7_75t_R _19114_ (.A(_13381_),
    .B(_13384_),
    .Y(_13385_));
 OR3x4_ASAP7_75t_R _19115_ (.A(_13374_),
    .B(_13379_),
    .C(_13385_),
    .Y(_13386_));
 NOR2x2_ASAP7_75t_R _19116_ (.A(_13373_),
    .B(_13386_),
    .Y(_13387_));
 INVx3_ASAP7_75t_R _19117_ (.A(_01552_),
    .Y(_13388_));
 BUFx6f_ASAP7_75t_R _19118_ (.A(_13388_),
    .Y(_13389_));
 BUFx6f_ASAP7_75t_R _19119_ (.A(_13389_),
    .Y(_13390_));
 INVx4_ASAP7_75t_R _19120_ (.A(_13382_),
    .Y(_13391_));
 INVx3_ASAP7_75t_R _19121_ (.A(_13383_),
    .Y(_13392_));
 AND2x2_ASAP7_75t_R _19122_ (.A(_13369_),
    .B(_13370_),
    .Y(_13393_));
 AND5x2_ASAP7_75t_R _19123_ (.A(_13391_),
    .B(_13392_),
    .C(_13376_),
    .D(_13381_),
    .E(_13393_),
    .Y(_13394_));
 BUFx6f_ASAP7_75t_R _19124_ (.A(_00404_),
    .Y(_13395_));
 NAND2x2_ASAP7_75t_R _19125_ (.A(net2000),
    .B(_00403_),
    .Y(_13396_));
 NOR2x2_ASAP7_75t_R _19126_ (.A(_13395_),
    .B(_13396_),
    .Y(_13397_));
 BUFx12f_ASAP7_75t_R _19127_ (.A(_13382_),
    .Y(_13398_));
 INVx5_ASAP7_75t_R _19128_ (.A(net2014),
    .Y(_13399_));
 AND2x2_ASAP7_75t_R _19129_ (.A(net2001),
    .B(_13376_),
    .Y(_13400_));
 NOR2x1_ASAP7_75t_R _19130_ (.A(_13382_),
    .B(_13376_),
    .Y(_13401_));
 AO31x2_ASAP7_75t_R _19131_ (.A1(_13398_),
    .A2(_13399_),
    .A3(_13400_),
    .B(_13401_),
    .Y(_13402_));
 OR2x4_ASAP7_75t_R _19132_ (.A(_00013_),
    .B(_13380_),
    .Y(_13403_));
 NAND2x1_ASAP7_75t_R _19133_ (.A(_13369_),
    .B(_13383_),
    .Y(_13404_));
 NOR2x1_ASAP7_75t_R _19134_ (.A(_13403_),
    .B(_13404_),
    .Y(_13405_));
 AOI22x1_ASAP7_75t_R _19135_ (.A1(_13394_),
    .A2(_13397_),
    .B1(_13402_),
    .B2(_13405_),
    .Y(_13406_));
 INVx3_ASAP7_75t_R _19136_ (.A(_01456_),
    .Y(_13407_));
 AND2x2_ASAP7_75t_R _19137_ (.A(_01776_),
    .B(_13407_),
    .Y(_13408_));
 OR2x4_ASAP7_75t_R _19138_ (.A(_13369_),
    .B(_13370_),
    .Y(_13409_));
 NAND2x1_ASAP7_75t_R _19139_ (.A(_13391_),
    .B(_13376_),
    .Y(_13410_));
 OR4x1_ASAP7_75t_R _19140_ (.A(_13408_),
    .B(_13409_),
    .C(_13403_),
    .D(_13410_),
    .Y(_13411_));
 BUFx4f_ASAP7_75t_R _19141_ (.A(_13411_),
    .Y(_13412_));
 NAND2x1_ASAP7_75t_R _19142_ (.A(_13361_),
    .B(_13363_),
    .Y(_13413_));
 BUFx6f_ASAP7_75t_R _19143_ (.A(_13413_),
    .Y(_13414_));
 AO21x2_ASAP7_75t_R _19144_ (.A1(_13406_),
    .A2(_13412_),
    .B(_13414_),
    .Y(_13415_));
 NAND2x1_ASAP7_75t_R _19145_ (.A(_13390_),
    .B(_13415_),
    .Y(_13416_));
 BUFx6f_ASAP7_75t_R _19146_ (.A(_00510_),
    .Y(_13417_));
 NAND2x1_ASAP7_75t_R _19147_ (.A(_13369_),
    .B(_13370_),
    .Y(_13418_));
 OR3x1_ASAP7_75t_R _19148_ (.A(_13395_),
    .B(_13418_),
    .C(_13396_),
    .Y(_13419_));
 OR4x2_ASAP7_75t_R _19149_ (.A(_13382_),
    .B(_13383_),
    .C(_13377_),
    .D(_13403_),
    .Y(_13420_));
 AO21x2_ASAP7_75t_R _19150_ (.A1(_13409_),
    .A2(_13419_),
    .B(_13420_),
    .Y(_13421_));
 BUFx4f_ASAP7_75t_R _19151_ (.A(_13381_),
    .Y(_13422_));
 AND3x2_ASAP7_75t_R _19152_ (.A(_13391_),
    .B(_13383_),
    .C(_13422_),
    .Y(_13423_));
 INVx1_ASAP7_75t_R _19153_ (.A(_18763_),
    .Y(_13424_));
 INVx2_ASAP7_75t_R _19154_ (.A(_13359_),
    .Y(_13425_));
 OA211x2_ASAP7_75t_R _19155_ (.A1(_13424_),
    .A2(_13357_),
    .B(_13425_),
    .C(_00399_),
    .Y(_13426_));
 NOR2x2_ASAP7_75t_R _19156_ (.A(_00399_),
    .B(_13362_),
    .Y(_13427_));
 AOI211x1_ASAP7_75t_R _19157_ (.A1(_13373_),
    .A2(_13423_),
    .B(_13426_),
    .C(_13427_),
    .Y(_13428_));
 AND2x2_ASAP7_75t_R _19158_ (.A(_13421_),
    .B(_13428_),
    .Y(_13429_));
 OR3x1_ASAP7_75t_R _19159_ (.A(_13417_),
    .B(_13415_),
    .C(_13429_),
    .Y(_13430_));
 OR2x2_ASAP7_75t_R _19160_ (.A(_13376_),
    .B(_13380_),
    .Y(_13431_));
 OR3x1_ASAP7_75t_R _19161_ (.A(_13375_),
    .B(net2016),
    .C(_13431_),
    .Y(_13432_));
 OR3x4_ASAP7_75t_R _19162_ (.A(net2020),
    .B(_13392_),
    .C(_13432_),
    .Y(_13433_));
 AND2x2_ASAP7_75t_R _19163_ (.A(_13381_),
    .B(_13384_),
    .Y(_13434_));
 AOI211x1_ASAP7_75t_R _19164_ (.A1(_13373_),
    .A2(_13434_),
    .B(_13426_),
    .C(_13427_),
    .Y(_13435_));
 NAND2x1_ASAP7_75t_R _19165_ (.A(_13433_),
    .B(_13435_),
    .Y(_13436_));
 AOI21x1_ASAP7_75t_R _19166_ (.A1(_13416_),
    .A2(_13430_),
    .B(_13436_),
    .Y(_13437_));
 BUFx4f_ASAP7_75t_R _19167_ (.A(_00031_),
    .Y(_13438_));
 INVx2_ASAP7_75t_R _19168_ (.A(_13438_),
    .Y(_13439_));
 NAND3x2_ASAP7_75t_R _19169_ (.B(_13406_),
    .C(_13412_),
    .Y(_13440_),
    .A(_13435_));
 AO211x2_ASAP7_75t_R _19170_ (.A1(_13373_),
    .A2(_13434_),
    .B(_13426_),
    .C(_13427_),
    .Y(_13441_));
 OA211x2_ASAP7_75t_R _19171_ (.A1(_13433_),
    .A2(_13441_),
    .B(_13421_),
    .C(_13428_),
    .Y(_13442_));
 BUFx3_ASAP7_75t_R _19172_ (.A(_13442_),
    .Y(_13443_));
 AND3x1_ASAP7_75t_R _19173_ (.A(_13439_),
    .B(_13440_),
    .C(_13443_),
    .Y(_13444_));
 INVx4_ASAP7_75t_R _19174_ (.A(_00366_),
    .Y(_13445_));
 BUFx6f_ASAP7_75t_R _19175_ (.A(_13445_),
    .Y(_13446_));
 BUFx6f_ASAP7_75t_R _19176_ (.A(_13446_),
    .Y(_13447_));
 BUFx4f_ASAP7_75t_R _19177_ (.A(_01551_),
    .Y(_13448_));
 INVx2_ASAP7_75t_R _19178_ (.A(_13448_),
    .Y(_13449_));
 BUFx6f_ASAP7_75t_R _19179_ (.A(_13449_),
    .Y(_13450_));
 BUFx6f_ASAP7_75t_R _19180_ (.A(_13450_),
    .Y(_13451_));
 INVx5_ASAP7_75t_R _19181_ (.A(_00367_),
    .Y(_13452_));
 BUFx6f_ASAP7_75t_R _19182_ (.A(_13452_),
    .Y(_13453_));
 BUFx10_ASAP7_75t_R _19183_ (.A(_13453_),
    .Y(_13454_));
 BUFx6f_ASAP7_75t_R _19184_ (.A(_01552_),
    .Y(_13455_));
 BUFx12f_ASAP7_75t_R _19185_ (.A(_13455_),
    .Y(_13456_));
 BUFx12f_ASAP7_75t_R _19186_ (.A(_13456_),
    .Y(_13457_));
 BUFx12f_ASAP7_75t_R _19187_ (.A(_13457_),
    .Y(_13458_));
 BUFx2_ASAP7_75t_R clone3 (.A(_13466_),
    .Y(net3));
 INVx1_ASAP7_75t_R _19189_ (.A(_00374_),
    .Y(_13460_));
 BUFx6f_ASAP7_75t_R _19190_ (.A(net2),
    .Y(_13461_));
 BUFx6f_ASAP7_75t_R _19191_ (.A(_13461_),
    .Y(_13462_));
 BUFx6f_ASAP7_75t_R _19192_ (.A(_13462_),
    .Y(_13463_));
 BUFx6f_ASAP7_75t_R _19193_ (.A(_13463_),
    .Y(_13464_));
 NAND2x1_ASAP7_75t_R _19194_ (.A(_13464_),
    .B(_00372_),
    .Y(_13465_));
 INVx2_ASAP7_75t_R _19195_ (.A(_00368_),
    .Y(_13466_));
 BUFx3_ASAP7_75t_R _19196_ (.A(_13466_),
    .Y(_13467_));
 BUFx3_ASAP7_75t_R _19197_ (.A(_13467_),
    .Y(_13468_));
 BUFx6f_ASAP7_75t_R _19198_ (.A(_13468_),
    .Y(_13469_));
 BUFx6f_ASAP7_75t_R _19199_ (.A(_13469_),
    .Y(_13470_));
 OA211x2_ASAP7_75t_R _19200_ (.A1(net12),
    .A2(_13460_),
    .B(_13465_),
    .C(net14),
    .Y(_13471_));
 BUFx6f_ASAP7_75t_R _19201_ (.A(_13462_),
    .Y(_13472_));
 BUFx3_ASAP7_75t_R _19202_ (.A(_13472_),
    .Y(_13473_));
 INVx1_ASAP7_75t_R _19203_ (.A(_00373_),
    .Y(_13474_));
 NAND2x1_ASAP7_75t_R _19204_ (.A(_13464_),
    .B(_00371_),
    .Y(_13475_));
 BUFx3_ASAP7_75t_R _19205_ (.A(_00368_),
    .Y(_13476_));
 BUFx4f_ASAP7_75t_R _19206_ (.A(_13476_),
    .Y(_13477_));
 BUFx6f_ASAP7_75t_R _19207_ (.A(_13477_),
    .Y(_13478_));
 BUFx16f_ASAP7_75t_R _19208_ (.A(_13478_),
    .Y(_13479_));
 OA211x2_ASAP7_75t_R _19209_ (.A1(_13473_),
    .A2(_13474_),
    .B(_13475_),
    .C(_13479_),
    .Y(_13480_));
 OR3x1_ASAP7_75t_R _19210_ (.A(_13454_),
    .B(_13471_),
    .C(_13480_),
    .Y(_13481_));
 BUFx6f_ASAP7_75t_R _19211_ (.A(_00367_),
    .Y(_13482_));
 BUFx6f_ASAP7_75t_R _19212_ (.A(_13482_),
    .Y(_13483_));
 BUFx10_ASAP7_75t_R _19213_ (.A(_13483_),
    .Y(_13484_));
 INVx1_ASAP7_75t_R _19214_ (.A(_00382_),
    .Y(_13485_));
 NAND2x1_ASAP7_75t_R _19215_ (.A(_13464_),
    .B(_00380_),
    .Y(_13486_));
 OA211x2_ASAP7_75t_R _19216_ (.A1(net12),
    .A2(_13485_),
    .B(_13486_),
    .C(net14),
    .Y(_13487_));
 INVx1_ASAP7_75t_R _19217_ (.A(_00381_),
    .Y(_13488_));
 NAND2x1_ASAP7_75t_R _19218_ (.A(_13464_),
    .B(_00379_),
    .Y(_13489_));
 BUFx6f_ASAP7_75t_R _19219_ (.A(_00368_),
    .Y(_13490_));
 BUFx6f_ASAP7_75t_R _19220_ (.A(_13490_),
    .Y(_13491_));
 BUFx6f_ASAP7_75t_R _19221_ (.A(_13491_),
    .Y(_13492_));
 OA211x2_ASAP7_75t_R _19222_ (.A1(_13473_),
    .A2(_13488_),
    .B(_13489_),
    .C(_13492_),
    .Y(_13493_));
 OR3x1_ASAP7_75t_R _19223_ (.A(_13484_),
    .B(_13487_),
    .C(_13493_),
    .Y(_13494_));
 AND3x1_ASAP7_75t_R _19224_ (.A(_13451_),
    .B(_13481_),
    .C(_13494_),
    .Y(_13495_));
 NAND2x2_ASAP7_75t_R _19225_ (.A(_13490_),
    .B(_13389_),
    .Y(_13496_));
 BUFx12_ASAP7_75t_R _19226_ (.A(_13496_),
    .Y(_13497_));
 AND2x2_ASAP7_75t_R _19227_ (.A(_13464_),
    .B(_01803_),
    .Y(_13498_));
 AO21x1_ASAP7_75t_R _19228_ (.A1(_00370_),
    .A2(_13390_),
    .B(_13498_),
    .Y(_13499_));
 OAI22x1_ASAP7_75t_R _19229_ (.A1(_00369_),
    .A2(_13497_),
    .B1(_13499_),
    .B2(_13479_),
    .Y(_13500_));
 INVx1_ASAP7_75t_R _19230_ (.A(_00378_),
    .Y(_13501_));
 BUFx6f_ASAP7_75t_R _19231_ (.A(_13457_),
    .Y(_13502_));
 NAND2x1_ASAP7_75t_R _19232_ (.A(_13502_),
    .B(_00376_),
    .Y(_13503_));
 OA211x2_ASAP7_75t_R _19233_ (.A1(_13473_),
    .A2(_13501_),
    .B(_13503_),
    .C(_13470_),
    .Y(_13504_));
 INVx1_ASAP7_75t_R _19234_ (.A(_00377_),
    .Y(_13505_));
 NAND2x1_ASAP7_75t_R _19235_ (.A(_13502_),
    .B(_00375_),
    .Y(_13506_));
 OA211x2_ASAP7_75t_R _19236_ (.A1(_13473_),
    .A2(_13505_),
    .B(_13506_),
    .C(_13492_),
    .Y(_13507_));
 OR3x1_ASAP7_75t_R _19237_ (.A(_13483_),
    .B(_13504_),
    .C(_13507_),
    .Y(_13508_));
 BUFx6f_ASAP7_75t_R _19238_ (.A(_13448_),
    .Y(_13509_));
 BUFx4f_ASAP7_75t_R _19239_ (.A(_13509_),
    .Y(_13510_));
 BUFx6f_ASAP7_75t_R _19240_ (.A(_13510_),
    .Y(_13511_));
 BUFx6f_ASAP7_75t_R _19241_ (.A(_13511_),
    .Y(_13512_));
 OA211x2_ASAP7_75t_R _19242_ (.A1(_13454_),
    .A2(_13500_),
    .B(_13508_),
    .C(_13512_),
    .Y(_13513_));
 OR3x4_ASAP7_75t_R _19243_ (.A(_13447_),
    .B(_13495_),
    .C(_13513_),
    .Y(_13514_));
 BUFx6f_ASAP7_75t_R _19244_ (.A(_00366_),
    .Y(_13515_));
 BUFx6f_ASAP7_75t_R _19245_ (.A(_13515_),
    .Y(_13516_));
 BUFx6f_ASAP7_75t_R _19246_ (.A(_13516_),
    .Y(_13517_));
 BUFx10_ASAP7_75t_R _19247_ (.A(_13517_),
    .Y(_13518_));
 INVx1_ASAP7_75t_R _19248_ (.A(_00390_),
    .Y(_13519_));
 NAND2x1_ASAP7_75t_R _19249_ (.A(_13464_),
    .B(_00388_),
    .Y(_13520_));
 OA211x2_ASAP7_75t_R _19250_ (.A1(net12),
    .A2(_13519_),
    .B(_13520_),
    .C(net14),
    .Y(_13521_));
 INVx2_ASAP7_75t_R _19251_ (.A(_00389_),
    .Y(_13522_));
 NAND2x1_ASAP7_75t_R _19252_ (.A(_13464_),
    .B(_00387_),
    .Y(_13523_));
 OA211x2_ASAP7_75t_R _19253_ (.A1(_13473_),
    .A2(_13522_),
    .B(_13523_),
    .C(_13492_),
    .Y(_13524_));
 OR3x1_ASAP7_75t_R _19254_ (.A(_13453_),
    .B(_13521_),
    .C(_13524_),
    .Y(_13525_));
 INVx2_ASAP7_75t_R _19255_ (.A(_00398_),
    .Y(_13526_));
 NAND2x1_ASAP7_75t_R _19256_ (.A(_13464_),
    .B(_00396_),
    .Y(_13527_));
 OA211x2_ASAP7_75t_R _19257_ (.A1(_13473_),
    .A2(_13526_),
    .B(_13527_),
    .C(net14),
    .Y(_13528_));
 INVx2_ASAP7_75t_R _19258_ (.A(_00397_),
    .Y(_13529_));
 NAND2x1_ASAP7_75t_R _19259_ (.A(_13502_),
    .B(_00395_),
    .Y(_13530_));
 OA211x2_ASAP7_75t_R _19260_ (.A1(_13473_),
    .A2(_13529_),
    .B(_13530_),
    .C(_13492_),
    .Y(_13531_));
 OR3x1_ASAP7_75t_R _19261_ (.A(_13483_),
    .B(_13528_),
    .C(_13531_),
    .Y(_13532_));
 AND3x1_ASAP7_75t_R _19262_ (.A(_13451_),
    .B(_13525_),
    .C(_13532_),
    .Y(_13533_));
 INVx1_ASAP7_75t_R _19263_ (.A(_00391_),
    .Y(_13534_));
 NOR2x1_ASAP7_75t_R _19264_ (.A(_13473_),
    .B(_00393_),
    .Y(_13535_));
 AO21x1_ASAP7_75t_R _19265_ (.A1(net12),
    .A2(_13534_),
    .B(_13535_),
    .Y(_13536_));
 INVx1_ASAP7_75t_R _19266_ (.A(_00394_),
    .Y(_13537_));
 NAND2x1_ASAP7_75t_R _19267_ (.A(_13464_),
    .B(_00392_),
    .Y(_13538_));
 OA211x2_ASAP7_75t_R _19268_ (.A1(net12),
    .A2(_13537_),
    .B(_13538_),
    .C(_13470_),
    .Y(_13539_));
 AO21x1_ASAP7_75t_R _19269_ (.A1(_13479_),
    .A2(_13536_),
    .B(_13539_),
    .Y(_13540_));
 INVx2_ASAP7_75t_R _19270_ (.A(_00386_),
    .Y(_13541_));
 NAND2x1_ASAP7_75t_R _19271_ (.A(_13502_),
    .B(_00384_),
    .Y(_13542_));
 OA211x2_ASAP7_75t_R _19272_ (.A1(_13473_),
    .A2(_13541_),
    .B(_13542_),
    .C(_13470_),
    .Y(_13543_));
 INVx2_ASAP7_75t_R _19273_ (.A(_00385_),
    .Y(_13544_));
 NAND2x1_ASAP7_75t_R _19274_ (.A(_13502_),
    .B(_00383_),
    .Y(_13545_));
 OA211x2_ASAP7_75t_R _19275_ (.A1(_13473_),
    .A2(_13544_),
    .B(_13545_),
    .C(_13492_),
    .Y(_13546_));
 OR3x1_ASAP7_75t_R _19276_ (.A(_13453_),
    .B(_13543_),
    .C(_13546_),
    .Y(_13547_));
 OA211x2_ASAP7_75t_R _19277_ (.A1(_13484_),
    .A2(_13540_),
    .B(_13547_),
    .C(_13512_),
    .Y(_13548_));
 OR3x4_ASAP7_75t_R _19278_ (.A(_13518_),
    .B(_13533_),
    .C(_13548_),
    .Y(_13549_));
 OR4x1_ASAP7_75t_R _19279_ (.A(net2014),
    .B(_13373_),
    .C(_13379_),
    .D(_13385_),
    .Y(_13550_));
 BUFx6f_ASAP7_75t_R _19280_ (.A(_13550_),
    .Y(_13551_));
 AO21x1_ASAP7_75t_R _19281_ (.A1(_13514_),
    .A2(_13549_),
    .B(_13551_),
    .Y(_13552_));
 OA31x2_ASAP7_75t_R _19282_ (.A1(_13387_),
    .A2(_13437_),
    .A3(_13444_),
    .B1(_13552_),
    .Y(_13553_));
 AND2x6_ASAP7_75t_R _19283_ (.A(_13367_),
    .B(_13553_),
    .Y(_18614_));
 BUFx4f_ASAP7_75t_R _19284_ (.A(_13369_),
    .Y(_13554_));
 INVx2_ASAP7_75t_R _19285_ (.A(_00013_),
    .Y(_13555_));
 NOR2x1_ASAP7_75t_R _19286_ (.A(_13376_),
    .B(_13380_),
    .Y(_13556_));
 BUFx4_ASAP7_75t_R clone51 (.A(net2014),
    .Y(net2013));
 AND3x1_ASAP7_75t_R _19288_ (.A(_13374_),
    .B(_13383_),
    .C(_13398_),
    .Y(_13558_));
 AND4x2_ASAP7_75t_R _19289_ (.A(_13558_),
    .B(_13555_),
    .C(_13556_),
    .D(_13554_),
    .Y(_13559_));
 BUFx4f_ASAP7_75t_R _19290_ (.A(_13395_),
    .Y(_13560_));
 BUFx4f_ASAP7_75t_R _19291_ (.A(_13560_),
    .Y(_13561_));
 INVx1_ASAP7_75t_R _19292_ (.A(_00403_),
    .Y(_13562_));
 BUFx6f_ASAP7_75t_R _19293_ (.A(_13562_),
    .Y(_13563_));
 AND2x2_ASAP7_75t_R _19294_ (.A(_13561_),
    .B(_13563_),
    .Y(_13564_));
 INVx2_ASAP7_75t_R _19295_ (.A(net2000),
    .Y(_13565_));
 BUFx6f_ASAP7_75t_R _19296_ (.A(_13565_),
    .Y(_13566_));
 BUFx6f_ASAP7_75t_R _19297_ (.A(_13566_),
    .Y(_13567_));
 BUFx6f_ASAP7_75t_R _19298_ (.A(_13408_),
    .Y(_13568_));
 BUFx4f_ASAP7_75t_R _19299_ (.A(_13376_),
    .Y(_13569_));
 AND4x2_ASAP7_75t_R _19300_ (.A(_13569_),
    .B(_13371_),
    .C(_13422_),
    .D(_13384_),
    .Y(_13570_));
 AND2x6_ASAP7_75t_R _19301_ (.A(_13568_),
    .B(_13570_),
    .Y(_13571_));
 INVx3_ASAP7_75t_R _19302_ (.A(_13395_),
    .Y(_13572_));
 BUFx4f_ASAP7_75t_R _19303_ (.A(_13572_),
    .Y(_13573_));
 BUFx4f_ASAP7_75t_R _19304_ (.A(_01546_),
    .Y(_13574_));
 BUFx4f_ASAP7_75t_R _19305_ (.A(_13574_),
    .Y(_13575_));
 BUFx4f_ASAP7_75t_R _19306_ (.A(_00402_),
    .Y(_13576_));
 BUFx6f_ASAP7_75t_R _19307_ (.A(_01547_),
    .Y(_13577_));
 BUFx10_ASAP7_75t_R _19308_ (.A(_01548_),
    .Y(_13578_));
 BUFx4f_ASAP7_75t_R _19309_ (.A(_01549_),
    .Y(_13579_));
 AND4x2_ASAP7_75t_R _19310_ (.A(_13576_),
    .B(_13577_),
    .C(_13578_),
    .D(_13579_),
    .Y(_13580_));
 AND2x4_ASAP7_75t_R _19311_ (.A(_13580_),
    .B(_13559_),
    .Y(_13581_));
 AND3x1_ASAP7_75t_R _19312_ (.A(_13573_),
    .B(_13575_),
    .C(_13581_),
    .Y(_13582_));
 OA22x2_ASAP7_75t_R _19313_ (.A1(_13567_),
    .A2(_13561_),
    .B1(_13582_),
    .B2(_13571_),
    .Y(_13583_));
 BUFx6f_ASAP7_75t_R _19314_ (.A(_00403_),
    .Y(_13584_));
 BUFx6f_ASAP7_75t_R _19315_ (.A(_13584_),
    .Y(_13585_));
 AND4x2_ASAP7_75t_R _19316_ (.A(_13554_),
    .B(_13555_),
    .C(_13384_),
    .D(_13556_),
    .Y(_13586_));
 AND2x2_ASAP7_75t_R _19317_ (.A(_13399_),
    .B(_13586_),
    .Y(_13587_));
 AND4x2_ASAP7_75t_R _19318_ (.A(_01547_),
    .B(_01548_),
    .C(_13579_),
    .D(_01550_),
    .Y(_13588_));
 BUFx6f_ASAP7_75t_R _19319_ (.A(_00405_),
    .Y(_13589_));
 AND2x2_ASAP7_75t_R _19320_ (.A(_13576_),
    .B(_13589_),
    .Y(_13590_));
 AND2x2_ASAP7_75t_R _19321_ (.A(_13585_),
    .B(_13575_),
    .Y(_13591_));
 BUFx12f_ASAP7_75t_R _19322_ (.A(_00401_),
    .Y(_13592_));
 BUFx10_ASAP7_75t_R _19323_ (.A(_13592_),
    .Y(_13593_));
 NOR2x2_ASAP7_75t_R _19324_ (.A(_13593_),
    .B(_13560_),
    .Y(_13594_));
 BUFx12f_ASAP7_75t_R _19325_ (.A(_13593_),
    .Y(_13595_));
 BUFx3_ASAP7_75t_R rebuffer46 (.A(_00227_),
    .Y(net2008));
 INVx1_ASAP7_75t_R _19327_ (.A(_13575_),
    .Y(_13597_));
 AND4x1_ASAP7_75t_R _19328_ (.A(_13597_),
    .B(_13561_),
    .C(_13585_),
    .D(_13595_),
    .Y(_13598_));
 AO221x1_ASAP7_75t_R _19329_ (.A1(_13575_),
    .A2(_13564_),
    .B1(_13591_),
    .B2(_13594_),
    .C(_13598_),
    .Y(_13599_));
 AND4x1_ASAP7_75t_R _19330_ (.A(_13587_),
    .B(_13588_),
    .C(_13590_),
    .D(_13599_),
    .Y(_13600_));
 AOI221x1_ASAP7_75t_R _19331_ (.A1(net2006),
    .A2(_13564_),
    .B1(_13583_),
    .B2(_13585_),
    .C(_13600_),
    .Y(_18777_));
 INVx1_ASAP7_75t_R _19332_ (.A(_18777_),
    .Y(_18781_));
 BUFx6f_ASAP7_75t_R _19333_ (.A(_01550_),
    .Y(_13601_));
 INVx2_ASAP7_75t_R _19334_ (.A(_13601_),
    .Y(_13602_));
 AND3x2_ASAP7_75t_R _19335_ (.A(_13593_),
    .B(_13560_),
    .C(_13585_),
    .Y(_13603_));
 AND3x1_ASAP7_75t_R _19336_ (.A(_13577_),
    .B(_13578_),
    .C(_13579_),
    .Y(_13604_));
 AND3x4_ASAP7_75t_R _19337_ (.A(_13576_),
    .B(_13589_),
    .C(_13574_),
    .Y(_13605_));
 AND2x2_ASAP7_75t_R _19338_ (.A(_13604_),
    .B(_13605_),
    .Y(_13606_));
 OA21x2_ASAP7_75t_R _19339_ (.A1(_13602_),
    .A2(_13603_),
    .B(_13606_),
    .Y(_13607_));
 NAND2x2_ASAP7_75t_R _19340_ (.A(_13588_),
    .B(_13590_),
    .Y(_13608_));
 NOR2x1_ASAP7_75t_R _19341_ (.A(_13592_),
    .B(_13574_),
    .Y(_13609_));
 AND3x1_ASAP7_75t_R _19342_ (.A(net2000),
    .B(_13584_),
    .C(_13574_),
    .Y(_13610_));
 OA21x2_ASAP7_75t_R _19343_ (.A1(_13609_),
    .A2(_13610_),
    .B(_13395_),
    .Y(_13611_));
 NAND2x1_ASAP7_75t_R _19344_ (.A(_13584_),
    .B(_13574_),
    .Y(_13612_));
 NOR2x1_ASAP7_75t_R _19345_ (.A(_13584_),
    .B(_13574_),
    .Y(_13613_));
 AO31x2_ASAP7_75t_R _19346_ (.A1(_13592_),
    .A2(_13572_),
    .A3(_13612_),
    .B(_13613_),
    .Y(_13614_));
 NOR3x2_ASAP7_75t_R _19347_ (.B(_13611_),
    .C(_13614_),
    .Y(_13615_),
    .A(_13608_));
 NOR2x1_ASAP7_75t_R _19348_ (.A(_13607_),
    .B(_13615_),
    .Y(_13616_));
 AND2x2_ASAP7_75t_R _19349_ (.A(_13566_),
    .B(_13560_),
    .Y(_13617_));
 AND3x1_ASAP7_75t_R _19350_ (.A(_13576_),
    .B(_13575_),
    .C(_13588_),
    .Y(_13618_));
 OA21x2_ASAP7_75t_R _19351_ (.A1(_13397_),
    .A2(_13617_),
    .B(_13618_),
    .Y(_13619_));
 OAI21x1_ASAP7_75t_R _19352_ (.A1(_13616_),
    .A2(_13619_),
    .B(_13587_),
    .Y(_13620_));
 NAND2x2_ASAP7_75t_R _19353_ (.A(_01776_),
    .B(_13407_),
    .Y(_13621_));
 BUFx4f_ASAP7_75t_R _19354_ (.A(_13621_),
    .Y(_13622_));
 NAND2x2_ASAP7_75t_R _19355_ (.A(_13382_),
    .B(_13383_),
    .Y(_13623_));
 OR4x2_ASAP7_75t_R _19356_ (.A(_13377_),
    .B(_13409_),
    .C(_13403_),
    .D(_13623_),
    .Y(_13624_));
 OR3x1_ASAP7_75t_R _19357_ (.A(_13573_),
    .B(_13622_),
    .C(_13624_),
    .Y(_13625_));
 NAND2x1_ASAP7_75t_R _19358_ (.A(_13573_),
    .B(net2006),
    .Y(_13626_));
 AO21x1_ASAP7_75t_R _19359_ (.A1(_13625_),
    .A2(_13626_),
    .B(_13567_),
    .Y(_13627_));
 AO21x1_ASAP7_75t_R _19360_ (.A1(_13398_),
    .A2(_13392_),
    .B(_13409_),
    .Y(_13628_));
 OR3x1_ASAP7_75t_R _19361_ (.A(_13398_),
    .B(_13383_),
    .C(_13418_),
    .Y(_13629_));
 NAND2x1_ASAP7_75t_R _19362_ (.A(_13569_),
    .B(_13422_),
    .Y(_13630_));
 AOI21x1_ASAP7_75t_R _19363_ (.A1(_13628_),
    .A2(_13629_),
    .B(_13630_),
    .Y(_13631_));
 AND4x1_ASAP7_75t_R _19364_ (.A(_13554_),
    .B(_13383_),
    .C(_13422_),
    .D(_13410_),
    .Y(_13632_));
 NAND2x1_ASAP7_75t_R _19365_ (.A(_13394_),
    .B(_13396_),
    .Y(_13633_));
 OA21x2_ASAP7_75t_R _19366_ (.A1(_13631_),
    .A2(_13632_),
    .B(_13633_),
    .Y(_13634_));
 AND2x2_ASAP7_75t_R _19367_ (.A(_13572_),
    .B(_13584_),
    .Y(_13635_));
 NAND2x2_ASAP7_75t_R _19368_ (.A(_13568_),
    .B(_13570_),
    .Y(_13636_));
 OA21x2_ASAP7_75t_R _19369_ (.A1(_13563_),
    .A2(_13580_),
    .B(_13573_),
    .Y(_13637_));
 NAND3x1_ASAP7_75t_R _19370_ (.A(_13382_),
    .B(_13383_),
    .C(net2014),
    .Y(_13638_));
 OR4x2_ASAP7_75t_R _19371_ (.A(_13375_),
    .B(net2015),
    .C(_13431_),
    .D(_13638_),
    .Y(_13639_));
 OA33x2_ASAP7_75t_R _19372_ (.A1(_13635_),
    .A2(_13636_),
    .A3(_13564_),
    .B1(_13637_),
    .B2(_13639_),
    .B3(_13595_),
    .Y(_13640_));
 AND4x2_ASAP7_75t_R _19373_ (.A(_13620_),
    .B(_13627_),
    .C(_13634_),
    .D(_13640_),
    .Y(_18779_));
 INVx3_ASAP7_75t_R _19374_ (.A(_01544_),
    .Y(\cs_registers_i.pc_id_i[1] ));
 INVx1_ASAP7_75t_R _19375_ (.A(_01532_),
    .Y(_13641_));
 BUFx4f_ASAP7_75t_R _19376_ (.A(_13414_),
    .Y(_13642_));
 AO21x1_ASAP7_75t_R _19377_ (.A1(_13375_),
    .A2(_13569_),
    .B(net2020),
    .Y(_13643_));
 AND3x1_ASAP7_75t_R _19378_ (.A(_13383_),
    .B(_13399_),
    .C(_13643_),
    .Y(_13644_));
 AND4x1_ASAP7_75t_R _19379_ (.A(_13391_),
    .B(_13392_),
    .C(_13569_),
    .D(_13374_),
    .Y(_13645_));
 OA21x2_ASAP7_75t_R _19380_ (.A1(_13384_),
    .A2(_13645_),
    .B(_13554_),
    .Y(_13646_));
 NOR2x2_ASAP7_75t_R _19381_ (.A(_13644_),
    .B(_13646_),
    .Y(_13647_));
 NAND3x2_ASAP7_75t_R _19382_ (.B(_13395_),
    .C(_13584_),
    .Y(_13648_),
    .A(net2005));
 AND2x2_ASAP7_75t_R _19383_ (.A(_13394_),
    .B(_13648_),
    .Y(_13649_));
 OR3x1_ASAP7_75t_R _19384_ (.A(_13554_),
    .B(_13569_),
    .C(_13374_),
    .Y(_13650_));
 OR3x1_ASAP7_75t_R _19385_ (.A(net2005),
    .B(_13623_),
    .C(_13650_),
    .Y(_13651_));
 NAND2x1_ASAP7_75t_R _19386_ (.A(_13422_),
    .B(_13651_),
    .Y(_13652_));
 AND3x1_ASAP7_75t_R _19387_ (.A(_13377_),
    .B(_13393_),
    .C(_13423_),
    .Y(_13653_));
 NAND2x1_ASAP7_75t_R _19388_ (.A(_13398_),
    .B(_13392_),
    .Y(_13654_));
 AND3x1_ASAP7_75t_R _19389_ (.A(_13569_),
    .B(_13371_),
    .C(_13422_),
    .Y(_13655_));
 OA211x2_ASAP7_75t_R _19390_ (.A1(_13392_),
    .A2(_13621_),
    .B(_13654_),
    .C(_13655_),
    .Y(_13656_));
 OR4x1_ASAP7_75t_R _19391_ (.A(_13649_),
    .B(_13652_),
    .C(_13653_),
    .D(_13656_),
    .Y(_13657_));
 BUFx4f_ASAP7_75t_R _19392_ (.A(_13657_),
    .Y(_13658_));
 OAI21x1_ASAP7_75t_R _19393_ (.A1(_13647_),
    .A2(_13658_),
    .B(_13366_),
    .Y(_13659_));
 BUFx10_ASAP7_75t_R _19394_ (.A(_13659_),
    .Y(_13660_));
 AO21x1_ASAP7_75t_R _19395_ (.A1(_13392_),
    .A2(_13393_),
    .B(_13371_),
    .Y(_13661_));
 AO21x1_ASAP7_75t_R _19396_ (.A1(_13377_),
    .A2(net2013),
    .B(net2020),
    .Y(_13662_));
 AO22x1_ASAP7_75t_R _19397_ (.A1(net2020),
    .A2(_13399_),
    .B1(_13662_),
    .B2(_13554_),
    .Y(_13663_));
 AO32x2_ASAP7_75t_R _19398_ (.A1(_13391_),
    .A2(_13569_),
    .A3(_13661_),
    .B1(_13663_),
    .B2(_13383_),
    .Y(_13664_));
 AND4x2_ASAP7_75t_R _19399_ (.A(_13365_),
    .B(_13422_),
    .C(_13633_),
    .D(_13651_),
    .Y(_13665_));
 AND2x2_ASAP7_75t_R _19400_ (.A(_13664_),
    .B(_13665_),
    .Y(_13666_));
 BUFx6f_ASAP7_75t_R _19401_ (.A(_13666_),
    .Y(_13667_));
 BUFx6f_ASAP7_75t_R _19402_ (.A(_00409_),
    .Y(_13668_));
 INVx3_ASAP7_75t_R _19403_ (.A(_13668_),
    .Y(_13669_));
 BUFx6f_ASAP7_75t_R _19404_ (.A(_13669_),
    .Y(_13670_));
 BUFx6f_ASAP7_75t_R _19405_ (.A(_00411_),
    .Y(_13671_));
 BUFx6f_ASAP7_75t_R _19406_ (.A(_13671_),
    .Y(_13672_));
 INVx2_ASAP7_75t_R _19407_ (.A(_13672_),
    .Y(_13673_));
 BUFx10_ASAP7_75t_R _19408_ (.A(_13673_),
    .Y(_13674_));
 INVx4_ASAP7_75t_R _19409_ (.A(_00410_),
    .Y(_13675_));
 BUFx10_ASAP7_75t_R _19410_ (.A(_13675_),
    .Y(_13676_));
 BUFx4f_ASAP7_75t_R _19411_ (.A(_00412_),
    .Y(_13677_));
 BUFx6f_ASAP7_75t_R _19412_ (.A(_13677_),
    .Y(_13678_));
 BUFx12f_ASAP7_75t_R _19413_ (.A(_13678_),
    .Y(_13679_));
 BUFx12f_ASAP7_75t_R _19414_ (.A(_13679_),
    .Y(_13680_));
 BUFx12f_ASAP7_75t_R _19415_ (.A(_13677_),
    .Y(_13681_));
 BUFx12f_ASAP7_75t_R _19416_ (.A(_13681_),
    .Y(_13682_));
 NAND2x1_ASAP7_75t_R _19417_ (.A(_00372_),
    .B(_13682_),
    .Y(_13683_));
 INVx1_ASAP7_75t_R _19418_ (.A(_00413_),
    .Y(_13684_));
 BUFx6f_ASAP7_75t_R _19419_ (.A(_13684_),
    .Y(_13685_));
 BUFx4f_ASAP7_75t_R _19420_ (.A(_13685_),
    .Y(_13686_));
 OA211x2_ASAP7_75t_R _19421_ (.A1(_13460_),
    .A2(_13680_),
    .B(_13683_),
    .C(_13686_),
    .Y(_13687_));
 BUFx10_ASAP7_75t_R _19422_ (.A(_13678_),
    .Y(_13688_));
 BUFx10_ASAP7_75t_R _19423_ (.A(_13688_),
    .Y(_13689_));
 BUFx12f_ASAP7_75t_R _19424_ (.A(_13681_),
    .Y(_13690_));
 NAND2x1_ASAP7_75t_R _19425_ (.A(_00371_),
    .B(_13690_),
    .Y(_13691_));
 BUFx10_ASAP7_75t_R _19426_ (.A(_00413_),
    .Y(_13692_));
 BUFx6f_ASAP7_75t_R _19427_ (.A(_13692_),
    .Y(_13693_));
 OA211x2_ASAP7_75t_R _19428_ (.A1(_13474_),
    .A2(_13689_),
    .B(_13691_),
    .C(_13693_),
    .Y(_13694_));
 OR3x1_ASAP7_75t_R _19429_ (.A(_13676_),
    .B(_13687_),
    .C(_13694_),
    .Y(_13695_));
 BUFx10_ASAP7_75t_R _19430_ (.A(_00410_),
    .Y(_13696_));
 NAND2x1_ASAP7_75t_R _19431_ (.A(_00380_),
    .B(_13690_),
    .Y(_13697_));
 OA211x2_ASAP7_75t_R _19432_ (.A1(_13485_),
    .A2(_13689_),
    .B(_13697_),
    .C(_13686_),
    .Y(_13698_));
 BUFx12_ASAP7_75t_R _19433_ (.A(_13678_),
    .Y(_13699_));
 BUFx10_ASAP7_75t_R _19434_ (.A(_13699_),
    .Y(_13700_));
 BUFx12_ASAP7_75t_R _19435_ (.A(_13681_),
    .Y(_13701_));
 NAND2x1_ASAP7_75t_R _19436_ (.A(_00379_),
    .B(_13701_),
    .Y(_13702_));
 OA211x2_ASAP7_75t_R _19437_ (.A1(_13488_),
    .A2(_13700_),
    .B(_13702_),
    .C(_13693_),
    .Y(_13703_));
 OR3x1_ASAP7_75t_R _19438_ (.A(_13696_),
    .B(_13698_),
    .C(_13703_),
    .Y(_13704_));
 AND3x1_ASAP7_75t_R _19439_ (.A(_13674_),
    .B(_13695_),
    .C(_13704_),
    .Y(_13705_));
 BUFx10_ASAP7_75t_R _19440_ (.A(_13675_),
    .Y(_13706_));
 BUFx6f_ASAP7_75t_R _19441_ (.A(_13706_),
    .Y(_13707_));
 INVx2_ASAP7_75t_R _19442_ (.A(_13677_),
    .Y(_13708_));
 BUFx6f_ASAP7_75t_R _19443_ (.A(_13708_),
    .Y(_13709_));
 NAND2x2_ASAP7_75t_R _19444_ (.A(_13692_),
    .B(_13709_),
    .Y(_13710_));
 BUFx12f_ASAP7_75t_R _19445_ (.A(_13681_),
    .Y(_13711_));
 AND2x2_ASAP7_75t_R _19446_ (.A(_13711_),
    .B(_01803_),
    .Y(_13712_));
 AO21x1_ASAP7_75t_R _19447_ (.A1(_00370_),
    .A2(_13709_),
    .B(_13712_),
    .Y(_13713_));
 BUFx6f_ASAP7_75t_R _19448_ (.A(_13692_),
    .Y(_13714_));
 BUFx10_ASAP7_75t_R _19449_ (.A(_13714_),
    .Y(_13715_));
 BUFx10_ASAP7_75t_R _19450_ (.A(_13715_),
    .Y(_13716_));
 OAI22x1_ASAP7_75t_R _19451_ (.A1(_00369_),
    .A2(_13710_),
    .B1(_13713_),
    .B2(_13716_),
    .Y(_13717_));
 BUFx6f_ASAP7_75t_R _19452_ (.A(_00410_),
    .Y(_13718_));
 BUFx6f_ASAP7_75t_R _19453_ (.A(_13677_),
    .Y(_13719_));
 BUFx12_ASAP7_75t_R _19454_ (.A(_13719_),
    .Y(_13720_));
 BUFx10_ASAP7_75t_R _19455_ (.A(_13720_),
    .Y(_13721_));
 BUFx10_ASAP7_75t_R _19456_ (.A(_13681_),
    .Y(_13722_));
 NAND2x1_ASAP7_75t_R _19457_ (.A(_00376_),
    .B(_13722_),
    .Y(_13723_));
 BUFx6f_ASAP7_75t_R _19458_ (.A(_13685_),
    .Y(_13724_));
 OA211x2_ASAP7_75t_R _19459_ (.A1(_13501_),
    .A2(_13721_),
    .B(_13723_),
    .C(_13724_),
    .Y(_13725_));
 BUFx12_ASAP7_75t_R _19460_ (.A(_13720_),
    .Y(_13726_));
 NAND2x1_ASAP7_75t_R _19461_ (.A(_00375_),
    .B(_13722_),
    .Y(_13727_));
 BUFx6f_ASAP7_75t_R _19462_ (.A(_13692_),
    .Y(_13728_));
 OA211x2_ASAP7_75t_R _19463_ (.A1(_13505_),
    .A2(_13726_),
    .B(_13727_),
    .C(_13728_),
    .Y(_13729_));
 OR3x1_ASAP7_75t_R _19464_ (.A(_13718_),
    .B(_13725_),
    .C(_13729_),
    .Y(_13730_));
 BUFx6f_ASAP7_75t_R _19465_ (.A(_13672_),
    .Y(_13731_));
 OA211x2_ASAP7_75t_R _19466_ (.A1(_13707_),
    .A2(_13717_),
    .B(_13730_),
    .C(_13731_),
    .Y(_13732_));
 OR3x4_ASAP7_75t_R _19467_ (.A(_13670_),
    .B(_13705_),
    .C(_13732_),
    .Y(_13733_));
 BUFx6f_ASAP7_75t_R _19468_ (.A(_13668_),
    .Y(_13734_));
 NAND2x1_ASAP7_75t_R _19469_ (.A(_00388_),
    .B(_13690_),
    .Y(_13735_));
 OA211x2_ASAP7_75t_R _19470_ (.A1(_13519_),
    .A2(_13689_),
    .B(_13735_),
    .C(_13686_),
    .Y(_13736_));
 NAND2x1_ASAP7_75t_R _19471_ (.A(_00387_),
    .B(_13701_),
    .Y(_13737_));
 OA211x2_ASAP7_75t_R _19472_ (.A1(_13522_),
    .A2(_13700_),
    .B(_13737_),
    .C(_13693_),
    .Y(_13738_));
 OR3x1_ASAP7_75t_R _19473_ (.A(_13706_),
    .B(_13736_),
    .C(_13738_),
    .Y(_13739_));
 NAND2x1_ASAP7_75t_R _19474_ (.A(_00396_),
    .B(_13690_),
    .Y(_13740_));
 OA211x2_ASAP7_75t_R _19475_ (.A1(_13526_),
    .A2(_13689_),
    .B(_13740_),
    .C(_13686_),
    .Y(_13741_));
 BUFx12_ASAP7_75t_R _19476_ (.A(_13681_),
    .Y(_13742_));
 NAND2x1_ASAP7_75t_R _19477_ (.A(_00395_),
    .B(_13742_),
    .Y(_13743_));
 BUFx6f_ASAP7_75t_R _19478_ (.A(_13692_),
    .Y(_13744_));
 OA211x2_ASAP7_75t_R _19479_ (.A1(_13529_),
    .A2(_13700_),
    .B(_13743_),
    .C(_13744_),
    .Y(_13745_));
 OR3x1_ASAP7_75t_R _19480_ (.A(_13696_),
    .B(_13741_),
    .C(_13745_),
    .Y(_13746_));
 AND3x1_ASAP7_75t_R _19481_ (.A(_13674_),
    .B(_13739_),
    .C(_13746_),
    .Y(_13747_));
 BUFx10_ASAP7_75t_R _19482_ (.A(_13718_),
    .Y(_13748_));
 BUFx12_ASAP7_75t_R _19483_ (.A(_13744_),
    .Y(_13749_));
 BUFx10_ASAP7_75t_R _19484_ (.A(_13722_),
    .Y(_13750_));
 BUFx12_ASAP7_75t_R _19485_ (.A(_13688_),
    .Y(_13751_));
 NOR2x1_ASAP7_75t_R _19486_ (.A(_00393_),
    .B(_13751_),
    .Y(_13752_));
 AO21x1_ASAP7_75t_R _19487_ (.A1(_13534_),
    .A2(_13750_),
    .B(_13752_),
    .Y(_13753_));
 BUFx12_ASAP7_75t_R _19488_ (.A(_13681_),
    .Y(_13754_));
 BUFx12f_ASAP7_75t_R _19489_ (.A(_13754_),
    .Y(_13755_));
 BUFx12f_ASAP7_75t_R _19490_ (.A(_13720_),
    .Y(_13756_));
 NAND2x1_ASAP7_75t_R _19491_ (.A(_00392_),
    .B(_13756_),
    .Y(_13757_));
 OA211x2_ASAP7_75t_R _19492_ (.A1(_13537_),
    .A2(_13755_),
    .B(_13757_),
    .C(_13686_),
    .Y(_13758_));
 AO21x1_ASAP7_75t_R _19493_ (.A1(_13749_),
    .A2(_13753_),
    .B(_13758_),
    .Y(_13759_));
 NAND2x1_ASAP7_75t_R _19494_ (.A(_00384_),
    .B(_13722_),
    .Y(_13760_));
 BUFx10_ASAP7_75t_R _19495_ (.A(_13685_),
    .Y(_13761_));
 OA211x2_ASAP7_75t_R _19496_ (.A1(_13541_),
    .A2(_13721_),
    .B(_13760_),
    .C(_13761_),
    .Y(_13762_));
 BUFx12f_ASAP7_75t_R _19497_ (.A(_13720_),
    .Y(_13763_));
 NAND2x1_ASAP7_75t_R _19498_ (.A(_00383_),
    .B(_13722_),
    .Y(_13764_));
 OA211x2_ASAP7_75t_R _19499_ (.A1(_13544_),
    .A2(_13763_),
    .B(_13764_),
    .C(_13728_),
    .Y(_13765_));
 OR3x1_ASAP7_75t_R _19500_ (.A(_13706_),
    .B(_13762_),
    .C(_13765_),
    .Y(_13766_));
 OA211x2_ASAP7_75t_R _19501_ (.A1(_13748_),
    .A2(_13759_),
    .B(_13766_),
    .C(_13731_),
    .Y(_13767_));
 OR3x4_ASAP7_75t_R _19502_ (.A(_13734_),
    .B(_13747_),
    .C(_13767_),
    .Y(_13768_));
 AND3x1_ASAP7_75t_R _19503_ (.A(_13667_),
    .B(_13733_),
    .C(_13768_),
    .Y(_13769_));
 OA21x2_ASAP7_75t_R _19504_ (.A1(_13647_),
    .A2(_13658_),
    .B(_13366_),
    .Y(_13770_));
 BUFx4f_ASAP7_75t_R _19505_ (.A(_13664_),
    .Y(_13771_));
 BUFx4f_ASAP7_75t_R _19506_ (.A(_13665_),
    .Y(_13772_));
 AND4x1_ASAP7_75t_R _19507_ (.A(_13377_),
    .B(_13371_),
    .C(_13422_),
    .D(_13384_),
    .Y(_13773_));
 BUFx6f_ASAP7_75t_R _19508_ (.A(_13773_),
    .Y(_13774_));
 AND2x2_ASAP7_75t_R _19509_ (.A(_13648_),
    .B(_13774_),
    .Y(_13775_));
 BUFx4f_ASAP7_75t_R _19510_ (.A(_13775_),
    .Y(_13776_));
 BUFx6f_ASAP7_75t_R _19511_ (.A(_13709_),
    .Y(_13777_));
 AO32x1_ASAP7_75t_R _19512_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(_13771_),
    .A3(_13772_),
    .B1(_13776_),
    .B2(_13777_),
    .Y(_13778_));
 AND2x2_ASAP7_75t_R _19513_ (.A(_13770_),
    .B(_13778_),
    .Y(_13779_));
 AO221x1_ASAP7_75t_R _19514_ (.A1(_13641_),
    .A2(_13642_),
    .B1(_13660_),
    .B2(_13769_),
    .C(_13779_),
    .Y(_13780_));
 BUFx6f_ASAP7_75t_R _19515_ (.A(_13780_),
    .Y(_18613_));
 INVx3_ASAP7_75t_R _19516_ (.A(_18613_),
    .Y(_18615_));
 AND3x2_ASAP7_75t_R _19517_ (.A(_13364_),
    .B(_13386_),
    .C(_13433_),
    .Y(_13781_));
 NAND2x2_ASAP7_75t_R _19518_ (.A(_13429_),
    .B(_13781_),
    .Y(_13782_));
 AND2x2_ASAP7_75t_R _19519_ (.A(_13479_),
    .B(_13415_),
    .Y(_13783_));
 AOI21x1_ASAP7_75t_R _19520_ (.A1(_13406_),
    .A2(_13412_),
    .B(_13414_),
    .Y(_13784_));
 AND2x2_ASAP7_75t_R _19521_ (.A(_00446_),
    .B(_13784_),
    .Y(_13785_));
 OR3x4_ASAP7_75t_R _19522_ (.A(_13782_),
    .B(_13783_),
    .C(_13785_),
    .Y(_13786_));
 NOR2x2_ASAP7_75t_R _19523_ (.A(_13414_),
    .B(_13551_),
    .Y(_13787_));
 BUFx6f_ASAP7_75t_R _19524_ (.A(_13787_),
    .Y(_13788_));
 AND2x2_ASAP7_75t_R _19525_ (.A(_13472_),
    .B(_01814_),
    .Y(_13789_));
 AO21x1_ASAP7_75t_R _19526_ (.A1(_13390_),
    .A2(_00417_),
    .B(_13789_),
    .Y(_13790_));
 OAI22x1_ASAP7_75t_R _19527_ (.A1(_00416_),
    .A2(_13497_),
    .B1(_13790_),
    .B2(_13479_),
    .Y(_13791_));
 INVx1_ASAP7_75t_R _19528_ (.A(_00425_),
    .Y(_13792_));
 NAND2x1_ASAP7_75t_R _19529_ (.A(_13463_),
    .B(_00423_),
    .Y(_13793_));
 BUFx4f_ASAP7_75t_R _19530_ (.A(_13467_),
    .Y(_13794_));
 BUFx6f_ASAP7_75t_R _19531_ (.A(_13794_),
    .Y(_13795_));
 OA211x2_ASAP7_75t_R _19532_ (.A1(_13458_),
    .A2(_13792_),
    .B(_13793_),
    .C(_13795_),
    .Y(_13796_));
 INVx2_ASAP7_75t_R _19533_ (.A(_00424_),
    .Y(_13797_));
 BUFx6f_ASAP7_75t_R _19534_ (.A(_01552_),
    .Y(_13798_));
 BUFx6f_ASAP7_75t_R _19535_ (.A(_13798_),
    .Y(_13799_));
 BUFx6f_ASAP7_75t_R _19536_ (.A(_13799_),
    .Y(_13800_));
 BUFx6f_ASAP7_75t_R _19537_ (.A(_13800_),
    .Y(_13801_));
 NAND2x1_ASAP7_75t_R _19538_ (.A(_13801_),
    .B(_00422_),
    .Y(_13802_));
 OA211x2_ASAP7_75t_R _19539_ (.A1(_13472_),
    .A2(_13797_),
    .B(_13802_),
    .C(_13478_),
    .Y(_13803_));
 OR3x1_ASAP7_75t_R _19540_ (.A(_13483_),
    .B(_13796_),
    .C(_13803_),
    .Y(_13804_));
 OA211x2_ASAP7_75t_R _19541_ (.A1(_13453_),
    .A2(_13791_),
    .B(_13804_),
    .C(_13512_),
    .Y(_13805_));
 INVx1_ASAP7_75t_R _19542_ (.A(_00421_),
    .Y(_13806_));
 NAND2x1_ASAP7_75t_R _19543_ (.A(_13472_),
    .B(_00419_),
    .Y(_13807_));
 OA211x2_ASAP7_75t_R _19544_ (.A1(_13502_),
    .A2(_13806_),
    .B(_13807_),
    .C(_13795_),
    .Y(_13808_));
 INVx1_ASAP7_75t_R _19545_ (.A(_00420_),
    .Y(_13809_));
 NAND2x1_ASAP7_75t_R _19546_ (.A(_13463_),
    .B(_00418_),
    .Y(_13810_));
 OA211x2_ASAP7_75t_R _19547_ (.A1(_13502_),
    .A2(_13809_),
    .B(_13810_),
    .C(_13492_),
    .Y(_13811_));
 OR3x1_ASAP7_75t_R _19548_ (.A(_13453_),
    .B(_13808_),
    .C(_13811_),
    .Y(_13812_));
 INVx1_ASAP7_75t_R _19549_ (.A(_00429_),
    .Y(_13813_));
 NAND2x1_ASAP7_75t_R _19550_ (.A(_13472_),
    .B(_00427_),
    .Y(_13814_));
 OA211x2_ASAP7_75t_R _19551_ (.A1(_13502_),
    .A2(_13813_),
    .B(_13814_),
    .C(_13795_),
    .Y(_13815_));
 INVx1_ASAP7_75t_R _19552_ (.A(_00428_),
    .Y(_13816_));
 NAND2x1_ASAP7_75t_R _19553_ (.A(_13463_),
    .B(_00426_),
    .Y(_13817_));
 OA211x2_ASAP7_75t_R _19554_ (.A1(net17),
    .A2(_13816_),
    .B(_13817_),
    .C(_13478_),
    .Y(_13818_));
 OR3x1_ASAP7_75t_R _19555_ (.A(_13483_),
    .B(_13815_),
    .C(_13818_),
    .Y(_13819_));
 AND3x1_ASAP7_75t_R _19556_ (.A(_13451_),
    .B(_13812_),
    .C(_13819_),
    .Y(_13820_));
 OR3x4_ASAP7_75t_R _19557_ (.A(_13447_),
    .B(_13805_),
    .C(_13820_),
    .Y(_13821_));
 INVx1_ASAP7_75t_R _19558_ (.A(_00437_),
    .Y(_13822_));
 NAND2x1_ASAP7_75t_R _19559_ (.A(_13463_),
    .B(_00435_),
    .Y(_13823_));
 OA211x2_ASAP7_75t_R _19560_ (.A1(net17),
    .A2(_13822_),
    .B(_13823_),
    .C(_13795_),
    .Y(_13824_));
 INVx1_ASAP7_75t_R _19561_ (.A(_00436_),
    .Y(_13825_));
 NAND2x1_ASAP7_75t_R _19562_ (.A(_13463_),
    .B(_00434_),
    .Y(_13826_));
 OA211x2_ASAP7_75t_R _19563_ (.A1(net17),
    .A2(_13825_),
    .B(_13826_),
    .C(_13478_),
    .Y(_13827_));
 OR3x1_ASAP7_75t_R _19564_ (.A(_13453_),
    .B(_13824_),
    .C(_13827_),
    .Y(_13828_));
 INVx2_ASAP7_75t_R _19565_ (.A(_00445_),
    .Y(_13829_));
 NAND2x1_ASAP7_75t_R _19566_ (.A(_13463_),
    .B(_00443_),
    .Y(_13830_));
 OA211x2_ASAP7_75t_R _19567_ (.A1(net17),
    .A2(_13829_),
    .B(_13830_),
    .C(_13795_),
    .Y(_13831_));
 INVx2_ASAP7_75t_R _19568_ (.A(_00444_),
    .Y(_13832_));
 NAND2x1_ASAP7_75t_R _19569_ (.A(_13463_),
    .B(_00442_),
    .Y(_13833_));
 OA211x2_ASAP7_75t_R _19570_ (.A1(net17),
    .A2(_13832_),
    .B(_13833_),
    .C(_13478_),
    .Y(_13834_));
 OR3x1_ASAP7_75t_R _19571_ (.A(_13483_),
    .B(_13831_),
    .C(_13834_),
    .Y(_13835_));
 AND3x1_ASAP7_75t_R _19572_ (.A(_13451_),
    .B(_13828_),
    .C(_13835_),
    .Y(_13836_));
 INVx1_ASAP7_75t_R _19573_ (.A(_00438_),
    .Y(_13837_));
 NOR2x1_ASAP7_75t_R _19574_ (.A(net12),
    .B(_00440_),
    .Y(_13838_));
 AO21x1_ASAP7_75t_R _19575_ (.A1(_13464_),
    .A2(_13837_),
    .B(_13838_),
    .Y(_13839_));
 INVx1_ASAP7_75t_R _19576_ (.A(_00441_),
    .Y(_13840_));
 NAND2x1_ASAP7_75t_R _19577_ (.A(_13472_),
    .B(_00439_),
    .Y(_13841_));
 OA211x2_ASAP7_75t_R _19578_ (.A1(_13502_),
    .A2(_13840_),
    .B(_13841_),
    .C(_13795_),
    .Y(_13842_));
 AO21x1_ASAP7_75t_R _19579_ (.A1(_13479_),
    .A2(_13839_),
    .B(_13842_),
    .Y(_13843_));
 INVx1_ASAP7_75t_R _19580_ (.A(_00433_),
    .Y(_13844_));
 NAND2x1_ASAP7_75t_R _19581_ (.A(_13801_),
    .B(_00431_),
    .Y(_13845_));
 OA211x2_ASAP7_75t_R _19582_ (.A1(_13472_),
    .A2(_13844_),
    .B(_13845_),
    .C(_13795_),
    .Y(_13846_));
 INVx1_ASAP7_75t_R _19583_ (.A(_00432_),
    .Y(_13847_));
 NAND2x1_ASAP7_75t_R _19584_ (.A(_13801_),
    .B(_00430_),
    .Y(_13848_));
 OA211x2_ASAP7_75t_R _19585_ (.A1(_13472_),
    .A2(_13847_),
    .B(_13848_),
    .C(_13478_),
    .Y(_13849_));
 OR3x1_ASAP7_75t_R _19586_ (.A(_13453_),
    .B(_13846_),
    .C(_13849_),
    .Y(_13850_));
 OA211x2_ASAP7_75t_R _19587_ (.A1(_13483_),
    .A2(_13843_),
    .B(_13850_),
    .C(_13512_),
    .Y(_13851_));
 OR3x4_ASAP7_75t_R _19588_ (.A(_13518_),
    .B(_13836_),
    .C(_13851_),
    .Y(_13852_));
 NAND3x2_ASAP7_75t_R _19589_ (.B(_13821_),
    .C(_13852_),
    .Y(_13853_),
    .A(_13788_));
 AND2x2_ASAP7_75t_R _19590_ (.A(_13786_),
    .B(_13853_),
    .Y(_13854_));
 INVx1_ASAP7_75t_R _19591_ (.A(_13854_),
    .Y(_13855_));
 BUFx4f_ASAP7_75t_R _19592_ (.A(_13855_),
    .Y(_18610_));
 BUFx6f_ASAP7_75t_R _19593_ (.A(_13854_),
    .Y(_18608_));
 BUFx12_ASAP7_75t_R _19594_ (.A(_13706_),
    .Y(_13856_));
 BUFx6f_ASAP7_75t_R _19595_ (.A(_13856_),
    .Y(_13857_));
 BUFx10_ASAP7_75t_R _19596_ (.A(_13710_),
    .Y(_13858_));
 BUFx6f_ASAP7_75t_R _19597_ (.A(_13709_),
    .Y(_13859_));
 BUFx12_ASAP7_75t_R _19598_ (.A(_13722_),
    .Y(_13860_));
 AND2x2_ASAP7_75t_R _19599_ (.A(_13860_),
    .B(_01814_),
    .Y(_13861_));
 AO21x1_ASAP7_75t_R _19600_ (.A1(_13859_),
    .A2(_00417_),
    .B(_13861_),
    .Y(_13862_));
 BUFx10_ASAP7_75t_R _19601_ (.A(_13749_),
    .Y(_13863_));
 OAI22x1_ASAP7_75t_R _19602_ (.A1(_00416_),
    .A2(_13858_),
    .B1(_13862_),
    .B2(_13863_),
    .Y(_13864_));
 BUFx6f_ASAP7_75t_R _19603_ (.A(_13701_),
    .Y(_13865_));
 BUFx12_ASAP7_75t_R _19604_ (.A(_13720_),
    .Y(_13866_));
 NAND2x1_ASAP7_75t_R _19605_ (.A(_13866_),
    .B(_00431_),
    .Y(_13867_));
 BUFx6f_ASAP7_75t_R _19606_ (.A(_13685_),
    .Y(_13868_));
 BUFx6f_ASAP7_75t_R _19607_ (.A(_13868_),
    .Y(_13869_));
 OA211x2_ASAP7_75t_R _19608_ (.A1(_13865_),
    .A2(_13844_),
    .B(_13867_),
    .C(_13869_),
    .Y(_13870_));
 BUFx6f_ASAP7_75t_R _19609_ (.A(_13742_),
    .Y(_13871_));
 BUFx12_ASAP7_75t_R _19610_ (.A(_13699_),
    .Y(_13872_));
 NAND2x1_ASAP7_75t_R _19611_ (.A(_13872_),
    .B(_00430_),
    .Y(_13873_));
 BUFx6f_ASAP7_75t_R _19612_ (.A(_13714_),
    .Y(_13874_));
 OA211x2_ASAP7_75t_R _19613_ (.A1(_13871_),
    .A2(_13847_),
    .B(_13873_),
    .C(_13874_),
    .Y(_13875_));
 OR3x1_ASAP7_75t_R _19614_ (.A(_13734_),
    .B(_13870_),
    .C(_13875_),
    .Y(_13876_));
 BUFx6f_ASAP7_75t_R _19615_ (.A(_13731_),
    .Y(_13877_));
 OA211x2_ASAP7_75t_R _19616_ (.A1(_13670_),
    .A2(_13864_),
    .B(_13876_),
    .C(_13877_),
    .Y(_13878_));
 BUFx6f_ASAP7_75t_R _19617_ (.A(_13674_),
    .Y(_13879_));
 BUFx16f_ASAP7_75t_R _19618_ (.A(_13720_),
    .Y(_13880_));
 BUFx6f_ASAP7_75t_R _19619_ (.A(_13880_),
    .Y(_13881_));
 BUFx12f_ASAP7_75t_R _19620_ (.A(_13679_),
    .Y(_13882_));
 NAND2x1_ASAP7_75t_R _19621_ (.A(_13882_),
    .B(_00419_),
    .Y(_13883_));
 BUFx6f_ASAP7_75t_R _19622_ (.A(_13761_),
    .Y(_13884_));
 OA211x2_ASAP7_75t_R _19623_ (.A1(_13881_),
    .A2(_13806_),
    .B(_13883_),
    .C(_13884_),
    .Y(_13885_));
 BUFx12_ASAP7_75t_R _19624_ (.A(_13720_),
    .Y(_13886_));
 BUFx6f_ASAP7_75t_R _19625_ (.A(_13886_),
    .Y(_13887_));
 BUFx12f_ASAP7_75t_R _19626_ (.A(_13679_),
    .Y(_13888_));
 NAND2x1_ASAP7_75t_R _19627_ (.A(_13888_),
    .B(_00418_),
    .Y(_13889_));
 BUFx6f_ASAP7_75t_R _19628_ (.A(_13728_),
    .Y(_13890_));
 OA211x2_ASAP7_75t_R _19629_ (.A1(_13887_),
    .A2(_13809_),
    .B(_13889_),
    .C(_13890_),
    .Y(_13891_));
 OR3x1_ASAP7_75t_R _19630_ (.A(_13670_),
    .B(_13885_),
    .C(_13891_),
    .Y(_13892_));
 NAND2x1_ASAP7_75t_R _19631_ (.A(_13882_),
    .B(_00435_),
    .Y(_13893_));
 OA211x2_ASAP7_75t_R _19632_ (.A1(_13881_),
    .A2(_13822_),
    .B(_13893_),
    .C(_13884_),
    .Y(_13894_));
 BUFx6f_ASAP7_75t_R _19633_ (.A(_13886_),
    .Y(_13895_));
 NAND2x1_ASAP7_75t_R _19634_ (.A(_13755_),
    .B(_00434_),
    .Y(_13896_));
 BUFx6f_ASAP7_75t_R _19635_ (.A(_13714_),
    .Y(_13897_));
 OA211x2_ASAP7_75t_R _19636_ (.A1(_13895_),
    .A2(_13825_),
    .B(_13896_),
    .C(_13897_),
    .Y(_13898_));
 OR3x1_ASAP7_75t_R _19637_ (.A(_13734_),
    .B(_13894_),
    .C(_13898_),
    .Y(_13899_));
 AND3x1_ASAP7_75t_R _19638_ (.A(_13879_),
    .B(_13892_),
    .C(_13899_),
    .Y(_13900_));
 OR3x4_ASAP7_75t_R _19639_ (.A(_13857_),
    .B(_13878_),
    .C(_13900_),
    .Y(_13901_));
 BUFx10_ASAP7_75t_R _19640_ (.A(_13718_),
    .Y(_13902_));
 BUFx6f_ASAP7_75t_R _19641_ (.A(_13902_),
    .Y(_13903_));
 BUFx10_ASAP7_75t_R _19642_ (.A(_13699_),
    .Y(_13904_));
 NAND2x1_ASAP7_75t_R _19643_ (.A(_13904_),
    .B(_00427_),
    .Y(_13905_));
 BUFx6f_ASAP7_75t_R _19644_ (.A(_13761_),
    .Y(_13906_));
 OA211x2_ASAP7_75t_R _19645_ (.A1(_13881_),
    .A2(_13813_),
    .B(_13905_),
    .C(_13906_),
    .Y(_13907_));
 NAND2x1_ASAP7_75t_R _19646_ (.A(_13882_),
    .B(_00426_),
    .Y(_13908_));
 OA211x2_ASAP7_75t_R _19647_ (.A1(_13881_),
    .A2(_13816_),
    .B(_13908_),
    .C(_13890_),
    .Y(_13909_));
 OR3x1_ASAP7_75t_R _19648_ (.A(_13670_),
    .B(_13907_),
    .C(_13909_),
    .Y(_13910_));
 NAND2x1_ASAP7_75t_R _19649_ (.A(_13904_),
    .B(_00443_),
    .Y(_13911_));
 OA211x2_ASAP7_75t_R _19650_ (.A1(_13881_),
    .A2(_13829_),
    .B(_13911_),
    .C(_13906_),
    .Y(_13912_));
 NAND2x1_ASAP7_75t_R _19651_ (.A(_13888_),
    .B(_00442_),
    .Y(_13913_));
 OA211x2_ASAP7_75t_R _19652_ (.A1(_13887_),
    .A2(_13832_),
    .B(_13913_),
    .C(_13890_),
    .Y(_13914_));
 OR3x1_ASAP7_75t_R _19653_ (.A(_13734_),
    .B(_13912_),
    .C(_13914_),
    .Y(_13915_));
 AND3x1_ASAP7_75t_R _19654_ (.A(_13879_),
    .B(_13910_),
    .C(_13915_),
    .Y(_13916_));
 BUFx6f_ASAP7_75t_R _19655_ (.A(_13728_),
    .Y(_13917_));
 BUFx10_ASAP7_75t_R _19656_ (.A(_13917_),
    .Y(_13918_));
 BUFx12f_ASAP7_75t_R _19657_ (.A(_13699_),
    .Y(_13919_));
 BUFx6f_ASAP7_75t_R _19658_ (.A(_13919_),
    .Y(_13920_));
 BUFx10_ASAP7_75t_R _19659_ (.A(_13682_),
    .Y(_13921_));
 NOR2x1_ASAP7_75t_R _19660_ (.A(_13921_),
    .B(_00440_),
    .Y(_13922_));
 AO21x1_ASAP7_75t_R _19661_ (.A1(_13920_),
    .A2(_13837_),
    .B(_13922_),
    .Y(_13923_));
 BUFx6f_ASAP7_75t_R _19662_ (.A(_13721_),
    .Y(_13924_));
 BUFx12_ASAP7_75t_R _19663_ (.A(_13679_),
    .Y(_13925_));
 NAND2x1_ASAP7_75t_R _19664_ (.A(_13925_),
    .B(_00439_),
    .Y(_13926_));
 BUFx6f_ASAP7_75t_R _19665_ (.A(_13761_),
    .Y(_13927_));
 OA211x2_ASAP7_75t_R _19666_ (.A1(_13924_),
    .A2(_13840_),
    .B(_13926_),
    .C(_13927_),
    .Y(_13928_));
 AO21x1_ASAP7_75t_R _19667_ (.A1(_13918_),
    .A2(_13923_),
    .B(_13928_),
    .Y(_13929_));
 BUFx6f_ASAP7_75t_R _19668_ (.A(_13742_),
    .Y(_13930_));
 NAND2x1_ASAP7_75t_R _19669_ (.A(_13872_),
    .B(_00423_),
    .Y(_13931_));
 BUFx6f_ASAP7_75t_R _19670_ (.A(_13868_),
    .Y(_13932_));
 OA211x2_ASAP7_75t_R _19671_ (.A1(_13930_),
    .A2(_13792_),
    .B(_13931_),
    .C(_13932_),
    .Y(_13933_));
 BUFx6f_ASAP7_75t_R _19672_ (.A(_13742_),
    .Y(_13934_));
 BUFx12_ASAP7_75t_R _19673_ (.A(_13688_),
    .Y(_13935_));
 NAND2x1_ASAP7_75t_R _19674_ (.A(_13935_),
    .B(_00422_),
    .Y(_13936_));
 BUFx6f_ASAP7_75t_R _19675_ (.A(_13714_),
    .Y(_13937_));
 OA211x2_ASAP7_75t_R _19676_ (.A1(_13934_),
    .A2(_13797_),
    .B(_13936_),
    .C(_13937_),
    .Y(_13938_));
 OR3x1_ASAP7_75t_R _19677_ (.A(_13670_),
    .B(_13933_),
    .C(_13938_),
    .Y(_13939_));
 OA211x2_ASAP7_75t_R _19678_ (.A1(_13734_),
    .A2(_13929_),
    .B(_13939_),
    .C(_13877_),
    .Y(_13940_));
 OR3x4_ASAP7_75t_R _19679_ (.A(_13903_),
    .B(_13916_),
    .C(_13940_),
    .Y(_13941_));
 NAND2x1_ASAP7_75t_R _19680_ (.A(_13771_),
    .B(_13772_),
    .Y(_13942_));
 AO21x1_ASAP7_75t_R _19681_ (.A1(_13901_),
    .A2(_13941_),
    .B(_13942_),
    .Y(_13943_));
 NAND2x1_ASAP7_75t_R _19682_ (.A(_01543_),
    .B(_13942_),
    .Y(_13944_));
 BUFx6f_ASAP7_75t_R _19683_ (.A(_13724_),
    .Y(_13945_));
 AND4x1_ASAP7_75t_R _19684_ (.A(_13945_),
    .B(_13770_),
    .C(_13942_),
    .D(_13776_),
    .Y(_13946_));
 AO31x2_ASAP7_75t_R _19685_ (.A1(_13660_),
    .A2(_13943_),
    .A3(_13944_),
    .B(_13946_),
    .Y(_18609_));
 INVx3_ASAP7_75t_R _19686_ (.A(_18609_),
    .Y(_18611_));
 XOR2x2_ASAP7_75t_R _19687_ (.A(_00415_),
    .B(_02229_),
    .Y(\alu_adder_result_ex[1] ));
 CKINVDCx10_ASAP7_75t_R _19688_ (.A(\alu_adder_result_ex[1] ),
    .Y(_18764_));
 BUFx10_ASAP7_75t_R _19689_ (.A(_13659_),
    .Y(_13947_));
 BUFx12_ASAP7_75t_R _19690_ (.A(_13710_),
    .Y(_13948_));
 AND2x2_ASAP7_75t_R _19691_ (.A(_13886_),
    .B(_01811_),
    .Y(_13949_));
 AO21x1_ASAP7_75t_R _19692_ (.A1(_13709_),
    .A2(_00450_),
    .B(_13949_),
    .Y(_13950_));
 OAI22x1_ASAP7_75t_R _19693_ (.A1(_00449_),
    .A2(_13948_),
    .B1(_13950_),
    .B2(_13716_),
    .Y(_13951_));
 BUFx12f_ASAP7_75t_R _19694_ (.A(_13688_),
    .Y(_13952_));
 INVx1_ASAP7_75t_R _19695_ (.A(_00466_),
    .Y(_13953_));
 NAND2x1_ASAP7_75t_R _19696_ (.A(_13754_),
    .B(_00464_),
    .Y(_13954_));
 OA211x2_ASAP7_75t_R _19697_ (.A1(_13952_),
    .A2(_13953_),
    .B(_13954_),
    .C(_13724_),
    .Y(_13955_));
 BUFx10_ASAP7_75t_R _19698_ (.A(_13688_),
    .Y(_13956_));
 INVx1_ASAP7_75t_R _19699_ (.A(_00465_),
    .Y(_13957_));
 NAND2x1_ASAP7_75t_R _19700_ (.A(_13754_),
    .B(_00463_),
    .Y(_13958_));
 OA211x2_ASAP7_75t_R _19701_ (.A1(_13956_),
    .A2(_13957_),
    .B(_13958_),
    .C(_13728_),
    .Y(_13959_));
 OR3x1_ASAP7_75t_R _19702_ (.A(_13668_),
    .B(_13955_),
    .C(_13959_),
    .Y(_13960_));
 BUFx4f_ASAP7_75t_R _19703_ (.A(_13731_),
    .Y(_13961_));
 OA211x2_ASAP7_75t_R _19704_ (.A1(_13670_),
    .A2(_13951_),
    .B(_13960_),
    .C(_13961_),
    .Y(_13962_));
 INVx1_ASAP7_75t_R _19705_ (.A(_00454_),
    .Y(_13963_));
 BUFx6f_ASAP7_75t_R _19706_ (.A(_13681_),
    .Y(_13964_));
 NAND2x1_ASAP7_75t_R _19707_ (.A(_13964_),
    .B(_00452_),
    .Y(_13965_));
 OA211x2_ASAP7_75t_R _19708_ (.A1(_13680_),
    .A2(_13963_),
    .B(_13965_),
    .C(_13686_),
    .Y(_13966_));
 INVx1_ASAP7_75t_R _19709_ (.A(_00453_),
    .Y(_13967_));
 NAND2x1_ASAP7_75t_R _19710_ (.A(_13964_),
    .B(_00451_),
    .Y(_13968_));
 OA211x2_ASAP7_75t_R _19711_ (.A1(_13689_),
    .A2(_13967_),
    .B(_13968_),
    .C(_13744_),
    .Y(_13969_));
 OR3x1_ASAP7_75t_R _19712_ (.A(_13669_),
    .B(_13966_),
    .C(_13969_),
    .Y(_13970_));
 INVx1_ASAP7_75t_R _19713_ (.A(_00470_),
    .Y(_13971_));
 NAND2x1_ASAP7_75t_R _19714_ (.A(_13964_),
    .B(_00468_),
    .Y(_13972_));
 OA211x2_ASAP7_75t_R _19715_ (.A1(_13689_),
    .A2(_13971_),
    .B(_13972_),
    .C(_13686_),
    .Y(_13973_));
 INVx1_ASAP7_75t_R _19716_ (.A(_00469_),
    .Y(_13974_));
 NAND2x1_ASAP7_75t_R _19717_ (.A(_13964_),
    .B(_00467_),
    .Y(_13975_));
 OA211x2_ASAP7_75t_R _19718_ (.A1(_13700_),
    .A2(_13974_),
    .B(_13975_),
    .C(_13744_),
    .Y(_13976_));
 OR3x1_ASAP7_75t_R _19719_ (.A(_13668_),
    .B(_13973_),
    .C(_13976_),
    .Y(_13977_));
 AND3x1_ASAP7_75t_R _19720_ (.A(_13674_),
    .B(_13970_),
    .C(_13977_),
    .Y(_13978_));
 OR3x4_ASAP7_75t_R _19721_ (.A(_13857_),
    .B(_13962_),
    .C(_13978_),
    .Y(_13979_));
 BUFx3_ASAP7_75t_R _19722_ (.A(_13671_),
    .Y(_13980_));
 BUFx4f_ASAP7_75t_R _19723_ (.A(_13980_),
    .Y(_13981_));
 INVx1_ASAP7_75t_R _19724_ (.A(_00462_),
    .Y(_13982_));
 NAND2x1_ASAP7_75t_R _19725_ (.A(_13981_),
    .B(_00458_),
    .Y(_13983_));
 OA211x2_ASAP7_75t_R _19726_ (.A1(_13981_),
    .A2(_13982_),
    .B(_13983_),
    .C(_13686_),
    .Y(_13984_));
 INVx1_ASAP7_75t_R _19727_ (.A(_00461_),
    .Y(_13985_));
 NAND2x1_ASAP7_75t_R _19728_ (.A(_13672_),
    .B(_00457_),
    .Y(_13986_));
 OA211x2_ASAP7_75t_R _19729_ (.A1(_13981_),
    .A2(_13985_),
    .B(_13986_),
    .C(_13693_),
    .Y(_13987_));
 OR3x1_ASAP7_75t_R _19730_ (.A(_13669_),
    .B(_13984_),
    .C(_13987_),
    .Y(_13988_));
 INVx2_ASAP7_75t_R _19731_ (.A(_00478_),
    .Y(_13989_));
 NAND2x1_ASAP7_75t_R _19732_ (.A(_13981_),
    .B(_00474_),
    .Y(_13990_));
 OA211x2_ASAP7_75t_R _19733_ (.A1(_13981_),
    .A2(_13989_),
    .B(_13990_),
    .C(_13686_),
    .Y(_13991_));
 INVx1_ASAP7_75t_R _19734_ (.A(_00477_),
    .Y(_13992_));
 NAND2x1_ASAP7_75t_R _19735_ (.A(_13672_),
    .B(_00473_),
    .Y(_13993_));
 OA211x2_ASAP7_75t_R _19736_ (.A1(_13981_),
    .A2(_13992_),
    .B(_13993_),
    .C(_13693_),
    .Y(_13994_));
 OR3x1_ASAP7_75t_R _19737_ (.A(_13734_),
    .B(_13991_),
    .C(_13994_),
    .Y(_13995_));
 AND3x1_ASAP7_75t_R _19738_ (.A(_13777_),
    .B(_13988_),
    .C(_13995_),
    .Y(_13996_));
 INVx1_ASAP7_75t_R _19739_ (.A(_00471_),
    .Y(_13997_));
 NOR2x1_ASAP7_75t_R _19740_ (.A(_13981_),
    .B(_00475_),
    .Y(_13998_));
 AO21x1_ASAP7_75t_R _19741_ (.A1(_13731_),
    .A2(_13997_),
    .B(_13998_),
    .Y(_13999_));
 INVx1_ASAP7_75t_R _19742_ (.A(_00476_),
    .Y(_14000_));
 NAND2x1_ASAP7_75t_R _19743_ (.A(_13981_),
    .B(_00472_),
    .Y(_14001_));
 OA211x2_ASAP7_75t_R _19744_ (.A1(_13731_),
    .A2(_14000_),
    .B(_14001_),
    .C(_13686_),
    .Y(_14002_));
 AO21x1_ASAP7_75t_R _19745_ (.A1(_13749_),
    .A2(_13999_),
    .B(_14002_),
    .Y(_14003_));
 INVx1_ASAP7_75t_R _19746_ (.A(_00460_),
    .Y(_14004_));
 NAND2x1_ASAP7_75t_R _19747_ (.A(_13672_),
    .B(_00456_),
    .Y(_14005_));
 OA211x2_ASAP7_75t_R _19748_ (.A1(_13981_),
    .A2(_14004_),
    .B(_14005_),
    .C(_13761_),
    .Y(_14006_));
 INVx1_ASAP7_75t_R _19749_ (.A(_00459_),
    .Y(_14007_));
 NAND2x1_ASAP7_75t_R _19750_ (.A(_13672_),
    .B(_00455_),
    .Y(_14008_));
 OA211x2_ASAP7_75t_R _19751_ (.A1(_13981_),
    .A2(_14007_),
    .B(_14008_),
    .C(_13728_),
    .Y(_14009_));
 OR3x1_ASAP7_75t_R _19752_ (.A(_13669_),
    .B(_14006_),
    .C(_14009_),
    .Y(_14010_));
 BUFx10_ASAP7_75t_R _19753_ (.A(_13680_),
    .Y(_14011_));
 OA211x2_ASAP7_75t_R _19754_ (.A1(_13734_),
    .A2(_14003_),
    .B(_14010_),
    .C(_14011_),
    .Y(_14012_));
 OR3x4_ASAP7_75t_R _19755_ (.A(_13903_),
    .B(_13996_),
    .C(_14012_),
    .Y(_14013_));
 INVx1_ASAP7_75t_R _19756_ (.A(_00044_),
    .Y(_14014_));
 OA211x2_ASAP7_75t_R _19757_ (.A1(_13647_),
    .A2(_13658_),
    .B(_14014_),
    .C(_13366_),
    .Y(_14015_));
 AO31x2_ASAP7_75t_R _19758_ (.A1(_13947_),
    .A2(_13979_),
    .A3(_14013_),
    .B(_14015_),
    .Y(_14016_));
 INVx1_ASAP7_75t_R _19759_ (.A(_01540_),
    .Y(_14017_));
 AO32x1_ASAP7_75t_R _19760_ (.A1(_13771_),
    .A2(_13772_),
    .A3(_14016_),
    .B1(_13642_),
    .B2(_14017_),
    .Y(_14018_));
 BUFx4f_ASAP7_75t_R _19761_ (.A(_14018_),
    .Y(_18667_));
 INVx4_ASAP7_75t_R _19762_ (.A(_18667_),
    .Y(_18669_));
 NAND2x2_ASAP7_75t_R _19763_ (.A(_13592_),
    .B(_13560_),
    .Y(_14019_));
 OA211x2_ASAP7_75t_R _19764_ (.A1(net2005),
    .A2(_13391_),
    .B(_13383_),
    .C(_13422_),
    .Y(_14020_));
 AOI22x1_ASAP7_75t_R _19765_ (.A1(_13423_),
    .A2(_14019_),
    .B1(_14020_),
    .B2(_13563_),
    .Y(_14021_));
 OR3x2_ASAP7_75t_R _19766_ (.A(_13377_),
    .B(_13409_),
    .C(_14021_),
    .Y(_14022_));
 OR4x1_ASAP7_75t_R _19767_ (.A(_13375_),
    .B(net2017),
    .C(_13623_),
    .D(_13431_),
    .Y(_14023_));
 OR3x2_ASAP7_75t_R _19768_ (.A(_13374_),
    .B(_14023_),
    .C(_13606_),
    .Y(_14024_));
 INVx1_ASAP7_75t_R _19769_ (.A(_13380_),
    .Y(_14025_));
 AND5x2_ASAP7_75t_R _19770_ (.A(_13554_),
    .B(_13555_),
    .C(_13376_),
    .D(_14025_),
    .E(_13384_),
    .Y(_14026_));
 NOR2x1_ASAP7_75t_R _19771_ (.A(_13395_),
    .B(_13584_),
    .Y(_14027_));
 OA22x2_ASAP7_75t_R _19772_ (.A1(_13562_),
    .A2(_13399_),
    .B1(_14027_),
    .B2(_13565_),
    .Y(_14028_));
 INVx2_ASAP7_75t_R _19773_ (.A(_01556_),
    .Y(_14029_));
 AOI221x1_ASAP7_75t_R _19774_ (.A1(_13394_),
    .A2(_13396_),
    .B1(_14026_),
    .B2(_14028_),
    .C(_14029_),
    .Y(_14030_));
 NAND2x1_ASAP7_75t_R _19775_ (.A(_13572_),
    .B(_13584_),
    .Y(_14031_));
 OA211x2_ASAP7_75t_R _19776_ (.A1(_13565_),
    .A2(_13575_),
    .B(_13588_),
    .C(_13590_),
    .Y(_14032_));
 OR3x1_ASAP7_75t_R _19777_ (.A(_14031_),
    .B(_13639_),
    .C(_14032_),
    .Y(_14033_));
 OA211x2_ASAP7_75t_R _19778_ (.A1(_13615_),
    .A2(_14024_),
    .B(_14030_),
    .C(_14033_),
    .Y(_14034_));
 BUFx4f_ASAP7_75t_R _19779_ (.A(_13476_),
    .Y(_14035_));
 BUFx6f_ASAP7_75t_R _19780_ (.A(_14035_),
    .Y(_14036_));
 NOR2x2_ASAP7_75t_R _19781_ (.A(_13577_),
    .B(_13578_),
    .Y(_14037_));
 AND2x6_ASAP7_75t_R _19782_ (.A(_13509_),
    .B(_13482_),
    .Y(_14038_));
 AND4x2_ASAP7_75t_R _19783_ (.A(_14036_),
    .B(_13390_),
    .C(_14037_),
    .D(_14038_),
    .Y(_14039_));
 BUFx6f_ASAP7_75t_R _19784_ (.A(_13509_),
    .Y(_14040_));
 BUFx6f_ASAP7_75t_R _19785_ (.A(_14040_),
    .Y(_14041_));
 NOR3x1_ASAP7_75t_R _19786_ (.A(_14036_),
    .B(_14041_),
    .C(_13578_),
    .Y(_14042_));
 BUFx6f_ASAP7_75t_R _19787_ (.A(_13448_),
    .Y(_14043_));
 BUFx6f_ASAP7_75t_R _19788_ (.A(_14043_),
    .Y(_14044_));
 AND2x2_ASAP7_75t_R _19789_ (.A(_14044_),
    .B(_13578_),
    .Y(_14045_));
 AND3x1_ASAP7_75t_R _19790_ (.A(net20),
    .B(_13482_),
    .C(_13577_),
    .Y(_14046_));
 OA21x2_ASAP7_75t_R _19791_ (.A1(_14042_),
    .A2(_14045_),
    .B(_14046_),
    .Y(_14047_));
 AND5x2_ASAP7_75t_R _19792_ (.A(_00413_),
    .B(_13677_),
    .C(_13671_),
    .D(_00410_),
    .E(_13668_),
    .Y(_14048_));
 BUFx6f_ASAP7_75t_R _19793_ (.A(_00034_),
    .Y(_14049_));
 BUFx4f_ASAP7_75t_R _19794_ (.A(_00037_),
    .Y(_14050_));
 AND3x4_ASAP7_75t_R _19795_ (.A(_14049_),
    .B(_14050_),
    .C(_00040_),
    .Y(_14051_));
 AND5x1_ASAP7_75t_R _19796_ (.A(net2005),
    .B(_00446_),
    .C(_13438_),
    .D(_14048_),
    .E(_14051_),
    .Y(_14052_));
 OAI21x1_ASAP7_75t_R _19797_ (.A1(_14039_),
    .A2(_14047_),
    .B(_14052_),
    .Y(_14053_));
 BUFx6f_ASAP7_75t_R _19798_ (.A(_13798_),
    .Y(_14054_));
 BUFx4f_ASAP7_75t_R _19799_ (.A(_14054_),
    .Y(_14055_));
 NAND2x2_ASAP7_75t_R _19800_ (.A(_14043_),
    .B(_13482_),
    .Y(_14056_));
 OR5x2_ASAP7_75t_R _19801_ (.A(_13794_),
    .B(_14055_),
    .C(_13577_),
    .D(_13578_),
    .E(_14056_),
    .Y(_14057_));
 INVx2_ASAP7_75t_R _19802_ (.A(_13576_),
    .Y(_14058_));
 INVx3_ASAP7_75t_R _19803_ (.A(_13589_),
    .Y(_14059_));
 BUFx6f_ASAP7_75t_R _19804_ (.A(_13515_),
    .Y(_14060_));
 OR4x1_ASAP7_75t_R _19805_ (.A(_14060_),
    .B(_13574_),
    .C(_13579_),
    .D(_13601_),
    .Y(_14061_));
 OR3x4_ASAP7_75t_R _19806_ (.A(_14058_),
    .B(_14059_),
    .C(_14061_),
    .Y(_14062_));
 BUFx6f_ASAP7_75t_R _19807_ (.A(_13515_),
    .Y(_14063_));
 AND3x2_ASAP7_75t_R _19808_ (.A(_14063_),
    .B(_13579_),
    .C(_13601_),
    .Y(_14064_));
 NAND2x2_ASAP7_75t_R _19809_ (.A(_13605_),
    .B(_14064_),
    .Y(_14065_));
 OA21x2_ASAP7_75t_R _19810_ (.A1(_14057_),
    .A2(_14062_),
    .B(_14065_),
    .Y(_14066_));
 AND3x1_ASAP7_75t_R _19811_ (.A(_13560_),
    .B(_13584_),
    .C(_13774_),
    .Y(_14067_));
 OAI21x1_ASAP7_75t_R _19812_ (.A1(_14053_),
    .A2(_14066_),
    .B(_14067_),
    .Y(_14068_));
 AND4x2_ASAP7_75t_R _19813_ (.A(_13775_),
    .B(_14022_),
    .C(_14034_),
    .D(_14068_),
    .Y(_14069_));
 BUFx6f_ASAP7_75t_R _19814_ (.A(_14069_),
    .Y(_14070_));
 BUFx6f_ASAP7_75t_R _19815_ (.A(_14070_),
    .Y(_14071_));
 AND2x2_ASAP7_75t_R _19816_ (.A(_18610_),
    .B(_14071_),
    .Y(_18855_));
 INVx1_ASAP7_75t_R _19817_ (.A(_18855_),
    .Y(_18856_));
 NAND2x2_ASAP7_75t_R _19818_ (.A(_18614_),
    .B(_14071_),
    .Y(_18854_));
 INVx1_ASAP7_75t_R _19819_ (.A(_18854_),
    .Y(_18858_));
 BUFx6f_ASAP7_75t_R _19820_ (.A(_13798_),
    .Y(_14072_));
 BUFx4f_ASAP7_75t_R _19821_ (.A(_14072_),
    .Y(_14073_));
 INVx1_ASAP7_75t_R _19822_ (.A(_00505_),
    .Y(_14074_));
 BUFx6f_ASAP7_75t_R _19823_ (.A(_13455_),
    .Y(_14075_));
 NAND2x1_ASAP7_75t_R _19824_ (.A(_14075_),
    .B(_00503_),
    .Y(_14076_));
 OA211x2_ASAP7_75t_R _19825_ (.A1(_14073_),
    .A2(_14074_),
    .B(_14076_),
    .C(_13468_),
    .Y(_14077_));
 INVx1_ASAP7_75t_R _19826_ (.A(_00504_),
    .Y(_14078_));
 BUFx6f_ASAP7_75t_R _19827_ (.A(_13455_),
    .Y(_14079_));
 NAND2x1_ASAP7_75t_R _19828_ (.A(_14079_),
    .B(_00502_),
    .Y(_14080_));
 OA211x2_ASAP7_75t_R _19829_ (.A1(_14073_),
    .A2(_14078_),
    .B(_14080_),
    .C(_14035_),
    .Y(_14081_));
 OR3x1_ASAP7_75t_R _19830_ (.A(_13450_),
    .B(_14077_),
    .C(_14081_),
    .Y(_14082_));
 INVx1_ASAP7_75t_R _19831_ (.A(_00509_),
    .Y(_14083_));
 NAND2x1_ASAP7_75t_R _19832_ (.A(_14075_),
    .B(_00507_),
    .Y(_14084_));
 OA211x2_ASAP7_75t_R _19833_ (.A1(_14073_),
    .A2(_14083_),
    .B(_14084_),
    .C(_13468_),
    .Y(_14085_));
 INVx1_ASAP7_75t_R _19834_ (.A(_00508_),
    .Y(_14086_));
 NAND2x1_ASAP7_75t_R _19835_ (.A(_14079_),
    .B(_00506_),
    .Y(_14087_));
 OA211x2_ASAP7_75t_R _19836_ (.A1(_13800_),
    .A2(_14086_),
    .B(_14087_),
    .C(_14035_),
    .Y(_14088_));
 OR3x1_ASAP7_75t_R _19837_ (.A(_13511_),
    .B(_14085_),
    .C(_14088_),
    .Y(_14089_));
 OR2x2_ASAP7_75t_R _19838_ (.A(_13482_),
    .B(_14060_),
    .Y(_14090_));
 AO21x1_ASAP7_75t_R _19839_ (.A1(_14082_),
    .A2(_14089_),
    .B(_14090_),
    .Y(_14091_));
 BUFx4f_ASAP7_75t_R _19840_ (.A(_14060_),
    .Y(_14092_));
 INVx1_ASAP7_75t_R _19841_ (.A(_00497_),
    .Y(_14093_));
 NAND2x1_ASAP7_75t_R _19842_ (.A(_14079_),
    .B(_00495_),
    .Y(_14094_));
 OA211x2_ASAP7_75t_R _19843_ (.A1(_13800_),
    .A2(_14093_),
    .B(_14094_),
    .C(_13468_),
    .Y(_14095_));
 INVx1_ASAP7_75t_R _19844_ (.A(_00496_),
    .Y(_14096_));
 BUFx6f_ASAP7_75t_R _19845_ (.A(_13455_),
    .Y(_14097_));
 NAND2x1_ASAP7_75t_R _19846_ (.A(_14097_),
    .B(_00494_),
    .Y(_14098_));
 OA211x2_ASAP7_75t_R _19847_ (.A1(_13800_),
    .A2(_14096_),
    .B(_14098_),
    .C(_14035_),
    .Y(_14099_));
 OR3x1_ASAP7_75t_R _19848_ (.A(_14092_),
    .B(_14095_),
    .C(_14099_),
    .Y(_14100_));
 INVx1_ASAP7_75t_R _19849_ (.A(_00480_),
    .Y(_14101_));
 AND2x4_ASAP7_75t_R _19850_ (.A(_13476_),
    .B(_13388_),
    .Y(_14102_));
 BUFx4f_ASAP7_75t_R _19851_ (.A(_13388_),
    .Y(_14103_));
 BUFx6f_ASAP7_75t_R _19852_ (.A(_13455_),
    .Y(_14104_));
 AND2x2_ASAP7_75t_R _19853_ (.A(_14104_),
    .B(_01792_),
    .Y(_14105_));
 AOI21x1_ASAP7_75t_R _19854_ (.A1(_14103_),
    .A2(_00481_),
    .B(_14105_),
    .Y(_14106_));
 AO221x1_ASAP7_75t_R _19855_ (.A1(_14101_),
    .A2(_14102_),
    .B1(_14106_),
    .B2(_13469_),
    .C(_13446_),
    .Y(_14107_));
 AO21x1_ASAP7_75t_R _19856_ (.A1(_14100_),
    .A2(_14107_),
    .B(_14056_),
    .Y(_14108_));
 OR3x4_ASAP7_75t_R _19857_ (.A(_14043_),
    .B(_13452_),
    .C(_13445_),
    .Y(_14109_));
 BUFx6f_ASAP7_75t_R _19858_ (.A(_14079_),
    .Y(_14110_));
 INVx1_ASAP7_75t_R _19859_ (.A(_00484_),
    .Y(_14111_));
 BUFx6f_ASAP7_75t_R _19860_ (.A(_13799_),
    .Y(_14112_));
 NAND2x1_ASAP7_75t_R _19861_ (.A(_14112_),
    .B(_00482_),
    .Y(_14113_));
 OA211x2_ASAP7_75t_R _19862_ (.A1(_14110_),
    .A2(_14111_),
    .B(_14113_),
    .C(_13477_),
    .Y(_14114_));
 INVx1_ASAP7_75t_R _19863_ (.A(_00485_),
    .Y(_14115_));
 NAND2x1_ASAP7_75t_R _19864_ (.A(_13800_),
    .B(_00483_),
    .Y(_14116_));
 BUFx4f_ASAP7_75t_R _19865_ (.A(_13467_),
    .Y(_14117_));
 OA211x2_ASAP7_75t_R _19866_ (.A1(_14110_),
    .A2(_14115_),
    .B(_14116_),
    .C(_14117_),
    .Y(_14118_));
 OR3x4_ASAP7_75t_R _19867_ (.A(_14040_),
    .B(_13452_),
    .C(_14060_),
    .Y(_14119_));
 INVx1_ASAP7_75t_R _19868_ (.A(_00500_),
    .Y(_14120_));
 NAND2x1_ASAP7_75t_R _19869_ (.A(_13800_),
    .B(_00498_),
    .Y(_14121_));
 OA211x2_ASAP7_75t_R _19870_ (.A1(_14110_),
    .A2(_14120_),
    .B(_14121_),
    .C(_13491_),
    .Y(_14122_));
 INVx1_ASAP7_75t_R _19871_ (.A(_00501_),
    .Y(_14123_));
 NAND2x1_ASAP7_75t_R _19872_ (.A(_13800_),
    .B(_00499_),
    .Y(_14124_));
 OA211x2_ASAP7_75t_R _19873_ (.A1(_14110_),
    .A2(_14123_),
    .B(_14124_),
    .C(_14117_),
    .Y(_14125_));
 OA33x2_ASAP7_75t_R _19874_ (.A1(_14109_),
    .A2(_14114_),
    .A3(_14118_),
    .B1(_14119_),
    .B2(_14122_),
    .B3(_14125_),
    .Y(_14126_));
 INVx1_ASAP7_75t_R _19875_ (.A(_00493_),
    .Y(_14127_));
 NOR2x2_ASAP7_75t_R _19876_ (.A(_13490_),
    .B(_14097_),
    .Y(_14128_));
 BUFx6f_ASAP7_75t_R _19877_ (.A(_13509_),
    .Y(_14129_));
 NAND2x1_ASAP7_75t_R _19878_ (.A(_14129_),
    .B(_00489_),
    .Y(_14130_));
 OA211x2_ASAP7_75t_R _19879_ (.A1(_14044_),
    .A2(_14127_),
    .B(_14128_),
    .C(_14130_),
    .Y(_14131_));
 NAND2x2_ASAP7_75t_R _19880_ (.A(_13452_),
    .B(_13516_),
    .Y(_14132_));
 INVx1_ASAP7_75t_R _19881_ (.A(_00490_),
    .Y(_14133_));
 AND2x2_ASAP7_75t_R _19882_ (.A(_13476_),
    .B(_14072_),
    .Y(_14134_));
 NAND2x1_ASAP7_75t_R _19883_ (.A(_14129_),
    .B(_00486_),
    .Y(_14135_));
 OA211x2_ASAP7_75t_R _19884_ (.A1(_14044_),
    .A2(_14133_),
    .B(_14134_),
    .C(_14135_),
    .Y(_14136_));
 BUFx4f_ASAP7_75t_R _19885_ (.A(_13466_),
    .Y(_14137_));
 AND2x2_ASAP7_75t_R _19886_ (.A(_14137_),
    .B(_14079_),
    .Y(_14138_));
 NAND2x1_ASAP7_75t_R _19887_ (.A(_13510_),
    .B(_00487_),
    .Y(_14139_));
 BUFx4f_ASAP7_75t_R _19888_ (.A(_13449_),
    .Y(_14140_));
 NAND2x1_ASAP7_75t_R _19889_ (.A(_14140_),
    .B(_00491_),
    .Y(_14141_));
 INVx1_ASAP7_75t_R _19890_ (.A(_00488_),
    .Y(_14142_));
 NOR2x1_ASAP7_75t_R _19891_ (.A(_14043_),
    .B(_00492_),
    .Y(_14143_));
 AO21x1_ASAP7_75t_R _19892_ (.A1(_14040_),
    .A2(_14142_),
    .B(_14143_),
    .Y(_14144_));
 AO32x1_ASAP7_75t_R _19893_ (.A1(_14138_),
    .A2(_14139_),
    .A3(_14141_),
    .B1(_14144_),
    .B2(_14102_),
    .Y(_14145_));
 OR4x1_ASAP7_75t_R _19894_ (.A(_14131_),
    .B(_14132_),
    .C(_14136_),
    .D(_14145_),
    .Y(_14146_));
 AND4x2_ASAP7_75t_R _19895_ (.A(_14091_),
    .B(_14108_),
    .C(_14126_),
    .D(_14146_),
    .Y(_14147_));
 BUFx6f_ASAP7_75t_R _19896_ (.A(_14147_),
    .Y(_14148_));
 OR2x2_ASAP7_75t_R _19897_ (.A(_13551_),
    .B(_14148_),
    .Y(_14149_));
 NAND2x2_ASAP7_75t_R _19898_ (.A(_13421_),
    .B(_13428_),
    .Y(_14150_));
 AND3x4_ASAP7_75t_R _19899_ (.A(_00510_),
    .B(_13784_),
    .C(_14150_),
    .Y(_14151_));
 AND4x2_ASAP7_75t_R _19900_ (.A(_13451_),
    .B(_13433_),
    .C(_13435_),
    .D(_13415_),
    .Y(_14152_));
 INVx5_ASAP7_75t_R _19901_ (.A(_14049_),
    .Y(_14153_));
 AND3x4_ASAP7_75t_R _19902_ (.A(_14153_),
    .B(_13440_),
    .C(_13443_),
    .Y(_14154_));
 OR4x1_ASAP7_75t_R _19903_ (.A(_13387_),
    .B(_14151_),
    .C(_14152_),
    .D(_14154_),
    .Y(_14155_));
 AO21x1_ASAP7_75t_R _19904_ (.A1(_14149_),
    .A2(_14155_),
    .B(_13414_),
    .Y(_14156_));
 BUFx4f_ASAP7_75t_R _19905_ (.A(_14156_),
    .Y(_18617_));
 INVx2_ASAP7_75t_R _19906_ (.A(_18617_),
    .Y(_18619_));
 AND2x2_ASAP7_75t_R _19907_ (.A(_13456_),
    .B(_01789_),
    .Y(_14157_));
 AO21x1_ASAP7_75t_R _19908_ (.A1(_14103_),
    .A2(_00512_),
    .B(_14157_),
    .Y(_14158_));
 OAI22x1_ASAP7_75t_R _19909_ (.A1(_00511_),
    .A2(_13497_),
    .B1(_14158_),
    .B2(_13478_),
    .Y(_14159_));
 BUFx6f_ASAP7_75t_R _19910_ (.A(_13799_),
    .Y(_14160_));
 INVx1_ASAP7_75t_R _19911_ (.A(_00528_),
    .Y(_14161_));
 NAND2x1_ASAP7_75t_R _19912_ (.A(_13461_),
    .B(_00526_),
    .Y(_14162_));
 OA211x2_ASAP7_75t_R _19913_ (.A1(_14160_),
    .A2(_14161_),
    .B(_14162_),
    .C(_13468_),
    .Y(_14163_));
 BUFx4f_ASAP7_75t_R _19914_ (.A(_13799_),
    .Y(_14164_));
 INVx1_ASAP7_75t_R _19915_ (.A(_00527_),
    .Y(_14165_));
 NAND2x1_ASAP7_75t_R _19916_ (.A(_13461_),
    .B(_00525_),
    .Y(_14166_));
 BUFx4f_ASAP7_75t_R _19917_ (.A(_13476_),
    .Y(_14167_));
 OA211x2_ASAP7_75t_R _19918_ (.A1(_14164_),
    .A2(_14165_),
    .B(_14166_),
    .C(_14167_),
    .Y(_14168_));
 OR3x1_ASAP7_75t_R _19919_ (.A(_14092_),
    .B(_14163_),
    .C(_14168_),
    .Y(_14169_));
 OA211x2_ASAP7_75t_R _19920_ (.A1(_13446_),
    .A2(_14159_),
    .B(_14169_),
    .C(_14038_),
    .Y(_14170_));
 NAND2x1_ASAP7_75t_R _19921_ (.A(_14041_),
    .B(_00533_),
    .Y(_14171_));
 NAND2x1_ASAP7_75t_R _19922_ (.A(_13450_),
    .B(_00537_),
    .Y(_14172_));
 AND2x2_ASAP7_75t_R _19923_ (.A(_14072_),
    .B(_13445_),
    .Y(_14173_));
 NOR2x1_ASAP7_75t_R _19924_ (.A(_13461_),
    .B(_14060_),
    .Y(_14174_));
 INVx1_ASAP7_75t_R _19925_ (.A(_00539_),
    .Y(_14175_));
 NAND2x1_ASAP7_75t_R _19926_ (.A(_14129_),
    .B(_00535_),
    .Y(_14176_));
 OA21x2_ASAP7_75t_R _19927_ (.A1(_14044_),
    .A2(_14175_),
    .B(_14176_),
    .Y(_14177_));
 AO32x1_ASAP7_75t_R _19928_ (.A1(_14171_),
    .A2(_14172_),
    .A3(_14173_),
    .B1(_14174_),
    .B2(_14177_),
    .Y(_14178_));
 NAND2x1_ASAP7_75t_R _19929_ (.A(_14044_),
    .B(_00517_),
    .Y(_14179_));
 NAND2x1_ASAP7_75t_R _19930_ (.A(_13450_),
    .B(_00521_),
    .Y(_14180_));
 AND2x2_ASAP7_75t_R _19931_ (.A(_14072_),
    .B(_13515_),
    .Y(_14181_));
 AND2x2_ASAP7_75t_R _19932_ (.A(_13388_),
    .B(_13515_),
    .Y(_14182_));
 INVx1_ASAP7_75t_R _19933_ (.A(_00523_),
    .Y(_14183_));
 NAND2x1_ASAP7_75t_R _19934_ (.A(_14129_),
    .B(_00519_),
    .Y(_14184_));
 OA21x2_ASAP7_75t_R _19935_ (.A1(_13510_),
    .A2(_14183_),
    .B(_14184_),
    .Y(_14185_));
 AO32x1_ASAP7_75t_R _19936_ (.A1(_14179_),
    .A2(_14180_),
    .A3(_14181_),
    .B1(_14182_),
    .B2(_14185_),
    .Y(_14186_));
 AND2x2_ASAP7_75t_R _19937_ (.A(_00368_),
    .B(_13452_),
    .Y(_14187_));
 OA21x2_ASAP7_75t_R _19938_ (.A1(_14178_),
    .A2(_14186_),
    .B(_14187_),
    .Y(_14188_));
 INVx1_ASAP7_75t_R _19939_ (.A(_00540_),
    .Y(_14189_));
 NAND2x1_ASAP7_75t_R _19940_ (.A(_14060_),
    .B(_00524_),
    .Y(_14190_));
 OA211x2_ASAP7_75t_R _19941_ (.A1(_14063_),
    .A2(_14189_),
    .B(_14190_),
    .C(_14140_),
    .Y(_14191_));
 INVx1_ASAP7_75t_R _19942_ (.A(_00536_),
    .Y(_14192_));
 NAND2x1_ASAP7_75t_R _19943_ (.A(_13515_),
    .B(_00520_),
    .Y(_14193_));
 OA211x2_ASAP7_75t_R _19944_ (.A1(_14063_),
    .A2(_14192_),
    .B(_14193_),
    .C(_14129_),
    .Y(_14194_));
 AND2x2_ASAP7_75t_R _19945_ (.A(_13452_),
    .B(_14128_),
    .Y(_14195_));
 OA21x2_ASAP7_75t_R _19946_ (.A1(_14191_),
    .A2(_14194_),
    .B(_14195_),
    .Y(_14196_));
 BUFx4f_ASAP7_75t_R _19947_ (.A(_01552_),
    .Y(_14197_));
 BUFx4f_ASAP7_75t_R _19948_ (.A(_14197_),
    .Y(_14198_));
 INVx1_ASAP7_75t_R _19949_ (.A(_00532_),
    .Y(_14199_));
 NAND2x1_ASAP7_75t_R _19950_ (.A(_14054_),
    .B(_00530_),
    .Y(_14200_));
 OA211x2_ASAP7_75t_R _19951_ (.A1(_14198_),
    .A2(_14199_),
    .B(_14200_),
    .C(_14137_),
    .Y(_14201_));
 INVx1_ASAP7_75t_R _19952_ (.A(_00531_),
    .Y(_14202_));
 NAND2x1_ASAP7_75t_R _19953_ (.A(_14054_),
    .B(_00529_),
    .Y(_14203_));
 OA211x2_ASAP7_75t_R _19954_ (.A1(_14198_),
    .A2(_14202_),
    .B(_14203_),
    .C(_14167_),
    .Y(_14204_));
 AND3x4_ASAP7_75t_R _19955_ (.A(_13449_),
    .B(_00367_),
    .C(_13445_),
    .Y(_14205_));
 OA21x2_ASAP7_75t_R _19956_ (.A1(_14201_),
    .A2(_14204_),
    .B(_14205_),
    .Y(_14206_));
 INVx1_ASAP7_75t_R _19957_ (.A(_00538_),
    .Y(_14207_));
 NAND2x1_ASAP7_75t_R _19958_ (.A(_13515_),
    .B(_00522_),
    .Y(_14208_));
 OA211x2_ASAP7_75t_R _19959_ (.A1(_14063_),
    .A2(_14207_),
    .B(_14208_),
    .C(_14140_),
    .Y(_14209_));
 INVx1_ASAP7_75t_R _19960_ (.A(_00534_),
    .Y(_14210_));
 NAND2x1_ASAP7_75t_R _19961_ (.A(_13515_),
    .B(_00518_),
    .Y(_14211_));
 OA211x2_ASAP7_75t_R _19962_ (.A1(_14063_),
    .A2(_14210_),
    .B(_14211_),
    .C(_14040_),
    .Y(_14212_));
 AND3x1_ASAP7_75t_R _19963_ (.A(_13468_),
    .B(_14112_),
    .C(_13452_),
    .Y(_14213_));
 OA21x2_ASAP7_75t_R _19964_ (.A1(_14209_),
    .A2(_14212_),
    .B(_14213_),
    .Y(_14214_));
 INVx1_ASAP7_75t_R _19965_ (.A(_00516_),
    .Y(_14215_));
 NAND2x1_ASAP7_75t_R _19966_ (.A(_14054_),
    .B(_00514_),
    .Y(_14216_));
 OA211x2_ASAP7_75t_R _19967_ (.A1(_13456_),
    .A2(_14215_),
    .B(_14216_),
    .C(_14137_),
    .Y(_14217_));
 INVx1_ASAP7_75t_R _19968_ (.A(_00515_),
    .Y(_14218_));
 NAND2x1_ASAP7_75t_R _19969_ (.A(_14054_),
    .B(_00513_),
    .Y(_14219_));
 OA211x2_ASAP7_75t_R _19970_ (.A1(_13456_),
    .A2(_14218_),
    .B(_14219_),
    .C(_14167_),
    .Y(_14220_));
 AND3x4_ASAP7_75t_R _19971_ (.A(_13449_),
    .B(_00367_),
    .C(_13515_),
    .Y(_14221_));
 OA21x2_ASAP7_75t_R _19972_ (.A1(_14217_),
    .A2(_14220_),
    .B(_14221_),
    .Y(_14222_));
 OR4x1_ASAP7_75t_R _19973_ (.A(_14196_),
    .B(_14206_),
    .C(_14214_),
    .D(_14222_),
    .Y(_14223_));
 OR3x2_ASAP7_75t_R _19974_ (.A(_14170_),
    .B(_14188_),
    .C(_14223_),
    .Y(_14224_));
 BUFx6f_ASAP7_75t_R _19975_ (.A(_14224_),
    .Y(_14225_));
 AND2x2_ASAP7_75t_R _19976_ (.A(_13415_),
    .B(_13781_),
    .Y(_14226_));
 INVx1_ASAP7_75t_R _19977_ (.A(_14050_),
    .Y(_14227_));
 AND3x1_ASAP7_75t_R _19978_ (.A(_14227_),
    .B(_13440_),
    .C(_13443_),
    .Y(_14228_));
 AOI221x1_ASAP7_75t_R _19979_ (.A1(_13788_),
    .A2(_14225_),
    .B1(_14226_),
    .B2(_13454_),
    .C(_14228_),
    .Y(_14229_));
 INVx2_ASAP7_75t_R _19980_ (.A(_14229_),
    .Y(_14230_));
 BUFx6f_ASAP7_75t_R _19981_ (.A(_14230_),
    .Y(_18623_));
 BUFx10_ASAP7_75t_R _19982_ (.A(_14229_),
    .Y(_18625_));
 BUFx6f_ASAP7_75t_R _19983_ (.A(_00040_),
    .Y(_14231_));
 INVx4_ASAP7_75t_R _19984_ (.A(_14231_),
    .Y(_14232_));
 AND2x2_ASAP7_75t_R _19985_ (.A(_13440_),
    .B(_13443_),
    .Y(_14233_));
 INVx1_ASAP7_75t_R _19986_ (.A(_00551_),
    .Y(_14234_));
 NOR2x1_ASAP7_75t_R _19987_ (.A(_13516_),
    .B(_00567_),
    .Y(_14235_));
 AO21x1_ASAP7_75t_R _19988_ (.A1(_13516_),
    .A2(_14234_),
    .B(_14235_),
    .Y(_14236_));
 INVx1_ASAP7_75t_R _19989_ (.A(_00569_),
    .Y(_14237_));
 NAND2x1_ASAP7_75t_R _19990_ (.A(_14060_),
    .B(_00553_),
    .Y(_14238_));
 OA211x2_ASAP7_75t_R _19991_ (.A1(_13516_),
    .A2(_14237_),
    .B(_14238_),
    .C(_14103_),
    .Y(_14239_));
 AO21x1_ASAP7_75t_R _19992_ (.A1(_13801_),
    .A2(_14236_),
    .B(_14239_),
    .Y(_14240_));
 INVx2_ASAP7_75t_R _19993_ (.A(_00570_),
    .Y(_14241_));
 NAND2x1_ASAP7_75t_R _19994_ (.A(_14060_),
    .B(_00554_),
    .Y(_14242_));
 OA211x2_ASAP7_75t_R _19995_ (.A1(_14063_),
    .A2(_14241_),
    .B(_14242_),
    .C(_13389_),
    .Y(_14243_));
 INVx1_ASAP7_75t_R _19996_ (.A(_00568_),
    .Y(_14244_));
 NAND2x1_ASAP7_75t_R _19997_ (.A(_14060_),
    .B(_00552_),
    .Y(_14245_));
 OA211x2_ASAP7_75t_R _19998_ (.A1(_14063_),
    .A2(_14244_),
    .B(_14245_),
    .C(_14198_),
    .Y(_14246_));
 OR3x1_ASAP7_75t_R _19999_ (.A(_14036_),
    .B(_14243_),
    .C(_14246_),
    .Y(_14247_));
 NOR2x1_ASAP7_75t_R _20000_ (.A(_13511_),
    .B(_13482_),
    .Y(_14248_));
 OA211x2_ASAP7_75t_R _20001_ (.A1(_13470_),
    .A2(_14240_),
    .B(_14247_),
    .C(_14248_),
    .Y(_14249_));
 AND2x2_ASAP7_75t_R _20002_ (.A(_13456_),
    .B(_01788_),
    .Y(_14250_));
 AO21x1_ASAP7_75t_R _20003_ (.A1(_14103_),
    .A2(_00542_),
    .B(_14250_),
    .Y(_14251_));
 OAI22x1_ASAP7_75t_R _20004_ (.A1(_00541_),
    .A2(_13497_),
    .B1(_14251_),
    .B2(_13478_),
    .Y(_14252_));
 INVx1_ASAP7_75t_R _20005_ (.A(_00558_),
    .Y(_14253_));
 NAND2x1_ASAP7_75t_R _20006_ (.A(_13461_),
    .B(_00556_),
    .Y(_14254_));
 OA211x2_ASAP7_75t_R _20007_ (.A1(_14164_),
    .A2(_14253_),
    .B(_14254_),
    .C(_14137_),
    .Y(_14255_));
 INVx1_ASAP7_75t_R _20008_ (.A(_00557_),
    .Y(_14256_));
 NAND2x1_ASAP7_75t_R _20009_ (.A(_14054_),
    .B(_00555_),
    .Y(_14257_));
 OA211x2_ASAP7_75t_R _20010_ (.A1(_14164_),
    .A2(_14256_),
    .B(_14257_),
    .C(_14167_),
    .Y(_14258_));
 OR3x1_ASAP7_75t_R _20011_ (.A(_14092_),
    .B(_14255_),
    .C(_14258_),
    .Y(_14259_));
 OA211x2_ASAP7_75t_R _20012_ (.A1(_13446_),
    .A2(_14252_),
    .B(_14259_),
    .C(_14038_),
    .Y(_14260_));
 AND2x2_ASAP7_75t_R _20013_ (.A(_13510_),
    .B(_13452_),
    .Y(_14261_));
 BUFx6f_ASAP7_75t_R _20014_ (.A(_14097_),
    .Y(_14262_));
 INVx1_ASAP7_75t_R _20015_ (.A(_00547_),
    .Y(_14263_));
 NOR2x1_ASAP7_75t_R _20016_ (.A(_14112_),
    .B(_00549_),
    .Y(_14264_));
 AO21x1_ASAP7_75t_R _20017_ (.A1(_14262_),
    .A2(_14263_),
    .B(_14264_),
    .Y(_14265_));
 INVx1_ASAP7_75t_R _20018_ (.A(_00550_),
    .Y(_14266_));
 BUFx6f_ASAP7_75t_R _20019_ (.A(net2),
    .Y(_14267_));
 NAND2x1_ASAP7_75t_R _20020_ (.A(_14267_),
    .B(_00548_),
    .Y(_14268_));
 OA211x2_ASAP7_75t_R _20021_ (.A1(_14055_),
    .A2(_14266_),
    .B(_14268_),
    .C(_13794_),
    .Y(_14269_));
 AO21x1_ASAP7_75t_R _20022_ (.A1(_14036_),
    .A2(_14265_),
    .B(_14269_),
    .Y(_14270_));
 INVx1_ASAP7_75t_R _20023_ (.A(_00543_),
    .Y(_14271_));
 NOR2x1_ASAP7_75t_R _20024_ (.A(_14112_),
    .B(_00545_),
    .Y(_14272_));
 AO21x1_ASAP7_75t_R _20025_ (.A1(_14262_),
    .A2(_14271_),
    .B(_14272_),
    .Y(_14273_));
 INVx1_ASAP7_75t_R _20026_ (.A(_00546_),
    .Y(_14274_));
 NAND2x1_ASAP7_75t_R _20027_ (.A(_14104_),
    .B(_00544_),
    .Y(_14275_));
 OA211x2_ASAP7_75t_R _20028_ (.A1(_14055_),
    .A2(_14274_),
    .B(_14275_),
    .C(_13794_),
    .Y(_14276_));
 AO21x1_ASAP7_75t_R _20029_ (.A1(_14036_),
    .A2(_14273_),
    .B(_14276_),
    .Y(_14277_));
 AO32x1_ASAP7_75t_R _20030_ (.A1(_13517_),
    .A2(_14261_),
    .A3(_14270_),
    .B1(_14277_),
    .B2(_14221_),
    .Y(_14278_));
 INVx1_ASAP7_75t_R _20031_ (.A(_00565_),
    .Y(_14279_));
 NAND2x1_ASAP7_75t_R _20032_ (.A(_14104_),
    .B(_00563_),
    .Y(_14280_));
 OA211x2_ASAP7_75t_R _20033_ (.A1(_14073_),
    .A2(_14279_),
    .B(_14280_),
    .C(_14035_),
    .Y(_14281_));
 INVx1_ASAP7_75t_R _20034_ (.A(_00566_),
    .Y(_14282_));
 NAND2x1_ASAP7_75t_R _20035_ (.A(_14104_),
    .B(_00564_),
    .Y(_14283_));
 OA211x2_ASAP7_75t_R _20036_ (.A1(_14073_),
    .A2(_14282_),
    .B(_14283_),
    .C(_13794_),
    .Y(_14284_));
 OA21x2_ASAP7_75t_R _20037_ (.A1(_14281_),
    .A2(_14284_),
    .B(_14261_),
    .Y(_14285_));
 INVx1_ASAP7_75t_R _20038_ (.A(_00561_),
    .Y(_14286_));
 NAND2x1_ASAP7_75t_R _20039_ (.A(_14104_),
    .B(_00559_),
    .Y(_14287_));
 OA211x2_ASAP7_75t_R _20040_ (.A1(_14073_),
    .A2(_14286_),
    .B(_14287_),
    .C(_14035_),
    .Y(_14288_));
 INVx1_ASAP7_75t_R _20041_ (.A(_00562_),
    .Y(_14289_));
 NAND2x1_ASAP7_75t_R _20042_ (.A(_14075_),
    .B(_00560_),
    .Y(_14290_));
 OA211x2_ASAP7_75t_R _20043_ (.A1(_14073_),
    .A2(_14289_),
    .B(_14290_),
    .C(_13794_),
    .Y(_14291_));
 AND2x2_ASAP7_75t_R _20044_ (.A(_14140_),
    .B(_13482_),
    .Y(_14292_));
 OA21x2_ASAP7_75t_R _20045_ (.A1(_14288_),
    .A2(_14291_),
    .B(_14292_),
    .Y(_14293_));
 OA21x2_ASAP7_75t_R _20046_ (.A1(_14285_),
    .A2(_14293_),
    .B(_13446_),
    .Y(_14294_));
 OR4x2_ASAP7_75t_R _20047_ (.A(_14249_),
    .B(_14260_),
    .C(_14278_),
    .D(_14294_),
    .Y(_14295_));
 AND3x1_ASAP7_75t_R _20048_ (.A(_13447_),
    .B(_13415_),
    .C(_13781_),
    .Y(_14296_));
 AOI221x1_ASAP7_75t_R _20049_ (.A1(_14232_),
    .A2(_14233_),
    .B1(_13788_),
    .B2(_14295_),
    .C(_14296_),
    .Y(_14297_));
 INVx4_ASAP7_75t_R _20050_ (.A(_14297_),
    .Y(_14298_));
 BUFx6f_ASAP7_75t_R _20051_ (.A(_14298_),
    .Y(_18629_));
 BUFx6f_ASAP7_75t_R _20052_ (.A(_14297_),
    .Y(_18627_));
 AND2x2_ASAP7_75t_R _20053_ (.A(_14070_),
    .B(_18629_),
    .Y(_18852_));
 BUFx4f_ASAP7_75t_R _20054_ (.A(_02306_),
    .Y(_14299_));
 BUFx4f_ASAP7_75t_R _20055_ (.A(_14299_),
    .Y(_14300_));
 OA21x2_ASAP7_75t_R _20056_ (.A1(_14151_),
    .A2(_14152_),
    .B(_13551_),
    .Y(_14301_));
 AO21x1_ASAP7_75t_R _20057_ (.A1(_13387_),
    .A2(_14148_),
    .B(_14154_),
    .Y(_14302_));
 BUFx4f_ASAP7_75t_R _20058_ (.A(_14227_),
    .Y(_14303_));
 AO31x2_ASAP7_75t_R _20059_ (.A1(_14303_),
    .A2(_13440_),
    .A3(_13443_),
    .B(_13414_),
    .Y(_14304_));
 AO221x2_ASAP7_75t_R _20060_ (.A1(_13788_),
    .A2(_14225_),
    .B1(_14226_),
    .B2(_13454_),
    .C(_14304_),
    .Y(_14305_));
 OA31x2_ASAP7_75t_R _20061_ (.A1(_14301_),
    .A2(_14302_),
    .A3(_14305_),
    .B1(_14069_),
    .Y(_14306_));
 BUFx3_ASAP7_75t_R _20062_ (.A(_14306_),
    .Y(_14307_));
 BUFx4f_ASAP7_75t_R _20063_ (.A(_14307_),
    .Y(_14308_));
 NOR2x2_ASAP7_75t_R _20064_ (.A(_14300_),
    .B(_14308_),
    .Y(_18853_));
 AND5x2_ASAP7_75t_R _20065_ (.A(_13554_),
    .B(_13555_),
    .C(_13383_),
    .D(_14025_),
    .E(_13401_),
    .Y(_14309_));
 AOI21x1_ASAP7_75t_R _20066_ (.A1(_13409_),
    .A2(_13419_),
    .B(_13420_),
    .Y(_14310_));
 AND2x2_ASAP7_75t_R _20067_ (.A(_13373_),
    .B(_13423_),
    .Y(_14311_));
 OR5x1_ASAP7_75t_R _20068_ (.A(_13414_),
    .B(_14309_),
    .C(_13441_),
    .D(_14310_),
    .E(_14311_),
    .Y(_14312_));
 NAND3x1_ASAP7_75t_R _20069_ (.A(_13365_),
    .B(_13406_),
    .C(_13412_),
    .Y(_14313_));
 AO21x2_ASAP7_75t_R _20070_ (.A1(_14312_),
    .A2(_14313_),
    .B(_13787_),
    .Y(_14314_));
 AND2x2_ASAP7_75t_R _20071_ (.A(_13456_),
    .B(_01787_),
    .Y(_14315_));
 AO21x1_ASAP7_75t_R _20072_ (.A1(_14103_),
    .A2(_00574_),
    .B(_14315_),
    .Y(_14316_));
 OAI22x1_ASAP7_75t_R _20073_ (.A1(_00573_),
    .A2(_13497_),
    .B1(_14316_),
    .B2(_14036_),
    .Y(_14317_));
 NAND2x1_ASAP7_75t_R _20074_ (.A(_13517_),
    .B(_14038_),
    .Y(_14318_));
 INVx1_ASAP7_75t_R _20075_ (.A(_00590_),
    .Y(_14319_));
 NAND2x1_ASAP7_75t_R _20076_ (.A(_13461_),
    .B(_00588_),
    .Y(_14320_));
 OA211x2_ASAP7_75t_R _20077_ (.A1(_14164_),
    .A2(_14319_),
    .B(_14320_),
    .C(_14137_),
    .Y(_14321_));
 INVx1_ASAP7_75t_R _20078_ (.A(_00589_),
    .Y(_14322_));
 NAND2x1_ASAP7_75t_R _20079_ (.A(_14054_),
    .B(_00587_),
    .Y(_14323_));
 OA211x2_ASAP7_75t_R _20080_ (.A1(_14198_),
    .A2(_14322_),
    .B(_14323_),
    .C(_14167_),
    .Y(_14324_));
 NAND2x1_ASAP7_75t_R _20081_ (.A(_13445_),
    .B(_14038_),
    .Y(_14325_));
 OR3x1_ASAP7_75t_R _20082_ (.A(_14321_),
    .B(_14324_),
    .C(_14325_),
    .Y(_14326_));
 INVx1_ASAP7_75t_R _20083_ (.A(_00578_),
    .Y(_14327_));
 NAND2x1_ASAP7_75t_R _20084_ (.A(_14072_),
    .B(_00576_),
    .Y(_14328_));
 OA211x2_ASAP7_75t_R _20085_ (.A1(_14104_),
    .A2(_14327_),
    .B(_14328_),
    .C(_14137_),
    .Y(_14329_));
 INVx1_ASAP7_75t_R _20086_ (.A(_00577_),
    .Y(_14330_));
 NAND2x1_ASAP7_75t_R _20087_ (.A(_14072_),
    .B(_00575_),
    .Y(_14331_));
 OA211x2_ASAP7_75t_R _20088_ (.A1(_14267_),
    .A2(_14330_),
    .B(_14331_),
    .C(_13490_),
    .Y(_14332_));
 INVx1_ASAP7_75t_R _20089_ (.A(_00594_),
    .Y(_14333_));
 NAND2x1_ASAP7_75t_R _20090_ (.A(_14072_),
    .B(_00592_),
    .Y(_14334_));
 OA211x2_ASAP7_75t_R _20091_ (.A1(_14267_),
    .A2(_14333_),
    .B(_14334_),
    .C(_14137_),
    .Y(_14335_));
 INVx1_ASAP7_75t_R _20092_ (.A(_00593_),
    .Y(_14336_));
 NAND2x1_ASAP7_75t_R _20093_ (.A(_14072_),
    .B(_00591_),
    .Y(_14337_));
 OA211x2_ASAP7_75t_R _20094_ (.A1(_14267_),
    .A2(_14336_),
    .B(_14337_),
    .C(_13490_),
    .Y(_14338_));
 OA33x2_ASAP7_75t_R _20095_ (.A1(_14109_),
    .A2(_14329_),
    .A3(_14332_),
    .B1(_14335_),
    .B2(_14338_),
    .B3(_14119_),
    .Y(_14339_));
 OA211x2_ASAP7_75t_R _20096_ (.A1(_14317_),
    .A2(_14318_),
    .B(_14326_),
    .C(_14339_),
    .Y(_14340_));
 INVx1_ASAP7_75t_R _20097_ (.A(_00602_),
    .Y(_14341_));
 NAND2x1_ASAP7_75t_R _20098_ (.A(_14040_),
    .B(_00598_),
    .Y(_14342_));
 OA211x2_ASAP7_75t_R _20099_ (.A1(_13510_),
    .A2(_14341_),
    .B(_14342_),
    .C(_13389_),
    .Y(_14343_));
 INVx1_ASAP7_75t_R _20100_ (.A(_00600_),
    .Y(_14344_));
 NAND2x1_ASAP7_75t_R _20101_ (.A(_14043_),
    .B(_00596_),
    .Y(_14345_));
 OA211x2_ASAP7_75t_R _20102_ (.A1(_14129_),
    .A2(_14344_),
    .B(_14345_),
    .C(_14164_),
    .Y(_14346_));
 OA21x2_ASAP7_75t_R _20103_ (.A1(_14343_),
    .A2(_14346_),
    .B(_13469_),
    .Y(_14347_));
 INVx1_ASAP7_75t_R _20104_ (.A(_00597_),
    .Y(_14348_));
 NOR2x1_ASAP7_75t_R _20105_ (.A(_14040_),
    .B(_00601_),
    .Y(_14349_));
 AO21x1_ASAP7_75t_R _20106_ (.A1(_14129_),
    .A2(_14348_),
    .B(_14349_),
    .Y(_14350_));
 OR2x2_ASAP7_75t_R _20107_ (.A(_14043_),
    .B(_00599_),
    .Y(_14351_));
 OAI21x1_ASAP7_75t_R _20108_ (.A1(_13450_),
    .A2(_00595_),
    .B(_14351_),
    .Y(_14352_));
 AO221x1_ASAP7_75t_R _20109_ (.A1(_14102_),
    .A2(_14350_),
    .B1(_14352_),
    .B2(_14134_),
    .C(_14090_),
    .Y(_14353_));
 INVx1_ASAP7_75t_R _20110_ (.A(_00586_),
    .Y(_14354_));
 BUFx6f_ASAP7_75t_R _20111_ (.A(_13798_),
    .Y(_14355_));
 NAND2x1_ASAP7_75t_R _20112_ (.A(_14355_),
    .B(_00584_),
    .Y(_14356_));
 OA211x2_ASAP7_75t_R _20113_ (.A1(_14079_),
    .A2(_14354_),
    .B(_14356_),
    .C(_13467_),
    .Y(_14357_));
 INVx1_ASAP7_75t_R _20114_ (.A(_00585_),
    .Y(_14358_));
 NAND2x1_ASAP7_75t_R _20115_ (.A(_13799_),
    .B(_00583_),
    .Y(_14359_));
 OA211x2_ASAP7_75t_R _20116_ (.A1(_14079_),
    .A2(_14358_),
    .B(_14359_),
    .C(_13490_),
    .Y(_14360_));
 OR4x1_ASAP7_75t_R _20117_ (.A(_14041_),
    .B(_14132_),
    .C(_14357_),
    .D(_14360_),
    .Y(_14361_));
 NAND2x1_ASAP7_75t_R _20118_ (.A(_14129_),
    .B(_13452_),
    .Y(_14362_));
 INVx1_ASAP7_75t_R _20119_ (.A(_00582_),
    .Y(_14363_));
 NAND2x1_ASAP7_75t_R _20120_ (.A(_13799_),
    .B(_00580_),
    .Y(_14364_));
 OA211x2_ASAP7_75t_R _20121_ (.A1(_14079_),
    .A2(_14363_),
    .B(_14364_),
    .C(_13467_),
    .Y(_14365_));
 INVx1_ASAP7_75t_R _20122_ (.A(_00581_),
    .Y(_14366_));
 NAND2x1_ASAP7_75t_R _20123_ (.A(_13799_),
    .B(_00579_),
    .Y(_14367_));
 OA211x2_ASAP7_75t_R _20124_ (.A1(_14097_),
    .A2(_14366_),
    .B(_14367_),
    .C(net4),
    .Y(_14368_));
 OR4x1_ASAP7_75t_R _20125_ (.A(_13445_),
    .B(_14362_),
    .C(_14365_),
    .D(_14368_),
    .Y(_14369_));
 OA211x2_ASAP7_75t_R _20126_ (.A1(_14347_),
    .A2(_14353_),
    .B(_14361_),
    .C(_14369_),
    .Y(_14370_));
 NAND2x2_ASAP7_75t_R _20127_ (.A(_14340_),
    .B(_14370_),
    .Y(_14371_));
 OR2x2_ASAP7_75t_R _20128_ (.A(_13413_),
    .B(_13551_),
    .Y(_14372_));
 BUFx6f_ASAP7_75t_R _20129_ (.A(_14372_),
    .Y(_14373_));
 OAI22x1_ASAP7_75t_R _20130_ (.A1(_13601_),
    .A2(_14314_),
    .B1(_14371_),
    .B2(_14373_),
    .Y(_18632_));
 INVx4_ASAP7_75t_R _20131_ (.A(_18632_),
    .Y(_18634_));
 AND3x1_ASAP7_75t_R _20132_ (.A(_14041_),
    .B(_13482_),
    .C(_14092_),
    .Y(_14374_));
 AND2x2_ASAP7_75t_R _20133_ (.A(_14054_),
    .B(_01786_),
    .Y(_14375_));
 AO21x1_ASAP7_75t_R _20134_ (.A1(_14103_),
    .A2(_00604_),
    .B(_14375_),
    .Y(_14376_));
 OA22x2_ASAP7_75t_R _20135_ (.A1(_00603_),
    .A2(_13496_),
    .B1(_14376_),
    .B2(_13491_),
    .Y(_14377_));
 INVx1_ASAP7_75t_R _20136_ (.A(_00620_),
    .Y(_14378_));
 NAND2x1_ASAP7_75t_R _20137_ (.A(_14097_),
    .B(_00618_),
    .Y(_14379_));
 OA211x2_ASAP7_75t_R _20138_ (.A1(_13800_),
    .A2(_14378_),
    .B(_14379_),
    .C(net16),
    .Y(_14380_));
 INVx1_ASAP7_75t_R _20139_ (.A(_00619_),
    .Y(_14381_));
 NAND2x1_ASAP7_75t_R _20140_ (.A(_14075_),
    .B(_00617_),
    .Y(_14382_));
 OA211x2_ASAP7_75t_R _20141_ (.A1(_14073_),
    .A2(_14381_),
    .B(_14382_),
    .C(_14035_),
    .Y(_14383_));
 NOR2x2_ASAP7_75t_R _20142_ (.A(_14380_),
    .B(_14383_),
    .Y(_14384_));
 AND2x2_ASAP7_75t_R _20143_ (.A(_13446_),
    .B(_14038_),
    .Y(_14385_));
 AND2x2_ASAP7_75t_R _20144_ (.A(_14197_),
    .B(_00622_),
    .Y(_14386_));
 AO211x2_ASAP7_75t_R _20145_ (.A1(_13389_),
    .A2(_00624_),
    .B(_14386_),
    .C(_14167_),
    .Y(_14387_));
 AND2x2_ASAP7_75t_R _20146_ (.A(_14197_),
    .B(_00621_),
    .Y(_14388_));
 AO211x2_ASAP7_75t_R _20147_ (.A1(_13389_),
    .A2(_00623_),
    .B(_14388_),
    .C(_14137_),
    .Y(_14389_));
 AND2x2_ASAP7_75t_R _20148_ (.A(_14197_),
    .B(_00606_),
    .Y(_14390_));
 AO211x2_ASAP7_75t_R _20149_ (.A1(_13389_),
    .A2(_00608_),
    .B(_14390_),
    .C(_14167_),
    .Y(_14391_));
 AND2x2_ASAP7_75t_R _20150_ (.A(_14197_),
    .B(_00605_),
    .Y(_14392_));
 AO211x2_ASAP7_75t_R _20151_ (.A1(_13389_),
    .A2(_00607_),
    .B(_14392_),
    .C(_14137_),
    .Y(_14393_));
 AO33x2_ASAP7_75t_R _20152_ (.A1(_14205_),
    .A2(_14387_),
    .A3(_14389_),
    .B1(_14391_),
    .B2(_14393_),
    .B3(_14221_),
    .Y(_14394_));
 AOI221x1_ASAP7_75t_R _20153_ (.A1(_14374_),
    .A2(_14377_),
    .B1(_14384_),
    .B2(_14385_),
    .C(_14394_),
    .Y(_14395_));
 INVx1_ASAP7_75t_R _20154_ (.A(_00631_),
    .Y(_14396_));
 NAND2x1_ASAP7_75t_R _20155_ (.A(_14355_),
    .B(_00629_),
    .Y(_14397_));
 OA211x2_ASAP7_75t_R _20156_ (.A1(_14075_),
    .A2(_14396_),
    .B(_14397_),
    .C(_14140_),
    .Y(_14398_));
 INVx1_ASAP7_75t_R _20157_ (.A(_00627_),
    .Y(_14399_));
 NAND2x1_ASAP7_75t_R _20158_ (.A(_14355_),
    .B(_00625_),
    .Y(_14400_));
 OA211x2_ASAP7_75t_R _20159_ (.A1(_14075_),
    .A2(_14399_),
    .B(_14400_),
    .C(_14043_),
    .Y(_14401_));
 OR3x1_ASAP7_75t_R _20160_ (.A(_14117_),
    .B(_14398_),
    .C(_14401_),
    .Y(_14402_));
 INVx1_ASAP7_75t_R _20161_ (.A(_00632_),
    .Y(_14403_));
 NAND2x1_ASAP7_75t_R _20162_ (.A(_14355_),
    .B(_00630_),
    .Y(_14404_));
 OA211x2_ASAP7_75t_R _20163_ (.A1(_14075_),
    .A2(_14403_),
    .B(_14404_),
    .C(_14140_),
    .Y(_14405_));
 INVx1_ASAP7_75t_R _20164_ (.A(_00628_),
    .Y(_14406_));
 NAND2x1_ASAP7_75t_R _20165_ (.A(_14355_),
    .B(_00626_),
    .Y(_14407_));
 OA211x2_ASAP7_75t_R _20166_ (.A1(_14079_),
    .A2(_14406_),
    .B(_14407_),
    .C(_14043_),
    .Y(_14408_));
 OR3x1_ASAP7_75t_R _20167_ (.A(_13491_),
    .B(_14405_),
    .C(_14408_),
    .Y(_14409_));
 AO21x1_ASAP7_75t_R _20168_ (.A1(_14402_),
    .A2(_14409_),
    .B(_14090_),
    .Y(_14410_));
 AND2x2_ASAP7_75t_R _20169_ (.A(_13453_),
    .B(_14092_),
    .Y(_14411_));
 AND2x2_ASAP7_75t_R _20170_ (.A(_14129_),
    .B(_00610_),
    .Y(_14412_));
 AOI21x1_ASAP7_75t_R _20171_ (.A1(_13450_),
    .A2(_00614_),
    .B(_14412_),
    .Y(_14413_));
 INVx1_ASAP7_75t_R _20172_ (.A(_00616_),
    .Y(_14414_));
 NAND2x1_ASAP7_75t_R _20173_ (.A(_14040_),
    .B(_00612_),
    .Y(_14415_));
 OA211x2_ASAP7_75t_R _20174_ (.A1(_13510_),
    .A2(_14414_),
    .B(_14128_),
    .C(_14415_),
    .Y(_14416_));
 AOI21x1_ASAP7_75t_R _20175_ (.A1(_14138_),
    .A2(_14413_),
    .B(_14416_),
    .Y(_14417_));
 INVx1_ASAP7_75t_R _20176_ (.A(_00615_),
    .Y(_14418_));
 NAND2x1_ASAP7_75t_R _20177_ (.A(_14129_),
    .B(_00611_),
    .Y(_14419_));
 OA21x2_ASAP7_75t_R _20178_ (.A1(_14044_),
    .A2(_14418_),
    .B(_14419_),
    .Y(_14420_));
 INVx1_ASAP7_75t_R _20179_ (.A(_00613_),
    .Y(_14421_));
 NAND2x1_ASAP7_75t_R _20180_ (.A(_14040_),
    .B(_00609_),
    .Y(_14422_));
 OA211x2_ASAP7_75t_R _20181_ (.A1(_13510_),
    .A2(_14421_),
    .B(_14134_),
    .C(_14422_),
    .Y(_14423_));
 AOI21x1_ASAP7_75t_R _20182_ (.A1(_14102_),
    .A2(_14420_),
    .B(_14423_),
    .Y(_14424_));
 NAND3x2_ASAP7_75t_R _20183_ (.B(_14417_),
    .C(_14424_),
    .Y(_14425_),
    .A(_14411_));
 AND3x4_ASAP7_75t_R _20184_ (.A(_14395_),
    .B(_14410_),
    .C(_14425_),
    .Y(_14426_));
 AND4x1_ASAP7_75t_R _20185_ (.A(_13433_),
    .B(_13435_),
    .C(_13421_),
    .D(_13428_),
    .Y(_14427_));
 AND3x1_ASAP7_75t_R _20186_ (.A(_13365_),
    .B(_13406_),
    .C(_13412_),
    .Y(_14428_));
 OA21x2_ASAP7_75t_R _20187_ (.A1(_14427_),
    .A2(_14428_),
    .B(_14373_),
    .Y(_14429_));
 AO32x1_ASAP7_75t_R _20188_ (.A1(_13365_),
    .A2(_13387_),
    .A3(_14426_),
    .B1(_14429_),
    .B2(_14059_),
    .Y(_14430_));
 BUFx3_ASAP7_75t_R _20189_ (.A(_14430_),
    .Y(_18638_));
 INVx1_ASAP7_75t_R _20190_ (.A(_18638_),
    .Y(_18640_));
 AND2x2_ASAP7_75t_R _20191_ (.A(_13456_),
    .B(_01785_),
    .Y(_14431_));
 AO21x1_ASAP7_75t_R _20192_ (.A1(_14103_),
    .A2(_00634_),
    .B(_14431_),
    .Y(_14432_));
 OAI22x1_ASAP7_75t_R _20193_ (.A1(_00633_),
    .A2(_13497_),
    .B1(_14432_),
    .B2(_14036_),
    .Y(_14433_));
 INVx1_ASAP7_75t_R _20194_ (.A(_00650_),
    .Y(_14434_));
 NAND2x1_ASAP7_75t_R _20195_ (.A(_14112_),
    .B(_00648_),
    .Y(_14435_));
 OA21x2_ASAP7_75t_R _20196_ (.A1(_13462_),
    .A2(_14434_),
    .B(_14435_),
    .Y(_14436_));
 INVx2_ASAP7_75t_R _20197_ (.A(_00649_),
    .Y(_14437_));
 NAND2x1_ASAP7_75t_R _20198_ (.A(_13456_),
    .B(_00647_),
    .Y(_14438_));
 OA211x2_ASAP7_75t_R _20199_ (.A1(_14055_),
    .A2(_14437_),
    .B(_14438_),
    .C(_14035_),
    .Y(_14439_));
 AO21x1_ASAP7_75t_R _20200_ (.A1(_13795_),
    .A2(_14436_),
    .B(_14439_),
    .Y(_14440_));
 INVx1_ASAP7_75t_R _20201_ (.A(_00654_),
    .Y(_14441_));
 NAND2x1_ASAP7_75t_R _20202_ (.A(_13461_),
    .B(_00652_),
    .Y(_14442_));
 OA211x2_ASAP7_75t_R _20203_ (.A1(_14164_),
    .A2(_14441_),
    .B(_14442_),
    .C(net16),
    .Y(_14443_));
 INVx1_ASAP7_75t_R _20204_ (.A(_00653_),
    .Y(_14444_));
 NAND2x1_ASAP7_75t_R _20205_ (.A(_13461_),
    .B(_00651_),
    .Y(_14445_));
 OA211x2_ASAP7_75t_R _20206_ (.A1(_14164_),
    .A2(_14444_),
    .B(_14445_),
    .C(_14167_),
    .Y(_14446_));
 INVx1_ASAP7_75t_R _20207_ (.A(_00638_),
    .Y(_14447_));
 NAND2x1_ASAP7_75t_R _20208_ (.A(_13461_),
    .B(_00636_),
    .Y(_14448_));
 OA211x2_ASAP7_75t_R _20209_ (.A1(_14160_),
    .A2(_14447_),
    .B(_14448_),
    .C(net16),
    .Y(_14449_));
 INVx1_ASAP7_75t_R _20210_ (.A(_00637_),
    .Y(_14450_));
 NAND2x1_ASAP7_75t_R _20211_ (.A(_14097_),
    .B(_00635_),
    .Y(_14451_));
 OA211x2_ASAP7_75t_R _20212_ (.A1(_14112_),
    .A2(_14450_),
    .B(_14451_),
    .C(_14167_),
    .Y(_14452_));
 OA33x2_ASAP7_75t_R _20213_ (.A1(_14119_),
    .A2(_14443_),
    .A3(_14446_),
    .B1(_14449_),
    .B2(_14452_),
    .B3(_14109_),
    .Y(_14453_));
 OA221x2_ASAP7_75t_R _20214_ (.A1(_14318_),
    .A2(_14433_),
    .B1(_14440_),
    .B2(_14325_),
    .C(_14453_),
    .Y(_14454_));
 INVx1_ASAP7_75t_R _20215_ (.A(_00645_),
    .Y(_14455_));
 NAND2x1_ASAP7_75t_R _20216_ (.A(_14267_),
    .B(_00643_),
    .Y(_14456_));
 OA211x2_ASAP7_75t_R _20217_ (.A1(_14055_),
    .A2(_14455_),
    .B(_14456_),
    .C(_14140_),
    .Y(_14457_));
 INVx1_ASAP7_75t_R _20218_ (.A(_00641_),
    .Y(_14458_));
 NAND2x1_ASAP7_75t_R _20219_ (.A(_14267_),
    .B(_00639_),
    .Y(_14459_));
 OA211x2_ASAP7_75t_R _20220_ (.A1(_14055_),
    .A2(_14458_),
    .B(_14459_),
    .C(_13510_),
    .Y(_14460_));
 OR3x1_ASAP7_75t_R _20221_ (.A(_13795_),
    .B(_14457_),
    .C(_14460_),
    .Y(_14461_));
 INVx1_ASAP7_75t_R _20222_ (.A(_00646_),
    .Y(_14462_));
 NAND2x1_ASAP7_75t_R _20223_ (.A(_14267_),
    .B(_00644_),
    .Y(_14463_));
 OA211x2_ASAP7_75t_R _20224_ (.A1(_14055_),
    .A2(_14462_),
    .B(_14463_),
    .C(_14140_),
    .Y(_14464_));
 INVx1_ASAP7_75t_R _20225_ (.A(_00642_),
    .Y(_14465_));
 NAND2x1_ASAP7_75t_R _20226_ (.A(_14267_),
    .B(_00640_),
    .Y(_14466_));
 OA211x2_ASAP7_75t_R _20227_ (.A1(_14055_),
    .A2(_14465_),
    .B(_14466_),
    .C(_13510_),
    .Y(_14467_));
 OR3x1_ASAP7_75t_R _20228_ (.A(_14036_),
    .B(_14464_),
    .C(_14467_),
    .Y(_14468_));
 AO21x1_ASAP7_75t_R _20229_ (.A1(_14461_),
    .A2(_14468_),
    .B(_14132_),
    .Y(_14469_));
 NOR2x2_ASAP7_75t_R _20230_ (.A(_13483_),
    .B(_13517_),
    .Y(_14470_));
 NAND2x1_ASAP7_75t_R _20231_ (.A(_13491_),
    .B(_13450_),
    .Y(_14471_));
 AND2x2_ASAP7_75t_R _20232_ (.A(_14198_),
    .B(_00659_),
    .Y(_14472_));
 AO21x1_ASAP7_75t_R _20233_ (.A1(_14103_),
    .A2(_00661_),
    .B(_14472_),
    .Y(_14473_));
 AND2x2_ASAP7_75t_R _20234_ (.A(_14198_),
    .B(_00660_),
    .Y(_14474_));
 AO21x1_ASAP7_75t_R _20235_ (.A1(_13390_),
    .A2(_00662_),
    .B(_14474_),
    .Y(_14475_));
 OR2x2_ASAP7_75t_R _20236_ (.A(_13477_),
    .B(_13510_),
    .Y(_14476_));
 OA22x2_ASAP7_75t_R _20237_ (.A1(_14471_),
    .A2(_14473_),
    .B1(_14475_),
    .B2(_14476_),
    .Y(_14477_));
 NAND2x1_ASAP7_75t_R _20238_ (.A(_13491_),
    .B(_14041_),
    .Y(_14478_));
 AND2x2_ASAP7_75t_R _20239_ (.A(_13456_),
    .B(_00655_),
    .Y(_14479_));
 AO21x1_ASAP7_75t_R _20240_ (.A1(_14103_),
    .A2(_00657_),
    .B(_14479_),
    .Y(_14480_));
 AND2x2_ASAP7_75t_R _20241_ (.A(_13456_),
    .B(_00656_),
    .Y(_14481_));
 AO21x1_ASAP7_75t_R _20242_ (.A1(_14103_),
    .A2(_00658_),
    .B(_14481_),
    .Y(_14482_));
 NAND2x1_ASAP7_75t_R _20243_ (.A(_13469_),
    .B(_14041_),
    .Y(_14483_));
 OA22x2_ASAP7_75t_R _20244_ (.A1(_14478_),
    .A2(_14480_),
    .B1(_14482_),
    .B2(_14483_),
    .Y(_14484_));
 NAND3x2_ASAP7_75t_R _20245_ (.B(_14477_),
    .C(_14484_),
    .Y(_14485_),
    .A(_14470_));
 AND3x4_ASAP7_75t_R _20246_ (.A(_14454_),
    .B(_14469_),
    .C(_14485_),
    .Y(_14486_));
 INVx1_ASAP7_75t_R _20247_ (.A(_13579_),
    .Y(_14487_));
 AO32x1_ASAP7_75t_R _20248_ (.A1(_13365_),
    .A2(_13387_),
    .A3(_14486_),
    .B1(_14429_),
    .B2(_14487_),
    .Y(_14488_));
 BUFx3_ASAP7_75t_R _20249_ (.A(_14488_),
    .Y(_18643_));
 INVx1_ASAP7_75t_R _20250_ (.A(_18643_),
    .Y(_18645_));
 AND2x2_ASAP7_75t_R _20251_ (.A(_14262_),
    .B(_01784_),
    .Y(_14489_));
 AO21x1_ASAP7_75t_R _20252_ (.A1(_13390_),
    .A2(_00664_),
    .B(_14489_),
    .Y(_14490_));
 OAI22x1_ASAP7_75t_R _20253_ (.A1(_00663_),
    .A2(_13497_),
    .B1(_14490_),
    .B2(_13492_),
    .Y(_14491_));
 INVx1_ASAP7_75t_R _20254_ (.A(_00680_),
    .Y(_14492_));
 NAND2x1_ASAP7_75t_R _20255_ (.A(_14112_),
    .B(_00678_),
    .Y(_14493_));
 OA211x2_ASAP7_75t_R _20256_ (.A1(_14110_),
    .A2(_14492_),
    .B(_14493_),
    .C(_14117_),
    .Y(_14494_));
 BUFx6f_ASAP7_75t_R _20257_ (.A(_14097_),
    .Y(_14495_));
 INVx1_ASAP7_75t_R _20258_ (.A(_00679_),
    .Y(_14496_));
 NAND2x1_ASAP7_75t_R _20259_ (.A(_14112_),
    .B(_00677_),
    .Y(_14497_));
 OA211x2_ASAP7_75t_R _20260_ (.A1(_14495_),
    .A2(_14496_),
    .B(_14497_),
    .C(_13477_),
    .Y(_14498_));
 OR3x1_ASAP7_75t_R _20261_ (.A(_13517_),
    .B(_14494_),
    .C(_14498_),
    .Y(_14499_));
 OA211x2_ASAP7_75t_R _20262_ (.A1(_13447_),
    .A2(_14491_),
    .B(_14499_),
    .C(_14038_),
    .Y(_14500_));
 INVx1_ASAP7_75t_R _20263_ (.A(_00689_),
    .Y(_14501_));
 NAND2x1_ASAP7_75t_R _20264_ (.A(_14041_),
    .B(_00685_),
    .Y(_14502_));
 OA21x2_ASAP7_75t_R _20265_ (.A1(_13511_),
    .A2(_14501_),
    .B(_14502_),
    .Y(_14503_));
 INVx1_ASAP7_75t_R _20266_ (.A(_00691_),
    .Y(_14504_));
 NAND2x1_ASAP7_75t_R _20267_ (.A(_14044_),
    .B(_00687_),
    .Y(_14505_));
 OA211x2_ASAP7_75t_R _20268_ (.A1(_14041_),
    .A2(_14504_),
    .B(_14174_),
    .C(_14505_),
    .Y(_14506_));
 AO21x1_ASAP7_75t_R _20269_ (.A1(_14173_),
    .A2(_14503_),
    .B(_14506_),
    .Y(_14507_));
 INVx2_ASAP7_75t_R _20270_ (.A(_00675_),
    .Y(_14508_));
 NAND2x1_ASAP7_75t_R _20271_ (.A(_14041_),
    .B(_00671_),
    .Y(_14509_));
 OA21x2_ASAP7_75t_R _20272_ (.A1(_13511_),
    .A2(_14508_),
    .B(_14509_),
    .Y(_14510_));
 INVx1_ASAP7_75t_R _20273_ (.A(_00673_),
    .Y(_14511_));
 NAND2x1_ASAP7_75t_R _20274_ (.A(_14044_),
    .B(_00669_),
    .Y(_14512_));
 OA211x2_ASAP7_75t_R _20275_ (.A1(_14041_),
    .A2(_14511_),
    .B(_14181_),
    .C(_14512_),
    .Y(_14513_));
 AO21x1_ASAP7_75t_R _20276_ (.A1(_14182_),
    .A2(_14510_),
    .B(_14513_),
    .Y(_14514_));
 OA21x2_ASAP7_75t_R _20277_ (.A1(_14507_),
    .A2(_14514_),
    .B(_14187_),
    .Y(_14515_));
 INVx2_ASAP7_75t_R _20278_ (.A(_00692_),
    .Y(_14516_));
 NAND2x1_ASAP7_75t_R _20279_ (.A(_13516_),
    .B(_00676_),
    .Y(_14517_));
 OA211x2_ASAP7_75t_R _20280_ (.A1(_14092_),
    .A2(_14516_),
    .B(_14517_),
    .C(_13450_),
    .Y(_14518_));
 INVx2_ASAP7_75t_R _20281_ (.A(_00688_),
    .Y(_14519_));
 NAND2x1_ASAP7_75t_R _20282_ (.A(_13516_),
    .B(_00672_),
    .Y(_14520_));
 OA211x2_ASAP7_75t_R _20283_ (.A1(_14092_),
    .A2(_14519_),
    .B(_14520_),
    .C(_14044_),
    .Y(_14521_));
 OA21x2_ASAP7_75t_R _20284_ (.A1(_14518_),
    .A2(_14521_),
    .B(_14195_),
    .Y(_14522_));
 INVx1_ASAP7_75t_R _20285_ (.A(_00684_),
    .Y(_14523_));
 NAND2x1_ASAP7_75t_R _20286_ (.A(_14112_),
    .B(_00682_),
    .Y(_14524_));
 OA211x2_ASAP7_75t_R _20287_ (.A1(_14110_),
    .A2(_14523_),
    .B(_14524_),
    .C(_14117_),
    .Y(_14525_));
 INVx1_ASAP7_75t_R _20288_ (.A(_00683_),
    .Y(_14526_));
 NAND2x1_ASAP7_75t_R _20289_ (.A(_14112_),
    .B(_00681_),
    .Y(_14527_));
 OA211x2_ASAP7_75t_R _20290_ (.A1(_14495_),
    .A2(_14526_),
    .B(_14527_),
    .C(_13477_),
    .Y(_14528_));
 OA21x2_ASAP7_75t_R _20291_ (.A1(_14525_),
    .A2(_14528_),
    .B(_14205_),
    .Y(_14529_));
 INVx1_ASAP7_75t_R _20292_ (.A(_00690_),
    .Y(_14530_));
 NAND2x1_ASAP7_75t_R _20293_ (.A(_14063_),
    .B(_00674_),
    .Y(_14531_));
 OA211x2_ASAP7_75t_R _20294_ (.A1(_13516_),
    .A2(_14530_),
    .B(_14531_),
    .C(_13450_),
    .Y(_14532_));
 INVx1_ASAP7_75t_R _20295_ (.A(_00686_),
    .Y(_14533_));
 NAND2x1_ASAP7_75t_R _20296_ (.A(_14063_),
    .B(_00670_),
    .Y(_14534_));
 OA211x2_ASAP7_75t_R _20297_ (.A1(_13516_),
    .A2(_14533_),
    .B(_14534_),
    .C(_14044_),
    .Y(_14535_));
 OA21x2_ASAP7_75t_R _20298_ (.A1(_14532_),
    .A2(_14535_),
    .B(_14213_),
    .Y(_14536_));
 INVx1_ASAP7_75t_R _20299_ (.A(_00668_),
    .Y(_14537_));
 NAND2x1_ASAP7_75t_R _20300_ (.A(_14160_),
    .B(_00666_),
    .Y(_14538_));
 OA211x2_ASAP7_75t_R _20301_ (.A1(_14495_),
    .A2(_14537_),
    .B(_14538_),
    .C(_14117_),
    .Y(_14539_));
 INVx1_ASAP7_75t_R _20302_ (.A(_00667_),
    .Y(_14540_));
 NAND2x1_ASAP7_75t_R _20303_ (.A(_14160_),
    .B(_00665_),
    .Y(_14541_));
 OA211x2_ASAP7_75t_R _20304_ (.A1(_14262_),
    .A2(_14540_),
    .B(_14541_),
    .C(_13477_),
    .Y(_14542_));
 OA21x2_ASAP7_75t_R _20305_ (.A1(_14539_),
    .A2(_14542_),
    .B(_14221_),
    .Y(_14543_));
 OR4x2_ASAP7_75t_R _20306_ (.A(_14522_),
    .B(_14529_),
    .C(_14536_),
    .D(_14543_),
    .Y(_14544_));
 OA31x2_ASAP7_75t_R _20307_ (.A1(_14500_),
    .A2(_14515_),
    .A3(_14544_),
    .B1(_13787_),
    .Y(_14545_));
 INVx2_ASAP7_75t_R _20308_ (.A(_13578_),
    .Y(_14546_));
 OA211x2_ASAP7_75t_R _20309_ (.A1(_14427_),
    .A2(_14428_),
    .B(_14546_),
    .C(_14373_),
    .Y(_14547_));
 OR2x2_ASAP7_75t_R _20310_ (.A(_14545_),
    .B(_14547_),
    .Y(_14548_));
 BUFx3_ASAP7_75t_R _20311_ (.A(_14548_),
    .Y(_18648_));
 INVx1_ASAP7_75t_R _20312_ (.A(_18648_),
    .Y(_18650_));
 AND2x2_ASAP7_75t_R _20313_ (.A(_14197_),
    .B(_01783_),
    .Y(_14549_));
 AO21x1_ASAP7_75t_R _20314_ (.A1(_13389_),
    .A2(_00694_),
    .B(_14549_),
    .Y(_14550_));
 OAI22x1_ASAP7_75t_R _20315_ (.A1(_00693_),
    .A2(_13496_),
    .B1(_14550_),
    .B2(_13491_),
    .Y(_14551_));
 INVx1_ASAP7_75t_R _20316_ (.A(_00710_),
    .Y(_14552_));
 NAND2x1_ASAP7_75t_R _20317_ (.A(_13798_),
    .B(_00708_),
    .Y(_14553_));
 OA211x2_ASAP7_75t_R _20318_ (.A1(_13799_),
    .A2(_14552_),
    .B(_14553_),
    .C(net3),
    .Y(_14554_));
 INVx1_ASAP7_75t_R _20319_ (.A(_00709_),
    .Y(_14555_));
 NAND2x1_ASAP7_75t_R _20320_ (.A(_13798_),
    .B(_00707_),
    .Y(_14556_));
 OA211x2_ASAP7_75t_R _20321_ (.A1(_13799_),
    .A2(_14555_),
    .B(_14556_),
    .C(net4),
    .Y(_14557_));
 OR3x1_ASAP7_75t_R _20322_ (.A(_13516_),
    .B(_14554_),
    .C(_14557_),
    .Y(_14558_));
 OA211x2_ASAP7_75t_R _20323_ (.A1(_13446_),
    .A2(_14551_),
    .B(_14558_),
    .C(_14038_),
    .Y(_14559_));
 NAND2x1_ASAP7_75t_R _20324_ (.A(_14040_),
    .B(_00716_),
    .Y(_14560_));
 NAND2x1_ASAP7_75t_R _20325_ (.A(_14140_),
    .B(_00720_),
    .Y(_14561_));
 INVx1_ASAP7_75t_R _20326_ (.A(_00722_),
    .Y(_14562_));
 NAND2x1_ASAP7_75t_R _20327_ (.A(_13509_),
    .B(_00718_),
    .Y(_14563_));
 OA21x2_ASAP7_75t_R _20328_ (.A1(_14043_),
    .A2(_14562_),
    .B(_14563_),
    .Y(_14564_));
 AO32x1_ASAP7_75t_R _20329_ (.A1(_14173_),
    .A2(_14560_),
    .A3(_14561_),
    .B1(_14564_),
    .B2(_14174_),
    .Y(_14565_));
 NAND2x1_ASAP7_75t_R _20330_ (.A(_14040_),
    .B(_00700_),
    .Y(_14566_));
 NAND2x1_ASAP7_75t_R _20331_ (.A(_14140_),
    .B(_00704_),
    .Y(_14567_));
 INVx1_ASAP7_75t_R _20332_ (.A(_00706_),
    .Y(_14568_));
 NAND2x1_ASAP7_75t_R _20333_ (.A(_13509_),
    .B(_00702_),
    .Y(_14569_));
 OA21x2_ASAP7_75t_R _20334_ (.A1(_14043_),
    .A2(_14568_),
    .B(_14569_),
    .Y(_14570_));
 AO32x1_ASAP7_75t_R _20335_ (.A1(_14181_),
    .A2(_14566_),
    .A3(_14567_),
    .B1(_14570_),
    .B2(_14182_),
    .Y(_14571_));
 OA211x2_ASAP7_75t_R _20336_ (.A1(_14565_),
    .A2(_14571_),
    .B(net11),
    .C(_13452_),
    .Y(_14572_));
 INVx2_ASAP7_75t_R _20337_ (.A(_00721_),
    .Y(_14573_));
 NAND2x1_ASAP7_75t_R _20338_ (.A(_13448_),
    .B(_00717_),
    .Y(_14574_));
 OA211x2_ASAP7_75t_R _20339_ (.A1(_13509_),
    .A2(_14573_),
    .B(_14574_),
    .C(_13388_),
    .Y(_14575_));
 INVx1_ASAP7_75t_R _20340_ (.A(_00719_),
    .Y(_14576_));
 NAND2x1_ASAP7_75t_R _20341_ (.A(_13448_),
    .B(_00715_),
    .Y(_14577_));
 OA211x2_ASAP7_75t_R _20342_ (.A1(_13509_),
    .A2(_14576_),
    .B(_14577_),
    .C(net2),
    .Y(_14578_));
 OA211x2_ASAP7_75t_R _20343_ (.A1(_14575_),
    .A2(_14578_),
    .B(_13445_),
    .C(_14187_),
    .Y(_14579_));
 INVx1_ASAP7_75t_R _20344_ (.A(_00705_),
    .Y(_14580_));
 NAND2x1_ASAP7_75t_R _20345_ (.A(_13448_),
    .B(_00701_),
    .Y(_14581_));
 OA211x2_ASAP7_75t_R _20346_ (.A1(_13509_),
    .A2(_14580_),
    .B(_14581_),
    .C(_13388_),
    .Y(_14582_));
 INVx1_ASAP7_75t_R _20347_ (.A(_00703_),
    .Y(_14583_));
 NAND2x1_ASAP7_75t_R _20348_ (.A(_13448_),
    .B(_00699_),
    .Y(_14584_));
 OA211x2_ASAP7_75t_R _20349_ (.A1(_13509_),
    .A2(_14583_),
    .B(_14584_),
    .C(net2),
    .Y(_14585_));
 OA211x2_ASAP7_75t_R _20350_ (.A1(_14582_),
    .A2(_14585_),
    .B(_14060_),
    .C(_14187_),
    .Y(_14586_));
 INVx1_ASAP7_75t_R _20351_ (.A(_00698_),
    .Y(_14587_));
 NAND2x1_ASAP7_75t_R _20352_ (.A(_13798_),
    .B(_00696_),
    .Y(_14588_));
 OA211x2_ASAP7_75t_R _20353_ (.A1(_14197_),
    .A2(_14587_),
    .B(_14588_),
    .C(net3),
    .Y(_14589_));
 INVx1_ASAP7_75t_R _20354_ (.A(_00697_),
    .Y(_14590_));
 NAND2x1_ASAP7_75t_R _20355_ (.A(_13798_),
    .B(_00695_),
    .Y(_14591_));
 OA211x2_ASAP7_75t_R _20356_ (.A1(_14197_),
    .A2(_14590_),
    .B(_14591_),
    .C(net4),
    .Y(_14592_));
 OA21x2_ASAP7_75t_R _20357_ (.A1(_14589_),
    .A2(_14592_),
    .B(_14221_),
    .Y(_14593_));
 INVx1_ASAP7_75t_R _20358_ (.A(_00714_),
    .Y(_14594_));
 NAND2x1_ASAP7_75t_R _20359_ (.A(_13798_),
    .B(_00712_),
    .Y(_14595_));
 OA211x2_ASAP7_75t_R _20360_ (.A1(_14197_),
    .A2(_14594_),
    .B(_14595_),
    .C(_13466_),
    .Y(_14596_));
 INVx1_ASAP7_75t_R _20361_ (.A(_00713_),
    .Y(_14597_));
 NAND2x1_ASAP7_75t_R _20362_ (.A(_13798_),
    .B(_00711_),
    .Y(_14598_));
 OA211x2_ASAP7_75t_R _20363_ (.A1(_14197_),
    .A2(_14597_),
    .B(_14598_),
    .C(net4),
    .Y(_14599_));
 OA21x2_ASAP7_75t_R _20364_ (.A1(_14596_),
    .A2(_14599_),
    .B(_14205_),
    .Y(_14600_));
 OR4x1_ASAP7_75t_R _20365_ (.A(_14579_),
    .B(_14586_),
    .C(_14593_),
    .D(_14600_),
    .Y(_14601_));
 OR3x2_ASAP7_75t_R _20366_ (.A(_14559_),
    .B(_14572_),
    .C(_14601_),
    .Y(_14602_));
 BUFx6f_ASAP7_75t_R _20367_ (.A(_14602_),
    .Y(_14603_));
 INVx1_ASAP7_75t_R _20368_ (.A(_13577_),
    .Y(_14604_));
 AO32x1_ASAP7_75t_R _20369_ (.A1(_13365_),
    .A2(_13387_),
    .A3(_14603_),
    .B1(_14429_),
    .B2(_14604_),
    .Y(_14605_));
 BUFx6f_ASAP7_75t_R _20370_ (.A(_14605_),
    .Y(_18652_));
 INVx3_ASAP7_75t_R _20371_ (.A(_18652_),
    .Y(_18654_));
 INVx1_ASAP7_75t_R _20372_ (.A(_00728_),
    .Y(_14606_));
 NAND2x1_ASAP7_75t_R _20373_ (.A(_14160_),
    .B(_00726_),
    .Y(_14607_));
 OA211x2_ASAP7_75t_R _20374_ (.A1(_14262_),
    .A2(_14606_),
    .B(_14607_),
    .C(_14117_),
    .Y(_14608_));
 INVx2_ASAP7_75t_R _20375_ (.A(_00727_),
    .Y(_14609_));
 NAND2x1_ASAP7_75t_R _20376_ (.A(_14160_),
    .B(_00725_),
    .Y(_14610_));
 OA211x2_ASAP7_75t_R _20377_ (.A1(_14262_),
    .A2(_14609_),
    .B(_14610_),
    .C(_13477_),
    .Y(_14611_));
 OA21x2_ASAP7_75t_R _20378_ (.A1(_14608_),
    .A2(_14611_),
    .B(_14292_),
    .Y(_14612_));
 INVx1_ASAP7_75t_R _20379_ (.A(_00732_),
    .Y(_14613_));
 NAND2x1_ASAP7_75t_R _20380_ (.A(_14160_),
    .B(_00730_),
    .Y(_14614_));
 OA211x2_ASAP7_75t_R _20381_ (.A1(_14262_),
    .A2(_14613_),
    .B(_14614_),
    .C(_14117_),
    .Y(_14615_));
 INVx2_ASAP7_75t_R _20382_ (.A(_00731_),
    .Y(_14616_));
 NAND2x1_ASAP7_75t_R _20383_ (.A(_14164_),
    .B(_00729_),
    .Y(_14617_));
 OA211x2_ASAP7_75t_R _20384_ (.A1(_14262_),
    .A2(_14616_),
    .B(_14617_),
    .C(_13477_),
    .Y(_14618_));
 OA21x2_ASAP7_75t_R _20385_ (.A1(_14615_),
    .A2(_14618_),
    .B(_14261_),
    .Y(_14619_));
 OA21x2_ASAP7_75t_R _20386_ (.A1(_14612_),
    .A2(_14619_),
    .B(_13517_),
    .Y(_14620_));
 INVx1_ASAP7_75t_R _20387_ (.A(_00744_),
    .Y(_14621_));
 NAND2x1_ASAP7_75t_R _20388_ (.A(_14198_),
    .B(_00742_),
    .Y(_14622_));
 OA211x2_ASAP7_75t_R _20389_ (.A1(_14262_),
    .A2(_14621_),
    .B(_14622_),
    .C(_13794_),
    .Y(_14623_));
 INVx2_ASAP7_75t_R _20390_ (.A(_00743_),
    .Y(_14624_));
 NAND2x1_ASAP7_75t_R _20391_ (.A(_14198_),
    .B(_00741_),
    .Y(_14625_));
 OA211x2_ASAP7_75t_R _20392_ (.A1(_13462_),
    .A2(_14624_),
    .B(_14625_),
    .C(_13477_),
    .Y(_14626_));
 OA21x2_ASAP7_75t_R _20393_ (.A1(_14623_),
    .A2(_14626_),
    .B(_14292_),
    .Y(_14627_));
 INVx1_ASAP7_75t_R _20394_ (.A(_00748_),
    .Y(_14628_));
 NAND2x1_ASAP7_75t_R _20395_ (.A(_14198_),
    .B(_00746_),
    .Y(_14629_));
 OA211x2_ASAP7_75t_R _20396_ (.A1(_13462_),
    .A2(_14628_),
    .B(_14629_),
    .C(_13794_),
    .Y(_14630_));
 INVx1_ASAP7_75t_R _20397_ (.A(_00747_),
    .Y(_14631_));
 NAND2x1_ASAP7_75t_R _20398_ (.A(_14198_),
    .B(_00745_),
    .Y(_14632_));
 OA211x2_ASAP7_75t_R _20399_ (.A1(_13462_),
    .A2(_14631_),
    .B(_14632_),
    .C(_13477_),
    .Y(_14633_));
 OA21x2_ASAP7_75t_R _20400_ (.A1(_14630_),
    .A2(_14633_),
    .B(_14261_),
    .Y(_14634_));
 OA21x2_ASAP7_75t_R _20401_ (.A1(_14627_),
    .A2(_14634_),
    .B(_13447_),
    .Y(_14635_));
 AND2x2_ASAP7_75t_R _20402_ (.A(net4),
    .B(_13445_),
    .Y(_14636_));
 INVx2_ASAP7_75t_R _20403_ (.A(_00751_),
    .Y(_14637_));
 NAND2x1_ASAP7_75t_R _20404_ (.A(_13462_),
    .B(_00749_),
    .Y(_14638_));
 OA21x2_ASAP7_75t_R _20405_ (.A1(_14110_),
    .A2(_14637_),
    .B(_14638_),
    .Y(_14639_));
 INVx2_ASAP7_75t_R _20406_ (.A(_00752_),
    .Y(_14640_));
 NOR2x1_ASAP7_75t_R _20407_ (.A(_13490_),
    .B(_14063_),
    .Y(_14641_));
 NAND2x1_ASAP7_75t_R _20408_ (.A(_14160_),
    .B(_00750_),
    .Y(_14642_));
 OA211x2_ASAP7_75t_R _20409_ (.A1(_14495_),
    .A2(_14640_),
    .B(_14641_),
    .C(_14642_),
    .Y(_14643_));
 AO21x1_ASAP7_75t_R _20410_ (.A1(_14636_),
    .A2(_14639_),
    .B(_14643_),
    .Y(_14644_));
 INVx1_ASAP7_75t_R _20411_ (.A(_00736_),
    .Y(_14645_));
 NAND2x1_ASAP7_75t_R _20412_ (.A(_13462_),
    .B(_00734_),
    .Y(_14646_));
 OA21x2_ASAP7_75t_R _20413_ (.A1(_14110_),
    .A2(_14645_),
    .B(_14646_),
    .Y(_14647_));
 AND2x2_ASAP7_75t_R _20414_ (.A(net3),
    .B(_13515_),
    .Y(_14648_));
 INVx2_ASAP7_75t_R _20415_ (.A(_00735_),
    .Y(_14649_));
 NAND2x1_ASAP7_75t_R _20416_ (.A(_14160_),
    .B(_00733_),
    .Y(_14650_));
 AND2x2_ASAP7_75t_R _20417_ (.A(_00368_),
    .B(_00366_),
    .Y(_14651_));
 OA211x2_ASAP7_75t_R _20418_ (.A1(_14495_),
    .A2(_14649_),
    .B(_14650_),
    .C(_14651_),
    .Y(_14652_));
 AO21x1_ASAP7_75t_R _20419_ (.A1(_14647_),
    .A2(_14648_),
    .B(_14652_),
    .Y(_14653_));
 OA21x2_ASAP7_75t_R _20420_ (.A1(_14644_),
    .A2(_14653_),
    .B(_14248_),
    .Y(_14654_));
 AND2x2_ASAP7_75t_R _20421_ (.A(_14160_),
    .B(_01813_),
    .Y(_14655_));
 AO21x1_ASAP7_75t_R _20422_ (.A1(_13390_),
    .A2(_00724_),
    .B(_14655_),
    .Y(_14656_));
 OAI22x1_ASAP7_75t_R _20423_ (.A1(_00723_),
    .A2(_13497_),
    .B1(_14656_),
    .B2(_13478_),
    .Y(_14657_));
 INVx1_ASAP7_75t_R _20424_ (.A(_00740_),
    .Y(_14658_));
 NAND2x1_ASAP7_75t_R _20425_ (.A(_14097_),
    .B(_00738_),
    .Y(_14659_));
 OA211x2_ASAP7_75t_R _20426_ (.A1(_13800_),
    .A2(_14658_),
    .B(_14659_),
    .C(net16),
    .Y(_14660_));
 INVx2_ASAP7_75t_R _20427_ (.A(_00739_),
    .Y(_14661_));
 NAND2x1_ASAP7_75t_R _20428_ (.A(_14097_),
    .B(_00737_),
    .Y(_14662_));
 OA211x2_ASAP7_75t_R _20429_ (.A1(_13800_),
    .A2(_14661_),
    .B(_14662_),
    .C(_14167_),
    .Y(_14663_));
 OR3x1_ASAP7_75t_R _20430_ (.A(_14092_),
    .B(_14660_),
    .C(_14663_),
    .Y(_14664_));
 OA211x2_ASAP7_75t_R _20431_ (.A1(_13446_),
    .A2(_14657_),
    .B(_14664_),
    .C(_14038_),
    .Y(_14665_));
 OR4x2_ASAP7_75t_R _20432_ (.A(_14620_),
    .B(_14635_),
    .C(_14654_),
    .D(_14665_),
    .Y(_14666_));
 AO32x2_ASAP7_75t_R _20433_ (.A1(_13366_),
    .A2(_13387_),
    .A3(_14666_),
    .B1(_14429_),
    .B2(_13597_),
    .Y(_14667_));
 BUFx4f_ASAP7_75t_R _20434_ (.A(_14667_),
    .Y(_14668_));
 INVx4_ASAP7_75t_R _20435_ (.A(_14668_),
    .Y(_18660_));
 INVx1_ASAP7_75t_R _20436_ (.A(_00757_),
    .Y(_14669_));
 NAND2x1_ASAP7_75t_R _20437_ (.A(_14075_),
    .B(_00755_),
    .Y(_14670_));
 OA211x2_ASAP7_75t_R _20438_ (.A1(_14073_),
    .A2(_14669_),
    .B(_14670_),
    .C(_14035_),
    .Y(_14671_));
 INVx1_ASAP7_75t_R _20439_ (.A(_00758_),
    .Y(_14672_));
 NAND2x1_ASAP7_75t_R _20440_ (.A(_14104_),
    .B(_00756_),
    .Y(_14673_));
 OA211x2_ASAP7_75t_R _20441_ (.A1(_14073_),
    .A2(_14672_),
    .B(_14673_),
    .C(_13794_),
    .Y(_14674_));
 INVx2_ASAP7_75t_R _20442_ (.A(_00773_),
    .Y(_14675_));
 NAND2x1_ASAP7_75t_R _20443_ (.A(_14267_),
    .B(_00771_),
    .Y(_14676_));
 OA211x2_ASAP7_75t_R _20444_ (.A1(_14055_),
    .A2(_14675_),
    .B(_14676_),
    .C(_14035_),
    .Y(_14677_));
 INVx1_ASAP7_75t_R _20445_ (.A(_00774_),
    .Y(_14678_));
 NAND2x1_ASAP7_75t_R _20446_ (.A(_14267_),
    .B(_00772_),
    .Y(_14679_));
 OA211x2_ASAP7_75t_R _20447_ (.A1(_14055_),
    .A2(_14678_),
    .B(_14679_),
    .C(_13794_),
    .Y(_14680_));
 OA33x2_ASAP7_75t_R _20448_ (.A1(_14109_),
    .A2(_14671_),
    .A3(_14674_),
    .B1(_14677_),
    .B2(_14680_),
    .B3(_14119_),
    .Y(_14681_));
 INVx1_ASAP7_75t_R _20449_ (.A(_00762_),
    .Y(_14682_));
 NAND2x1_ASAP7_75t_R _20450_ (.A(_14072_),
    .B(_00760_),
    .Y(_14683_));
 OA211x2_ASAP7_75t_R _20451_ (.A1(_14104_),
    .A2(_14682_),
    .B(_14683_),
    .C(_14137_),
    .Y(_14684_));
 INVx2_ASAP7_75t_R _20452_ (.A(_00761_),
    .Y(_14685_));
 NAND2x1_ASAP7_75t_R _20453_ (.A(_14355_),
    .B(_00759_),
    .Y(_14686_));
 OA211x2_ASAP7_75t_R _20454_ (.A1(_14104_),
    .A2(_14685_),
    .B(_14686_),
    .C(_13490_),
    .Y(_14687_));
 OR3x1_ASAP7_75t_R _20455_ (.A(_13446_),
    .B(_14684_),
    .C(_14687_),
    .Y(_14688_));
 INVx1_ASAP7_75t_R _20456_ (.A(_00778_),
    .Y(_14689_));
 NAND2x1_ASAP7_75t_R _20457_ (.A(_14355_),
    .B(_00776_),
    .Y(_14690_));
 OA211x2_ASAP7_75t_R _20458_ (.A1(_14104_),
    .A2(_14689_),
    .B(_14690_),
    .C(net3),
    .Y(_14691_));
 INVx2_ASAP7_75t_R _20459_ (.A(_00777_),
    .Y(_14692_));
 NAND2x1_ASAP7_75t_R _20460_ (.A(_14355_),
    .B(_00775_),
    .Y(_14693_));
 OA211x2_ASAP7_75t_R _20461_ (.A1(_14075_),
    .A2(_14692_),
    .B(_14693_),
    .C(_13490_),
    .Y(_14694_));
 OR3x1_ASAP7_75t_R _20462_ (.A(_14092_),
    .B(_14691_),
    .C(_14694_),
    .Y(_14695_));
 AO21x1_ASAP7_75t_R _20463_ (.A1(_14688_),
    .A2(_14695_),
    .B(_14362_),
    .Y(_14696_));
 INVx1_ASAP7_75t_R _20464_ (.A(_00782_),
    .Y(_14697_));
 NAND2x1_ASAP7_75t_R _20465_ (.A(_14355_),
    .B(_00780_),
    .Y(_14698_));
 OA21x2_ASAP7_75t_R _20466_ (.A1(_14097_),
    .A2(_14697_),
    .B(_14698_),
    .Y(_14699_));
 INVx2_ASAP7_75t_R _20467_ (.A(_00765_),
    .Y(_14700_));
 NAND2x1_ASAP7_75t_R _20468_ (.A(net2),
    .B(_00763_),
    .Y(_14701_));
 OA211x2_ASAP7_75t_R _20469_ (.A1(_14054_),
    .A2(_14700_),
    .B(_14651_),
    .C(_14701_),
    .Y(_14702_));
 AO21x1_ASAP7_75t_R _20470_ (.A1(_14641_),
    .A2(_14699_),
    .B(_14702_),
    .Y(_14703_));
 INVx2_ASAP7_75t_R _20471_ (.A(_00781_),
    .Y(_14704_));
 NAND2x1_ASAP7_75t_R _20472_ (.A(_13461_),
    .B(_00779_),
    .Y(_14705_));
 OA211x2_ASAP7_75t_R _20473_ (.A1(_14164_),
    .A2(_14704_),
    .B(_14636_),
    .C(_14705_),
    .Y(_14706_));
 INVx1_ASAP7_75t_R _20474_ (.A(_00766_),
    .Y(_14707_));
 NAND2x1_ASAP7_75t_R _20475_ (.A(_14054_),
    .B(_00764_),
    .Y(_14708_));
 OA211x2_ASAP7_75t_R _20476_ (.A1(_14164_),
    .A2(_14707_),
    .B(_14648_),
    .C(_14708_),
    .Y(_14709_));
 OR5x1_ASAP7_75t_R _20477_ (.A(_13511_),
    .B(_13482_),
    .C(_14703_),
    .D(_14706_),
    .E(_14709_),
    .Y(_14710_));
 INVx1_ASAP7_75t_R _20478_ (.A(_00770_),
    .Y(_14711_));
 NAND2x1_ASAP7_75t_R _20479_ (.A(_14355_),
    .B(_00768_),
    .Y(_14712_));
 OA211x2_ASAP7_75t_R _20480_ (.A1(_14075_),
    .A2(_14711_),
    .B(_14712_),
    .C(net3),
    .Y(_14713_));
 INVx1_ASAP7_75t_R _20481_ (.A(_00769_),
    .Y(_14714_));
 NAND2x1_ASAP7_75t_R _20482_ (.A(_13799_),
    .B(_00767_),
    .Y(_14715_));
 OA211x2_ASAP7_75t_R _20483_ (.A1(_14079_),
    .A2(_14714_),
    .B(_14715_),
    .C(_13490_),
    .Y(_14716_));
 OR3x1_ASAP7_75t_R _20484_ (.A(_14092_),
    .B(_14713_),
    .C(_14716_),
    .Y(_14717_));
 INVx1_ASAP7_75t_R _20485_ (.A(_00753_),
    .Y(_14718_));
 AND2x2_ASAP7_75t_R _20486_ (.A(_14072_),
    .B(_01812_),
    .Y(_14719_));
 AOI21x1_ASAP7_75t_R _20487_ (.A1(_13389_),
    .A2(_00754_),
    .B(_14719_),
    .Y(_14720_));
 AO221x1_ASAP7_75t_R _20488_ (.A1(_14718_),
    .A2(_14102_),
    .B1(_14720_),
    .B2(_14117_),
    .C(_13445_),
    .Y(_14721_));
 AO21x1_ASAP7_75t_R _20489_ (.A1(_14717_),
    .A2(_14721_),
    .B(_14056_),
    .Y(_14722_));
 AND4x2_ASAP7_75t_R _20490_ (.A(_14681_),
    .B(_14696_),
    .C(_14710_),
    .D(_14722_),
    .Y(_14723_));
 AND2x2_ASAP7_75t_R _20491_ (.A(net14),
    .B(_14150_),
    .Y(_14724_));
 AND4x1_ASAP7_75t_R _20492_ (.A(_14058_),
    .B(_13365_),
    .C(_13386_),
    .D(_13433_),
    .Y(_14725_));
 INVx4_ASAP7_75t_R _20493_ (.A(_00446_),
    .Y(_14726_));
 AND4x1_ASAP7_75t_R _20494_ (.A(_14726_),
    .B(_13365_),
    .C(_13373_),
    .D(_13434_),
    .Y(_14727_));
 OA21x2_ASAP7_75t_R _20495_ (.A1(_14725_),
    .A2(_14727_),
    .B(_13429_),
    .Y(_14728_));
 AOI221x1_ASAP7_75t_R _20496_ (.A1(_13788_),
    .A2(_14723_),
    .B1(_14724_),
    .B2(_14226_),
    .C(_14728_),
    .Y(_18665_));
 INVx2_ASAP7_75t_R _20497_ (.A(_18665_),
    .Y(_14729_));
 BUFx6f_ASAP7_75t_R _20498_ (.A(_14729_),
    .Y(_18663_));
 OR3x2_ASAP7_75t_R _20499_ (.A(_13403_),
    .B(_13623_),
    .C(_13650_),
    .Y(_14730_));
 AO21x1_ASAP7_75t_R _20500_ (.A1(_13563_),
    .A2(_14048_),
    .B(_13561_),
    .Y(_14731_));
 OR2x4_ASAP7_75t_R _20501_ (.A(_14730_),
    .B(_14731_),
    .Y(_18862_));
 INVx1_ASAP7_75t_R _20502_ (.A(_18862_),
    .Y(_18863_));
 BUFx12_ASAP7_75t_R _20503_ (.A(_13674_),
    .Y(_14732_));
 BUFx6f_ASAP7_75t_R _20504_ (.A(_13670_),
    .Y(_14733_));
 OR5x1_ASAP7_75t_R _20505_ (.A(_13945_),
    .B(_13777_),
    .C(_14732_),
    .D(_13857_),
    .E(_14733_),
    .Y(_14734_));
 AND3x2_ASAP7_75t_R _20506_ (.A(_13563_),
    .B(_13774_),
    .C(_14734_),
    .Y(_14735_));
 BUFx3_ASAP7_75t_R _20507_ (.A(_14735_),
    .Y(_14736_));
 INVx1_ASAP7_75t_R _20508_ (.A(_14736_),
    .Y(_18865_));
 BUFx10_ASAP7_75t_R _20509_ (.A(_13659_),
    .Y(_14737_));
 BUFx10_ASAP7_75t_R _20510_ (.A(_13670_),
    .Y(_14738_));
 BUFx10_ASAP7_75t_R _20511_ (.A(_13675_),
    .Y(_14739_));
 BUFx6f_ASAP7_75t_R _20512_ (.A(_14739_),
    .Y(_14740_));
 BUFx12_ASAP7_75t_R _20513_ (.A(_13710_),
    .Y(_14741_));
 BUFx6f_ASAP7_75t_R _20514_ (.A(_13709_),
    .Y(_14742_));
 BUFx12_ASAP7_75t_R _20515_ (.A(_13679_),
    .Y(_14743_));
 AND2x2_ASAP7_75t_R _20516_ (.A(_14743_),
    .B(_01812_),
    .Y(_14744_));
 AO21x1_ASAP7_75t_R _20517_ (.A1(_14742_),
    .A2(_00754_),
    .B(_14744_),
    .Y(_14745_));
 BUFx10_ASAP7_75t_R _20518_ (.A(_13749_),
    .Y(_14746_));
 OAI22x1_ASAP7_75t_R _20519_ (.A1(_00753_),
    .A2(_14741_),
    .B1(_14745_),
    .B2(_14746_),
    .Y(_14747_));
 BUFx10_ASAP7_75t_R _20520_ (.A(_13718_),
    .Y(_14748_));
 BUFx10_ASAP7_75t_R _20521_ (.A(_13754_),
    .Y(_14749_));
 NAND2x1_ASAP7_75t_R _20522_ (.A(_13711_),
    .B(_00760_),
    .Y(_14750_));
 BUFx6f_ASAP7_75t_R _20523_ (.A(_13685_),
    .Y(_14751_));
 OA211x2_ASAP7_75t_R _20524_ (.A1(_14749_),
    .A2(_14682_),
    .B(_14750_),
    .C(_14751_),
    .Y(_14752_));
 NAND2x1_ASAP7_75t_R _20525_ (.A(_13711_),
    .B(_00759_),
    .Y(_14753_));
 BUFx6f_ASAP7_75t_R _20526_ (.A(_13692_),
    .Y(_14754_));
 OA211x2_ASAP7_75t_R _20527_ (.A1(_14749_),
    .A2(_14685_),
    .B(_14753_),
    .C(_14754_),
    .Y(_14755_));
 OR3x1_ASAP7_75t_R _20528_ (.A(_14748_),
    .B(_14752_),
    .C(_14755_),
    .Y(_14756_));
 BUFx6f_ASAP7_75t_R _20529_ (.A(_13731_),
    .Y(_14757_));
 OA211x2_ASAP7_75t_R _20530_ (.A1(_14740_),
    .A2(_14747_),
    .B(_14756_),
    .C(_14757_),
    .Y(_14758_));
 BUFx10_ASAP7_75t_R _20531_ (.A(_13674_),
    .Y(_14759_));
 BUFx6f_ASAP7_75t_R _20532_ (.A(_13675_),
    .Y(_14760_));
 BUFx6f_ASAP7_75t_R _20533_ (.A(_13742_),
    .Y(_14761_));
 NAND2x1_ASAP7_75t_R _20534_ (.A(_13866_),
    .B(_00756_),
    .Y(_14762_));
 OA211x2_ASAP7_75t_R _20535_ (.A1(_14761_),
    .A2(_14672_),
    .B(_14762_),
    .C(_13869_),
    .Y(_14763_));
 BUFx12_ASAP7_75t_R _20536_ (.A(_13688_),
    .Y(_14764_));
 NAND2x1_ASAP7_75t_R _20537_ (.A(_14764_),
    .B(_00755_),
    .Y(_14765_));
 OA211x2_ASAP7_75t_R _20538_ (.A1(_13865_),
    .A2(_14669_),
    .B(_14765_),
    .C(_13874_),
    .Y(_14766_));
 OR3x1_ASAP7_75t_R _20539_ (.A(_14760_),
    .B(_14763_),
    .C(_14766_),
    .Y(_14767_));
 BUFx6f_ASAP7_75t_R _20540_ (.A(_13718_),
    .Y(_14768_));
 NAND2x1_ASAP7_75t_R _20541_ (.A(_13866_),
    .B(_00764_),
    .Y(_14769_));
 OA211x2_ASAP7_75t_R _20542_ (.A1(_14761_),
    .A2(_14707_),
    .B(_14769_),
    .C(_13869_),
    .Y(_14770_));
 NAND2x1_ASAP7_75t_R _20543_ (.A(_14764_),
    .B(_00763_),
    .Y(_14771_));
 OA211x2_ASAP7_75t_R _20544_ (.A1(_13871_),
    .A2(_14700_),
    .B(_14771_),
    .C(_13874_),
    .Y(_14772_));
 OR3x1_ASAP7_75t_R _20545_ (.A(_14768_),
    .B(_14770_),
    .C(_14772_),
    .Y(_14773_));
 AND3x1_ASAP7_75t_R _20546_ (.A(_14759_),
    .B(_14767_),
    .C(_14773_),
    .Y(_14774_));
 OR3x4_ASAP7_75t_R _20547_ (.A(_14738_),
    .B(_14758_),
    .C(_14774_),
    .Y(_14775_));
 BUFx6f_ASAP7_75t_R _20548_ (.A(_13734_),
    .Y(_14776_));
 BUFx10_ASAP7_75t_R _20549_ (.A(_13706_),
    .Y(_14777_));
 BUFx12f_ASAP7_75t_R _20550_ (.A(_13688_),
    .Y(_14778_));
 NAND2x1_ASAP7_75t_R _20551_ (.A(_14778_),
    .B(_00772_),
    .Y(_14779_));
 BUFx6f_ASAP7_75t_R _20552_ (.A(_13868_),
    .Y(_14780_));
 OA211x2_ASAP7_75t_R _20553_ (.A1(_14761_),
    .A2(_14678_),
    .B(_14779_),
    .C(_14780_),
    .Y(_14781_));
 NAND2x1_ASAP7_75t_R _20554_ (.A(_13866_),
    .B(_00771_),
    .Y(_14782_));
 OA211x2_ASAP7_75t_R _20555_ (.A1(_14761_),
    .A2(_14675_),
    .B(_14782_),
    .C(_13874_),
    .Y(_14783_));
 OR3x1_ASAP7_75t_R _20556_ (.A(_14777_),
    .B(_14781_),
    .C(_14783_),
    .Y(_14784_));
 NAND2x1_ASAP7_75t_R _20557_ (.A(_14778_),
    .B(_00780_),
    .Y(_14785_));
 OA211x2_ASAP7_75t_R _20558_ (.A1(_14761_),
    .A2(_14697_),
    .B(_14785_),
    .C(_13869_),
    .Y(_14786_));
 NAND2x1_ASAP7_75t_R _20559_ (.A(_13866_),
    .B(_00779_),
    .Y(_14787_));
 OA211x2_ASAP7_75t_R _20560_ (.A1(_13865_),
    .A2(_14704_),
    .B(_14787_),
    .C(_13874_),
    .Y(_14788_));
 OR3x1_ASAP7_75t_R _20561_ (.A(_14768_),
    .B(_14786_),
    .C(_14788_),
    .Y(_14789_));
 AND3x1_ASAP7_75t_R _20562_ (.A(_14759_),
    .B(_14784_),
    .C(_14789_),
    .Y(_14790_));
 BUFx6f_ASAP7_75t_R _20563_ (.A(_13731_),
    .Y(_14791_));
 NAND2x1_ASAP7_75t_R _20564_ (.A(_13866_),
    .B(_00768_),
    .Y(_14792_));
 OA211x2_ASAP7_75t_R _20565_ (.A1(_14761_),
    .A2(_14711_),
    .B(_14792_),
    .C(_13869_),
    .Y(_14793_));
 NAND2x1_ASAP7_75t_R _20566_ (.A(_14764_),
    .B(_00767_),
    .Y(_14794_));
 OA211x2_ASAP7_75t_R _20567_ (.A1(_13865_),
    .A2(_14714_),
    .B(_14794_),
    .C(_13874_),
    .Y(_14795_));
 OR3x1_ASAP7_75t_R _20568_ (.A(_14760_),
    .B(_14793_),
    .C(_14795_),
    .Y(_14796_));
 NAND2x1_ASAP7_75t_R _20569_ (.A(_14764_),
    .B(_00776_),
    .Y(_14797_));
 OA211x2_ASAP7_75t_R _20570_ (.A1(_13865_),
    .A2(_14689_),
    .B(_14797_),
    .C(_13869_),
    .Y(_14798_));
 NAND2x1_ASAP7_75t_R _20571_ (.A(_13872_),
    .B(_00775_),
    .Y(_14799_));
 OA211x2_ASAP7_75t_R _20572_ (.A1(_13871_),
    .A2(_14692_),
    .B(_14799_),
    .C(_13874_),
    .Y(_14800_));
 OR3x1_ASAP7_75t_R _20573_ (.A(_14768_),
    .B(_14798_),
    .C(_14800_),
    .Y(_14801_));
 AND3x1_ASAP7_75t_R _20574_ (.A(_14791_),
    .B(_14796_),
    .C(_14801_),
    .Y(_14802_));
 OR3x4_ASAP7_75t_R _20575_ (.A(_14776_),
    .B(_14790_),
    .C(_14802_),
    .Y(_14803_));
 BUFx3_ASAP7_75t_R _20576_ (.A(_13647_),
    .Y(_14804_));
 BUFx3_ASAP7_75t_R _20577_ (.A(_13658_),
    .Y(_14805_));
 INVx2_ASAP7_75t_R _20578_ (.A(_00042_),
    .Y(_14806_));
 BUFx2_ASAP7_75t_R _20579_ (.A(_13366_),
    .Y(_14807_));
 OA211x2_ASAP7_75t_R _20580_ (.A1(_14804_),
    .A2(_14805_),
    .B(_14806_),
    .C(_14807_),
    .Y(_14808_));
 AO31x2_ASAP7_75t_R _20581_ (.A1(_14737_),
    .A2(_14775_),
    .A3(_14803_),
    .B(_14808_),
    .Y(_14809_));
 NOR2x1_ASAP7_75t_R _20582_ (.A(_01541_),
    .B(_13367_),
    .Y(_14810_));
 AO21x1_ASAP7_75t_R _20583_ (.A1(_13667_),
    .A2(_14809_),
    .B(_14810_),
    .Y(_14811_));
 BUFx4f_ASAP7_75t_R _20584_ (.A(_14811_),
    .Y(_18662_));
 INVx4_ASAP7_75t_R _20585_ (.A(_18662_),
    .Y(_18664_));
 INVx1_ASAP7_75t_R _20586_ (.A(_02135_),
    .Y(\cs_registers_i.mhpmcounter[2][1] ));
 INVx1_ASAP7_75t_R _20587_ (.A(_02198_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[1] ));
 BUFx3_ASAP7_75t_R _20588_ (.A(_02082_),
    .Y(_14812_));
 INVx1_ASAP7_75t_R _20589_ (.A(_14812_),
    .Y(\cs_registers_i.priv_lvl_q[0] ));
 INVx3_ASAP7_75t_R _20590_ (.A(_00012_),
    .Y(\cs_registers_i.pc_id_i[2] ));
 NOR2x1_ASAP7_75t_R _20591_ (.A(_01521_),
    .B(_13667_),
    .Y(_14813_));
 BUFx6f_ASAP7_75t_R _20592_ (.A(_13670_),
    .Y(_14814_));
 BUFx10_ASAP7_75t_R _20593_ (.A(_13706_),
    .Y(_14815_));
 BUFx12_ASAP7_75t_R _20594_ (.A(_13688_),
    .Y(_14816_));
 AND2x2_ASAP7_75t_R _20595_ (.A(_14816_),
    .B(_01792_),
    .Y(_14817_));
 AO21x1_ASAP7_75t_R _20596_ (.A1(_13709_),
    .A2(_00481_),
    .B(_14817_),
    .Y(_14818_));
 OAI22x1_ASAP7_75t_R _20597_ (.A1(_00480_),
    .A2(_13948_),
    .B1(_14818_),
    .B2(_13716_),
    .Y(_14819_));
 BUFx10_ASAP7_75t_R _20598_ (.A(_13688_),
    .Y(_14820_));
 INVx1_ASAP7_75t_R _20599_ (.A(_00489_),
    .Y(_14821_));
 BUFx10_ASAP7_75t_R _20600_ (.A(_13681_),
    .Y(_14822_));
 NAND2x1_ASAP7_75t_R _20601_ (.A(_14822_),
    .B(_00487_),
    .Y(_14823_));
 OA211x2_ASAP7_75t_R _20602_ (.A1(_14820_),
    .A2(_14821_),
    .B(_14823_),
    .C(_13724_),
    .Y(_14824_));
 NAND2x1_ASAP7_75t_R _20603_ (.A(_14822_),
    .B(_00486_),
    .Y(_14825_));
 OA211x2_ASAP7_75t_R _20604_ (.A1(_14820_),
    .A2(_14142_),
    .B(_14825_),
    .C(_13744_),
    .Y(_14826_));
 OR3x1_ASAP7_75t_R _20605_ (.A(_13696_),
    .B(_14824_),
    .C(_14826_),
    .Y(_14827_));
 OA211x2_ASAP7_75t_R _20606_ (.A1(_14815_),
    .A2(_14819_),
    .B(_14827_),
    .C(_13961_),
    .Y(_14828_));
 NOR2x1_ASAP7_75t_R _20607_ (.A(_13919_),
    .B(_00492_),
    .Y(_14829_));
 AO21x1_ASAP7_75t_R _20608_ (.A1(_13921_),
    .A2(_14133_),
    .B(_14829_),
    .Y(_14830_));
 BUFx10_ASAP7_75t_R _20609_ (.A(_13679_),
    .Y(_14831_));
 NAND2x1_ASAP7_75t_R _20610_ (.A(_13711_),
    .B(_00491_),
    .Y(_14832_));
 OA211x2_ASAP7_75t_R _20611_ (.A1(_14831_),
    .A2(_14127_),
    .B(_14832_),
    .C(_14751_),
    .Y(_14833_));
 AO21x1_ASAP7_75t_R _20612_ (.A1(_13749_),
    .A2(_14830_),
    .B(_14833_),
    .Y(_14834_));
 NAND2x1_ASAP7_75t_R _20613_ (.A(_14822_),
    .B(_00483_),
    .Y(_14835_));
 OA211x2_ASAP7_75t_R _20614_ (.A1(_14820_),
    .A2(_14115_),
    .B(_14835_),
    .C(_13724_),
    .Y(_14836_));
 NAND2x1_ASAP7_75t_R _20615_ (.A(_14822_),
    .B(_00482_),
    .Y(_14837_));
 OA211x2_ASAP7_75t_R _20616_ (.A1(_13751_),
    .A2(_14111_),
    .B(_14837_),
    .C(_13744_),
    .Y(_14838_));
 OR3x1_ASAP7_75t_R _20617_ (.A(_13706_),
    .B(_14836_),
    .C(_14838_),
    .Y(_14839_));
 OA211x2_ASAP7_75t_R _20618_ (.A1(_13748_),
    .A2(_14834_),
    .B(_14839_),
    .C(_13674_),
    .Y(_14840_));
 OR3x4_ASAP7_75t_R _20619_ (.A(_14814_),
    .B(_14828_),
    .C(_14840_),
    .Y(_14841_));
 BUFx6f_ASAP7_75t_R _20620_ (.A(_13734_),
    .Y(_14842_));
 BUFx10_ASAP7_75t_R _20621_ (.A(_13673_),
    .Y(_14843_));
 BUFx10_ASAP7_75t_R _20622_ (.A(_13679_),
    .Y(_14844_));
 NAND2x1_ASAP7_75t_R _20623_ (.A(_13756_),
    .B(_00499_),
    .Y(_14845_));
 BUFx6f_ASAP7_75t_R _20624_ (.A(_13685_),
    .Y(_14846_));
 OA211x2_ASAP7_75t_R _20625_ (.A1(_14844_),
    .A2(_14123_),
    .B(_14845_),
    .C(_14846_),
    .Y(_14847_));
 BUFx12f_ASAP7_75t_R _20626_ (.A(_13754_),
    .Y(_14848_));
 NAND2x1_ASAP7_75t_R _20627_ (.A(_13756_),
    .B(_00498_),
    .Y(_14849_));
 BUFx10_ASAP7_75t_R _20628_ (.A(_13692_),
    .Y(_14850_));
 OA211x2_ASAP7_75t_R _20629_ (.A1(_14848_),
    .A2(_14120_),
    .B(_14849_),
    .C(_14850_),
    .Y(_14851_));
 OR3x1_ASAP7_75t_R _20630_ (.A(_13676_),
    .B(_14847_),
    .C(_14851_),
    .Y(_14852_));
 BUFx10_ASAP7_75t_R _20631_ (.A(_13718_),
    .Y(_14853_));
 BUFx12f_ASAP7_75t_R _20632_ (.A(_13754_),
    .Y(_14854_));
 NAND2x1_ASAP7_75t_R _20633_ (.A(_13756_),
    .B(_00507_),
    .Y(_14855_));
 OA211x2_ASAP7_75t_R _20634_ (.A1(_14854_),
    .A2(_14083_),
    .B(_14855_),
    .C(_14846_),
    .Y(_14856_));
 BUFx10_ASAP7_75t_R _20635_ (.A(_13699_),
    .Y(_14857_));
 BUFx12_ASAP7_75t_R _20636_ (.A(_13681_),
    .Y(_14858_));
 NAND2x1_ASAP7_75t_R _20637_ (.A(_14858_),
    .B(_00506_),
    .Y(_14859_));
 OA211x2_ASAP7_75t_R _20638_ (.A1(_14857_),
    .A2(_14086_),
    .B(_14859_),
    .C(_14850_),
    .Y(_14860_));
 OR3x1_ASAP7_75t_R _20639_ (.A(_14853_),
    .B(_14856_),
    .C(_14860_),
    .Y(_14861_));
 AND3x1_ASAP7_75t_R _20640_ (.A(_14843_),
    .B(_14852_),
    .C(_14861_),
    .Y(_14862_));
 BUFx6f_ASAP7_75t_R _20641_ (.A(_13731_),
    .Y(_14863_));
 NAND2x1_ASAP7_75t_R _20642_ (.A(_13756_),
    .B(_00495_),
    .Y(_14864_));
 OA211x2_ASAP7_75t_R _20643_ (.A1(_14848_),
    .A2(_14093_),
    .B(_14864_),
    .C(_14846_),
    .Y(_14865_));
 NAND2x1_ASAP7_75t_R _20644_ (.A(_14858_),
    .B(_00494_),
    .Y(_14866_));
 BUFx6f_ASAP7_75t_R _20645_ (.A(_13692_),
    .Y(_14867_));
 OA211x2_ASAP7_75t_R _20646_ (.A1(_13925_),
    .A2(_14096_),
    .B(_14866_),
    .C(_14867_),
    .Y(_14868_));
 OR3x1_ASAP7_75t_R _20647_ (.A(_13676_),
    .B(_14865_),
    .C(_14868_),
    .Y(_14869_));
 NAND2x1_ASAP7_75t_R _20648_ (.A(_14858_),
    .B(_00503_),
    .Y(_14870_));
 OA211x2_ASAP7_75t_R _20649_ (.A1(_14857_),
    .A2(_14074_),
    .B(_14870_),
    .C(_14846_),
    .Y(_14871_));
 BUFx12f_ASAP7_75t_R _20650_ (.A(_13679_),
    .Y(_14872_));
 NAND2x1_ASAP7_75t_R _20651_ (.A(_14858_),
    .B(_00502_),
    .Y(_14873_));
 OA211x2_ASAP7_75t_R _20652_ (.A1(_14872_),
    .A2(_14078_),
    .B(_14873_),
    .C(_14867_),
    .Y(_14874_));
 OR3x1_ASAP7_75t_R _20653_ (.A(_14853_),
    .B(_14871_),
    .C(_14874_),
    .Y(_14875_));
 AND3x1_ASAP7_75t_R _20654_ (.A(_14863_),
    .B(_14869_),
    .C(_14875_),
    .Y(_14876_));
 OR3x4_ASAP7_75t_R _20655_ (.A(_14842_),
    .B(_14862_),
    .C(_14876_),
    .Y(_14877_));
 AND3x1_ASAP7_75t_R _20656_ (.A(_13667_),
    .B(_14841_),
    .C(_14877_),
    .Y(_14878_));
 AND3x1_ASAP7_75t_R _20657_ (.A(\cs_registers_i.pc_id_i[2] ),
    .B(_13771_),
    .C(_13772_),
    .Y(_14879_));
 AND2x2_ASAP7_75t_R _20658_ (.A(_13391_),
    .B(_13569_),
    .Y(_14880_));
 AOI22x1_ASAP7_75t_R _20659_ (.A1(_13383_),
    .A2(_13663_),
    .B1(_13661_),
    .B2(_14880_),
    .Y(_14881_));
 AND2x2_ASAP7_75t_R _20660_ (.A(_13394_),
    .B(_13396_),
    .Y(_14882_));
 OR3x1_ASAP7_75t_R _20661_ (.A(_13414_),
    .B(_14882_),
    .C(_13652_),
    .Y(_14883_));
 OA211x2_ASAP7_75t_R _20662_ (.A1(_14881_),
    .A2(_14883_),
    .B(_13776_),
    .C(_14732_),
    .Y(_14884_));
 OR3x1_ASAP7_75t_R _20663_ (.A(_13947_),
    .B(_14879_),
    .C(_14884_),
    .Y(_14885_));
 OA31x2_ASAP7_75t_R _20664_ (.A1(_13770_),
    .A2(_14813_),
    .A3(_14878_),
    .B1(_14885_),
    .Y(_14886_));
 BUFx6f_ASAP7_75t_R _20665_ (.A(_14886_),
    .Y(_18618_));
 INVx1_ASAP7_75t_R _20666_ (.A(_18618_),
    .Y(_18620_));
 OR2x2_ASAP7_75t_R _20667_ (.A(_13615_),
    .B(_14024_),
    .Y(_14887_));
 AND4x1_ASAP7_75t_R _20668_ (.A(_13593_),
    .B(_13560_),
    .C(_13563_),
    .D(_13606_),
    .Y(_14888_));
 OA31x2_ASAP7_75t_R _20669_ (.A1(_13608_),
    .A2(_13611_),
    .A3(_13614_),
    .B1(_14019_),
    .Y(_14889_));
 AND3x1_ASAP7_75t_R _20670_ (.A(_13399_),
    .B(_13601_),
    .C(_13586_),
    .Y(_14890_));
 OAI21x1_ASAP7_75t_R _20671_ (.A1(_14888_),
    .A2(_14889_),
    .B(_14890_),
    .Y(_14891_));
 AO21x1_ASAP7_75t_R _20672_ (.A1(_13628_),
    .A2(_13629_),
    .B(_13630_),
    .Y(_14892_));
 OR3x1_ASAP7_75t_R _20673_ (.A(_13403_),
    .B(_14880_),
    .C(_13404_),
    .Y(_14893_));
 NAND2x2_ASAP7_75t_R _20674_ (.A(net2005),
    .B(_13563_),
    .Y(_14894_));
 OR4x1_ASAP7_75t_R _20675_ (.A(_13592_),
    .B(_13395_),
    .C(_13563_),
    .D(_13580_),
    .Y(_14895_));
 NAND2x1_ASAP7_75t_R _20676_ (.A(_14894_),
    .B(_14895_),
    .Y(_14896_));
 AOI221x1_ASAP7_75t_R _20677_ (.A1(_14892_),
    .A2(_14893_),
    .B1(_14896_),
    .B2(_13559_),
    .C(_14882_),
    .Y(_14897_));
 AND3x4_ASAP7_75t_R _20678_ (.A(_14887_),
    .B(_14891_),
    .C(_14897_),
    .Y(_14898_));
 NAND2x1_ASAP7_75t_R _20679_ (.A(_13559_),
    .B(_13580_),
    .Y(_14899_));
 NAND3x1_ASAP7_75t_R _20680_ (.A(_13399_),
    .B(_13586_),
    .C(_14032_),
    .Y(_14900_));
 OR3x2_ASAP7_75t_R _20681_ (.A(_13565_),
    .B(_13368_),
    .C(net2019),
    .Y(_14901_));
 OR5x2_ASAP7_75t_R _20682_ (.A(_13375_),
    .B(_13565_),
    .C(net2017),
    .D(_13431_),
    .E(_13638_),
    .Y(_14902_));
 OA21x2_ASAP7_75t_R _20683_ (.A1(_13624_),
    .A2(_14901_),
    .B(_14902_),
    .Y(_14903_));
 AO31x2_ASAP7_75t_R _20684_ (.A1(_14899_),
    .A2(_14900_),
    .A3(_14903_),
    .B(_14031_),
    .Y(_14904_));
 AND5x1_ASAP7_75t_R _20685_ (.A(_13566_),
    .B(_13576_),
    .C(_13589_),
    .D(_13575_),
    .E(_13588_),
    .Y(_14905_));
 OA211x2_ASAP7_75t_R _20686_ (.A1(net2013),
    .A2(_14905_),
    .B(_14027_),
    .C(_13586_),
    .Y(_14906_));
 AOI21x1_ASAP7_75t_R _20687_ (.A1(_13571_),
    .A2(_13594_),
    .B(_14906_),
    .Y(_14907_));
 AND3x1_ASAP7_75t_R _20688_ (.A(_13584_),
    .B(_02296_),
    .C(_14019_),
    .Y(_14908_));
 AO31x2_ASAP7_75t_R _20689_ (.A1(_14904_),
    .A2(_14907_),
    .A3(_14908_),
    .B(_13636_),
    .Y(_14909_));
 AND3x1_ASAP7_75t_R _20690_ (.A(_13399_),
    .B(_13586_),
    .C(_14032_),
    .Y(_14910_));
 OAI21x1_ASAP7_75t_R _20691_ (.A1(_13624_),
    .A2(_14901_),
    .B(_14902_),
    .Y(_14911_));
 OA31x2_ASAP7_75t_R _20692_ (.A1(_13581_),
    .A2(_14910_),
    .A3(_14911_),
    .B1(_13635_),
    .Y(_14912_));
 AO21x1_ASAP7_75t_R _20693_ (.A1(_13571_),
    .A2(_13594_),
    .B(_14906_),
    .Y(_14913_));
 OR4x2_ASAP7_75t_R _20694_ (.A(_00406_),
    .B(_13571_),
    .C(_14912_),
    .D(_14913_),
    .Y(_14914_));
 NOR2x1_ASAP7_75t_R _20695_ (.A(_13615_),
    .B(_14024_),
    .Y(_14915_));
 NOR2x1_ASAP7_75t_R _20696_ (.A(_13636_),
    .B(_14894_),
    .Y(_14916_));
 OA21x2_ASAP7_75t_R _20697_ (.A1(_14888_),
    .A2(_14889_),
    .B(_14890_),
    .Y(_14917_));
 AO221x1_ASAP7_75t_R _20698_ (.A1(_14892_),
    .A2(_14893_),
    .B1(_14896_),
    .B2(_13559_),
    .C(_14882_),
    .Y(_14918_));
 OR4x2_ASAP7_75t_R _20699_ (.A(_14915_),
    .B(_14916_),
    .C(_14917_),
    .D(_14918_),
    .Y(_14919_));
 INVx3_ASAP7_75t_R _20700_ (.A(net1974),
    .Y(_14920_));
 AO32x1_ASAP7_75t_R _20701_ (.A1(_14898_),
    .A2(_14914_),
    .A3(_14909_),
    .B1(_14919_),
    .B2(_14920_),
    .Y(_14921_));
 BUFx6f_ASAP7_75t_R _20702_ (.A(_14921_),
    .Y(_14922_));
 NAND2x2_ASAP7_75t_R _20703_ (.A(_13604_),
    .B(_13605_),
    .Y(_14923_));
 OR4x2_ASAP7_75t_R _20704_ (.A(net2013),
    .B(_13601_),
    .C(_14023_),
    .D(_14923_),
    .Y(_14924_));
 BUFx10_ASAP7_75t_R _20705_ (.A(_14924_),
    .Y(_14925_));
 NAND2x2_ASAP7_75t_R _20706_ (.A(_14922_),
    .B(_14925_),
    .Y(_17344_));
 NOR2x1_ASAP7_75t_R _20707_ (.A(_01518_),
    .B(_13667_),
    .Y(_14926_));
 AND2x2_ASAP7_75t_R _20708_ (.A(_13726_),
    .B(_01789_),
    .Y(_14927_));
 AO21x1_ASAP7_75t_R _20709_ (.A1(_13709_),
    .A2(_00512_),
    .B(_14927_),
    .Y(_14928_));
 OAI22x1_ASAP7_75t_R _20710_ (.A1(_00511_),
    .A2(_13948_),
    .B1(_14928_),
    .B2(_13716_),
    .Y(_14929_));
 INVx1_ASAP7_75t_R _20711_ (.A(_00520_),
    .Y(_14930_));
 NAND2x1_ASAP7_75t_R _20712_ (.A(_14822_),
    .B(_00518_),
    .Y(_14931_));
 OA211x2_ASAP7_75t_R _20713_ (.A1(_14778_),
    .A2(_14930_),
    .B(_14931_),
    .C(_13724_),
    .Y(_14932_));
 INVx1_ASAP7_75t_R _20714_ (.A(_00519_),
    .Y(_14933_));
 NAND2x1_ASAP7_75t_R _20715_ (.A(_14822_),
    .B(_00517_),
    .Y(_14934_));
 OA211x2_ASAP7_75t_R _20716_ (.A1(_13866_),
    .A2(_14933_),
    .B(_14934_),
    .C(_13744_),
    .Y(_14935_));
 OR3x1_ASAP7_75t_R _20717_ (.A(_13696_),
    .B(_14932_),
    .C(_14935_),
    .Y(_14936_));
 OA211x2_ASAP7_75t_R _20718_ (.A1(_14815_),
    .A2(_14929_),
    .B(_14936_),
    .C(_13961_),
    .Y(_14937_));
 BUFx12_ASAP7_75t_R _20719_ (.A(_13699_),
    .Y(_14938_));
 NAND2x1_ASAP7_75t_R _20720_ (.A(_13682_),
    .B(_00514_),
    .Y(_14939_));
 BUFx6f_ASAP7_75t_R _20721_ (.A(_13685_),
    .Y(_14940_));
 OA211x2_ASAP7_75t_R _20722_ (.A1(_14938_),
    .A2(_14215_),
    .B(_14939_),
    .C(_14940_),
    .Y(_14941_));
 NAND2x1_ASAP7_75t_R _20723_ (.A(_13701_),
    .B(_00513_),
    .Y(_14942_));
 OA211x2_ASAP7_75t_R _20724_ (.A1(_13904_),
    .A2(_14218_),
    .B(_14942_),
    .C(_14867_),
    .Y(_14943_));
 OR3x1_ASAP7_75t_R _20725_ (.A(_13676_),
    .B(_14941_),
    .C(_14943_),
    .Y(_14944_));
 BUFx12f_ASAP7_75t_R _20726_ (.A(_13699_),
    .Y(_14945_));
 INVx1_ASAP7_75t_R _20727_ (.A(_00524_),
    .Y(_14946_));
 NAND2x1_ASAP7_75t_R _20728_ (.A(_13690_),
    .B(_00522_),
    .Y(_14947_));
 OA211x2_ASAP7_75t_R _20729_ (.A1(_14945_),
    .A2(_14946_),
    .B(_14947_),
    .C(_14940_),
    .Y(_14948_));
 NAND2x1_ASAP7_75t_R _20730_ (.A(_13701_),
    .B(_00521_),
    .Y(_14949_));
 OA211x2_ASAP7_75t_R _20731_ (.A1(_13904_),
    .A2(_14183_),
    .B(_14949_),
    .C(_13693_),
    .Y(_14950_));
 OR3x1_ASAP7_75t_R _20732_ (.A(_13696_),
    .B(_14948_),
    .C(_14950_),
    .Y(_14951_));
 AND3x1_ASAP7_75t_R _20733_ (.A(_14843_),
    .B(_14944_),
    .C(_14951_),
    .Y(_14952_));
 OR3x4_ASAP7_75t_R _20734_ (.A(_14814_),
    .B(_14937_),
    .C(_14952_),
    .Y(_14953_));
 NAND2x1_ASAP7_75t_R _20735_ (.A(_13682_),
    .B(_00530_),
    .Y(_14954_));
 OA211x2_ASAP7_75t_R _20736_ (.A1(_14938_),
    .A2(_14199_),
    .B(_14954_),
    .C(_14940_),
    .Y(_14955_));
 NAND2x1_ASAP7_75t_R _20737_ (.A(_13701_),
    .B(_00529_),
    .Y(_14956_));
 OA211x2_ASAP7_75t_R _20738_ (.A1(_13904_),
    .A2(_14202_),
    .B(_14956_),
    .C(_14867_),
    .Y(_14957_));
 OR3x1_ASAP7_75t_R _20739_ (.A(_13676_),
    .B(_14955_),
    .C(_14957_),
    .Y(_14958_));
 NAND2x1_ASAP7_75t_R _20740_ (.A(_13690_),
    .B(_00538_),
    .Y(_14959_));
 OA211x2_ASAP7_75t_R _20741_ (.A1(_14945_),
    .A2(_14189_),
    .B(_14959_),
    .C(_14940_),
    .Y(_14960_));
 NAND2x1_ASAP7_75t_R _20742_ (.A(_13701_),
    .B(_00537_),
    .Y(_14961_));
 OA211x2_ASAP7_75t_R _20743_ (.A1(_13904_),
    .A2(_14175_),
    .B(_14961_),
    .C(_13693_),
    .Y(_14962_));
 OR3x1_ASAP7_75t_R _20744_ (.A(_13696_),
    .B(_14960_),
    .C(_14962_),
    .Y(_14963_));
 AND3x1_ASAP7_75t_R _20745_ (.A(_14843_),
    .B(_14958_),
    .C(_14963_),
    .Y(_14964_));
 NAND2x1_ASAP7_75t_R _20746_ (.A(_13701_),
    .B(_00526_),
    .Y(_14965_));
 OA211x2_ASAP7_75t_R _20747_ (.A1(_13904_),
    .A2(_14161_),
    .B(_14965_),
    .C(_14940_),
    .Y(_14966_));
 NAND2x1_ASAP7_75t_R _20748_ (.A(_13742_),
    .B(_00525_),
    .Y(_14967_));
 OA211x2_ASAP7_75t_R _20749_ (.A1(_13882_),
    .A2(_14165_),
    .B(_14967_),
    .C(_13693_),
    .Y(_14968_));
 OR3x1_ASAP7_75t_R _20750_ (.A(_13676_),
    .B(_14966_),
    .C(_14968_),
    .Y(_14969_));
 NAND2x1_ASAP7_75t_R _20751_ (.A(_13701_),
    .B(_00534_),
    .Y(_14970_));
 OA211x2_ASAP7_75t_R _20752_ (.A1(_13904_),
    .A2(_14192_),
    .B(_14970_),
    .C(_14940_),
    .Y(_14971_));
 INVx1_ASAP7_75t_R _20753_ (.A(_00535_),
    .Y(_14972_));
 NAND2x1_ASAP7_75t_R _20754_ (.A(_13742_),
    .B(_00533_),
    .Y(_14973_));
 OA211x2_ASAP7_75t_R _20755_ (.A1(_13888_),
    .A2(_14972_),
    .B(_14973_),
    .C(_13693_),
    .Y(_14974_));
 OR3x1_ASAP7_75t_R _20756_ (.A(_13696_),
    .B(_14971_),
    .C(_14974_),
    .Y(_14975_));
 AND3x1_ASAP7_75t_R _20757_ (.A(_14863_),
    .B(_14969_),
    .C(_14975_),
    .Y(_14976_));
 OR3x4_ASAP7_75t_R _20758_ (.A(_14842_),
    .B(_14964_),
    .C(_14976_),
    .Y(_14977_));
 AND3x1_ASAP7_75t_R _20759_ (.A(_13667_),
    .B(_14953_),
    .C(_14977_),
    .Y(_14978_));
 INVx1_ASAP7_75t_R _20760_ (.A(_00020_),
    .Y(_14979_));
 AND3x1_ASAP7_75t_R _20761_ (.A(_14979_),
    .B(_13664_),
    .C(_13665_),
    .Y(_14980_));
 OA211x2_ASAP7_75t_R _20762_ (.A1(_14881_),
    .A2(_14883_),
    .B(_13776_),
    .C(_13857_),
    .Y(_14981_));
 OR3x1_ASAP7_75t_R _20763_ (.A(_13659_),
    .B(_14980_),
    .C(_14981_),
    .Y(_14982_));
 OA31x2_ASAP7_75t_R _20764_ (.A1(_13770_),
    .A2(_14926_),
    .A3(_14978_),
    .B1(_14982_),
    .Y(_14983_));
 BUFx4f_ASAP7_75t_R _20765_ (.A(_14983_),
    .Y(_18622_));
 INVx1_ASAP7_75t_R _20766_ (.A(_18622_),
    .Y(_18624_));
 NOR2x1_ASAP7_75t_R _20767_ (.A(_01517_),
    .B(_13667_),
    .Y(_14984_));
 BUFx12_ASAP7_75t_R _20768_ (.A(_13675_),
    .Y(_14985_));
 BUFx4f_ASAP7_75t_R _20769_ (.A(_14985_),
    .Y(_14986_));
 BUFx10_ASAP7_75t_R _20770_ (.A(_13964_),
    .Y(_14987_));
 AND2x2_ASAP7_75t_R _20771_ (.A(_14987_),
    .B(_01788_),
    .Y(_14988_));
 AO21x1_ASAP7_75t_R _20772_ (.A1(_13859_),
    .A2(_00542_),
    .B(_14988_),
    .Y(_14989_));
 BUFx10_ASAP7_75t_R _20773_ (.A(_13749_),
    .Y(_14990_));
 OAI22x1_ASAP7_75t_R _20774_ (.A1(_00541_),
    .A2(_13858_),
    .B1(_14989_),
    .B2(_14990_),
    .Y(_14991_));
 BUFx6f_ASAP7_75t_R _20775_ (.A(_14858_),
    .Y(_14992_));
 BUFx10_ASAP7_75t_R _20776_ (.A(_13699_),
    .Y(_14993_));
 NAND2x1_ASAP7_75t_R _20777_ (.A(_14993_),
    .B(_00548_),
    .Y(_14994_));
 BUFx6f_ASAP7_75t_R _20778_ (.A(_13868_),
    .Y(_14995_));
 OA211x2_ASAP7_75t_R _20779_ (.A1(_14992_),
    .A2(_14266_),
    .B(_14994_),
    .C(_14995_),
    .Y(_14996_));
 INVx1_ASAP7_75t_R _20780_ (.A(_00549_),
    .Y(_14997_));
 NAND2x1_ASAP7_75t_R _20781_ (.A(_13751_),
    .B(_00547_),
    .Y(_14998_));
 OA211x2_ASAP7_75t_R _20782_ (.A1(_13921_),
    .A2(_14997_),
    .B(_14998_),
    .C(_13715_),
    .Y(_14999_));
 OR3x2_ASAP7_75t_R _20783_ (.A(_13902_),
    .B(_14996_),
    .C(_14999_),
    .Y(_15000_));
 OA211x2_ASAP7_75t_R _20784_ (.A1(_14986_),
    .A2(_14991_),
    .B(_15000_),
    .C(_14791_),
    .Y(_15001_));
 BUFx10_ASAP7_75t_R _20785_ (.A(_13674_),
    .Y(_15002_));
 NAND2x1_ASAP7_75t_R _20786_ (.A(_14857_),
    .B(_00544_),
    .Y(_15003_));
 BUFx6f_ASAP7_75t_R _20787_ (.A(_13761_),
    .Y(_15004_));
 OA211x2_ASAP7_75t_R _20788_ (.A1(_13924_),
    .A2(_14274_),
    .B(_15003_),
    .C(_15004_),
    .Y(_15005_));
 BUFx6f_ASAP7_75t_R _20789_ (.A(_13763_),
    .Y(_15006_));
 INVx1_ASAP7_75t_R _20790_ (.A(_00545_),
    .Y(_15007_));
 NAND2x1_ASAP7_75t_R _20791_ (.A(_14743_),
    .B(_00543_),
    .Y(_15008_));
 BUFx6f_ASAP7_75t_R _20792_ (.A(_13728_),
    .Y(_15009_));
 OA211x2_ASAP7_75t_R _20793_ (.A1(_15006_),
    .A2(_15007_),
    .B(_15008_),
    .C(_15009_),
    .Y(_15010_));
 OR3x1_ASAP7_75t_R _20794_ (.A(_13707_),
    .B(_15005_),
    .C(_15010_),
    .Y(_15011_));
 BUFx10_ASAP7_75t_R _20795_ (.A(_13718_),
    .Y(_15012_));
 BUFx6f_ASAP7_75t_R _20796_ (.A(_13726_),
    .Y(_15013_));
 INVx1_ASAP7_75t_R _20797_ (.A(_00554_),
    .Y(_15014_));
 NAND2x1_ASAP7_75t_R _20798_ (.A(_13925_),
    .B(_00552_),
    .Y(_15015_));
 OA211x2_ASAP7_75t_R _20799_ (.A1(_15013_),
    .A2(_15014_),
    .B(_15015_),
    .C(_13927_),
    .Y(_15016_));
 BUFx6f_ASAP7_75t_R _20800_ (.A(_13763_),
    .Y(_15017_));
 INVx1_ASAP7_75t_R _20801_ (.A(_00553_),
    .Y(_15018_));
 BUFx12f_ASAP7_75t_R _20802_ (.A(_13754_),
    .Y(_15019_));
 NAND2x1_ASAP7_75t_R _20803_ (.A(_15019_),
    .B(_00551_),
    .Y(_15020_));
 OA211x2_ASAP7_75t_R _20804_ (.A1(_15017_),
    .A2(_15018_),
    .B(_15020_),
    .C(_13917_),
    .Y(_15021_));
 OR3x1_ASAP7_75t_R _20805_ (.A(_15012_),
    .B(_15016_),
    .C(_15021_),
    .Y(_15022_));
 AND3x2_ASAP7_75t_R _20806_ (.A(_15002_),
    .B(_15011_),
    .C(_15022_),
    .Y(_15023_));
 OR3x2_ASAP7_75t_R _20807_ (.A(_14733_),
    .B(_15001_),
    .C(_15023_),
    .Y(_15024_));
 BUFx10_ASAP7_75t_R _20808_ (.A(_13734_),
    .Y(_15025_));
 NAND2x1_ASAP7_75t_R _20809_ (.A(_14857_),
    .B(_00560_),
    .Y(_15026_));
 OA211x2_ASAP7_75t_R _20810_ (.A1(_13924_),
    .A2(_14289_),
    .B(_15026_),
    .C(_15004_),
    .Y(_15027_));
 NAND2x1_ASAP7_75t_R _20811_ (.A(_14872_),
    .B(_00559_),
    .Y(_15028_));
 OA211x2_ASAP7_75t_R _20812_ (.A1(_15006_),
    .A2(_14286_),
    .B(_15028_),
    .C(_15009_),
    .Y(_15029_));
 OR3x1_ASAP7_75t_R _20813_ (.A(_13707_),
    .B(_15027_),
    .C(_15029_),
    .Y(_15030_));
 BUFx6f_ASAP7_75t_R _20814_ (.A(_13718_),
    .Y(_15031_));
 NAND2x1_ASAP7_75t_R _20815_ (.A(_13925_),
    .B(_00568_),
    .Y(_15032_));
 OA211x2_ASAP7_75t_R _20816_ (.A1(_15013_),
    .A2(_14241_),
    .B(_15032_),
    .C(_13927_),
    .Y(_15033_));
 NAND2x1_ASAP7_75t_R _20817_ (.A(_15019_),
    .B(_00567_),
    .Y(_15034_));
 OA211x2_ASAP7_75t_R _20818_ (.A1(_15017_),
    .A2(_14237_),
    .B(_15034_),
    .C(_15009_),
    .Y(_15035_));
 OR3x1_ASAP7_75t_R _20819_ (.A(_15031_),
    .B(_15033_),
    .C(_15035_),
    .Y(_15036_));
 AND3x1_ASAP7_75t_R _20820_ (.A(_15002_),
    .B(_15030_),
    .C(_15036_),
    .Y(_15037_));
 BUFx6f_ASAP7_75t_R _20821_ (.A(_13731_),
    .Y(_15038_));
 BUFx10_ASAP7_75t_R _20822_ (.A(_13706_),
    .Y(_15039_));
 NAND2x1_ASAP7_75t_R _20823_ (.A(_14743_),
    .B(_00556_),
    .Y(_15040_));
 OA211x2_ASAP7_75t_R _20824_ (.A1(_15006_),
    .A2(_14253_),
    .B(_15040_),
    .C(_13927_),
    .Y(_15041_));
 BUFx6f_ASAP7_75t_R _20825_ (.A(_13880_),
    .Y(_15042_));
 NAND2x1_ASAP7_75t_R _20826_ (.A(_14938_),
    .B(_00555_),
    .Y(_15043_));
 OA211x2_ASAP7_75t_R _20827_ (.A1(_15042_),
    .A2(_14256_),
    .B(_15043_),
    .C(_13917_),
    .Y(_15044_));
 OR3x1_ASAP7_75t_R _20828_ (.A(_15039_),
    .B(_15041_),
    .C(_15044_),
    .Y(_15045_));
 NAND2x1_ASAP7_75t_R _20829_ (.A(_15019_),
    .B(_00564_),
    .Y(_15046_));
 OA211x2_ASAP7_75t_R _20830_ (.A1(_15017_),
    .A2(_14282_),
    .B(_15046_),
    .C(_13906_),
    .Y(_15047_));
 NAND2x1_ASAP7_75t_R _20831_ (.A(_14938_),
    .B(_00563_),
    .Y(_15048_));
 OA211x2_ASAP7_75t_R _20832_ (.A1(_15042_),
    .A2(_14279_),
    .B(_15048_),
    .C(_13917_),
    .Y(_15049_));
 OR3x1_ASAP7_75t_R _20833_ (.A(_15012_),
    .B(_15047_),
    .C(_15049_),
    .Y(_15050_));
 AND3x1_ASAP7_75t_R _20834_ (.A(_15038_),
    .B(_15045_),
    .C(_15050_),
    .Y(_15051_));
 OR3x4_ASAP7_75t_R _20835_ (.A(_15025_),
    .B(_15037_),
    .C(_15051_),
    .Y(_15052_));
 AND3x1_ASAP7_75t_R _20836_ (.A(_13667_),
    .B(_15024_),
    .C(_15052_),
    .Y(_15053_));
 INVx2_ASAP7_75t_R _20837_ (.A(_00023_),
    .Y(_15054_));
 AND3x1_ASAP7_75t_R _20838_ (.A(_15054_),
    .B(_13771_),
    .C(_13772_),
    .Y(_15055_));
 OA211x2_ASAP7_75t_R _20839_ (.A1(_14881_),
    .A2(_14883_),
    .B(_13776_),
    .C(_14738_),
    .Y(_15056_));
 OR3x1_ASAP7_75t_R _20840_ (.A(_14737_),
    .B(_15055_),
    .C(_15056_),
    .Y(_15057_));
 OA31x2_ASAP7_75t_R _20841_ (.A1(_13770_),
    .A2(_14984_),
    .A3(_15053_),
    .B1(_15057_),
    .Y(_15058_));
 BUFx6f_ASAP7_75t_R _20842_ (.A(_15058_),
    .Y(_18630_));
 INVx1_ASAP7_75t_R _20843_ (.A(_18630_),
    .Y(_18628_));
 BUFx3_ASAP7_75t_R _20844_ (.A(_13771_),
    .Y(_15059_));
 BUFx3_ASAP7_75t_R _20845_ (.A(_13772_),
    .Y(_15060_));
 BUFx6f_ASAP7_75t_R _20846_ (.A(_13754_),
    .Y(_15061_));
 AND2x2_ASAP7_75t_R _20847_ (.A(_15061_),
    .B(_01787_),
    .Y(_15062_));
 AO21x1_ASAP7_75t_R _20848_ (.A1(_13859_),
    .A2(_00574_),
    .B(_15062_),
    .Y(_15063_));
 OAI22x1_ASAP7_75t_R _20849_ (.A1(_00573_),
    .A2(_14741_),
    .B1(_15063_),
    .B2(_13863_),
    .Y(_15064_));
 NAND2x1_ASAP7_75t_R _20850_ (.A(_13872_),
    .B(_00580_),
    .Y(_15065_));
 OA211x2_ASAP7_75t_R _20851_ (.A1(_13871_),
    .A2(_14363_),
    .B(_15065_),
    .C(_13932_),
    .Y(_15066_));
 BUFx12_ASAP7_75t_R _20852_ (.A(_13688_),
    .Y(_15067_));
 NAND2x1_ASAP7_75t_R _20853_ (.A(_15067_),
    .B(_00579_),
    .Y(_15068_));
 OA211x2_ASAP7_75t_R _20854_ (.A1(_13930_),
    .A2(_14366_),
    .B(_15068_),
    .C(_13937_),
    .Y(_15069_));
 OR3x2_ASAP7_75t_R _20855_ (.A(_14768_),
    .B(_15066_),
    .C(_15069_),
    .Y(_15070_));
 OA211x2_ASAP7_75t_R _20856_ (.A1(_14986_),
    .A2(_15064_),
    .B(_15070_),
    .C(_13877_),
    .Y(_15071_));
 NAND2x1_ASAP7_75t_R _20857_ (.A(_13888_),
    .B(_00576_),
    .Y(_15072_));
 OA211x2_ASAP7_75t_R _20858_ (.A1(_13887_),
    .A2(_14327_),
    .B(_15072_),
    .C(_13884_),
    .Y(_15073_));
 BUFx6f_ASAP7_75t_R _20859_ (.A(_13886_),
    .Y(_15074_));
 BUFx12f_ASAP7_75t_R _20860_ (.A(_13679_),
    .Y(_15075_));
 NAND2x1_ASAP7_75t_R _20861_ (.A(_15075_),
    .B(_00575_),
    .Y(_15076_));
 OA211x2_ASAP7_75t_R _20862_ (.A1(_15074_),
    .A2(_14330_),
    .B(_15076_),
    .C(_13897_),
    .Y(_15077_));
 OR3x1_ASAP7_75t_R _20863_ (.A(_13856_),
    .B(_15073_),
    .C(_15077_),
    .Y(_15078_));
 BUFx12_ASAP7_75t_R _20864_ (.A(_13718_),
    .Y(_15079_));
 NAND2x1_ASAP7_75t_R _20865_ (.A(_13755_),
    .B(_00584_),
    .Y(_15080_));
 BUFx6f_ASAP7_75t_R _20866_ (.A(_13761_),
    .Y(_15081_));
 OA211x2_ASAP7_75t_R _20867_ (.A1(_13895_),
    .A2(_14354_),
    .B(_15080_),
    .C(_15081_),
    .Y(_15082_));
 NAND2x1_ASAP7_75t_R _20868_ (.A(_15075_),
    .B(_00583_),
    .Y(_15083_));
 OA211x2_ASAP7_75t_R _20869_ (.A1(_15074_),
    .A2(_14358_),
    .B(_15083_),
    .C(_13897_),
    .Y(_15084_));
 OR3x1_ASAP7_75t_R _20870_ (.A(_15079_),
    .B(_15082_),
    .C(_15084_),
    .Y(_15085_));
 AND3x2_ASAP7_75t_R _20871_ (.A(_13879_),
    .B(_15078_),
    .C(_15085_),
    .Y(_15086_));
 OR3x4_ASAP7_75t_R _20872_ (.A(_14738_),
    .B(_15071_),
    .C(_15086_),
    .Y(_15087_));
 NAND2x1_ASAP7_75t_R _20873_ (.A(_13882_),
    .B(_00592_),
    .Y(_15088_));
 OA211x2_ASAP7_75t_R _20874_ (.A1(_13881_),
    .A2(_14333_),
    .B(_15088_),
    .C(_13884_),
    .Y(_15089_));
 NAND2x1_ASAP7_75t_R _20875_ (.A(_13755_),
    .B(_00591_),
    .Y(_15090_));
 OA211x2_ASAP7_75t_R _20876_ (.A1(_13895_),
    .A2(_14336_),
    .B(_15090_),
    .C(_13890_),
    .Y(_15091_));
 OR3x1_ASAP7_75t_R _20877_ (.A(_15039_),
    .B(_15089_),
    .C(_15091_),
    .Y(_15092_));
 NAND2x1_ASAP7_75t_R _20878_ (.A(_13888_),
    .B(_00600_),
    .Y(_15093_));
 OA211x2_ASAP7_75t_R _20879_ (.A1(_13887_),
    .A2(_14341_),
    .B(_15093_),
    .C(_13884_),
    .Y(_15094_));
 INVx1_ASAP7_75t_R _20880_ (.A(_00601_),
    .Y(_15095_));
 NAND2x1_ASAP7_75t_R _20881_ (.A(_15075_),
    .B(_00599_),
    .Y(_15096_));
 OA211x2_ASAP7_75t_R _20882_ (.A1(_13895_),
    .A2(_15095_),
    .B(_15096_),
    .C(_13897_),
    .Y(_15097_));
 OR3x1_ASAP7_75t_R _20883_ (.A(_15012_),
    .B(_15094_),
    .C(_15097_),
    .Y(_15098_));
 AND3x1_ASAP7_75t_R _20884_ (.A(_13879_),
    .B(_15092_),
    .C(_15098_),
    .Y(_15099_));
 NAND2x1_ASAP7_75t_R _20885_ (.A(_13755_),
    .B(_00588_),
    .Y(_15100_));
 OA211x2_ASAP7_75t_R _20886_ (.A1(_13895_),
    .A2(_14319_),
    .B(_15100_),
    .C(_15081_),
    .Y(_15101_));
 NAND2x1_ASAP7_75t_R _20887_ (.A(_13680_),
    .B(_00587_),
    .Y(_15102_));
 OA211x2_ASAP7_75t_R _20888_ (.A1(_15074_),
    .A2(_14322_),
    .B(_15102_),
    .C(_13897_),
    .Y(_15103_));
 OR3x1_ASAP7_75t_R _20889_ (.A(_13856_),
    .B(_15101_),
    .C(_15103_),
    .Y(_15104_));
 INVx1_ASAP7_75t_R _20890_ (.A(_00598_),
    .Y(_15105_));
 NAND2x1_ASAP7_75t_R _20891_ (.A(_15075_),
    .B(_00596_),
    .Y(_15106_));
 OA211x2_ASAP7_75t_R _20892_ (.A1(_13895_),
    .A2(_15105_),
    .B(_15106_),
    .C(_15081_),
    .Y(_15107_));
 NAND2x1_ASAP7_75t_R _20893_ (.A(_13680_),
    .B(_00595_),
    .Y(_15108_));
 BUFx6f_ASAP7_75t_R _20894_ (.A(_13714_),
    .Y(_15109_));
 OA211x2_ASAP7_75t_R _20895_ (.A1(_15074_),
    .A2(_14348_),
    .B(_15108_),
    .C(_15109_),
    .Y(_15110_));
 OR3x1_ASAP7_75t_R _20896_ (.A(_15079_),
    .B(_15107_),
    .C(_15110_),
    .Y(_15111_));
 AND3x1_ASAP7_75t_R _20897_ (.A(_15038_),
    .B(_15104_),
    .C(_15111_),
    .Y(_15112_));
 OR3x4_ASAP7_75t_R _20898_ (.A(_14776_),
    .B(_15099_),
    .C(_15112_),
    .Y(_15113_));
 BUFx3_ASAP7_75t_R _20899_ (.A(_13647_),
    .Y(_15114_));
 BUFx3_ASAP7_75t_R _20900_ (.A(_13658_),
    .Y(_15115_));
 INVx2_ASAP7_75t_R _20901_ (.A(_00026_),
    .Y(_15116_));
 OA211x2_ASAP7_75t_R _20902_ (.A1(_15114_),
    .A2(_15115_),
    .B(_15116_),
    .C(_14807_),
    .Y(_15117_));
 AO31x2_ASAP7_75t_R _20903_ (.A1(_14737_),
    .A2(_15087_),
    .A3(_15113_),
    .B(_15117_),
    .Y(_15118_));
 BUFx3_ASAP7_75t_R _20904_ (.A(_13642_),
    .Y(_15119_));
 INVx1_ASAP7_75t_R _20905_ (.A(_01516_),
    .Y(_15120_));
 AO32x1_ASAP7_75t_R _20906_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_15118_),
    .B1(_15119_),
    .B2(_15120_),
    .Y(_15121_));
 BUFx6f_ASAP7_75t_R _20907_ (.A(_15121_),
    .Y(_18633_));
 INVx1_ASAP7_75t_R _20908_ (.A(_18633_),
    .Y(_18635_));
 AND2x2_ASAP7_75t_R _20909_ (.A(_14749_),
    .B(_01786_),
    .Y(_15122_));
 AO21x1_ASAP7_75t_R _20910_ (.A1(_13859_),
    .A2(_00604_),
    .B(_15122_),
    .Y(_15123_));
 OAI22x1_ASAP7_75t_R _20911_ (.A1(_00603_),
    .A2(_14741_),
    .B1(_15123_),
    .B2(_13863_),
    .Y(_15124_));
 BUFx10_ASAP7_75t_R _20912_ (.A(_13718_),
    .Y(_15125_));
 BUFx10_ASAP7_75t_R _20913_ (.A(_14822_),
    .Y(_15126_));
 INVx1_ASAP7_75t_R _20914_ (.A(_00612_),
    .Y(_15127_));
 NAND2x1_ASAP7_75t_R _20915_ (.A(_13956_),
    .B(_00610_),
    .Y(_15128_));
 BUFx6f_ASAP7_75t_R _20916_ (.A(_13868_),
    .Y(_15129_));
 OA211x2_ASAP7_75t_R _20917_ (.A1(_15126_),
    .A2(_15127_),
    .B(_15128_),
    .C(_15129_),
    .Y(_15130_));
 BUFx6f_ASAP7_75t_R _20918_ (.A(_13722_),
    .Y(_15131_));
 INVx1_ASAP7_75t_R _20919_ (.A(_00611_),
    .Y(_15132_));
 NAND2x1_ASAP7_75t_R _20920_ (.A(_13721_),
    .B(_00609_),
    .Y(_15133_));
 BUFx6f_ASAP7_75t_R _20921_ (.A(_13714_),
    .Y(_15134_));
 OA211x2_ASAP7_75t_R _20922_ (.A1(_15131_),
    .A2(_15132_),
    .B(_15133_),
    .C(_15134_),
    .Y(_15135_));
 OR3x1_ASAP7_75t_R _20923_ (.A(_15125_),
    .B(_15130_),
    .C(_15135_),
    .Y(_15136_));
 OA211x2_ASAP7_75t_R _20924_ (.A1(_14986_),
    .A2(_15124_),
    .B(_15136_),
    .C(_14757_),
    .Y(_15137_));
 BUFx10_ASAP7_75t_R _20925_ (.A(_13711_),
    .Y(_15138_));
 INVx1_ASAP7_75t_R _20926_ (.A(_00608_),
    .Y(_15139_));
 NAND2x1_ASAP7_75t_R _20927_ (.A(_13700_),
    .B(_00606_),
    .Y(_15140_));
 BUFx6f_ASAP7_75t_R _20928_ (.A(_13761_),
    .Y(_15141_));
 OA211x2_ASAP7_75t_R _20929_ (.A1(_15138_),
    .A2(_15139_),
    .B(_15140_),
    .C(_15141_),
    .Y(_15142_));
 BUFx10_ASAP7_75t_R _20930_ (.A(_13742_),
    .Y(_15143_));
 INVx1_ASAP7_75t_R _20931_ (.A(_00607_),
    .Y(_15144_));
 NAND2x1_ASAP7_75t_R _20932_ (.A(_13919_),
    .B(_00605_),
    .Y(_15145_));
 OA211x2_ASAP7_75t_R _20933_ (.A1(_15143_),
    .A2(_15144_),
    .B(_15145_),
    .C(_15109_),
    .Y(_15146_));
 OR3x1_ASAP7_75t_R _20934_ (.A(_13856_),
    .B(_15142_),
    .C(_15146_),
    .Y(_15147_));
 NAND2x1_ASAP7_75t_R _20935_ (.A(_13700_),
    .B(_00614_),
    .Y(_15148_));
 OA211x2_ASAP7_75t_R _20936_ (.A1(_15143_),
    .A2(_14414_),
    .B(_15148_),
    .C(_15141_),
    .Y(_15149_));
 NAND2x1_ASAP7_75t_R _20937_ (.A(_13919_),
    .B(_00613_),
    .Y(_15150_));
 OA211x2_ASAP7_75t_R _20938_ (.A1(_15143_),
    .A2(_14418_),
    .B(_15150_),
    .C(_15109_),
    .Y(_15151_));
 OR3x1_ASAP7_75t_R _20939_ (.A(_15079_),
    .B(_15149_),
    .C(_15151_),
    .Y(_15152_));
 AND3x2_ASAP7_75t_R _20940_ (.A(_14759_),
    .B(_15147_),
    .C(_15152_),
    .Y(_15153_));
 OR3x4_ASAP7_75t_R _20941_ (.A(_14738_),
    .B(_15137_),
    .C(_15153_),
    .Y(_15154_));
 INVx1_ASAP7_75t_R _20942_ (.A(_00624_),
    .Y(_15155_));
 NAND2x1_ASAP7_75t_R _20943_ (.A(_13689_),
    .B(_00622_),
    .Y(_15156_));
 OA211x2_ASAP7_75t_R _20944_ (.A1(_15138_),
    .A2(_15155_),
    .B(_15156_),
    .C(_15081_),
    .Y(_15157_));
 INVx1_ASAP7_75t_R _20945_ (.A(_00623_),
    .Y(_15158_));
 NAND2x1_ASAP7_75t_R _20946_ (.A(_13700_),
    .B(_00621_),
    .Y(_15159_));
 OA211x2_ASAP7_75t_R _20947_ (.A1(_15138_),
    .A2(_15158_),
    .B(_15159_),
    .C(_15109_),
    .Y(_15160_));
 OR3x1_ASAP7_75t_R _20948_ (.A(_13856_),
    .B(_15157_),
    .C(_15160_),
    .Y(_15161_));
 NAND2x1_ASAP7_75t_R _20949_ (.A(_13689_),
    .B(_00630_),
    .Y(_15162_));
 OA211x2_ASAP7_75t_R _20950_ (.A1(_15138_),
    .A2(_14403_),
    .B(_15162_),
    .C(_15141_),
    .Y(_15163_));
 NAND2x1_ASAP7_75t_R _20951_ (.A(_13700_),
    .B(_00629_),
    .Y(_15164_));
 OA211x2_ASAP7_75t_R _20952_ (.A1(_15138_),
    .A2(_14396_),
    .B(_15164_),
    .C(_15109_),
    .Y(_15165_));
 OR3x1_ASAP7_75t_R _20953_ (.A(_15079_),
    .B(_15163_),
    .C(_15165_),
    .Y(_15166_));
 AND3x1_ASAP7_75t_R _20954_ (.A(_14759_),
    .B(_15161_),
    .C(_15166_),
    .Y(_15167_));
 NAND2x1_ASAP7_75t_R _20955_ (.A(_13700_),
    .B(_00618_),
    .Y(_15168_));
 OA211x2_ASAP7_75t_R _20956_ (.A1(_15138_),
    .A2(_14378_),
    .B(_15168_),
    .C(_15141_),
    .Y(_15169_));
 NAND2x1_ASAP7_75t_R _20957_ (.A(_13919_),
    .B(_00617_),
    .Y(_15170_));
 OA211x2_ASAP7_75t_R _20958_ (.A1(_15143_),
    .A2(_14381_),
    .B(_15170_),
    .C(_15109_),
    .Y(_15171_));
 OR3x1_ASAP7_75t_R _20959_ (.A(_13856_),
    .B(_15169_),
    .C(_15171_),
    .Y(_15172_));
 NAND2x1_ASAP7_75t_R _20960_ (.A(_13700_),
    .B(_00626_),
    .Y(_15173_));
 OA211x2_ASAP7_75t_R _20961_ (.A1(_15143_),
    .A2(_14406_),
    .B(_15173_),
    .C(_15141_),
    .Y(_15174_));
 NAND2x1_ASAP7_75t_R _20962_ (.A(_13919_),
    .B(_00625_),
    .Y(_15175_));
 OA211x2_ASAP7_75t_R _20963_ (.A1(_15143_),
    .A2(_14399_),
    .B(_15175_),
    .C(_15109_),
    .Y(_15176_));
 OR3x1_ASAP7_75t_R _20964_ (.A(_15079_),
    .B(_15174_),
    .C(_15176_),
    .Y(_15177_));
 AND3x1_ASAP7_75t_R _20965_ (.A(_15038_),
    .B(_15172_),
    .C(_15177_),
    .Y(_15178_));
 OR3x4_ASAP7_75t_R _20966_ (.A(_14776_),
    .B(_15167_),
    .C(_15178_),
    .Y(_15179_));
 INVx1_ASAP7_75t_R _20967_ (.A(_00028_),
    .Y(_15180_));
 OA211x2_ASAP7_75t_R _20968_ (.A1(_15114_),
    .A2(_15115_),
    .B(_15180_),
    .C(_14807_),
    .Y(_15181_));
 AO31x2_ASAP7_75t_R _20969_ (.A1(_13660_),
    .A2(_15154_),
    .A3(_15179_),
    .B(_15181_),
    .Y(_15182_));
 INVx1_ASAP7_75t_R _20970_ (.A(_01515_),
    .Y(_15183_));
 AO32x1_ASAP7_75t_R _20971_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_15182_),
    .B1(_15119_),
    .B2(_15183_),
    .Y(_15184_));
 BUFx6f_ASAP7_75t_R _20972_ (.A(_15184_),
    .Y(_18637_));
 INVx1_ASAP7_75t_R _20973_ (.A(_18637_),
    .Y(_18639_));
 AND2x2_ASAP7_75t_R _20974_ (.A(_15126_),
    .B(_01785_),
    .Y(_15185_));
 AO21x1_ASAP7_75t_R _20975_ (.A1(_13859_),
    .A2(_00634_),
    .B(_15185_),
    .Y(_15186_));
 OAI22x1_ASAP7_75t_R _20976_ (.A1(_00633_),
    .A2(_13858_),
    .B1(_15186_),
    .B2(_14990_),
    .Y(_15187_));
 NAND2x1_ASAP7_75t_R _20977_ (.A(_14993_),
    .B(_00640_),
    .Y(_15188_));
 OA211x2_ASAP7_75t_R _20978_ (.A1(_14992_),
    .A2(_14465_),
    .B(_15188_),
    .C(_14780_),
    .Y(_15189_));
 BUFx12f_ASAP7_75t_R _20979_ (.A(_13699_),
    .Y(_15190_));
 NAND2x1_ASAP7_75t_R _20980_ (.A(_15190_),
    .B(_00639_),
    .Y(_15191_));
 OA211x2_ASAP7_75t_R _20981_ (.A1(_13921_),
    .A2(_14458_),
    .B(_15191_),
    .C(_13715_),
    .Y(_15192_));
 OR3x2_ASAP7_75t_R _20982_ (.A(_13902_),
    .B(_15189_),
    .C(_15192_),
    .Y(_15193_));
 OA211x2_ASAP7_75t_R _20983_ (.A1(_14986_),
    .A2(_15187_),
    .B(_15193_),
    .C(_14791_),
    .Y(_15194_));
 NAND2x1_ASAP7_75t_R _20984_ (.A(_13925_),
    .B(_00636_),
    .Y(_15195_));
 OA211x2_ASAP7_75t_R _20985_ (.A1(_13924_),
    .A2(_14447_),
    .B(_15195_),
    .C(_13927_),
    .Y(_15196_));
 NAND2x1_ASAP7_75t_R _20986_ (.A(_14743_),
    .B(_00635_),
    .Y(_15197_));
 OA211x2_ASAP7_75t_R _20987_ (.A1(_15006_),
    .A2(_14450_),
    .B(_15197_),
    .C(_15009_),
    .Y(_15198_));
 OR3x1_ASAP7_75t_R _20988_ (.A(_15039_),
    .B(_15196_),
    .C(_15198_),
    .Y(_15199_));
 NAND2x1_ASAP7_75t_R _20989_ (.A(_14872_),
    .B(_00644_),
    .Y(_15200_));
 OA211x2_ASAP7_75t_R _20990_ (.A1(_15013_),
    .A2(_14462_),
    .B(_15200_),
    .C(_13927_),
    .Y(_15201_));
 NAND2x1_ASAP7_75t_R _20991_ (.A(_15019_),
    .B(_00643_),
    .Y(_15202_));
 OA211x2_ASAP7_75t_R _20992_ (.A1(_15017_),
    .A2(_14455_),
    .B(_15202_),
    .C(_13917_),
    .Y(_15203_));
 OR3x1_ASAP7_75t_R _20993_ (.A(_15012_),
    .B(_15201_),
    .C(_15203_),
    .Y(_15204_));
 AND3x2_ASAP7_75t_R _20994_ (.A(_15002_),
    .B(_15199_),
    .C(_15204_),
    .Y(_15205_));
 OR3x4_ASAP7_75t_R _20995_ (.A(_14733_),
    .B(_15194_),
    .C(_15205_),
    .Y(_15206_));
 BUFx6f_ASAP7_75t_R _20996_ (.A(_13721_),
    .Y(_15207_));
 NAND2x1_ASAP7_75t_R _20997_ (.A(_14848_),
    .B(_00652_),
    .Y(_15208_));
 OA211x2_ASAP7_75t_R _20998_ (.A1(_15207_),
    .A2(_14441_),
    .B(_15208_),
    .C(_15004_),
    .Y(_15209_));
 NAND2x1_ASAP7_75t_R _20999_ (.A(_14872_),
    .B(_00651_),
    .Y(_15210_));
 OA211x2_ASAP7_75t_R _21000_ (.A1(_15013_),
    .A2(_14444_),
    .B(_15210_),
    .C(_15009_),
    .Y(_15211_));
 OR3x1_ASAP7_75t_R _21001_ (.A(_13707_),
    .B(_15209_),
    .C(_15211_),
    .Y(_15212_));
 INVx1_ASAP7_75t_R _21002_ (.A(_00662_),
    .Y(_15213_));
 NAND2x1_ASAP7_75t_R _21003_ (.A(_14857_),
    .B(_00660_),
    .Y(_15214_));
 OA211x2_ASAP7_75t_R _21004_ (.A1(_13924_),
    .A2(_15213_),
    .B(_15214_),
    .C(_15004_),
    .Y(_15215_));
 INVx1_ASAP7_75t_R _21005_ (.A(_00661_),
    .Y(_15216_));
 NAND2x1_ASAP7_75t_R _21006_ (.A(_14743_),
    .B(_00659_),
    .Y(_15217_));
 OA211x2_ASAP7_75t_R _21007_ (.A1(_15006_),
    .A2(_15216_),
    .B(_15217_),
    .C(_15009_),
    .Y(_15218_));
 OR3x1_ASAP7_75t_R _21008_ (.A(_15031_),
    .B(_15215_),
    .C(_15218_),
    .Y(_15219_));
 AND3x1_ASAP7_75t_R _21009_ (.A(_15002_),
    .B(_15212_),
    .C(_15219_),
    .Y(_15220_));
 NAND2x1_ASAP7_75t_R _21010_ (.A(_14872_),
    .B(_00648_),
    .Y(_15221_));
 OA211x2_ASAP7_75t_R _21011_ (.A1(_15006_),
    .A2(_14434_),
    .B(_15221_),
    .C(_13927_),
    .Y(_15222_));
 NAND2x1_ASAP7_75t_R _21012_ (.A(_15019_),
    .B(_00647_),
    .Y(_15223_));
 OA211x2_ASAP7_75t_R _21013_ (.A1(_15017_),
    .A2(_14437_),
    .B(_15223_),
    .C(_13917_),
    .Y(_15224_));
 OR3x1_ASAP7_75t_R _21014_ (.A(_15039_),
    .B(_15222_),
    .C(_15224_),
    .Y(_15225_));
 INVx1_ASAP7_75t_R _21015_ (.A(_00658_),
    .Y(_15226_));
 NAND2x1_ASAP7_75t_R _21016_ (.A(_14743_),
    .B(_00656_),
    .Y(_15227_));
 OA211x2_ASAP7_75t_R _21017_ (.A1(_15006_),
    .A2(_15226_),
    .B(_15227_),
    .C(_13906_),
    .Y(_15228_));
 INVx1_ASAP7_75t_R _21018_ (.A(_00657_),
    .Y(_15229_));
 NAND2x1_ASAP7_75t_R _21019_ (.A(_14938_),
    .B(_00655_),
    .Y(_15230_));
 OA211x2_ASAP7_75t_R _21020_ (.A1(_15042_),
    .A2(_15229_),
    .B(_15230_),
    .C(_13917_),
    .Y(_15231_));
 OR3x1_ASAP7_75t_R _21021_ (.A(_15012_),
    .B(_15228_),
    .C(_15231_),
    .Y(_15232_));
 AND3x1_ASAP7_75t_R _21022_ (.A(_15038_),
    .B(_15225_),
    .C(_15232_),
    .Y(_15233_));
 OR3x4_ASAP7_75t_R _21023_ (.A(_15025_),
    .B(_15220_),
    .C(_15233_),
    .Y(_15234_));
 INVx2_ASAP7_75t_R _21024_ (.A(_00030_),
    .Y(_15235_));
 OA211x2_ASAP7_75t_R _21025_ (.A1(_15114_),
    .A2(_15115_),
    .B(_15235_),
    .C(_14807_),
    .Y(_15236_));
 AO31x2_ASAP7_75t_R _21026_ (.A1(_13660_),
    .A2(_15206_),
    .A3(_15234_),
    .B(_15236_),
    .Y(_15237_));
 INVx1_ASAP7_75t_R _21027_ (.A(_01514_),
    .Y(_15238_));
 AO32x1_ASAP7_75t_R _21028_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_15237_),
    .B1(_15119_),
    .B2(_15238_),
    .Y(_15239_));
 BUFx6f_ASAP7_75t_R _21029_ (.A(_15239_),
    .Y(_18642_));
 INVx1_ASAP7_75t_R _21030_ (.A(_18642_),
    .Y(_18644_));
 OA211x2_ASAP7_75t_R _21031_ (.A1(_00415_),
    .A2(_02229_),
    .B(_00797_),
    .C(_00794_),
    .Y(_15240_));
 AO21x1_ASAP7_75t_R _21032_ (.A1(_00793_),
    .A2(_00797_),
    .B(_00796_),
    .Y(_15241_));
 AND3x1_ASAP7_75t_R _21033_ (.A(_00800_),
    .B(_00803_),
    .C(_00806_),
    .Y(_15242_));
 OA21x2_ASAP7_75t_R _21034_ (.A1(_15240_),
    .A2(_15241_),
    .B(_15242_),
    .Y(_15243_));
 AO21x1_ASAP7_75t_R _21035_ (.A1(_00799_),
    .A2(_00803_),
    .B(_00802_),
    .Y(_15244_));
 AO21x1_ASAP7_75t_R _21036_ (.A1(_00806_),
    .A2(_15244_),
    .B(_00805_),
    .Y(_15245_));
 OA21x2_ASAP7_75t_R _21037_ (.A1(_15243_),
    .A2(_15245_),
    .B(_00808_),
    .Y(_15246_));
 XNOR2x2_ASAP7_75t_R _21038_ (.A(_02298_),
    .B(_15246_),
    .Y(_15247_));
 INVx5_ASAP7_75t_R _21039_ (.A(_15247_),
    .Y(\alu_adder_result_ex[7] ));
 OR3x4_ASAP7_75t_R _21040_ (.A(_14915_),
    .B(_14917_),
    .C(_14918_),
    .Y(_15248_));
 INVx1_ASAP7_75t_R _21041_ (.A(_14908_),
    .Y(_15249_));
 OA31x2_ASAP7_75t_R _21042_ (.A1(_14912_),
    .A2(_14913_),
    .A3(_15249_),
    .B1(_13571_),
    .Y(_15250_));
 INVx2_ASAP7_75t_R _21043_ (.A(_00406_),
    .Y(_15251_));
 AND4x2_ASAP7_75t_R _21044_ (.A(_15251_),
    .B(_13636_),
    .C(_14904_),
    .D(_14907_),
    .Y(_15252_));
 OA21x2_ASAP7_75t_R _21045_ (.A1(_00797_),
    .A2(_00796_),
    .B(_00800_),
    .Y(_15253_));
 OR2x2_ASAP7_75t_R _21046_ (.A(_00799_),
    .B(_00802_),
    .Y(_15254_));
 OA21x2_ASAP7_75t_R _21047_ (.A1(_00803_),
    .A2(_00802_),
    .B(_00806_),
    .Y(_15255_));
 OA21x2_ASAP7_75t_R _21048_ (.A1(_15253_),
    .A2(_15254_),
    .B(_15255_),
    .Y(_15256_));
 OA21x2_ASAP7_75t_R _21049_ (.A1(_00415_),
    .A2(_00448_),
    .B(_00794_),
    .Y(_15257_));
 NAND3x2_ASAP7_75t_R _21050_ (.B(_15256_),
    .C(_15257_),
    .Y(_15258_),
    .A(_14925_));
 OR4x1_ASAP7_75t_R _21051_ (.A(_15248_),
    .B(_15250_),
    .C(_15252_),
    .D(_15258_),
    .Y(_15259_));
 BUFx3_ASAP7_75t_R _21052_ (.A(_15259_),
    .Y(_15260_));
 OR3x1_ASAP7_75t_R _21053_ (.A(_13621_),
    .B(_13624_),
    .C(_14894_),
    .Y(_15261_));
 AND4x2_ASAP7_75t_R _21054_ (.A(_14887_),
    .B(_15261_),
    .C(_14891_),
    .D(_14897_),
    .Y(_15262_));
 OR2x2_ASAP7_75t_R _21055_ (.A(_00415_),
    .B(_02297_),
    .Y(_15263_));
 OR3x1_ASAP7_75t_R _21056_ (.A(net1991),
    .B(_00796_),
    .C(_15254_),
    .Y(_15264_));
 AO21x1_ASAP7_75t_R _21057_ (.A1(_15257_),
    .A2(_15263_),
    .B(_15264_),
    .Y(_15265_));
 AND2x2_ASAP7_75t_R _21058_ (.A(_15256_),
    .B(_15265_),
    .Y(_15266_));
 INVx1_ASAP7_75t_R _21059_ (.A(_15266_),
    .Y(_15267_));
 OA31x2_ASAP7_75t_R _21060_ (.A1(net1975),
    .A2(_15262_),
    .A3(_15258_),
    .B1(_15267_),
    .Y(_15268_));
 INVx1_ASAP7_75t_R _21061_ (.A(net1982),
    .Y(_15269_));
 AOI21x1_ASAP7_75t_R _21062_ (.A1(_15260_),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15270_));
 AND3x1_ASAP7_75t_R _21063_ (.A(_15269_),
    .B(_15260_),
    .C(_15268_),
    .Y(_15271_));
 OR2x6_ASAP7_75t_R _21064_ (.A(_15270_),
    .B(_15271_),
    .Y(_15272_));
 INVx3_ASAP7_75t_R _21065_ (.A(_15272_),
    .Y(\alu_adder_result_ex[6] ));
 BUFx4f_ASAP7_75t_R _21066_ (.A(_13771_),
    .Y(_15273_));
 BUFx3_ASAP7_75t_R _21067_ (.A(_13772_),
    .Y(_15274_));
 AND2x2_ASAP7_75t_R _21068_ (.A(_13888_),
    .B(_01784_),
    .Y(_15275_));
 AO21x1_ASAP7_75t_R _21069_ (.A1(_14742_),
    .A2(_00664_),
    .B(_15275_),
    .Y(_15276_));
 OAI22x1_ASAP7_75t_R _21070_ (.A1(_00663_),
    .A2(_13948_),
    .B1(_15276_),
    .B2(_14746_),
    .Y(_15277_));
 BUFx10_ASAP7_75t_R _21071_ (.A(_13679_),
    .Y(_15278_));
 INVx1_ASAP7_75t_R _21072_ (.A(_00672_),
    .Y(_15279_));
 BUFx12f_ASAP7_75t_R _21073_ (.A(_13720_),
    .Y(_15280_));
 NAND2x1_ASAP7_75t_R _21074_ (.A(_15280_),
    .B(_00670_),
    .Y(_15281_));
 BUFx6f_ASAP7_75t_R _21075_ (.A(_13685_),
    .Y(_15282_));
 OA211x2_ASAP7_75t_R _21076_ (.A1(_15278_),
    .A2(_15279_),
    .B(_15281_),
    .C(_15282_),
    .Y(_15283_));
 INVx1_ASAP7_75t_R _21077_ (.A(_00671_),
    .Y(_15284_));
 NAND2x1_ASAP7_75t_R _21078_ (.A(_15280_),
    .B(_00669_),
    .Y(_15285_));
 OA211x2_ASAP7_75t_R _21079_ (.A1(_15278_),
    .A2(_15284_),
    .B(_15285_),
    .C(_14850_),
    .Y(_15286_));
 OR3x1_ASAP7_75t_R _21080_ (.A(_14853_),
    .B(_15283_),
    .C(_15286_),
    .Y(_15287_));
 OA211x2_ASAP7_75t_R _21081_ (.A1(_14740_),
    .A2(_15277_),
    .B(_15287_),
    .C(_14863_),
    .Y(_15288_));
 BUFx10_ASAP7_75t_R _21082_ (.A(_13674_),
    .Y(_15289_));
 BUFx6f_ASAP7_75t_R _21083_ (.A(_13964_),
    .Y(_15290_));
 NAND2x1_ASAP7_75t_R _21084_ (.A(_14816_),
    .B(_00666_),
    .Y(_15291_));
 OA211x2_ASAP7_75t_R _21085_ (.A1(_15290_),
    .A2(_14537_),
    .B(_15291_),
    .C(_15129_),
    .Y(_15292_));
 NAND2x1_ASAP7_75t_R _21086_ (.A(_13956_),
    .B(_00665_),
    .Y(_15293_));
 OA211x2_ASAP7_75t_R _21087_ (.A1(_14987_),
    .A2(_14540_),
    .B(_15293_),
    .C(_15134_),
    .Y(_15294_));
 OR3x1_ASAP7_75t_R _21088_ (.A(_14985_),
    .B(_15292_),
    .C(_15294_),
    .Y(_15295_));
 INVx1_ASAP7_75t_R _21089_ (.A(_00676_),
    .Y(_15296_));
 NAND2x1_ASAP7_75t_R _21090_ (.A(_13952_),
    .B(_00674_),
    .Y(_15297_));
 OA211x2_ASAP7_75t_R _21091_ (.A1(_15290_),
    .A2(_15296_),
    .B(_15297_),
    .C(_15129_),
    .Y(_15298_));
 NAND2x1_ASAP7_75t_R _21092_ (.A(_13956_),
    .B(_00673_),
    .Y(_15299_));
 OA211x2_ASAP7_75t_R _21093_ (.A1(_14987_),
    .A2(_14508_),
    .B(_15299_),
    .C(_15134_),
    .Y(_15300_));
 OR3x1_ASAP7_75t_R _21094_ (.A(_15125_),
    .B(_15298_),
    .C(_15300_),
    .Y(_15301_));
 AND3x1_ASAP7_75t_R _21095_ (.A(_15289_),
    .B(_15295_),
    .C(_15301_),
    .Y(_15302_));
 OR3x4_ASAP7_75t_R _21096_ (.A(_14814_),
    .B(_15288_),
    .C(_15302_),
    .Y(_15303_));
 NAND2x1_ASAP7_75t_R _21097_ (.A(_13935_),
    .B(_00682_),
    .Y(_15304_));
 BUFx6f_ASAP7_75t_R _21098_ (.A(_13868_),
    .Y(_15305_));
 OA211x2_ASAP7_75t_R _21099_ (.A1(_13934_),
    .A2(_14523_),
    .B(_15304_),
    .C(_15305_),
    .Y(_15306_));
 BUFx6f_ASAP7_75t_R _21100_ (.A(_13742_),
    .Y(_15307_));
 NAND2x1_ASAP7_75t_R _21101_ (.A(_14816_),
    .B(_00681_),
    .Y(_15308_));
 BUFx6f_ASAP7_75t_R _21102_ (.A(_13714_),
    .Y(_15309_));
 OA211x2_ASAP7_75t_R _21103_ (.A1(_15307_),
    .A2(_14526_),
    .B(_15308_),
    .C(_15309_),
    .Y(_15310_));
 OR3x1_ASAP7_75t_R _21104_ (.A(_14760_),
    .B(_15306_),
    .C(_15310_),
    .Y(_15311_));
 NAND2x1_ASAP7_75t_R _21105_ (.A(_13935_),
    .B(_00690_),
    .Y(_15312_));
 OA211x2_ASAP7_75t_R _21106_ (.A1(_15307_),
    .A2(_14516_),
    .B(_15312_),
    .C(_15305_),
    .Y(_15313_));
 NAND2x1_ASAP7_75t_R _21107_ (.A(_13952_),
    .B(_00689_),
    .Y(_15314_));
 OA211x2_ASAP7_75t_R _21108_ (.A1(_15290_),
    .A2(_14504_),
    .B(_15314_),
    .C(_15309_),
    .Y(_15315_));
 OR3x1_ASAP7_75t_R _21109_ (.A(_15125_),
    .B(_15313_),
    .C(_15315_),
    .Y(_15316_));
 AND3x1_ASAP7_75t_R _21110_ (.A(_15289_),
    .B(_15311_),
    .C(_15316_),
    .Y(_15317_));
 BUFx6f_ASAP7_75t_R _21111_ (.A(_14853_),
    .Y(_15318_));
 BUFx6f_ASAP7_75t_R _21112_ (.A(_13721_),
    .Y(_15319_));
 INVx1_ASAP7_75t_R _21113_ (.A(_00685_),
    .Y(_15320_));
 NOR2x1_ASAP7_75t_R _21114_ (.A(_14749_),
    .B(_00687_),
    .Y(_15321_));
 AO21x1_ASAP7_75t_R _21115_ (.A1(_15319_),
    .A2(_15320_),
    .B(_15321_),
    .Y(_15322_));
 NAND2x1_ASAP7_75t_R _21116_ (.A(_14778_),
    .B(_00686_),
    .Y(_15323_));
 OA211x2_ASAP7_75t_R _21117_ (.A1(_14761_),
    .A2(_14519_),
    .B(_15323_),
    .C(_13869_),
    .Y(_15324_));
 AO21x1_ASAP7_75t_R _21118_ (.A1(_13716_),
    .A2(_15322_),
    .B(_15324_),
    .Y(_15325_));
 NAND2x1_ASAP7_75t_R _21119_ (.A(_15280_),
    .B(_00678_),
    .Y(_15326_));
 OA211x2_ASAP7_75t_R _21120_ (.A1(_15278_),
    .A2(_14492_),
    .B(_15326_),
    .C(_15282_),
    .Y(_15327_));
 NAND2x1_ASAP7_75t_R _21121_ (.A(_13756_),
    .B(_00677_),
    .Y(_15328_));
 OA211x2_ASAP7_75t_R _21122_ (.A1(_14844_),
    .A2(_14496_),
    .B(_15328_),
    .C(_14850_),
    .Y(_15329_));
 OR3x1_ASAP7_75t_R _21123_ (.A(_14739_),
    .B(_15327_),
    .C(_15329_),
    .Y(_15330_));
 OA211x2_ASAP7_75t_R _21124_ (.A1(_15318_),
    .A2(_15325_),
    .B(_15330_),
    .C(_14863_),
    .Y(_15331_));
 OR3x4_ASAP7_75t_R _21125_ (.A(_14842_),
    .B(_15317_),
    .C(_15331_),
    .Y(_15332_));
 INVx1_ASAP7_75t_R _21126_ (.A(_00033_),
    .Y(_15333_));
 BUFx4f_ASAP7_75t_R _21127_ (.A(_13366_),
    .Y(_15334_));
 OA211x2_ASAP7_75t_R _21128_ (.A1(_14804_),
    .A2(_14805_),
    .B(_15333_),
    .C(_15334_),
    .Y(_15335_));
 AO31x2_ASAP7_75t_R _21129_ (.A1(_14737_),
    .A2(_15303_),
    .A3(_15332_),
    .B(_15335_),
    .Y(_15336_));
 BUFx3_ASAP7_75t_R _21130_ (.A(_13642_),
    .Y(_15337_));
 INVx1_ASAP7_75t_R _21131_ (.A(_01513_),
    .Y(_15338_));
 AO32x1_ASAP7_75t_R _21132_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_15336_),
    .B1(_15337_),
    .B2(_15338_),
    .Y(_15339_));
 BUFx6f_ASAP7_75t_R _21133_ (.A(_15339_),
    .Y(_18647_));
 INVx1_ASAP7_75t_R _21134_ (.A(_18647_),
    .Y(_18649_));
 AND2x2_ASAP7_75t_R _21135_ (.A(_13680_),
    .B(_01783_),
    .Y(_15340_));
 AO21x1_ASAP7_75t_R _21136_ (.A1(_14742_),
    .A2(_00694_),
    .B(_15340_),
    .Y(_15341_));
 OAI22x1_ASAP7_75t_R _21137_ (.A1(_00693_),
    .A2(_13948_),
    .B1(_15341_),
    .B2(_13918_),
    .Y(_15342_));
 INVx1_ASAP7_75t_R _21138_ (.A(_00702_),
    .Y(_15343_));
 NAND2x1_ASAP7_75t_R _21139_ (.A(_14858_),
    .B(_00700_),
    .Y(_15344_));
 OA211x2_ASAP7_75t_R _21140_ (.A1(_14848_),
    .A2(_15343_),
    .B(_15344_),
    .C(_14846_),
    .Y(_15345_));
 INVx1_ASAP7_75t_R _21141_ (.A(_00701_),
    .Y(_15346_));
 NAND2x1_ASAP7_75t_R _21142_ (.A(_14858_),
    .B(_00699_),
    .Y(_15347_));
 OA211x2_ASAP7_75t_R _21143_ (.A1(_13925_),
    .A2(_15346_),
    .B(_15347_),
    .C(_14867_),
    .Y(_15348_));
 OR3x1_ASAP7_75t_R _21144_ (.A(_14853_),
    .B(_15345_),
    .C(_15348_),
    .Y(_15349_));
 OA211x2_ASAP7_75t_R _21145_ (.A1(_14740_),
    .A2(_15342_),
    .B(_15349_),
    .C(_13961_),
    .Y(_15350_));
 NAND2x1_ASAP7_75t_R _21146_ (.A(_13726_),
    .B(_00696_),
    .Y(_15351_));
 BUFx6f_ASAP7_75t_R _21147_ (.A(_13868_),
    .Y(_15352_));
 OA211x2_ASAP7_75t_R _21148_ (.A1(_15131_),
    .A2(_14587_),
    .B(_15351_),
    .C(_15352_),
    .Y(_15353_));
 NAND2x1_ASAP7_75t_R _21149_ (.A(_13763_),
    .B(_00695_),
    .Y(_15354_));
 BUFx6f_ASAP7_75t_R _21150_ (.A(_13692_),
    .Y(_15355_));
 OA211x2_ASAP7_75t_R _21151_ (.A1(_13750_),
    .A2(_14590_),
    .B(_15354_),
    .C(_15355_),
    .Y(_15356_));
 OR3x1_ASAP7_75t_R _21152_ (.A(_14985_),
    .B(_15353_),
    .C(_15356_),
    .Y(_15357_));
 BUFx6f_ASAP7_75t_R _21153_ (.A(_13722_),
    .Y(_15358_));
 NAND2x1_ASAP7_75t_R _21154_ (.A(_13726_),
    .B(_00704_),
    .Y(_15359_));
 OA211x2_ASAP7_75t_R _21155_ (.A1(_15358_),
    .A2(_14568_),
    .B(_15359_),
    .C(_15352_),
    .Y(_15360_));
 NAND2x1_ASAP7_75t_R _21156_ (.A(_13763_),
    .B(_00703_),
    .Y(_15361_));
 OA211x2_ASAP7_75t_R _21157_ (.A1(_13860_),
    .A2(_14580_),
    .B(_15361_),
    .C(_15355_),
    .Y(_15362_));
 OR3x1_ASAP7_75t_R _21158_ (.A(_14748_),
    .B(_15360_),
    .C(_15362_),
    .Y(_15363_));
 AND3x1_ASAP7_75t_R _21159_ (.A(_14843_),
    .B(_15357_),
    .C(_15363_),
    .Y(_15364_));
 OR3x4_ASAP7_75t_R _21160_ (.A(_14814_),
    .B(_15350_),
    .C(_15364_),
    .Y(_15365_));
 NAND2x1_ASAP7_75t_R _21161_ (.A(_13721_),
    .B(_00712_),
    .Y(_15366_));
 OA211x2_ASAP7_75t_R _21162_ (.A1(_15131_),
    .A2(_14594_),
    .B(_15366_),
    .C(_15352_),
    .Y(_15367_));
 NAND2x1_ASAP7_75t_R _21163_ (.A(_13726_),
    .B(_00711_),
    .Y(_15368_));
 OA211x2_ASAP7_75t_R _21164_ (.A1(_15358_),
    .A2(_14597_),
    .B(_15368_),
    .C(_15134_),
    .Y(_15369_));
 OR3x1_ASAP7_75t_R _21165_ (.A(_14985_),
    .B(_15367_),
    .C(_15369_),
    .Y(_15370_));
 NAND2x1_ASAP7_75t_R _21166_ (.A(_13721_),
    .B(_00720_),
    .Y(_15371_));
 OA211x2_ASAP7_75t_R _21167_ (.A1(_15131_),
    .A2(_14562_),
    .B(_15371_),
    .C(_15352_),
    .Y(_15372_));
 NAND2x1_ASAP7_75t_R _21168_ (.A(_13763_),
    .B(_00719_),
    .Y(_15373_));
 OA211x2_ASAP7_75t_R _21169_ (.A1(_13750_),
    .A2(_14573_),
    .B(_15373_),
    .C(_15355_),
    .Y(_15374_));
 OR3x1_ASAP7_75t_R _21170_ (.A(_15125_),
    .B(_15372_),
    .C(_15374_),
    .Y(_15375_));
 AND3x1_ASAP7_75t_R _21171_ (.A(_14843_),
    .B(_15370_),
    .C(_15375_),
    .Y(_15376_));
 NAND2x1_ASAP7_75t_R _21172_ (.A(_13726_),
    .B(_00708_),
    .Y(_15377_));
 OA211x2_ASAP7_75t_R _21173_ (.A1(_15358_),
    .A2(_14552_),
    .B(_15377_),
    .C(_15352_),
    .Y(_15378_));
 NAND2x1_ASAP7_75t_R _21174_ (.A(_13880_),
    .B(_00707_),
    .Y(_15379_));
 OA211x2_ASAP7_75t_R _21175_ (.A1(_13860_),
    .A2(_14555_),
    .B(_15379_),
    .C(_15355_),
    .Y(_15380_));
 OR3x1_ASAP7_75t_R _21176_ (.A(_14739_),
    .B(_15378_),
    .C(_15380_),
    .Y(_15381_));
 INVx1_ASAP7_75t_R _21177_ (.A(_00718_),
    .Y(_15382_));
 NAND2x1_ASAP7_75t_R _21178_ (.A(_13763_),
    .B(_00716_),
    .Y(_15383_));
 OA211x2_ASAP7_75t_R _21179_ (.A1(_13750_),
    .A2(_15382_),
    .B(_15383_),
    .C(_15352_),
    .Y(_15384_));
 INVx1_ASAP7_75t_R _21180_ (.A(_00717_),
    .Y(_15385_));
 NAND2x1_ASAP7_75t_R _21181_ (.A(_13880_),
    .B(_00715_),
    .Y(_15386_));
 OA211x2_ASAP7_75t_R _21182_ (.A1(_13860_),
    .A2(_15385_),
    .B(_15386_),
    .C(_15355_),
    .Y(_15387_));
 OR3x1_ASAP7_75t_R _21183_ (.A(_14748_),
    .B(_15384_),
    .C(_15387_),
    .Y(_15388_));
 AND3x1_ASAP7_75t_R _21184_ (.A(_13877_),
    .B(_15381_),
    .C(_15388_),
    .Y(_15389_));
 OR3x4_ASAP7_75t_R _21185_ (.A(_14842_),
    .B(_15376_),
    .C(_15389_),
    .Y(_15390_));
 INVx1_ASAP7_75t_R _21186_ (.A(_00036_),
    .Y(_15391_));
 OA211x2_ASAP7_75t_R _21187_ (.A1(_14804_),
    .A2(_14805_),
    .B(_15391_),
    .C(_14807_),
    .Y(_15392_));
 AO31x2_ASAP7_75t_R _21188_ (.A1(_14737_),
    .A2(_15365_),
    .A3(_15390_),
    .B(_15392_),
    .Y(_15393_));
 INVx1_ASAP7_75t_R _21189_ (.A(_01512_),
    .Y(_15394_));
 AO32x1_ASAP7_75t_R _21190_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_15393_),
    .B1(_15337_),
    .B2(_15394_),
    .Y(_15395_));
 BUFx6f_ASAP7_75t_R _21191_ (.A(_15395_),
    .Y(_18653_));
 INVx1_ASAP7_75t_R _21192_ (.A(_18653_),
    .Y(_18655_));
 OR2x2_ASAP7_75t_R _21193_ (.A(net1981),
    .B(_02298_),
    .Y(_15396_));
 AO21x1_ASAP7_75t_R _21194_ (.A1(_00806_),
    .A2(_15244_),
    .B(_15396_),
    .Y(_15397_));
 OA21x2_ASAP7_75t_R _21195_ (.A1(_00808_),
    .A2(_02298_),
    .B(_00811_),
    .Y(_15398_));
 OA21x2_ASAP7_75t_R _21196_ (.A1(_15243_),
    .A2(_15397_),
    .B(_15398_),
    .Y(_15399_));
 OA21x2_ASAP7_75t_R _21197_ (.A1(_00810_),
    .A2(_15399_),
    .B(_00814_),
    .Y(_15400_));
 XOR2x2_ASAP7_75t_R _21198_ (.A(_00813_),
    .B(_15400_),
    .Y(\alu_adder_result_ex[9] ));
 OR2x2_ASAP7_75t_R _21199_ (.A(_15254_),
    .B(_15396_),
    .Y(_15401_));
 OA21x2_ASAP7_75t_R _21200_ (.A1(net1991),
    .A2(_15257_),
    .B(_00797_),
    .Y(_15402_));
 OR3x4_ASAP7_75t_R _21201_ (.A(net1992),
    .B(_00796_),
    .C(_15263_),
    .Y(_15403_));
 OA211x2_ASAP7_75t_R _21202_ (.A1(_00796_),
    .A2(_15402_),
    .B(_15403_),
    .C(_00800_),
    .Y(_15404_));
 OA21x2_ASAP7_75t_R _21203_ (.A1(_15255_),
    .A2(_15396_),
    .B(_15398_),
    .Y(_15405_));
 OA21x2_ASAP7_75t_R _21204_ (.A1(_15401_),
    .A2(_15404_),
    .B(_15405_),
    .Y(_15406_));
 INVx1_ASAP7_75t_R _21205_ (.A(_15406_),
    .Y(_15407_));
 OA21x2_ASAP7_75t_R _21206_ (.A1(_00796_),
    .A2(_15402_),
    .B(_00800_),
    .Y(_15408_));
 OR2x2_ASAP7_75t_R _21207_ (.A(_15254_),
    .B(_15408_),
    .Y(_15409_));
 NAND3x1_ASAP7_75t_R _21208_ (.A(_14925_),
    .B(_15405_),
    .C(_15409_),
    .Y(_15410_));
 OR3x1_ASAP7_75t_R _21209_ (.A(net1973),
    .B(_15262_),
    .C(_15410_),
    .Y(_15411_));
 OR4x1_ASAP7_75t_R _21210_ (.A(_15248_),
    .B(_15250_),
    .C(_15252_),
    .D(_15410_),
    .Y(_15412_));
 INVx1_ASAP7_75t_R _21211_ (.A(net1980),
    .Y(_15413_));
 AO31x2_ASAP7_75t_R _21212_ (.A1(_15407_),
    .A2(_15411_),
    .A3(_15412_),
    .B(_15413_),
    .Y(_15414_));
 AND3x1_ASAP7_75t_R _21213_ (.A(_14925_),
    .B(_15405_),
    .C(_15409_),
    .Y(_15415_));
 AO211x2_ASAP7_75t_R _21214_ (.A1(net2003),
    .A2(_15415_),
    .B(_15406_),
    .C(net1980),
    .Y(_15416_));
 NAND2x2_ASAP7_75t_R _21215_ (.A(_15414_),
    .B(_15416_),
    .Y(_15417_));
 INVx2_ASAP7_75t_R _21216_ (.A(_15417_),
    .Y(\alu_adder_result_ex[8] ));
 AND2x2_ASAP7_75t_R _21217_ (.A(_14945_),
    .B(_01813_),
    .Y(_15418_));
 AO21x1_ASAP7_75t_R _21218_ (.A1(_14742_),
    .A2(_00724_),
    .B(_15418_),
    .Y(_15419_));
 OAI22x1_ASAP7_75t_R _21219_ (.A1(_00723_),
    .A2(_14741_),
    .B1(_15419_),
    .B2(_14746_),
    .Y(_15420_));
 NAND2x1_ASAP7_75t_R _21220_ (.A(_13711_),
    .B(_00730_),
    .Y(_15421_));
 OA211x2_ASAP7_75t_R _21221_ (.A1(_14831_),
    .A2(_14613_),
    .B(_15421_),
    .C(_15282_),
    .Y(_15422_));
 BUFx6f_ASAP7_75t_R _21222_ (.A(_13754_),
    .Y(_15423_));
 BUFx12_ASAP7_75t_R _21223_ (.A(_13720_),
    .Y(_15424_));
 NAND2x1_ASAP7_75t_R _21224_ (.A(_15424_),
    .B(_00729_),
    .Y(_15425_));
 OA211x2_ASAP7_75t_R _21225_ (.A1(_15423_),
    .A2(_14616_),
    .B(_15425_),
    .C(_14754_),
    .Y(_15426_));
 OR3x1_ASAP7_75t_R _21226_ (.A(_14748_),
    .B(_15422_),
    .C(_15426_),
    .Y(_15427_));
 OA211x2_ASAP7_75t_R _21227_ (.A1(_14740_),
    .A2(_15420_),
    .B(_15427_),
    .C(_14863_),
    .Y(_15428_));
 NAND2x1_ASAP7_75t_R _21228_ (.A(_13872_),
    .B(_00726_),
    .Y(_15429_));
 OA211x2_ASAP7_75t_R _21229_ (.A1(_13871_),
    .A2(_14606_),
    .B(_15429_),
    .C(_13932_),
    .Y(_15430_));
 NAND2x1_ASAP7_75t_R _21230_ (.A(_15067_),
    .B(_00725_),
    .Y(_15431_));
 OA211x2_ASAP7_75t_R _21231_ (.A1(_13934_),
    .A2(_14609_),
    .B(_15431_),
    .C(_13937_),
    .Y(_15432_));
 OR3x1_ASAP7_75t_R _21232_ (.A(_14760_),
    .B(_15430_),
    .C(_15432_),
    .Y(_15433_));
 NAND2x1_ASAP7_75t_R _21233_ (.A(_15067_),
    .B(_00734_),
    .Y(_15434_));
 OA211x2_ASAP7_75t_R _21234_ (.A1(_13930_),
    .A2(_14645_),
    .B(_15434_),
    .C(_15305_),
    .Y(_15435_));
 NAND2x1_ASAP7_75t_R _21235_ (.A(_13935_),
    .B(_00733_),
    .Y(_15436_));
 OA211x2_ASAP7_75t_R _21236_ (.A1(_13934_),
    .A2(_14649_),
    .B(_15436_),
    .C(_15309_),
    .Y(_15437_));
 OR3x1_ASAP7_75t_R _21237_ (.A(_14768_),
    .B(_15435_),
    .C(_15437_),
    .Y(_15438_));
 AND3x1_ASAP7_75t_R _21238_ (.A(_15289_),
    .B(_15433_),
    .C(_15438_),
    .Y(_15439_));
 OR3x4_ASAP7_75t_R _21239_ (.A(_14814_),
    .B(_15428_),
    .C(_15439_),
    .Y(_15440_));
 NAND2x1_ASAP7_75t_R _21240_ (.A(_13872_),
    .B(_00742_),
    .Y(_15441_));
 OA211x2_ASAP7_75t_R _21241_ (.A1(_13871_),
    .A2(_14621_),
    .B(_15441_),
    .C(_13932_),
    .Y(_15442_));
 NAND2x1_ASAP7_75t_R _21242_ (.A(_15067_),
    .B(_00741_),
    .Y(_15443_));
 OA211x2_ASAP7_75t_R _21243_ (.A1(_13930_),
    .A2(_14624_),
    .B(_15443_),
    .C(_13937_),
    .Y(_15444_));
 OR3x1_ASAP7_75t_R _21244_ (.A(_14760_),
    .B(_15442_),
    .C(_15444_),
    .Y(_15445_));
 NAND2x1_ASAP7_75t_R _21245_ (.A(_15067_),
    .B(_00750_),
    .Y(_15446_));
 OA211x2_ASAP7_75t_R _21246_ (.A1(_13930_),
    .A2(_14640_),
    .B(_15446_),
    .C(_15305_),
    .Y(_15447_));
 NAND2x1_ASAP7_75t_R _21247_ (.A(_13935_),
    .B(_00749_),
    .Y(_15448_));
 OA211x2_ASAP7_75t_R _21248_ (.A1(_13934_),
    .A2(_14637_),
    .B(_15448_),
    .C(_13937_),
    .Y(_15449_));
 OR3x1_ASAP7_75t_R _21249_ (.A(_14768_),
    .B(_15447_),
    .C(_15449_),
    .Y(_15450_));
 AND3x1_ASAP7_75t_R _21250_ (.A(_15289_),
    .B(_15445_),
    .C(_15450_),
    .Y(_15451_));
 NAND2x1_ASAP7_75t_R _21251_ (.A(_13935_),
    .B(_00738_),
    .Y(_15452_));
 OA211x2_ASAP7_75t_R _21252_ (.A1(_13934_),
    .A2(_14658_),
    .B(_15452_),
    .C(_15305_),
    .Y(_15453_));
 NAND2x1_ASAP7_75t_R _21253_ (.A(_14816_),
    .B(_00737_),
    .Y(_15454_));
 OA211x2_ASAP7_75t_R _21254_ (.A1(_15307_),
    .A2(_14661_),
    .B(_15454_),
    .C(_15309_),
    .Y(_15455_));
 OR3x1_ASAP7_75t_R _21255_ (.A(_14760_),
    .B(_15453_),
    .C(_15455_),
    .Y(_15456_));
 NAND2x1_ASAP7_75t_R _21256_ (.A(_13935_),
    .B(_00746_),
    .Y(_15457_));
 OA211x2_ASAP7_75t_R _21257_ (.A1(_13934_),
    .A2(_14628_),
    .B(_15457_),
    .C(_15305_),
    .Y(_15458_));
 NAND2x1_ASAP7_75t_R _21258_ (.A(_14816_),
    .B(_00745_),
    .Y(_15459_));
 OA211x2_ASAP7_75t_R _21259_ (.A1(_15290_),
    .A2(_14631_),
    .B(_15459_),
    .C(_15309_),
    .Y(_15460_));
 OR3x1_ASAP7_75t_R _21260_ (.A(_15125_),
    .B(_15458_),
    .C(_15460_),
    .Y(_15461_));
 AND3x1_ASAP7_75t_R _21261_ (.A(_14791_),
    .B(_15456_),
    .C(_15461_),
    .Y(_15462_));
 OR3x4_ASAP7_75t_R _21262_ (.A(_14842_),
    .B(_15451_),
    .C(_15462_),
    .Y(_15463_));
 INVx1_ASAP7_75t_R _21263_ (.A(_00039_),
    .Y(_15464_));
 OA211x2_ASAP7_75t_R _21264_ (.A1(_14804_),
    .A2(_14805_),
    .B(_15464_),
    .C(_15334_),
    .Y(_15465_));
 AO31x2_ASAP7_75t_R _21265_ (.A1(_13947_),
    .A2(_15440_),
    .A3(_15463_),
    .B(_15465_),
    .Y(_15466_));
 INVx1_ASAP7_75t_R _21266_ (.A(_01542_),
    .Y(_15467_));
 AO32x1_ASAP7_75t_R _21267_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_15466_),
    .B1(_15337_),
    .B2(_15467_),
    .Y(_15468_));
 BUFx6f_ASAP7_75t_R _21268_ (.A(_15468_),
    .Y(_18657_));
 INVx2_ASAP7_75t_R _21269_ (.A(_18657_),
    .Y(_18659_));
 BUFx3_ASAP7_75t_R _21270_ (.A(_00819_),
    .Y(_15469_));
 BUFx3_ASAP7_75t_R _21271_ (.A(_00816_),
    .Y(_15470_));
 OR4x2_ASAP7_75t_R _21272_ (.A(_00805_),
    .B(_00810_),
    .C(_00813_),
    .D(_02298_),
    .Y(_15471_));
 AO21x1_ASAP7_75t_R _21273_ (.A1(_00806_),
    .A2(_15244_),
    .B(_15471_),
    .Y(_15472_));
 OR2x2_ASAP7_75t_R _21274_ (.A(net1979),
    .B(net1989),
    .Y(_15473_));
 OR2x2_ASAP7_75t_R _21275_ (.A(_00814_),
    .B(net1989),
    .Y(_15474_));
 OA211x2_ASAP7_75t_R _21276_ (.A1(_15398_),
    .A2(_15473_),
    .B(_15474_),
    .C(_00817_),
    .Y(_15475_));
 OA21x2_ASAP7_75t_R _21277_ (.A1(_15243_),
    .A2(_15472_),
    .B(_15475_),
    .Y(_15476_));
 OA21x2_ASAP7_75t_R _21278_ (.A1(_15470_),
    .A2(_15476_),
    .B(_00820_),
    .Y(_15477_));
 XOR2x2_ASAP7_75t_R _21279_ (.A(_15469_),
    .B(_15477_),
    .Y(\alu_adder_result_ex[11] ));
 OA21x2_ASAP7_75t_R _21280_ (.A1(_15398_),
    .A2(_15473_),
    .B(_15474_),
    .Y(_15478_));
 NAND2x1_ASAP7_75t_R _21281_ (.A(_00817_),
    .B(_15478_),
    .Y(_15479_));
 INVx1_ASAP7_75t_R _21282_ (.A(_15470_),
    .Y(_15480_));
 AND3x1_ASAP7_75t_R _21283_ (.A(_15480_),
    .B(_15471_),
    .C(_15475_),
    .Y(_15481_));
 AND3x1_ASAP7_75t_R _21284_ (.A(_15480_),
    .B(_15266_),
    .C(_15475_),
    .Y(_15482_));
 AOI211x1_ASAP7_75t_R _21285_ (.A1(_15470_),
    .A2(_15479_),
    .B(_15481_),
    .C(_15482_),
    .Y(_15483_));
 AND3x2_ASAP7_75t_R _21286_ (.A(_14925_),
    .B(_15256_),
    .C(_15257_),
    .Y(_15484_));
 AND4x2_ASAP7_75t_R _21287_ (.A(_14898_),
    .B(_14909_),
    .C(_14914_),
    .D(_15484_),
    .Y(_15485_));
 AND3x1_ASAP7_75t_R _21288_ (.A(_14920_),
    .B(_14919_),
    .C(_15484_),
    .Y(_15486_));
 AND2x2_ASAP7_75t_R _21289_ (.A(_15480_),
    .B(_15475_),
    .Y(_15487_));
 OAI21x1_ASAP7_75t_R _21290_ (.A1(_15485_),
    .A2(_15486_),
    .B(_15487_),
    .Y(_15488_));
 OR5x2_ASAP7_75t_R _21291_ (.A(_15480_),
    .B(_15266_),
    .C(_15485_),
    .D(_15486_),
    .E(_15471_),
    .Y(_15489_));
 NAND3x2_ASAP7_75t_R _21292_ (.B(_15488_),
    .C(_15489_),
    .Y(\alu_adder_result_ex[10] ),
    .A(_15483_));
 BUFx3_ASAP7_75t_R _21293_ (.A(_14373_),
    .Y(_15490_));
 BUFx3_ASAP7_75t_R _21294_ (.A(_15490_),
    .Y(_15491_));
 AND3x1_ASAP7_75t_R _21295_ (.A(_13406_),
    .B(_13412_),
    .C(_14150_),
    .Y(_15492_));
 OA21x2_ASAP7_75t_R _21296_ (.A1(_13436_),
    .A2(_15492_),
    .B(_13435_),
    .Y(_15493_));
 AND2x4_ASAP7_75t_R _21297_ (.A(_14058_),
    .B(_13443_),
    .Y(_15494_));
 AO21x1_ASAP7_75t_R _21298_ (.A1(_13572_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_15495_));
 BUFx4f_ASAP7_75t_R _21299_ (.A(_13788_),
    .Y(_15496_));
 BUFx4f_ASAP7_75t_R _21300_ (.A(_13447_),
    .Y(_15497_));
 BUFx6f_ASAP7_75t_R _21301_ (.A(_13454_),
    .Y(_15498_));
 BUFx6f_ASAP7_75t_R _21302_ (.A(_15498_),
    .Y(_15499_));
 BUFx16f_ASAP7_75t_R _21303_ (.A(_13497_),
    .Y(_15500_));
 BUFx3_ASAP7_75t_R clone2 (.A(_01552_),
    .Y(net2));
 BUFx6f_ASAP7_75t_R _21305_ (.A(_13390_),
    .Y(_15502_));
 BUFx12f_ASAP7_75t_R _21306_ (.A(_13458_),
    .Y(_15503_));
 BUFx6f_ASAP7_75t_R _21307_ (.A(_15503_),
    .Y(_15504_));
 BUFx6f_ASAP7_75t_R _21308_ (.A(_15504_),
    .Y(_15505_));
 AND2x2_ASAP7_75t_R _21309_ (.A(_15505_),
    .B(_01811_),
    .Y(_15506_));
 AO21x1_ASAP7_75t_R _21310_ (.A1(_15502_),
    .A2(_00450_),
    .B(_15506_),
    .Y(_15507_));
 BUFx3_ASAP7_75t_R clone8 (.A(_09647_),
    .Y(net8));
 BUFx4f_ASAP7_75t_R _21312_ (.A(_13479_),
    .Y(_15509_));
 BUFx12_ASAP7_75t_R _21313_ (.A(_15509_),
    .Y(_15510_));
 OAI22x1_ASAP7_75t_R _21314_ (.A1(_00449_),
    .A2(_15500_),
    .B1(_15507_),
    .B2(_15510_),
    .Y(_15511_));
 BUFx6f_ASAP7_75t_R _21315_ (.A(_13484_),
    .Y(_15512_));
 BUFx6f_ASAP7_75t_R _21316_ (.A(net5),
    .Y(_15513_));
 INVx1_ASAP7_75t_R _21317_ (.A(_00458_),
    .Y(_15514_));
 BUFx12f_ASAP7_75t_R _21318_ (.A(_13458_),
    .Y(_15515_));
 BUFx10_ASAP7_75t_R _21319_ (.A(_15515_),
    .Y(_15516_));
 NAND2x1_ASAP7_75t_R _21320_ (.A(_15516_),
    .B(_00456_),
    .Y(_15517_));
 BUFx12f_ASAP7_75t_R _21321_ (.A(_13470_),
    .Y(_15518_));
 BUFx6f_ASAP7_75t_R _21322_ (.A(net10),
    .Y(_15519_));
 OA211x2_ASAP7_75t_R _21323_ (.A1(_15513_),
    .A2(_15514_),
    .B(_15517_),
    .C(_15519_),
    .Y(_15520_));
 INVx1_ASAP7_75t_R _21324_ (.A(_00457_),
    .Y(_15521_));
 NAND2x1_ASAP7_75t_R _21325_ (.A(_15516_),
    .B(_00455_),
    .Y(_15522_));
 BUFx4f_ASAP7_75t_R _21326_ (.A(_13479_),
    .Y(_15523_));
 OA211x2_ASAP7_75t_R _21327_ (.A1(_15513_),
    .A2(_15521_),
    .B(_15522_),
    .C(_15523_),
    .Y(_15524_));
 OR3x1_ASAP7_75t_R _21328_ (.A(_15512_),
    .B(_15520_),
    .C(_15524_),
    .Y(_15525_));
 BUFx4f_ASAP7_75t_R _21329_ (.A(_13512_),
    .Y(_15526_));
 OA211x2_ASAP7_75t_R _21330_ (.A1(_15499_),
    .A2(_15511_),
    .B(_15525_),
    .C(_15526_),
    .Y(_15527_));
 BUFx6f_ASAP7_75t_R _21331_ (.A(_13451_),
    .Y(_15528_));
 BUFx10_ASAP7_75t_R _21332_ (.A(_15528_),
    .Y(_15529_));
 BUFx6f_ASAP7_75t_R _21333_ (.A(_13454_),
    .Y(_15530_));
 BUFx6f_ASAP7_75t_R _21334_ (.A(_15530_),
    .Y(_15531_));
 BUFx10_ASAP7_75t_R _21335_ (.A(_15503_),
    .Y(_15532_));
 BUFx6f_ASAP7_75t_R _21336_ (.A(_15532_),
    .Y(_15533_));
 BUFx6f_ASAP7_75t_R _21337_ (.A(_13458_),
    .Y(_15534_));
 BUFx10_ASAP7_75t_R _21338_ (.A(_15534_),
    .Y(_15535_));
 NAND2x1_ASAP7_75t_R _21339_ (.A(_15535_),
    .B(_00452_),
    .Y(_15536_));
 BUFx6f_ASAP7_75t_R _21340_ (.A(_15518_),
    .Y(_15537_));
 BUFx6f_ASAP7_75t_R _21341_ (.A(_15537_),
    .Y(_15538_));
 OA211x2_ASAP7_75t_R _21342_ (.A1(_15533_),
    .A2(_13963_),
    .B(_15536_),
    .C(_15538_),
    .Y(_15539_));
 BUFx4f_ASAP7_75t_R _21343_ (.A(_15532_),
    .Y(_15540_));
 BUFx6f_ASAP7_75t_R _21344_ (.A(_13458_),
    .Y(_15541_));
 BUFx6f_ASAP7_75t_R _21345_ (.A(_15541_),
    .Y(_15542_));
 NAND2x1_ASAP7_75t_R _21346_ (.A(_15542_),
    .B(_00451_),
    .Y(_15543_));
 BUFx4f_ASAP7_75t_R _21347_ (.A(_13479_),
    .Y(_15544_));
 OA211x2_ASAP7_75t_R _21348_ (.A1(_15540_),
    .A2(_13967_),
    .B(_15543_),
    .C(_15544_),
    .Y(_15545_));
 OR3x1_ASAP7_75t_R _21349_ (.A(_15531_),
    .B(_15539_),
    .C(_15545_),
    .Y(_15546_));
 BUFx6f_ASAP7_75t_R _21350_ (.A(_13484_),
    .Y(_15547_));
 NAND2x1_ASAP7_75t_R _21351_ (.A(_15535_),
    .B(_00460_),
    .Y(_15548_));
 OA211x2_ASAP7_75t_R _21352_ (.A1(_15533_),
    .A2(_13982_),
    .B(_15548_),
    .C(_15538_),
    .Y(_15549_));
 NAND2x1_ASAP7_75t_R _21353_ (.A(_15542_),
    .B(_00459_),
    .Y(_15550_));
 OA211x2_ASAP7_75t_R _21354_ (.A1(_15540_),
    .A2(_13985_),
    .B(_15550_),
    .C(_15544_),
    .Y(_15551_));
 OR3x1_ASAP7_75t_R _21355_ (.A(_15547_),
    .B(_15549_),
    .C(_15551_),
    .Y(_15552_));
 AND3x1_ASAP7_75t_R _21356_ (.A(_15529_),
    .B(_15546_),
    .C(_15552_),
    .Y(_15553_));
 OR3x4_ASAP7_75t_R _21357_ (.A(_15497_),
    .B(_15527_),
    .C(_15553_),
    .Y(_15554_));
 BUFx10_ASAP7_75t_R _21358_ (.A(_13518_),
    .Y(_15555_));
 NAND2x1_ASAP7_75t_R _21359_ (.A(_15535_),
    .B(_00468_),
    .Y(_15556_));
 OA211x2_ASAP7_75t_R _21360_ (.A1(_15533_),
    .A2(_13971_),
    .B(_15556_),
    .C(_15538_),
    .Y(_15557_));
 NAND2x1_ASAP7_75t_R _21361_ (.A(_15542_),
    .B(_00467_),
    .Y(_15558_));
 OA211x2_ASAP7_75t_R _21362_ (.A1(_15533_),
    .A2(_13974_),
    .B(_15558_),
    .C(_15544_),
    .Y(_15559_));
 OR3x1_ASAP7_75t_R _21363_ (.A(_15531_),
    .B(_15557_),
    .C(_15559_),
    .Y(_15560_));
 NAND2x1_ASAP7_75t_R _21364_ (.A(_15535_),
    .B(_00476_),
    .Y(_15561_));
 OA211x2_ASAP7_75t_R _21365_ (.A1(_15533_),
    .A2(_13989_),
    .B(_15561_),
    .C(_15538_),
    .Y(_15562_));
 NAND2x1_ASAP7_75t_R _21366_ (.A(_15542_),
    .B(_00475_),
    .Y(_15563_));
 OA211x2_ASAP7_75t_R _21367_ (.A1(_15540_),
    .A2(_13992_),
    .B(_15563_),
    .C(_15544_),
    .Y(_15564_));
 OR3x1_ASAP7_75t_R _21368_ (.A(_15547_),
    .B(_15562_),
    .C(_15564_),
    .Y(_15565_));
 AND3x1_ASAP7_75t_R _21369_ (.A(_15529_),
    .B(_15560_),
    .C(_15565_),
    .Y(_15566_));
 BUFx6f_ASAP7_75t_R _21370_ (.A(_13484_),
    .Y(_15567_));
 BUFx6f_ASAP7_75t_R _21371_ (.A(_15567_),
    .Y(_15568_));
 BUFx6f_ASAP7_75t_R _21372_ (.A(_15509_),
    .Y(_15569_));
 BUFx6f_ASAP7_75t_R _21373_ (.A(_15534_),
    .Y(_15570_));
 BUFx4f_ASAP7_75t_R _21374_ (.A(_15570_),
    .Y(_15571_));
 BUFx10_ASAP7_75t_R _21375_ (.A(_15503_),
    .Y(_15572_));
 BUFx4f_ASAP7_75t_R _21376_ (.A(_15572_),
    .Y(_15573_));
 NOR2x1_ASAP7_75t_R _21377_ (.A(_15573_),
    .B(_00473_),
    .Y(_15574_));
 AO21x1_ASAP7_75t_R _21378_ (.A1(_15571_),
    .A2(_13997_),
    .B(_15574_),
    .Y(_15575_));
 BUFx6f_ASAP7_75t_R _21379_ (.A(_15503_),
    .Y(_15576_));
 BUFx6f_ASAP7_75t_R _21380_ (.A(_15576_),
    .Y(_15577_));
 INVx1_ASAP7_75t_R _21381_ (.A(_00474_),
    .Y(_15578_));
 BUFx6f_ASAP7_75t_R _21382_ (.A(_15534_),
    .Y(_15579_));
 NAND2x1_ASAP7_75t_R _21383_ (.A(_15579_),
    .B(_00472_),
    .Y(_15580_));
 BUFx4f_ASAP7_75t_R _21384_ (.A(_15537_),
    .Y(_15581_));
 OA211x2_ASAP7_75t_R _21385_ (.A1(_15577_),
    .A2(_15578_),
    .B(_15580_),
    .C(_15581_),
    .Y(_15582_));
 AO21x1_ASAP7_75t_R _21386_ (.A1(_15569_),
    .A2(_15575_),
    .B(_15582_),
    .Y(_15583_));
 NAND2x1_ASAP7_75t_R _21387_ (.A(_15516_),
    .B(_00464_),
    .Y(_15584_));
 OA211x2_ASAP7_75t_R _21388_ (.A1(_15513_),
    .A2(_13953_),
    .B(_15584_),
    .C(_15519_),
    .Y(_15585_));
 BUFx16f_ASAP7_75t_R _21389_ (.A(_15503_),
    .Y(_15586_));
 BUFx6f_ASAP7_75t_R _21390_ (.A(_15586_),
    .Y(_15587_));
 NAND2x1_ASAP7_75t_R _21391_ (.A(_15516_),
    .B(_00463_),
    .Y(_15588_));
 OA211x2_ASAP7_75t_R _21392_ (.A1(_15587_),
    .A2(_13957_),
    .B(_15588_),
    .C(_15523_),
    .Y(_15589_));
 OR3x1_ASAP7_75t_R _21393_ (.A(_15498_),
    .B(_15585_),
    .C(_15589_),
    .Y(_15590_));
 OA211x2_ASAP7_75t_R _21394_ (.A1(_15568_),
    .A2(_15583_),
    .B(_15590_),
    .C(_15526_),
    .Y(_15591_));
 OR3x4_ASAP7_75t_R _21395_ (.A(_15555_),
    .B(_15566_),
    .C(_15591_),
    .Y(_15592_));
 AND3x1_ASAP7_75t_R _21396_ (.A(_15496_),
    .B(_15554_),
    .C(_15592_),
    .Y(_15593_));
 AO21x2_ASAP7_75t_R _21397_ (.A1(_15491_),
    .A2(_15495_),
    .B(_15593_),
    .Y(_18668_));
 BUFx6f_ASAP7_75t_R _21398_ (.A(_15504_),
    .Y(_15594_));
 AND2x2_ASAP7_75t_R _21399_ (.A(_15594_),
    .B(_01810_),
    .Y(_15595_));
 AO21x1_ASAP7_75t_R _21400_ (.A1(_15502_),
    .A2(_00825_),
    .B(_15595_),
    .Y(_15596_));
 OAI22x1_ASAP7_75t_R _21401_ (.A1(_00824_),
    .A2(_15500_),
    .B1(_15596_),
    .B2(_15569_),
    .Y(_15597_));
 INVx1_ASAP7_75t_R _21402_ (.A(_00833_),
    .Y(_15598_));
 NAND2x1_ASAP7_75t_R _21403_ (.A(_15516_),
    .B(_00831_),
    .Y(_15599_));
 OA211x2_ASAP7_75t_R _21404_ (.A1(_15513_),
    .A2(_15598_),
    .B(_15599_),
    .C(_15519_),
    .Y(_15600_));
 INVx2_ASAP7_75t_R _21405_ (.A(_00832_),
    .Y(_15601_));
 BUFx12f_ASAP7_75t_R _21406_ (.A(_15515_),
    .Y(_15602_));
 NAND2x1_ASAP7_75t_R _21407_ (.A(_15602_),
    .B(_00830_),
    .Y(_15603_));
 OA211x2_ASAP7_75t_R _21408_ (.A1(_15587_),
    .A2(_15601_),
    .B(_15603_),
    .C(_15523_),
    .Y(_15604_));
 OR3x1_ASAP7_75t_R _21409_ (.A(_15512_),
    .B(_15600_),
    .C(_15604_),
    .Y(_15605_));
 OA211x2_ASAP7_75t_R _21410_ (.A1(_15499_),
    .A2(_15597_),
    .B(_15605_),
    .C(_15526_),
    .Y(_15606_));
 BUFx6f_ASAP7_75t_R _21411_ (.A(_13451_),
    .Y(_15607_));
 BUFx6f_ASAP7_75t_R _21412_ (.A(_13454_),
    .Y(_15608_));
 BUFx12f_ASAP7_75t_R _21413_ (.A(_15515_),
    .Y(_15609_));
 BUFx4f_ASAP7_75t_R _21414_ (.A(_15609_),
    .Y(_15610_));
 INVx1_ASAP7_75t_R _21415_ (.A(_00829_),
    .Y(_15611_));
 BUFx6f_ASAP7_75t_R _21416_ (.A(_15534_),
    .Y(_15612_));
 NAND2x1_ASAP7_75t_R _21417_ (.A(_15612_),
    .B(_00827_),
    .Y(_15613_));
 BUFx3_ASAP7_75t_R _21418_ (.A(_15537_),
    .Y(_15614_));
 OA211x2_ASAP7_75t_R _21419_ (.A1(_15610_),
    .A2(_15611_),
    .B(_15613_),
    .C(net145),
    .Y(_15615_));
 INVx1_ASAP7_75t_R _21420_ (.A(_00828_),
    .Y(_15616_));
 BUFx6f_ASAP7_75t_R _21421_ (.A(_15534_),
    .Y(_15617_));
 NAND2x1_ASAP7_75t_R _21422_ (.A(_15617_),
    .B(_00826_),
    .Y(_15618_));
 BUFx3_ASAP7_75t_R _21423_ (.A(_13479_),
    .Y(_15619_));
 OA211x2_ASAP7_75t_R _21424_ (.A1(_15610_),
    .A2(_15616_),
    .B(_15618_),
    .C(_15619_),
    .Y(_15620_));
 OR3x1_ASAP7_75t_R _21425_ (.A(_15608_),
    .B(_15615_),
    .C(_15620_),
    .Y(_15621_));
 INVx2_ASAP7_75t_R _21426_ (.A(_00837_),
    .Y(_15622_));
 NAND2x1_ASAP7_75t_R _21427_ (.A(_15617_),
    .B(_00835_),
    .Y(_15623_));
 OA211x2_ASAP7_75t_R _21428_ (.A1(_15610_),
    .A2(_15622_),
    .B(_15623_),
    .C(net145),
    .Y(_15624_));
 BUFx6f_ASAP7_75t_R _21429_ (.A(_15572_),
    .Y(_15625_));
 INVx2_ASAP7_75t_R _21430_ (.A(_00836_),
    .Y(_15626_));
 BUFx6f_ASAP7_75t_R _21431_ (.A(_15515_),
    .Y(_15627_));
 NAND2x1_ASAP7_75t_R _21432_ (.A(_15627_),
    .B(_00834_),
    .Y(_15628_));
 OA211x2_ASAP7_75t_R _21433_ (.A1(_15625_),
    .A2(_15626_),
    .B(_15628_),
    .C(_15619_),
    .Y(_15629_));
 OR3x1_ASAP7_75t_R _21434_ (.A(_15547_),
    .B(_15624_),
    .C(_15629_),
    .Y(_15630_));
 AND3x1_ASAP7_75t_R _21435_ (.A(_15607_),
    .B(_15621_),
    .C(_15630_),
    .Y(_15631_));
 OR3x4_ASAP7_75t_R _21436_ (.A(_15497_),
    .B(_15606_),
    .C(_15631_),
    .Y(_15632_));
 INVx2_ASAP7_75t_R _21437_ (.A(_00845_),
    .Y(_15633_));
 NAND2x1_ASAP7_75t_R _21438_ (.A(_15612_),
    .B(_00843_),
    .Y(_15634_));
 OA211x2_ASAP7_75t_R _21439_ (.A1(_15540_),
    .A2(_15633_),
    .B(_15634_),
    .C(net145),
    .Y(_15635_));
 INVx2_ASAP7_75t_R _21440_ (.A(_00844_),
    .Y(_15636_));
 NAND2x1_ASAP7_75t_R _21441_ (.A(_15617_),
    .B(_00842_),
    .Y(_15637_));
 OA211x2_ASAP7_75t_R _21442_ (.A1(_15610_),
    .A2(_15636_),
    .B(_15637_),
    .C(_15544_),
    .Y(_15638_));
 OR3x1_ASAP7_75t_R _21443_ (.A(_15608_),
    .B(_15635_),
    .C(_15638_),
    .Y(_15639_));
 INVx2_ASAP7_75t_R _21444_ (.A(_00853_),
    .Y(_15640_));
 NAND2x1_ASAP7_75t_R _21445_ (.A(_15612_),
    .B(_00851_),
    .Y(_15641_));
 OA211x2_ASAP7_75t_R _21446_ (.A1(_15610_),
    .A2(_15640_),
    .B(_15641_),
    .C(net145),
    .Y(_15642_));
 INVx2_ASAP7_75t_R _21447_ (.A(_00852_),
    .Y(_15643_));
 NAND2x1_ASAP7_75t_R _21448_ (.A(_15617_),
    .B(_00850_),
    .Y(_15644_));
 OA211x2_ASAP7_75t_R _21449_ (.A1(_15610_),
    .A2(_15643_),
    .B(_15644_),
    .C(_15619_),
    .Y(_15645_));
 OR3x1_ASAP7_75t_R _21450_ (.A(_15547_),
    .B(_15642_),
    .C(_15645_),
    .Y(_15646_));
 AND3x1_ASAP7_75t_R _21451_ (.A(_15607_),
    .B(_15639_),
    .C(_15646_),
    .Y(_15647_));
 BUFx6f_ASAP7_75t_R _21452_ (.A(_13479_),
    .Y(_15648_));
 BUFx6f_ASAP7_75t_R _21453_ (.A(_15648_),
    .Y(_15649_));
 INVx1_ASAP7_75t_R _21454_ (.A(_00846_),
    .Y(_15650_));
 BUFx6f_ASAP7_75t_R _21455_ (.A(net15),
    .Y(_15651_));
 BUFx6f_ASAP7_75t_R _21456_ (.A(_15651_),
    .Y(_15652_));
 NOR2x1_ASAP7_75t_R _21457_ (.A(_15652_),
    .B(_00848_),
    .Y(_15653_));
 AO21x1_ASAP7_75t_R _21458_ (.A1(_15571_),
    .A2(_15650_),
    .B(_15653_),
    .Y(_15654_));
 INVx1_ASAP7_75t_R _21459_ (.A(_00849_),
    .Y(_15655_));
 BUFx6f_ASAP7_75t_R _21460_ (.A(_15534_),
    .Y(_15656_));
 NAND2x1_ASAP7_75t_R _21461_ (.A(_15656_),
    .B(_00847_),
    .Y(_15657_));
 OA211x2_ASAP7_75t_R _21462_ (.A1(_15577_),
    .A2(_15655_),
    .B(_15657_),
    .C(_15538_),
    .Y(_15658_));
 AO21x1_ASAP7_75t_R _21463_ (.A1(_15649_),
    .A2(_15654_),
    .B(_15658_),
    .Y(_15659_));
 INVx1_ASAP7_75t_R _21464_ (.A(_00841_),
    .Y(_15660_));
 NAND2x1_ASAP7_75t_R _21465_ (.A(_15602_),
    .B(_00839_),
    .Y(_15661_));
 OA211x2_ASAP7_75t_R _21466_ (.A1(_15587_),
    .A2(_15660_),
    .B(_15661_),
    .C(_15519_),
    .Y(_15662_));
 BUFx3_ASAP7_75t_R clone7 (.A(_09647_),
    .Y(net7));
 INVx2_ASAP7_75t_R _21468_ (.A(_00840_),
    .Y(_15664_));
 BUFx6f_ASAP7_75t_R _21469_ (.A(_15515_),
    .Y(_15665_));
 NAND2x1_ASAP7_75t_R _21470_ (.A(_15665_),
    .B(_00838_),
    .Y(_15666_));
 OA211x2_ASAP7_75t_R _21471_ (.A1(net5),
    .A2(_15664_),
    .B(_15666_),
    .C(_15523_),
    .Y(_15667_));
 OR3x1_ASAP7_75t_R _21472_ (.A(_15498_),
    .B(_15662_),
    .C(_15667_),
    .Y(_15668_));
 OA211x2_ASAP7_75t_R _21473_ (.A1(_15568_),
    .A2(_15659_),
    .B(_15668_),
    .C(_15526_),
    .Y(_15669_));
 OR3x2_ASAP7_75t_R _21474_ (.A(_15555_),
    .B(_15647_),
    .C(_15669_),
    .Y(_15670_));
 AND2x2_ASAP7_75t_R _21475_ (.A(_15632_),
    .B(_15670_),
    .Y(_15671_));
 AO21x1_ASAP7_75t_R _21476_ (.A1(_13563_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_15672_));
 AND2x2_ASAP7_75t_R _21477_ (.A(_15491_),
    .B(_15672_),
    .Y(_15673_));
 AO21x2_ASAP7_75t_R _21478_ (.A1(_15496_),
    .A2(_15671_),
    .B(_15673_),
    .Y(_18673_));
 AND2x2_ASAP7_75t_R _21479_ (.A(_15290_),
    .B(_01810_),
    .Y(_15674_));
 AO21x1_ASAP7_75t_R _21480_ (.A1(_13777_),
    .A2(_00825_),
    .B(_15674_),
    .Y(_15675_));
 OAI22x1_ASAP7_75t_R _21481_ (.A1(_00824_),
    .A2(_13858_),
    .B1(_15675_),
    .B2(_14990_),
    .Y(_15676_));
 BUFx6f_ASAP7_75t_R _21482_ (.A(_14858_),
    .Y(_15677_));
 NAND2x1_ASAP7_75t_R _21483_ (.A(_14820_),
    .B(_00831_),
    .Y(_15678_));
 OA211x2_ASAP7_75t_R _21484_ (.A1(_15677_),
    .A2(_15598_),
    .B(_15678_),
    .C(_14995_),
    .Y(_15679_));
 NAND2x1_ASAP7_75t_R _21485_ (.A(_14993_),
    .B(_00830_),
    .Y(_15680_));
 BUFx6f_ASAP7_75t_R _21486_ (.A(_13714_),
    .Y(_15681_));
 OA211x2_ASAP7_75t_R _21487_ (.A1(_14992_),
    .A2(_15601_),
    .B(_15680_),
    .C(_15681_),
    .Y(_15682_));
 OR3x2_ASAP7_75t_R _21488_ (.A(_13902_),
    .B(_15679_),
    .C(_15682_),
    .Y(_15683_));
 OA211x2_ASAP7_75t_R _21489_ (.A1(_14986_),
    .A2(_15676_),
    .B(_15683_),
    .C(_14791_),
    .Y(_15684_));
 NAND2x1_ASAP7_75t_R _21490_ (.A(_14854_),
    .B(_00827_),
    .Y(_15685_));
 BUFx4f_ASAP7_75t_R _21491_ (.A(_13761_),
    .Y(_15686_));
 OA211x2_ASAP7_75t_R _21492_ (.A1(_15319_),
    .A2(_15611_),
    .B(_15685_),
    .C(_15686_),
    .Y(_15687_));
 NAND2x1_ASAP7_75t_R _21493_ (.A(_14857_),
    .B(_00826_),
    .Y(_15688_));
 BUFx4f_ASAP7_75t_R _21494_ (.A(_13728_),
    .Y(_15689_));
 OA211x2_ASAP7_75t_R _21495_ (.A1(_13924_),
    .A2(_15616_),
    .B(_15688_),
    .C(_15689_),
    .Y(_15690_));
 OR3x1_ASAP7_75t_R _21496_ (.A(_13707_),
    .B(_15687_),
    .C(_15690_),
    .Y(_15691_));
 NAND2x1_ASAP7_75t_R _21497_ (.A(_14848_),
    .B(_00835_),
    .Y(_15692_));
 OA211x2_ASAP7_75t_R _21498_ (.A1(_15207_),
    .A2(_15622_),
    .B(_15692_),
    .C(_15004_),
    .Y(_15693_));
 NAND2x1_ASAP7_75t_R _21499_ (.A(_13925_),
    .B(_00834_),
    .Y(_15694_));
 OA211x2_ASAP7_75t_R _21500_ (.A1(_15013_),
    .A2(_15626_),
    .B(_15694_),
    .C(_15689_),
    .Y(_15695_));
 OR3x1_ASAP7_75t_R _21501_ (.A(_15031_),
    .B(_15693_),
    .C(_15695_),
    .Y(_15696_));
 AND3x2_ASAP7_75t_R _21502_ (.A(_15002_),
    .B(_15691_),
    .C(_15696_),
    .Y(_15697_));
 OR3x4_ASAP7_75t_R _21503_ (.A(_14733_),
    .B(_15684_),
    .C(_15697_),
    .Y(_15698_));
 NAND2x1_ASAP7_75t_R _21504_ (.A(_14844_),
    .B(_00843_),
    .Y(_15699_));
 OA211x2_ASAP7_75t_R _21505_ (.A1(_15319_),
    .A2(_15633_),
    .B(_15699_),
    .C(_15686_),
    .Y(_15700_));
 NAND2x1_ASAP7_75t_R _21506_ (.A(_14854_),
    .B(_00842_),
    .Y(_15701_));
 OA211x2_ASAP7_75t_R _21507_ (.A1(_15207_),
    .A2(_15636_),
    .B(_15701_),
    .C(_15689_),
    .Y(_15702_));
 OR3x1_ASAP7_75t_R _21508_ (.A(_13707_),
    .B(_15700_),
    .C(_15702_),
    .Y(_15703_));
 NAND2x1_ASAP7_75t_R _21509_ (.A(_14844_),
    .B(_00851_),
    .Y(_15704_));
 OA211x2_ASAP7_75t_R _21510_ (.A1(_15319_),
    .A2(_15640_),
    .B(_15704_),
    .C(_15686_),
    .Y(_15705_));
 NAND2x1_ASAP7_75t_R _21511_ (.A(_14848_),
    .B(_00850_),
    .Y(_15706_));
 OA211x2_ASAP7_75t_R _21512_ (.A1(_15207_),
    .A2(_15643_),
    .B(_15706_),
    .C(_15689_),
    .Y(_15707_));
 OR3x1_ASAP7_75t_R _21513_ (.A(_15031_),
    .B(_15705_),
    .C(_15707_),
    .Y(_15708_));
 AND3x1_ASAP7_75t_R _21514_ (.A(_15002_),
    .B(_15703_),
    .C(_15708_),
    .Y(_15709_));
 NOR2x1_ASAP7_75t_R _21515_ (.A(_15143_),
    .B(_00848_),
    .Y(_15710_));
 AO21x1_ASAP7_75t_R _21516_ (.A1(_14011_),
    .A2(_15650_),
    .B(_15710_),
    .Y(_15711_));
 BUFx6f_ASAP7_75t_R _21517_ (.A(_13886_),
    .Y(_15712_));
 NAND2x1_ASAP7_75t_R _21518_ (.A(_14831_),
    .B(_00847_),
    .Y(_15713_));
 OA211x2_ASAP7_75t_R _21519_ (.A1(_15712_),
    .A2(_15655_),
    .B(_15713_),
    .C(_15686_),
    .Y(_15714_));
 AO21x1_ASAP7_75t_R _21520_ (.A1(_14746_),
    .A2(_15711_),
    .B(_15714_),
    .Y(_15715_));
 NAND2x1_ASAP7_75t_R _21521_ (.A(_14993_),
    .B(_00839_),
    .Y(_15716_));
 OA211x2_ASAP7_75t_R _21522_ (.A1(_14992_),
    .A2(_15660_),
    .B(_15716_),
    .C(_14780_),
    .Y(_15717_));
 BUFx6f_ASAP7_75t_R _21523_ (.A(_13690_),
    .Y(_15718_));
 NAND2x1_ASAP7_75t_R _21524_ (.A(_15190_),
    .B(_00838_),
    .Y(_15719_));
 OA211x2_ASAP7_75t_R _21525_ (.A1(_15718_),
    .A2(_15664_),
    .B(_15719_),
    .C(_13715_),
    .Y(_15720_));
 OR3x1_ASAP7_75t_R _21526_ (.A(_14777_),
    .B(_15717_),
    .C(_15720_),
    .Y(_15721_));
 OA211x2_ASAP7_75t_R _21527_ (.A1(_13903_),
    .A2(_15715_),
    .B(_15721_),
    .C(_14791_),
    .Y(_15722_));
 OR3x4_ASAP7_75t_R _21528_ (.A(_15025_),
    .B(_15709_),
    .C(_15722_),
    .Y(_15723_));
 INVx1_ASAP7_75t_R _21529_ (.A(_00046_),
    .Y(_15724_));
 OA211x2_ASAP7_75t_R _21530_ (.A1(_15114_),
    .A2(_15115_),
    .B(_15724_),
    .C(_14807_),
    .Y(_15725_));
 AO31x2_ASAP7_75t_R _21531_ (.A1(_13660_),
    .A2(_15698_),
    .A3(_15723_),
    .B(_15725_),
    .Y(_15726_));
 INVx1_ASAP7_75t_R _21532_ (.A(_01539_),
    .Y(_15727_));
 AO32x1_ASAP7_75t_R _21533_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_15726_),
    .B1(_15119_),
    .B2(_15727_),
    .Y(_15728_));
 BUFx6f_ASAP7_75t_R _21534_ (.A(_15728_),
    .Y(_18672_));
 INVx1_ASAP7_75t_R _21535_ (.A(_18672_),
    .Y(_18674_));
 OA21x2_ASAP7_75t_R _21536_ (.A1(_00820_),
    .A2(_15469_),
    .B(_00823_),
    .Y(_15729_));
 OR3x1_ASAP7_75t_R _21537_ (.A(_15470_),
    .B(_15469_),
    .C(_15476_),
    .Y(_15730_));
 AO21x1_ASAP7_75t_R _21538_ (.A1(_15729_),
    .A2(_15730_),
    .B(_00822_),
    .Y(_15731_));
 AND2x2_ASAP7_75t_R _21539_ (.A(_00856_),
    .B(_15731_),
    .Y(_15732_));
 XNOR2x2_ASAP7_75t_R _21540_ (.A(net1988),
    .B(_15732_),
    .Y(_15733_));
 CKINVDCx6p67_ASAP7_75t_R _21541_ (.A(_15733_),
    .Y(\alu_adder_result_ex[13] ));
 INVx1_ASAP7_75t_R _21542_ (.A(net1978),
    .Y(_15734_));
 OR4x1_ASAP7_75t_R _21543_ (.A(_15470_),
    .B(_15469_),
    .C(_15406_),
    .D(_15473_),
    .Y(_15735_));
 OR2x2_ASAP7_75t_R _21544_ (.A(_15734_),
    .B(_15735_),
    .Y(_15736_));
 AO21x2_ASAP7_75t_R _21545_ (.A1(net2003),
    .A2(_15415_),
    .B(_15736_),
    .Y(_15737_));
 OA21x2_ASAP7_75t_R _21546_ (.A1(_00814_),
    .A2(net1989),
    .B(_00817_),
    .Y(_15738_));
 OA21x2_ASAP7_75t_R _21547_ (.A1(_15470_),
    .A2(_15738_),
    .B(_00820_),
    .Y(_15739_));
 OA21x2_ASAP7_75t_R _21548_ (.A1(_15469_),
    .A2(_15739_),
    .B(_00823_),
    .Y(_15740_));
 AND2x2_ASAP7_75t_R _21549_ (.A(_15734_),
    .B(_15740_),
    .Y(_15741_));
 AND2x2_ASAP7_75t_R _21550_ (.A(_15415_),
    .B(_15741_),
    .Y(_15742_));
 NOR2x1_ASAP7_75t_R _21551_ (.A(_15734_),
    .B(_15740_),
    .Y(_15743_));
 AOI221x1_ASAP7_75t_R _21552_ (.A1(_15735_),
    .A2(_15741_),
    .B1(_15742_),
    .B2(net2003),
    .C(_15743_),
    .Y(_15744_));
 NAND2x2_ASAP7_75t_R _21553_ (.A(_15737_),
    .B(_15744_),
    .Y(\alu_adder_result_ex[12] ));
 BUFx12_ASAP7_75t_R _21554_ (.A(_13447_),
    .Y(_15745_));
 BUFx4f_ASAP7_75t_R _21555_ (.A(_13512_),
    .Y(_15746_));
 BUFx6f_ASAP7_75t_R _21556_ (.A(_15746_),
    .Y(_15747_));
 BUFx10_ASAP7_75t_R _21557_ (.A(_15503_),
    .Y(_15748_));
 BUFx4f_ASAP7_75t_R _21558_ (.A(_15748_),
    .Y(_15749_));
 AND2x2_ASAP7_75t_R _21559_ (.A(_15749_),
    .B(_01809_),
    .Y(_15750_));
 AO21x1_ASAP7_75t_R _21560_ (.A1(_15502_),
    .A2(_00858_),
    .B(_15750_),
    .Y(_15751_));
 OAI22x1_ASAP7_75t_R _21561_ (.A1(_00857_),
    .A2(_15500_),
    .B1(_15751_),
    .B2(_15510_),
    .Y(_15752_));
 BUFx6f_ASAP7_75t_R _21562_ (.A(_13484_),
    .Y(_15753_));
 BUFx2_ASAP7_75t_R clone6 (.A(_09579_),
    .Y(net6));
 INVx1_ASAP7_75t_R _21564_ (.A(_00866_),
    .Y(_15755_));
 BUFx6f_ASAP7_75t_R _21565_ (.A(_15541_),
    .Y(_15756_));
 NAND2x1_ASAP7_75t_R _21566_ (.A(_15756_),
    .B(_00864_),
    .Y(_15757_));
 BUFx3_ASAP7_75t_R _21567_ (.A(net18),
    .Y(_15758_));
 OA211x2_ASAP7_75t_R _21568_ (.A1(_15602_),
    .A2(_15755_),
    .B(_15757_),
    .C(net19),
    .Y(_15759_));
 INVx1_ASAP7_75t_R _21569_ (.A(_00865_),
    .Y(_15760_));
 NAND2x1_ASAP7_75t_R _21570_ (.A(_15756_),
    .B(_00863_),
    .Y(_15761_));
 OA211x2_ASAP7_75t_R _21571_ (.A1(_15602_),
    .A2(_15760_),
    .B(_15761_),
    .C(_15509_),
    .Y(_15762_));
 OR3x1_ASAP7_75t_R _21572_ (.A(_15753_),
    .B(_15759_),
    .C(_15762_),
    .Y(_15763_));
 OA21x2_ASAP7_75t_R _21573_ (.A1(_15499_),
    .A2(_15752_),
    .B(_15763_),
    .Y(_15764_));
 BUFx6f_ASAP7_75t_R _21574_ (.A(_15576_),
    .Y(_15765_));
 INVx1_ASAP7_75t_R _21575_ (.A(_00862_),
    .Y(_15766_));
 BUFx6f_ASAP7_75t_R _21576_ (.A(_15534_),
    .Y(_15767_));
 NAND2x1_ASAP7_75t_R _21577_ (.A(_15767_),
    .B(_00860_),
    .Y(_15768_));
 OA211x2_ASAP7_75t_R _21578_ (.A1(_15765_),
    .A2(_15766_),
    .B(_15768_),
    .C(_15581_),
    .Y(_15769_));
 INVx1_ASAP7_75t_R _21579_ (.A(_00861_),
    .Y(_15770_));
 NAND2x1_ASAP7_75t_R _21580_ (.A(_15579_),
    .B(_00859_),
    .Y(_15771_));
 OA211x2_ASAP7_75t_R _21581_ (.A1(_15765_),
    .A2(_15770_),
    .B(_15771_),
    .C(_15648_),
    .Y(_15772_));
 OR3x1_ASAP7_75t_R _21582_ (.A(_15531_),
    .B(_15769_),
    .C(_15772_),
    .Y(_15773_));
 INVx1_ASAP7_75t_R _21583_ (.A(_00870_),
    .Y(_15774_));
 NAND2x1_ASAP7_75t_R _21584_ (.A(_15767_),
    .B(_00868_),
    .Y(_15775_));
 OA211x2_ASAP7_75t_R _21585_ (.A1(_15765_),
    .A2(_15774_),
    .B(_15775_),
    .C(_15581_),
    .Y(_15776_));
 INVx1_ASAP7_75t_R _21586_ (.A(_00869_),
    .Y(_15777_));
 NAND2x1_ASAP7_75t_R _21587_ (.A(_15579_),
    .B(_00867_),
    .Y(_15778_));
 OA211x2_ASAP7_75t_R _21588_ (.A1(_15577_),
    .A2(_15777_),
    .B(_15778_),
    .C(_15648_),
    .Y(_15779_));
 OR3x1_ASAP7_75t_R _21589_ (.A(_15753_),
    .B(_15776_),
    .C(_15779_),
    .Y(_15780_));
 AND3x1_ASAP7_75t_R _21590_ (.A(_15529_),
    .B(_15773_),
    .C(_15780_),
    .Y(_15781_));
 AO21x1_ASAP7_75t_R _21591_ (.A1(_15747_),
    .A2(_15764_),
    .B(_15781_),
    .Y(_15782_));
 INVx2_ASAP7_75t_R _21592_ (.A(_00878_),
    .Y(_15783_));
 NAND2x1_ASAP7_75t_R _21593_ (.A(_15617_),
    .B(_00876_),
    .Y(_15784_));
 OA211x2_ASAP7_75t_R _21594_ (.A1(_15610_),
    .A2(_15783_),
    .B(_15784_),
    .C(_15614_),
    .Y(_15785_));
 INVx2_ASAP7_75t_R _21595_ (.A(_00877_),
    .Y(_15786_));
 NAND2x1_ASAP7_75t_R _21596_ (.A(_15627_),
    .B(_00875_),
    .Y(_15787_));
 OA211x2_ASAP7_75t_R _21597_ (.A1(_15625_),
    .A2(_15786_),
    .B(_15787_),
    .C(_15619_),
    .Y(_15788_));
 OR3x1_ASAP7_75t_R _21598_ (.A(_15608_),
    .B(_15785_),
    .C(_15788_),
    .Y(_15789_));
 INVx1_ASAP7_75t_R _21599_ (.A(_00886_),
    .Y(_15790_));
 NAND2x1_ASAP7_75t_R _21600_ (.A(_15627_),
    .B(_00884_),
    .Y(_15791_));
 OA211x2_ASAP7_75t_R _21601_ (.A1(_15625_),
    .A2(_15790_),
    .B(_15791_),
    .C(_15614_),
    .Y(_15792_));
 INVx2_ASAP7_75t_R _21602_ (.A(_00885_),
    .Y(_15793_));
 NAND2x1_ASAP7_75t_R _21603_ (.A(_15627_),
    .B(_00883_),
    .Y(_15794_));
 OA211x2_ASAP7_75t_R _21604_ (.A1(_15625_),
    .A2(_15793_),
    .B(_15794_),
    .C(_15619_),
    .Y(_15795_));
 OR3x1_ASAP7_75t_R _21605_ (.A(_15547_),
    .B(_15792_),
    .C(_15795_),
    .Y(_15796_));
 AND3x1_ASAP7_75t_R _21606_ (.A(_15607_),
    .B(_15789_),
    .C(_15796_),
    .Y(_15797_));
 INVx1_ASAP7_75t_R _21607_ (.A(_00879_),
    .Y(_15798_));
 NOR2x1_ASAP7_75t_R _21608_ (.A(_15513_),
    .B(_00881_),
    .Y(_15799_));
 AO21x1_ASAP7_75t_R _21609_ (.A1(_15571_),
    .A2(_15798_),
    .B(_15799_),
    .Y(_15800_));
 INVx1_ASAP7_75t_R _21610_ (.A(_00882_),
    .Y(_15801_));
 NAND2x1_ASAP7_75t_R _21611_ (.A(_15535_),
    .B(_00880_),
    .Y(_15802_));
 OA211x2_ASAP7_75t_R _21612_ (.A1(_15533_),
    .A2(_15801_),
    .B(_15802_),
    .C(_15538_),
    .Y(_15803_));
 AO21x1_ASAP7_75t_R _21613_ (.A1(_15649_),
    .A2(_15800_),
    .B(_15803_),
    .Y(_15804_));
 INVx1_ASAP7_75t_R _21614_ (.A(_00874_),
    .Y(_15805_));
 NAND2x1_ASAP7_75t_R _21615_ (.A(_15665_),
    .B(_00872_),
    .Y(_15806_));
 BUFx4f_ASAP7_75t_R _21616_ (.A(_15518_),
    .Y(_15807_));
 OA211x2_ASAP7_75t_R _21617_ (.A1(net5),
    .A2(_15805_),
    .B(_15806_),
    .C(_15807_),
    .Y(_15808_));
 INVx1_ASAP7_75t_R _21618_ (.A(_00873_),
    .Y(_15809_));
 NAND2x1_ASAP7_75t_R _21619_ (.A(_15665_),
    .B(_00871_),
    .Y(_15810_));
 BUFx6f_ASAP7_75t_R _21620_ (.A(_13479_),
    .Y(_15811_));
 OA211x2_ASAP7_75t_R _21621_ (.A1(net5),
    .A2(_15809_),
    .B(_15810_),
    .C(_15811_),
    .Y(_15812_));
 OR3x1_ASAP7_75t_R _21622_ (.A(_15498_),
    .B(_15808_),
    .C(_15812_),
    .Y(_15813_));
 OA211x2_ASAP7_75t_R _21623_ (.A1(_15568_),
    .A2(_15804_),
    .B(_15813_),
    .C(_15526_),
    .Y(_15814_));
 OR3x1_ASAP7_75t_R _21624_ (.A(_15555_),
    .B(_15797_),
    .C(_15814_),
    .Y(_15815_));
 OA21x2_ASAP7_75t_R _21625_ (.A1(_15745_),
    .A2(_15782_),
    .B(_15815_),
    .Y(_15816_));
 AO21x1_ASAP7_75t_R _21626_ (.A1(_13567_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_15817_));
 AND2x2_ASAP7_75t_R _21627_ (.A(_15491_),
    .B(_15817_),
    .Y(_15818_));
 AO21x2_ASAP7_75t_R _21628_ (.A1(_15496_),
    .A2(_15816_),
    .B(_15818_),
    .Y(_18679_));
 AND2x2_ASAP7_75t_R _21629_ (.A(_15290_),
    .B(_01809_),
    .Y(_15819_));
 AO21x1_ASAP7_75t_R _21630_ (.A1(_13777_),
    .A2(_00858_),
    .B(_15819_),
    .Y(_15820_));
 OAI22x1_ASAP7_75t_R _21631_ (.A1(_00857_),
    .A2(_13858_),
    .B1(_15820_),
    .B2(_14990_),
    .Y(_15821_));
 NAND2x1_ASAP7_75t_R _21632_ (.A(_14820_),
    .B(_00864_),
    .Y(_15822_));
 OA211x2_ASAP7_75t_R _21633_ (.A1(_15677_),
    .A2(_15755_),
    .B(_15822_),
    .C(_14995_),
    .Y(_15823_));
 NAND2x1_ASAP7_75t_R _21634_ (.A(_14993_),
    .B(_00863_),
    .Y(_15824_));
 OA211x2_ASAP7_75t_R _21635_ (.A1(_15677_),
    .A2(_15760_),
    .B(_15824_),
    .C(_15681_),
    .Y(_15825_));
 OR3x2_ASAP7_75t_R _21636_ (.A(_15079_),
    .B(_15823_),
    .C(_15825_),
    .Y(_15826_));
 OA211x2_ASAP7_75t_R _21637_ (.A1(_13857_),
    .A2(_15821_),
    .B(_15826_),
    .C(_14791_),
    .Y(_15827_));
 NAND2x1_ASAP7_75t_R _21638_ (.A(_14844_),
    .B(_00860_),
    .Y(_15828_));
 OA211x2_ASAP7_75t_R _21639_ (.A1(_15319_),
    .A2(_15766_),
    .B(_15828_),
    .C(_15686_),
    .Y(_15829_));
 NAND2x1_ASAP7_75t_R _21640_ (.A(_14848_),
    .B(_00859_),
    .Y(_15830_));
 OA211x2_ASAP7_75t_R _21641_ (.A1(_15207_),
    .A2(_15770_),
    .B(_15830_),
    .C(_15689_),
    .Y(_15831_));
 OR3x1_ASAP7_75t_R _21642_ (.A(_13707_),
    .B(_15829_),
    .C(_15831_),
    .Y(_15832_));
 NAND2x1_ASAP7_75t_R _21643_ (.A(_14854_),
    .B(_00868_),
    .Y(_15833_));
 OA211x2_ASAP7_75t_R _21644_ (.A1(_15319_),
    .A2(_15774_),
    .B(_15833_),
    .C(_15004_),
    .Y(_15834_));
 NAND2x1_ASAP7_75t_R _21645_ (.A(_14857_),
    .B(_00867_),
    .Y(_15835_));
 OA211x2_ASAP7_75t_R _21646_ (.A1(_13924_),
    .A2(_15777_),
    .B(_15835_),
    .C(_15689_),
    .Y(_15836_));
 OR3x1_ASAP7_75t_R _21647_ (.A(_15031_),
    .B(_15834_),
    .C(_15836_),
    .Y(_15837_));
 AND3x2_ASAP7_75t_R _21648_ (.A(_15002_),
    .B(_15832_),
    .C(_15837_),
    .Y(_15838_));
 OR3x4_ASAP7_75t_R _21649_ (.A(_14733_),
    .B(_15827_),
    .C(_15838_),
    .Y(_15839_));
 NAND2x1_ASAP7_75t_R _21650_ (.A(_14844_),
    .B(_00876_),
    .Y(_15840_));
 OA211x2_ASAP7_75t_R _21651_ (.A1(_15712_),
    .A2(_15783_),
    .B(_15840_),
    .C(_15686_),
    .Y(_15841_));
 NAND2x1_ASAP7_75t_R _21652_ (.A(_14854_),
    .B(_00875_),
    .Y(_15842_));
 OA211x2_ASAP7_75t_R _21653_ (.A1(_15319_),
    .A2(_15786_),
    .B(_15842_),
    .C(_15689_),
    .Y(_15843_));
 OR3x1_ASAP7_75t_R _21654_ (.A(_13707_),
    .B(_15841_),
    .C(_15843_),
    .Y(_15844_));
 NAND2x1_ASAP7_75t_R _21655_ (.A(_14844_),
    .B(_00884_),
    .Y(_15845_));
 OA211x2_ASAP7_75t_R _21656_ (.A1(_15319_),
    .A2(_15790_),
    .B(_15845_),
    .C(_15686_),
    .Y(_15846_));
 NAND2x1_ASAP7_75t_R _21657_ (.A(_14854_),
    .B(_00883_),
    .Y(_15847_));
 OA211x2_ASAP7_75t_R _21658_ (.A1(_15207_),
    .A2(_15793_),
    .B(_15847_),
    .C(_15689_),
    .Y(_15848_));
 OR3x1_ASAP7_75t_R _21659_ (.A(_15031_),
    .B(_15846_),
    .C(_15848_),
    .Y(_15849_));
 AND3x1_ASAP7_75t_R _21660_ (.A(_15002_),
    .B(_15844_),
    .C(_15849_),
    .Y(_15850_));
 NOR2x1_ASAP7_75t_R _21661_ (.A(_15143_),
    .B(_00881_),
    .Y(_15851_));
 AO21x1_ASAP7_75t_R _21662_ (.A1(_14011_),
    .A2(_15798_),
    .B(_15851_),
    .Y(_15852_));
 NAND2x1_ASAP7_75t_R _21663_ (.A(_14831_),
    .B(_00880_),
    .Y(_15853_));
 BUFx4f_ASAP7_75t_R _21664_ (.A(_13761_),
    .Y(_15854_));
 OA211x2_ASAP7_75t_R _21665_ (.A1(_15712_),
    .A2(_15801_),
    .B(_15853_),
    .C(_15854_),
    .Y(_15855_));
 AO21x1_ASAP7_75t_R _21666_ (.A1(_14746_),
    .A2(_15852_),
    .B(_15855_),
    .Y(_15856_));
 NAND2x1_ASAP7_75t_R _21667_ (.A(_14993_),
    .B(_00872_),
    .Y(_15857_));
 OA211x2_ASAP7_75t_R _21668_ (.A1(_14992_),
    .A2(_15805_),
    .B(_15857_),
    .C(_14995_),
    .Y(_15858_));
 NAND2x1_ASAP7_75t_R _21669_ (.A(_13751_),
    .B(_00871_),
    .Y(_15859_));
 OA211x2_ASAP7_75t_R _21670_ (.A1(_13921_),
    .A2(_15809_),
    .B(_15859_),
    .C(_13715_),
    .Y(_15860_));
 OR3x2_ASAP7_75t_R _21671_ (.A(_14777_),
    .B(_15858_),
    .C(_15860_),
    .Y(_15861_));
 OA211x2_ASAP7_75t_R _21672_ (.A1(_13903_),
    .A2(_15856_),
    .B(_15861_),
    .C(_14791_),
    .Y(_15862_));
 OR3x4_ASAP7_75t_R _21673_ (.A(_15025_),
    .B(_15850_),
    .C(_15862_),
    .Y(_15863_));
 INVx1_ASAP7_75t_R _21674_ (.A(_00048_),
    .Y(_15864_));
 OA211x2_ASAP7_75t_R _21675_ (.A1(_15114_),
    .A2(_15115_),
    .B(_15864_),
    .C(_13367_),
    .Y(_15865_));
 AO31x2_ASAP7_75t_R _21676_ (.A1(_13660_),
    .A2(_15839_),
    .A3(_15863_),
    .B(_15865_),
    .Y(_15866_));
 INVx1_ASAP7_75t_R _21677_ (.A(_01538_),
    .Y(_15867_));
 AO32x1_ASAP7_75t_R _21678_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_15866_),
    .B1(_15119_),
    .B2(_15867_),
    .Y(_15868_));
 BUFx6f_ASAP7_75t_R _21679_ (.A(_15868_),
    .Y(_18680_));
 INVx1_ASAP7_75t_R _21680_ (.A(_18680_),
    .Y(_18678_));
 BUFx6f_ASAP7_75t_R _21681_ (.A(_13454_),
    .Y(_15869_));
 BUFx4f_ASAP7_75t_R _21682_ (.A(_15869_),
    .Y(_15870_));
 BUFx4f_ASAP7_75t_R _21683_ (.A(_13390_),
    .Y(_15871_));
 BUFx6f_ASAP7_75t_R _21684_ (.A(_15515_),
    .Y(_15872_));
 AND2x2_ASAP7_75t_R _21685_ (.A(_15872_),
    .B(_01808_),
    .Y(_15873_));
 AO21x1_ASAP7_75t_R _21686_ (.A1(_15871_),
    .A2(_00891_),
    .B(_15873_),
    .Y(_15874_));
 OAI22x1_ASAP7_75t_R _21687_ (.A1(_00890_),
    .A2(_15500_),
    .B1(_15874_),
    .B2(_15649_),
    .Y(_15875_));
 BUFx6f_ASAP7_75t_R _21688_ (.A(_13484_),
    .Y(_15876_));
 INVx1_ASAP7_75t_R _21689_ (.A(_00899_),
    .Y(_15877_));
 NAND2x1_ASAP7_75t_R _21690_ (.A(_15572_),
    .B(_00897_),
    .Y(_15878_));
 BUFx4f_ASAP7_75t_R _21691_ (.A(net10),
    .Y(_15879_));
 OA211x2_ASAP7_75t_R _21692_ (.A1(_15612_),
    .A2(_15877_),
    .B(_15878_),
    .C(_15879_),
    .Y(_15880_));
 INVx1_ASAP7_75t_R _21693_ (.A(_00898_),
    .Y(_15881_));
 NAND2x1_ASAP7_75t_R _21694_ (.A(_15586_),
    .B(_00896_),
    .Y(_15882_));
 BUFx4f_ASAP7_75t_R _21695_ (.A(_13479_),
    .Y(_15883_));
 OA211x2_ASAP7_75t_R _21696_ (.A1(_15617_),
    .A2(_15881_),
    .B(_15882_),
    .C(_15883_),
    .Y(_15884_));
 OR3x1_ASAP7_75t_R _21697_ (.A(_15876_),
    .B(_15880_),
    .C(_15884_),
    .Y(_15885_));
 OA211x2_ASAP7_75t_R _21698_ (.A1(_15870_),
    .A2(_15875_),
    .B(_15885_),
    .C(_15746_),
    .Y(_15886_));
 BUFx6f_ASAP7_75t_R _21699_ (.A(_13451_),
    .Y(_15887_));
 BUFx4f_ASAP7_75t_R _21700_ (.A(_13454_),
    .Y(_15888_));
 BUFx6f_ASAP7_75t_R _21701_ (.A(_15504_),
    .Y(_15889_));
 INVx1_ASAP7_75t_R _21702_ (.A(_00895_),
    .Y(_15890_));
 BUFx12f_ASAP7_75t_R _21703_ (.A(_15515_),
    .Y(_15891_));
 NAND2x1_ASAP7_75t_R _21704_ (.A(_15891_),
    .B(_00893_),
    .Y(_15892_));
 BUFx6f_ASAP7_75t_R _21705_ (.A(_15518_),
    .Y(_15893_));
 OA211x2_ASAP7_75t_R _21706_ (.A1(_15889_),
    .A2(_15890_),
    .B(_15892_),
    .C(_15893_),
    .Y(_15894_));
 BUFx6f_ASAP7_75t_R _21707_ (.A(_15504_),
    .Y(_15895_));
 INVx1_ASAP7_75t_R _21708_ (.A(_00894_),
    .Y(_15896_));
 BUFx6f_ASAP7_75t_R _21709_ (.A(net15),
    .Y(_15897_));
 NAND2x1_ASAP7_75t_R _21710_ (.A(_15897_),
    .B(_00892_),
    .Y(_15898_));
 BUFx3_ASAP7_75t_R _21711_ (.A(_13479_),
    .Y(_15899_));
 OA211x2_ASAP7_75t_R _21712_ (.A1(_15895_),
    .A2(_15896_),
    .B(_15898_),
    .C(_15899_),
    .Y(_15900_));
 OR3x1_ASAP7_75t_R _21713_ (.A(_15888_),
    .B(_15894_),
    .C(_15900_),
    .Y(_15901_));
 BUFx6f_ASAP7_75t_R _21714_ (.A(_13484_),
    .Y(_15902_));
 INVx1_ASAP7_75t_R _21715_ (.A(_00903_),
    .Y(_15903_));
 NAND2x1_ASAP7_75t_R _21716_ (.A(_15609_),
    .B(_00901_),
    .Y(_15904_));
 OA211x2_ASAP7_75t_R _21717_ (.A1(_15895_),
    .A2(_15903_),
    .B(_15904_),
    .C(_15893_),
    .Y(_15905_));
 INVx1_ASAP7_75t_R _21718_ (.A(_00902_),
    .Y(_15906_));
 NAND2x1_ASAP7_75t_R _21719_ (.A(_15897_),
    .B(_00900_),
    .Y(_15907_));
 OA211x2_ASAP7_75t_R _21720_ (.A1(_15756_),
    .A2(_15906_),
    .B(_15907_),
    .C(_15899_),
    .Y(_15908_));
 OR3x1_ASAP7_75t_R _21721_ (.A(_15902_),
    .B(_15905_),
    .C(_15908_),
    .Y(_15909_));
 AND3x2_ASAP7_75t_R _21722_ (.A(_15887_),
    .B(_15901_),
    .C(_15909_),
    .Y(_15910_));
 OR3x4_ASAP7_75t_R _21723_ (.A(_15497_),
    .B(_15886_),
    .C(_15910_),
    .Y(_15911_));
 BUFx4f_ASAP7_75t_R _21724_ (.A(_13518_),
    .Y(_15912_));
 INVx1_ASAP7_75t_R _21725_ (.A(_00911_),
    .Y(_15913_));
 NAND2x1_ASAP7_75t_R _21726_ (.A(_15891_),
    .B(_00909_),
    .Y(_15914_));
 OA211x2_ASAP7_75t_R _21727_ (.A1(_15889_),
    .A2(_15913_),
    .B(_15914_),
    .C(_15893_),
    .Y(_15915_));
 INVx1_ASAP7_75t_R _21728_ (.A(_00910_),
    .Y(_15916_));
 NAND2x1_ASAP7_75t_R _21729_ (.A(_15609_),
    .B(_00908_),
    .Y(_15917_));
 BUFx4f_ASAP7_75t_R _21730_ (.A(_13479_),
    .Y(_15918_));
 OA211x2_ASAP7_75t_R _21731_ (.A1(_15895_),
    .A2(_15916_),
    .B(_15917_),
    .C(_15918_),
    .Y(_15919_));
 OR3x1_ASAP7_75t_R _21732_ (.A(_15888_),
    .B(_15915_),
    .C(_15919_),
    .Y(_15920_));
 INVx1_ASAP7_75t_R _21733_ (.A(_00919_),
    .Y(_15921_));
 NAND2x1_ASAP7_75t_R _21734_ (.A(_15891_),
    .B(_00917_),
    .Y(_15922_));
 OA211x2_ASAP7_75t_R _21735_ (.A1(_15889_),
    .A2(_15921_),
    .B(_15922_),
    .C(_15893_),
    .Y(_15923_));
 INVx1_ASAP7_75t_R _21736_ (.A(_00918_),
    .Y(_15924_));
 NAND2x1_ASAP7_75t_R _21737_ (.A(_15609_),
    .B(_00916_),
    .Y(_15925_));
 OA211x2_ASAP7_75t_R _21738_ (.A1(_15895_),
    .A2(_15924_),
    .B(_15925_),
    .C(_15899_),
    .Y(_15926_));
 OR3x1_ASAP7_75t_R _21739_ (.A(_15902_),
    .B(_15923_),
    .C(_15926_),
    .Y(_15927_));
 AND3x1_ASAP7_75t_R _21740_ (.A(_15887_),
    .B(_15920_),
    .C(_15927_),
    .Y(_15928_));
 BUFx4f_ASAP7_75t_R _21741_ (.A(_15876_),
    .Y(_15929_));
 BUFx4f_ASAP7_75t_R _21742_ (.A(_13479_),
    .Y(_15930_));
 BUFx4f_ASAP7_75t_R _21743_ (.A(_15930_),
    .Y(_15931_));
 INVx2_ASAP7_75t_R _21744_ (.A(_00912_),
    .Y(_15932_));
 NOR2x1_ASAP7_75t_R _21745_ (.A(_15535_),
    .B(_00914_),
    .Y(_15933_));
 AO21x1_ASAP7_75t_R _21746_ (.A1(_15625_),
    .A2(_15932_),
    .B(_15933_),
    .Y(_15934_));
 INVx1_ASAP7_75t_R _21747_ (.A(_00915_),
    .Y(_15935_));
 BUFx12f_ASAP7_75t_R _21748_ (.A(_15515_),
    .Y(_15936_));
 NAND2x1_ASAP7_75t_R _21749_ (.A(_15936_),
    .B(_00913_),
    .Y(_15937_));
 OA211x2_ASAP7_75t_R _21750_ (.A1(_15594_),
    .A2(_15935_),
    .B(_15937_),
    .C(_15807_),
    .Y(_15938_));
 AO21x1_ASAP7_75t_R _21751_ (.A1(_15931_),
    .A2(_15934_),
    .B(_15938_),
    .Y(_15939_));
 INVx1_ASAP7_75t_R _21752_ (.A(_00907_),
    .Y(_15940_));
 NAND2x1_ASAP7_75t_R _21753_ (.A(_15586_),
    .B(_00905_),
    .Y(_15941_));
 OA211x2_ASAP7_75t_R _21754_ (.A1(_15627_),
    .A2(_15940_),
    .B(_15941_),
    .C(_15879_),
    .Y(_15942_));
 INVx2_ASAP7_75t_R _21755_ (.A(_00906_),
    .Y(_15943_));
 NAND2x1_ASAP7_75t_R _21756_ (.A(_15651_),
    .B(_00904_),
    .Y(_15944_));
 BUFx4f_ASAP7_75t_R _21757_ (.A(_13479_),
    .Y(_15945_));
 OA211x2_ASAP7_75t_R _21758_ (.A1(_15627_),
    .A2(_15943_),
    .B(_15944_),
    .C(_15945_),
    .Y(_15946_));
 OR3x1_ASAP7_75t_R _21759_ (.A(_15530_),
    .B(_15942_),
    .C(_15946_),
    .Y(_15947_));
 OA211x2_ASAP7_75t_R _21760_ (.A1(_15929_),
    .A2(_15939_),
    .B(_15947_),
    .C(_15746_),
    .Y(_15948_));
 OR3x2_ASAP7_75t_R _21761_ (.A(_15912_),
    .B(_15928_),
    .C(_15948_),
    .Y(_15949_));
 AND2x4_ASAP7_75t_R _21762_ (.A(_15911_),
    .B(_15949_),
    .Y(_15950_));
 AO21x1_ASAP7_75t_R _21763_ (.A1(_13945_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_15951_));
 AND2x2_ASAP7_75t_R _21764_ (.A(_15491_),
    .B(_15951_),
    .Y(_15952_));
 AO21x2_ASAP7_75t_R _21765_ (.A1(_15496_),
    .A2(_15950_),
    .B(_15952_),
    .Y(_18684_));
 BUFx3_ASAP7_75t_R _21766_ (.A(_13667_),
    .Y(_15953_));
 BUFx6f_ASAP7_75t_R _21767_ (.A(_13756_),
    .Y(_15954_));
 AND2x2_ASAP7_75t_R _21768_ (.A(_15954_),
    .B(_01808_),
    .Y(_15955_));
 AO21x1_ASAP7_75t_R _21769_ (.A1(_13777_),
    .A2(_00891_),
    .B(_15955_),
    .Y(_15956_));
 OAI22x1_ASAP7_75t_R _21770_ (.A1(_00890_),
    .A2(_13858_),
    .B1(_15956_),
    .B2(_14990_),
    .Y(_15957_));
 NAND2x1_ASAP7_75t_R _21771_ (.A(_13882_),
    .B(_00897_),
    .Y(_15958_));
 OA211x2_ASAP7_75t_R _21772_ (.A1(_13881_),
    .A2(_15877_),
    .B(_15958_),
    .C(_13884_),
    .Y(_15959_));
 NAND2x1_ASAP7_75t_R _21773_ (.A(_13888_),
    .B(_00896_),
    .Y(_15960_));
 OA211x2_ASAP7_75t_R _21774_ (.A1(_13887_),
    .A2(_15881_),
    .B(_15960_),
    .C(_13890_),
    .Y(_15961_));
 OR3x2_ASAP7_75t_R _21775_ (.A(_15012_),
    .B(_15959_),
    .C(_15961_),
    .Y(_15962_));
 OA211x2_ASAP7_75t_R _21776_ (.A1(_13857_),
    .A2(_15957_),
    .B(_15962_),
    .C(_15038_),
    .Y(_15963_));
 BUFx4f_ASAP7_75t_R _21777_ (.A(_13751_),
    .Y(_15964_));
 NAND2x1_ASAP7_75t_R _21778_ (.A(_15061_),
    .B(_00893_),
    .Y(_15965_));
 OA211x2_ASAP7_75t_R _21779_ (.A1(_15964_),
    .A2(_15890_),
    .B(_15965_),
    .C(_15854_),
    .Y(_15966_));
 BUFx6f_ASAP7_75t_R _21780_ (.A(_13722_),
    .Y(_15967_));
 NAND2x1_ASAP7_75t_R _21781_ (.A(_15967_),
    .B(_00892_),
    .Y(_15968_));
 BUFx6f_ASAP7_75t_R _21782_ (.A(_13728_),
    .Y(_15969_));
 OA211x2_ASAP7_75t_R _21783_ (.A1(_15964_),
    .A2(_15896_),
    .B(_15968_),
    .C(_15969_),
    .Y(_15970_));
 OR3x1_ASAP7_75t_R _21784_ (.A(_14815_),
    .B(_15966_),
    .C(_15970_),
    .Y(_15971_));
 NAND2x1_ASAP7_75t_R _21785_ (.A(_15967_),
    .B(_00901_),
    .Y(_15972_));
 OA211x2_ASAP7_75t_R _21786_ (.A1(_15964_),
    .A2(_15903_),
    .B(_15972_),
    .C(_15854_),
    .Y(_15973_));
 NAND2x1_ASAP7_75t_R _21787_ (.A(_15967_),
    .B(_00900_),
    .Y(_15974_));
 OA211x2_ASAP7_75t_R _21788_ (.A1(_15964_),
    .A2(_15906_),
    .B(_15974_),
    .C(_15969_),
    .Y(_15975_));
 OR3x1_ASAP7_75t_R _21789_ (.A(_13748_),
    .B(_15973_),
    .C(_15975_),
    .Y(_15976_));
 AND3x2_ASAP7_75t_R _21790_ (.A(_14732_),
    .B(_15971_),
    .C(_15976_),
    .Y(_15977_));
 OR3x4_ASAP7_75t_R _21791_ (.A(_14733_),
    .B(_15963_),
    .C(_15977_),
    .Y(_15978_));
 NAND2x1_ASAP7_75t_R _21792_ (.A(_15061_),
    .B(_00909_),
    .Y(_15979_));
 OA211x2_ASAP7_75t_R _21793_ (.A1(_15964_),
    .A2(_15913_),
    .B(_15979_),
    .C(_15854_),
    .Y(_15980_));
 NAND2x1_ASAP7_75t_R _21794_ (.A(_15967_),
    .B(_00908_),
    .Y(_15981_));
 OA211x2_ASAP7_75t_R _21795_ (.A1(_15964_),
    .A2(_15916_),
    .B(_15981_),
    .C(_15969_),
    .Y(_15982_));
 OR3x1_ASAP7_75t_R _21796_ (.A(_14815_),
    .B(_15980_),
    .C(_15982_),
    .Y(_15983_));
 NAND2x1_ASAP7_75t_R _21797_ (.A(_15967_),
    .B(_00917_),
    .Y(_15984_));
 OA211x2_ASAP7_75t_R _21798_ (.A1(_15964_),
    .A2(_15921_),
    .B(_15984_),
    .C(_15854_),
    .Y(_15985_));
 NAND2x1_ASAP7_75t_R _21799_ (.A(_15967_),
    .B(_00916_),
    .Y(_15986_));
 OA211x2_ASAP7_75t_R _21800_ (.A1(_15964_),
    .A2(_15924_),
    .B(_15986_),
    .C(_15969_),
    .Y(_15987_));
 OR3x1_ASAP7_75t_R _21801_ (.A(_13748_),
    .B(_15985_),
    .C(_15987_),
    .Y(_15988_));
 AND3x2_ASAP7_75t_R _21802_ (.A(_14732_),
    .B(_15983_),
    .C(_15988_),
    .Y(_15989_));
 NOR2x1_ASAP7_75t_R _21803_ (.A(_15042_),
    .B(_00914_),
    .Y(_15990_));
 AO21x1_ASAP7_75t_R _21804_ (.A1(_14011_),
    .A2(_15932_),
    .B(_15990_),
    .Y(_15991_));
 BUFx6f_ASAP7_75t_R _21805_ (.A(_13919_),
    .Y(_15992_));
 NAND2x1_ASAP7_75t_R _21806_ (.A(_13750_),
    .B(_00913_),
    .Y(_15993_));
 OA211x2_ASAP7_75t_R _21807_ (.A1(_15992_),
    .A2(_15935_),
    .B(_15993_),
    .C(_15854_),
    .Y(_15994_));
 AO21x1_ASAP7_75t_R _21808_ (.A1(_13863_),
    .A2(_15991_),
    .B(_15994_),
    .Y(_15995_));
 NAND2x1_ASAP7_75t_R _21809_ (.A(_15075_),
    .B(_00905_),
    .Y(_15996_));
 OA211x2_ASAP7_75t_R _21810_ (.A1(_15074_),
    .A2(_15940_),
    .B(_15996_),
    .C(_15081_),
    .Y(_15997_));
 NAND2x1_ASAP7_75t_R _21811_ (.A(_13680_),
    .B(_00904_),
    .Y(_15998_));
 OA211x2_ASAP7_75t_R _21812_ (.A1(_15138_),
    .A2(_15943_),
    .B(_15998_),
    .C(_15109_),
    .Y(_15999_));
 OR3x1_ASAP7_75t_R _21813_ (.A(_13856_),
    .B(_15997_),
    .C(_15999_),
    .Y(_16000_));
 OA211x2_ASAP7_75t_R _21814_ (.A1(_13903_),
    .A2(_15995_),
    .B(_16000_),
    .C(_14791_),
    .Y(_16001_));
 OR3x4_ASAP7_75t_R _21815_ (.A(_15025_),
    .B(_15989_),
    .C(_16001_),
    .Y(_16002_));
 INVx2_ASAP7_75t_R _21816_ (.A(_00050_),
    .Y(_16003_));
 OA211x2_ASAP7_75t_R _21817_ (.A1(_15114_),
    .A2(_15115_),
    .B(_16003_),
    .C(_13367_),
    .Y(_16004_));
 AO31x2_ASAP7_75t_R _21818_ (.A1(_13660_),
    .A2(_15978_),
    .A3(_16002_),
    .B(_16004_),
    .Y(_16005_));
 INVx1_ASAP7_75t_R _21819_ (.A(_01537_),
    .Y(_16006_));
 AND2x2_ASAP7_75t_R _21820_ (.A(_16006_),
    .B(_13642_),
    .Y(_16007_));
 AO21x1_ASAP7_75t_R _21821_ (.A1(_15953_),
    .A2(_16005_),
    .B(_16007_),
    .Y(_16008_));
 BUFx4f_ASAP7_75t_R _21822_ (.A(_16008_),
    .Y(_18685_));
 INVx1_ASAP7_75t_R _21823_ (.A(_18685_),
    .Y(_18683_));
 BUFx4f_ASAP7_75t_R _21824_ (.A(_00888_),
    .Y(_16009_));
 OR4x2_ASAP7_75t_R _21825_ (.A(_15470_),
    .B(_15469_),
    .C(net1983),
    .D(net1976),
    .Y(_16010_));
 OA21x2_ASAP7_75t_R _21826_ (.A1(_15243_),
    .A2(_15472_),
    .B(_15478_),
    .Y(_16011_));
 OA21x2_ASAP7_75t_R _21827_ (.A1(_00817_),
    .A2(_15470_),
    .B(_00820_),
    .Y(_16012_));
 OR4x1_ASAP7_75t_R _21828_ (.A(_15469_),
    .B(net1976),
    .C(net1983),
    .D(_16012_),
    .Y(_16013_));
 OA211x2_ASAP7_75t_R _21829_ (.A1(_16010_),
    .A2(_16011_),
    .B(_16013_),
    .C(_00889_),
    .Y(_16014_));
 OA21x2_ASAP7_75t_R _21830_ (.A1(_00823_),
    .A2(_00822_),
    .B(_00856_),
    .Y(_16015_));
 OR3x1_ASAP7_75t_R _21831_ (.A(net1987),
    .B(_00888_),
    .C(_16015_),
    .Y(_16016_));
 OA211x2_ASAP7_75t_R _21832_ (.A1(_16009_),
    .A2(_16014_),
    .B(_16016_),
    .C(_00922_),
    .Y(_16017_));
 XOR2x2_ASAP7_75t_R _21833_ (.A(net2028),
    .B(_16017_),
    .Y(\alu_adder_result_ex[15] ));
 NAND2x1_ASAP7_75t_R _21834_ (.A(_15260_),
    .B(_15268_),
    .Y(_16018_));
 AO21x1_ASAP7_75t_R _21835_ (.A1(_15471_),
    .A2(_15475_),
    .B(_16010_),
    .Y(_16019_));
 OA21x2_ASAP7_75t_R _21836_ (.A1(net1976),
    .A2(_15729_),
    .B(_00856_),
    .Y(_16020_));
 OA21x2_ASAP7_75t_R _21837_ (.A1(net1984),
    .A2(_16020_),
    .B(_00889_),
    .Y(_16021_));
 NAND2x1_ASAP7_75t_R _21838_ (.A(_16019_),
    .B(_16021_),
    .Y(_16022_));
 XNOR2x1_ASAP7_75t_R _21839_ (.B(_16022_),
    .Y(_16023_),
    .A(_16009_));
 OR2x2_ASAP7_75t_R _21840_ (.A(_15475_),
    .B(_16010_),
    .Y(_16024_));
 NAND2x1_ASAP7_75t_R _21841_ (.A(_16021_),
    .B(_16024_),
    .Y(_16025_));
 XNOR2x1_ASAP7_75t_R _21842_ (.B(_16025_),
    .Y(_16026_),
    .A(_16009_));
 AO21x1_ASAP7_75t_R _21843_ (.A1(_15260_),
    .A2(_15268_),
    .B(_16026_),
    .Y(_16027_));
 OAI21x1_ASAP7_75t_R _21844_ (.A1(_16018_),
    .A2(_16023_),
    .B(_16027_),
    .Y(_16028_));
 INVx3_ASAP7_75t_R _21845_ (.A(_16028_),
    .Y(\alu_adder_result_ex[14] ));
 BUFx6f_ASAP7_75t_R _21846_ (.A(_15515_),
    .Y(_16029_));
 AND2x2_ASAP7_75t_R _21847_ (.A(_16029_),
    .B(_01807_),
    .Y(_16030_));
 AO21x1_ASAP7_75t_R _21848_ (.A1(_15871_),
    .A2(_00924_),
    .B(_16030_),
    .Y(_16031_));
 OAI22x1_ASAP7_75t_R _21849_ (.A1(_00923_),
    .A2(_15500_),
    .B1(_16031_),
    .B2(_15931_),
    .Y(_16032_));
 INVx1_ASAP7_75t_R _21850_ (.A(_00932_),
    .Y(_16033_));
 NAND2x1_ASAP7_75t_R _21851_ (.A(_15586_),
    .B(_00930_),
    .Y(_16034_));
 OA211x2_ASAP7_75t_R _21852_ (.A1(_15627_),
    .A2(_16033_),
    .B(_16034_),
    .C(_15879_),
    .Y(_16035_));
 BUFx4f_ASAP7_75t_R _21853_ (.A(_15534_),
    .Y(_16036_));
 INVx2_ASAP7_75t_R _21854_ (.A(_00931_),
    .Y(_16037_));
 NAND2x1_ASAP7_75t_R _21855_ (.A(_15651_),
    .B(_00929_),
    .Y(_16038_));
 OA211x2_ASAP7_75t_R _21856_ (.A1(_16036_),
    .A2(_16037_),
    .B(_16038_),
    .C(_15945_),
    .Y(_16039_));
 OR3x1_ASAP7_75t_R _21857_ (.A(_15876_),
    .B(_16035_),
    .C(_16039_),
    .Y(_16040_));
 OA211x2_ASAP7_75t_R _21858_ (.A1(_15531_),
    .A2(_16032_),
    .B(_16040_),
    .C(_15746_),
    .Y(_16041_));
 INVx2_ASAP7_75t_R _21859_ (.A(_00928_),
    .Y(_16042_));
 NAND2x1_ASAP7_75t_R _21860_ (.A(_15897_),
    .B(_00926_),
    .Y(_16043_));
 BUFx4f_ASAP7_75t_R _21861_ (.A(_15518_),
    .Y(_16044_));
 OA211x2_ASAP7_75t_R _21862_ (.A1(_15756_),
    .A2(_16042_),
    .B(_16043_),
    .C(_16044_),
    .Y(_16045_));
 BUFx6f_ASAP7_75t_R _21863_ (.A(_15541_),
    .Y(_16046_));
 INVx2_ASAP7_75t_R _21864_ (.A(_00927_),
    .Y(_16047_));
 BUFx6f_ASAP7_75t_R _21865_ (.A(net15),
    .Y(_16048_));
 NAND2x1_ASAP7_75t_R _21866_ (.A(_16048_),
    .B(_00925_),
    .Y(_16049_));
 OA211x2_ASAP7_75t_R _21867_ (.A1(_16046_),
    .A2(_16047_),
    .B(_16049_),
    .C(_15930_),
    .Y(_16050_));
 OR3x1_ASAP7_75t_R _21868_ (.A(_15869_),
    .B(_16045_),
    .C(_16050_),
    .Y(_16051_));
 INVx1_ASAP7_75t_R _21869_ (.A(_00936_),
    .Y(_16052_));
 NAND2x1_ASAP7_75t_R _21870_ (.A(_15897_),
    .B(_00934_),
    .Y(_16053_));
 OA211x2_ASAP7_75t_R _21871_ (.A1(_15756_),
    .A2(_16052_),
    .B(_16053_),
    .C(_16044_),
    .Y(_16054_));
 INVx1_ASAP7_75t_R _21872_ (.A(_00935_),
    .Y(_16055_));
 NAND2x1_ASAP7_75t_R _21873_ (.A(_16048_),
    .B(_00933_),
    .Y(_16056_));
 OA211x2_ASAP7_75t_R _21874_ (.A1(_16046_),
    .A2(_16055_),
    .B(_16056_),
    .C(_15930_),
    .Y(_16057_));
 OR3x1_ASAP7_75t_R _21875_ (.A(_15902_),
    .B(_16054_),
    .C(_16057_),
    .Y(_16058_));
 AND3x1_ASAP7_75t_R _21876_ (.A(_15528_),
    .B(_16051_),
    .C(_16058_),
    .Y(_16059_));
 OR3x4_ASAP7_75t_R _21877_ (.A(_15497_),
    .B(_16041_),
    .C(_16059_),
    .Y(_16060_));
 INVx2_ASAP7_75t_R _21878_ (.A(_00944_),
    .Y(_16061_));
 NAND2x1_ASAP7_75t_R _21879_ (.A(_15897_),
    .B(_00942_),
    .Y(_16062_));
 OA211x2_ASAP7_75t_R _21880_ (.A1(_15895_),
    .A2(_16061_),
    .B(_16062_),
    .C(_15893_),
    .Y(_16063_));
 INVx2_ASAP7_75t_R _21881_ (.A(_00943_),
    .Y(_16064_));
 NAND2x1_ASAP7_75t_R _21882_ (.A(_16048_),
    .B(_00941_),
    .Y(_16065_));
 OA211x2_ASAP7_75t_R _21883_ (.A1(_15756_),
    .A2(_16064_),
    .B(_16065_),
    .C(_15899_),
    .Y(_16066_));
 OR3x1_ASAP7_75t_R _21884_ (.A(_15869_),
    .B(_16063_),
    .C(_16066_),
    .Y(_16067_));
 INVx2_ASAP7_75t_R _21885_ (.A(_00952_),
    .Y(_16068_));
 NAND2x1_ASAP7_75t_R _21886_ (.A(_15897_),
    .B(_00950_),
    .Y(_16069_));
 OA211x2_ASAP7_75t_R _21887_ (.A1(_15756_),
    .A2(_16068_),
    .B(_16069_),
    .C(_16044_),
    .Y(_16070_));
 INVx3_ASAP7_75t_R _21888_ (.A(_00951_),
    .Y(_16071_));
 NAND2x1_ASAP7_75t_R _21889_ (.A(_16048_),
    .B(_00949_),
    .Y(_16072_));
 OA211x2_ASAP7_75t_R _21890_ (.A1(_16046_),
    .A2(_16071_),
    .B(_16072_),
    .C(_15899_),
    .Y(_16073_));
 OR3x1_ASAP7_75t_R _21891_ (.A(_15902_),
    .B(_16070_),
    .C(_16073_),
    .Y(_16074_));
 AND3x1_ASAP7_75t_R _21892_ (.A(_15528_),
    .B(_16067_),
    .C(_16074_),
    .Y(_16075_));
 INVx1_ASAP7_75t_R _21893_ (.A(_00945_),
    .Y(_16076_));
 NOR2x1_ASAP7_75t_R _21894_ (.A(_15542_),
    .B(_00947_),
    .Y(_16077_));
 AO21x1_ASAP7_75t_R _21895_ (.A1(_15749_),
    .A2(_16076_),
    .B(_16077_),
    .Y(_16078_));
 BUFx12f_ASAP7_75t_R _21896_ (.A(_15504_),
    .Y(_16079_));
 INVx2_ASAP7_75t_R _21897_ (.A(_00948_),
    .Y(_16080_));
 NAND2x1_ASAP7_75t_R _21898_ (.A(_15532_),
    .B(_00946_),
    .Y(_16081_));
 BUFx4f_ASAP7_75t_R _21899_ (.A(_15518_),
    .Y(_16082_));
 OA211x2_ASAP7_75t_R _21900_ (.A1(_16079_),
    .A2(_16080_),
    .B(_16081_),
    .C(_16082_),
    .Y(_16083_));
 AO21x1_ASAP7_75t_R _21901_ (.A1(_15931_),
    .A2(_16078_),
    .B(_16083_),
    .Y(_16084_));
 INVx2_ASAP7_75t_R _21902_ (.A(_00940_),
    .Y(_16085_));
 NAND2x1_ASAP7_75t_R _21903_ (.A(_15651_),
    .B(_00938_),
    .Y(_16086_));
 OA211x2_ASAP7_75t_R _21904_ (.A1(_16036_),
    .A2(_16085_),
    .B(_16086_),
    .C(_15879_),
    .Y(_16087_));
 INVx2_ASAP7_75t_R _21905_ (.A(_00939_),
    .Y(_16088_));
 NAND2x1_ASAP7_75t_R _21906_ (.A(_15651_),
    .B(_00937_),
    .Y(_16089_));
 OA211x2_ASAP7_75t_R _21907_ (.A1(_15570_),
    .A2(_16088_),
    .B(_16089_),
    .C(_15945_),
    .Y(_16090_));
 OR3x1_ASAP7_75t_R _21908_ (.A(_15530_),
    .B(_16087_),
    .C(_16090_),
    .Y(_16091_));
 OA211x2_ASAP7_75t_R _21909_ (.A1(_15929_),
    .A2(_16084_),
    .B(_16091_),
    .C(_15746_),
    .Y(_16092_));
 OR3x4_ASAP7_75t_R _21910_ (.A(_15912_),
    .B(_16075_),
    .C(_16092_),
    .Y(_16093_));
 AND2x4_ASAP7_75t_R _21911_ (.A(_16060_),
    .B(_16093_),
    .Y(_16094_));
 AO21x1_ASAP7_75t_R _21912_ (.A1(_13777_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_16095_));
 AND2x2_ASAP7_75t_R _21913_ (.A(_15491_),
    .B(_16095_),
    .Y(_16096_));
 AO21x2_ASAP7_75t_R _21914_ (.A1(_15496_),
    .A2(_16094_),
    .B(_16096_),
    .Y(_18688_));
 AND2x2_ASAP7_75t_R _21915_ (.A(_13882_),
    .B(_01807_),
    .Y(_16097_));
 AO21x1_ASAP7_75t_R _21916_ (.A1(_14742_),
    .A2(_00924_),
    .B(_16097_),
    .Y(_16098_));
 OAI22x1_ASAP7_75t_R _21917_ (.A1(_00923_),
    .A2(_13948_),
    .B1(_16098_),
    .B2(_14746_),
    .Y(_16099_));
 NAND2x1_ASAP7_75t_R _21918_ (.A(_15424_),
    .B(_00930_),
    .Y(_16100_));
 OA211x2_ASAP7_75t_R _21919_ (.A1(_15423_),
    .A2(_16033_),
    .B(_16100_),
    .C(_15282_),
    .Y(_16101_));
 NAND2x1_ASAP7_75t_R _21920_ (.A(_15280_),
    .B(_00929_),
    .Y(_16102_));
 OA211x2_ASAP7_75t_R _21921_ (.A1(_15278_),
    .A2(_16037_),
    .B(_16102_),
    .C(_14850_),
    .Y(_16103_));
 OR3x1_ASAP7_75t_R _21922_ (.A(_14853_),
    .B(_16101_),
    .C(_16103_),
    .Y(_16104_));
 OA211x2_ASAP7_75t_R _21923_ (.A1(_14740_),
    .A2(_16099_),
    .B(_16104_),
    .C(_14863_),
    .Y(_16105_));
 NAND2x1_ASAP7_75t_R _21924_ (.A(_14816_),
    .B(_00926_),
    .Y(_16106_));
 OA211x2_ASAP7_75t_R _21925_ (.A1(_15307_),
    .A2(_16042_),
    .B(_16106_),
    .C(_15305_),
    .Y(_16107_));
 NAND2x1_ASAP7_75t_R _21926_ (.A(_13952_),
    .B(_00925_),
    .Y(_16108_));
 OA211x2_ASAP7_75t_R _21927_ (.A1(_15290_),
    .A2(_16047_),
    .B(_16108_),
    .C(_15309_),
    .Y(_16109_));
 OR3x1_ASAP7_75t_R _21928_ (.A(_14985_),
    .B(_16107_),
    .C(_16109_),
    .Y(_16110_));
 NAND2x1_ASAP7_75t_R _21929_ (.A(_14816_),
    .B(_00934_),
    .Y(_16111_));
 OA211x2_ASAP7_75t_R _21930_ (.A1(_15307_),
    .A2(_16052_),
    .B(_16111_),
    .C(_15129_),
    .Y(_16112_));
 NAND2x1_ASAP7_75t_R _21931_ (.A(_13952_),
    .B(_00933_),
    .Y(_16113_));
 OA211x2_ASAP7_75t_R _21932_ (.A1(_14987_),
    .A2(_16055_),
    .B(_16113_),
    .C(_15134_),
    .Y(_16114_));
 OR3x1_ASAP7_75t_R _21933_ (.A(_15125_),
    .B(_16112_),
    .C(_16114_),
    .Y(_16115_));
 AND3x1_ASAP7_75t_R _21934_ (.A(_15289_),
    .B(_16110_),
    .C(_16115_),
    .Y(_16116_));
 OR3x4_ASAP7_75t_R _21935_ (.A(_14814_),
    .B(_16105_),
    .C(_16116_),
    .Y(_16117_));
 NAND2x1_ASAP7_75t_R _21936_ (.A(_13935_),
    .B(_00942_),
    .Y(_16118_));
 OA211x2_ASAP7_75t_R _21937_ (.A1(_15307_),
    .A2(_16061_),
    .B(_16118_),
    .C(_15305_),
    .Y(_16119_));
 NAND2x1_ASAP7_75t_R _21938_ (.A(_13952_),
    .B(_00941_),
    .Y(_16120_));
 OA211x2_ASAP7_75t_R _21939_ (.A1(_15290_),
    .A2(_16064_),
    .B(_16120_),
    .C(_15309_),
    .Y(_16121_));
 OR3x1_ASAP7_75t_R _21940_ (.A(_14760_),
    .B(_16119_),
    .C(_16121_),
    .Y(_16122_));
 NAND2x1_ASAP7_75t_R _21941_ (.A(_14816_),
    .B(_00950_),
    .Y(_16123_));
 OA211x2_ASAP7_75t_R _21942_ (.A1(_15307_),
    .A2(_16068_),
    .B(_16123_),
    .C(_15129_),
    .Y(_16124_));
 NAND2x1_ASAP7_75t_R _21943_ (.A(_13952_),
    .B(_00949_),
    .Y(_16125_));
 OA211x2_ASAP7_75t_R _21944_ (.A1(_15290_),
    .A2(_16071_),
    .B(_16125_),
    .C(_15309_),
    .Y(_16126_));
 OR3x1_ASAP7_75t_R _21945_ (.A(_15125_),
    .B(_16124_),
    .C(_16126_),
    .Y(_16127_));
 AND3x1_ASAP7_75t_R _21946_ (.A(_15289_),
    .B(_16122_),
    .C(_16127_),
    .Y(_16128_));
 NOR2x1_ASAP7_75t_R _21947_ (.A(_14749_),
    .B(_00947_),
    .Y(_16129_));
 AO21x1_ASAP7_75t_R _21948_ (.A1(_15319_),
    .A2(_16076_),
    .B(_16129_),
    .Y(_16130_));
 NAND2x1_ASAP7_75t_R _21949_ (.A(_14778_),
    .B(_00946_),
    .Y(_16131_));
 OA211x2_ASAP7_75t_R _21950_ (.A1(_14761_),
    .A2(_16080_),
    .B(_16131_),
    .C(_13869_),
    .Y(_16132_));
 AO21x1_ASAP7_75t_R _21951_ (.A1(_13716_),
    .A2(_16130_),
    .B(_16132_),
    .Y(_16133_));
 NAND2x1_ASAP7_75t_R _21952_ (.A(_15280_),
    .B(_00938_),
    .Y(_16134_));
 OA211x2_ASAP7_75t_R _21953_ (.A1(_15278_),
    .A2(_16085_),
    .B(_16134_),
    .C(_14846_),
    .Y(_16135_));
 NAND2x1_ASAP7_75t_R _21954_ (.A(_13756_),
    .B(_00937_),
    .Y(_16136_));
 OA211x2_ASAP7_75t_R _21955_ (.A1(_14844_),
    .A2(_16088_),
    .B(_16136_),
    .C(_14850_),
    .Y(_16137_));
 OR3x1_ASAP7_75t_R _21956_ (.A(_14739_),
    .B(_16135_),
    .C(_16137_),
    .Y(_16138_));
 OA211x2_ASAP7_75t_R _21957_ (.A1(_15318_),
    .A2(_16133_),
    .B(_16138_),
    .C(_14863_),
    .Y(_16139_));
 OR3x4_ASAP7_75t_R _21958_ (.A(_14842_),
    .B(_16128_),
    .C(_16139_),
    .Y(_16140_));
 INVx1_ASAP7_75t_R _21959_ (.A(_00051_),
    .Y(_16141_));
 OA211x2_ASAP7_75t_R _21960_ (.A1(_13647_),
    .A2(_13658_),
    .B(_16141_),
    .C(_15334_),
    .Y(_16142_));
 AO31x2_ASAP7_75t_R _21961_ (.A1(_13947_),
    .A2(_16117_),
    .A3(_16140_),
    .B(_16142_),
    .Y(_16143_));
 INVx1_ASAP7_75t_R _21962_ (.A(_01536_),
    .Y(_16144_));
 AO32x1_ASAP7_75t_R _21963_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_16143_),
    .B1(_15337_),
    .B2(_16144_),
    .Y(_16145_));
 BUFx6f_ASAP7_75t_R _21964_ (.A(_16145_),
    .Y(_18687_));
 INVx1_ASAP7_75t_R _21965_ (.A(_18687_),
    .Y(_18689_));
 AND2x2_ASAP7_75t_R _21966_ (.A(_16036_),
    .B(_01806_),
    .Y(_16146_));
 AO21x1_ASAP7_75t_R _21967_ (.A1(_15871_),
    .A2(_00957_),
    .B(_16146_),
    .Y(_16147_));
 OAI22x1_ASAP7_75t_R _21968_ (.A1(_00956_),
    .A2(_15500_),
    .B1(_16147_),
    .B2(_15649_),
    .Y(_16148_));
 BUFx6f_ASAP7_75t_R _21969_ (.A(_15534_),
    .Y(_16149_));
 INVx1_ASAP7_75t_R _21970_ (.A(_00965_),
    .Y(_16150_));
 BUFx10_ASAP7_75t_R _21971_ (.A(net15),
    .Y(_16151_));
 NAND2x1_ASAP7_75t_R _21972_ (.A(_16151_),
    .B(_00963_),
    .Y(_16152_));
 BUFx6f_ASAP7_75t_R _21973_ (.A(net10),
    .Y(_16153_));
 OA211x2_ASAP7_75t_R _21974_ (.A1(_16149_),
    .A2(_16150_),
    .B(_16152_),
    .C(_16153_),
    .Y(_16154_));
 INVx1_ASAP7_75t_R _21975_ (.A(_00964_),
    .Y(_16155_));
 NAND2x1_ASAP7_75t_R _21976_ (.A(_16151_),
    .B(_00962_),
    .Y(_16156_));
 OA211x2_ASAP7_75t_R _21977_ (.A1(_15656_),
    .A2(_16155_),
    .B(_16156_),
    .C(_15883_),
    .Y(_16157_));
 OR3x1_ASAP7_75t_R _21978_ (.A(_15876_),
    .B(_16154_),
    .C(_16157_),
    .Y(_16158_));
 BUFx3_ASAP7_75t_R _21979_ (.A(_13512_),
    .Y(_16159_));
 OA211x2_ASAP7_75t_R _21980_ (.A1(_15870_),
    .A2(_16148_),
    .B(_16158_),
    .C(_16159_),
    .Y(_16160_));
 BUFx6f_ASAP7_75t_R _21981_ (.A(_15541_),
    .Y(_16161_));
 INVx1_ASAP7_75t_R _21982_ (.A(_00961_),
    .Y(_16162_));
 NAND2x1_ASAP7_75t_R _21983_ (.A(_15576_),
    .B(_00959_),
    .Y(_16163_));
 OA211x2_ASAP7_75t_R _21984_ (.A1(_16161_),
    .A2(_16162_),
    .B(_16163_),
    .C(_15807_),
    .Y(_16164_));
 INVx2_ASAP7_75t_R _21985_ (.A(_00960_),
    .Y(_16165_));
 NAND2x1_ASAP7_75t_R _21986_ (.A(_15936_),
    .B(_00958_),
    .Y(_16166_));
 OA211x2_ASAP7_75t_R _21987_ (.A1(_15505_),
    .A2(_16165_),
    .B(_16166_),
    .C(_15811_),
    .Y(_16167_));
 OR3x1_ASAP7_75t_R _21988_ (.A(_15888_),
    .B(_16164_),
    .C(_16167_),
    .Y(_16168_));
 INVx1_ASAP7_75t_R _21989_ (.A(_00969_),
    .Y(_16169_));
 NAND2x1_ASAP7_75t_R _21990_ (.A(_15576_),
    .B(_00967_),
    .Y(_16170_));
 OA211x2_ASAP7_75t_R _21991_ (.A1(_15505_),
    .A2(_16169_),
    .B(_16170_),
    .C(_15807_),
    .Y(_16171_));
 INVx1_ASAP7_75t_R _21992_ (.A(_00968_),
    .Y(_16172_));
 NAND2x1_ASAP7_75t_R _21993_ (.A(_15936_),
    .B(_00966_),
    .Y(_16173_));
 OA211x2_ASAP7_75t_R _21994_ (.A1(_15594_),
    .A2(_16172_),
    .B(_16173_),
    .C(_15811_),
    .Y(_16174_));
 OR3x1_ASAP7_75t_R _21995_ (.A(_15567_),
    .B(_16171_),
    .C(_16174_),
    .Y(_16175_));
 AND3x1_ASAP7_75t_R _21996_ (.A(_15887_),
    .B(_16168_),
    .C(_16175_),
    .Y(_16176_));
 OR3x4_ASAP7_75t_R _21997_ (.A(_15497_),
    .B(_16160_),
    .C(_16176_),
    .Y(_16177_));
 INVx1_ASAP7_75t_R _21998_ (.A(_00977_),
    .Y(_16178_));
 NAND2x1_ASAP7_75t_R _21999_ (.A(_15576_),
    .B(_00975_),
    .Y(_16179_));
 OA211x2_ASAP7_75t_R _22000_ (.A1(_16161_),
    .A2(_16178_),
    .B(_16179_),
    .C(_15807_),
    .Y(_16180_));
 INVx1_ASAP7_75t_R _22001_ (.A(_00976_),
    .Y(_16181_));
 NAND2x1_ASAP7_75t_R _22002_ (.A(_15576_),
    .B(_00974_),
    .Y(_16182_));
 OA211x2_ASAP7_75t_R _22003_ (.A1(_15505_),
    .A2(_16181_),
    .B(_16182_),
    .C(_15811_),
    .Y(_16183_));
 OR3x1_ASAP7_75t_R _22004_ (.A(_15498_),
    .B(_16180_),
    .C(_16183_),
    .Y(_16184_));
 INVx1_ASAP7_75t_R _22005_ (.A(_00985_),
    .Y(_16185_));
 NAND2x1_ASAP7_75t_R _22006_ (.A(_15576_),
    .B(_00983_),
    .Y(_16186_));
 OA211x2_ASAP7_75t_R _22007_ (.A1(_16161_),
    .A2(_16185_),
    .B(_16186_),
    .C(_15807_),
    .Y(_16187_));
 INVx1_ASAP7_75t_R _22008_ (.A(_00984_),
    .Y(_16188_));
 NAND2x1_ASAP7_75t_R _22009_ (.A(_15576_),
    .B(_00982_),
    .Y(_16189_));
 OA211x2_ASAP7_75t_R _22010_ (.A1(_15505_),
    .A2(_16188_),
    .B(_16189_),
    .C(_15811_),
    .Y(_16190_));
 OR3x1_ASAP7_75t_R _22011_ (.A(_15567_),
    .B(_16187_),
    .C(_16190_),
    .Y(_16191_));
 AND3x1_ASAP7_75t_R _22012_ (.A(_15887_),
    .B(_16184_),
    .C(_16191_),
    .Y(_16192_));
 INVx2_ASAP7_75t_R _22013_ (.A(_00978_),
    .Y(_16193_));
 NOR2x1_ASAP7_75t_R _22014_ (.A(_15767_),
    .B(_00980_),
    .Y(_16194_));
 AO21x1_ASAP7_75t_R _22015_ (.A1(_15533_),
    .A2(_16193_),
    .B(_16194_),
    .Y(_16195_));
 INVx1_ASAP7_75t_R _22016_ (.A(_00981_),
    .Y(_16196_));
 NAND2x1_ASAP7_75t_R _22017_ (.A(_15602_),
    .B(_00979_),
    .Y(_16197_));
 OA211x2_ASAP7_75t_R _22018_ (.A1(_15587_),
    .A2(_16196_),
    .B(_16197_),
    .C(_15519_),
    .Y(_16198_));
 AO21x1_ASAP7_75t_R _22019_ (.A1(_15931_),
    .A2(_16195_),
    .B(_16198_),
    .Y(_16199_));
 INVx1_ASAP7_75t_R _22020_ (.A(_00973_),
    .Y(_16200_));
 NAND2x1_ASAP7_75t_R _22021_ (.A(_15572_),
    .B(_00971_),
    .Y(_16201_));
 OA211x2_ASAP7_75t_R _22022_ (.A1(_15656_),
    .A2(_16200_),
    .B(_16201_),
    .C(_16153_),
    .Y(_16202_));
 INVx1_ASAP7_75t_R _22023_ (.A(_00972_),
    .Y(_16203_));
 NAND2x1_ASAP7_75t_R _22024_ (.A(_15572_),
    .B(_00970_),
    .Y(_16204_));
 OA211x2_ASAP7_75t_R _22025_ (.A1(_15535_),
    .A2(_16203_),
    .B(_16204_),
    .C(_15883_),
    .Y(_16205_));
 OR3x1_ASAP7_75t_R _22026_ (.A(_15869_),
    .B(_16202_),
    .C(_16205_),
    .Y(_16206_));
 OA211x2_ASAP7_75t_R _22027_ (.A1(_15929_),
    .A2(_16199_),
    .B(_16206_),
    .C(_16159_),
    .Y(_16207_));
 OR3x2_ASAP7_75t_R _22028_ (.A(_15912_),
    .B(_16192_),
    .C(_16207_),
    .Y(_16208_));
 AND2x4_ASAP7_75t_R _22029_ (.A(_16177_),
    .B(_16208_),
    .Y(_16209_));
 AO21x1_ASAP7_75t_R _22030_ (.A1(_14732_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_16210_));
 AND2x2_ASAP7_75t_R _22031_ (.A(_15491_),
    .B(_16210_),
    .Y(_16211_));
 AO21x2_ASAP7_75t_R _22032_ (.A1(_15496_),
    .A2(_16209_),
    .B(_16211_),
    .Y(_18693_));
 AND2x2_ASAP7_75t_R _22033_ (.A(_15075_),
    .B(_01806_),
    .Y(_16212_));
 AO21x1_ASAP7_75t_R _22034_ (.A1(_14742_),
    .A2(_00957_),
    .B(_16212_),
    .Y(_16213_));
 OAI22x1_ASAP7_75t_R _22035_ (.A1(_00956_),
    .A2(_13948_),
    .B1(_16213_),
    .B2(_13918_),
    .Y(_16214_));
 NAND2x1_ASAP7_75t_R _22036_ (.A(_15280_),
    .B(_00963_),
    .Y(_16215_));
 OA211x2_ASAP7_75t_R _22037_ (.A1(_15278_),
    .A2(_16150_),
    .B(_16215_),
    .C(_15282_),
    .Y(_16216_));
 NAND2x1_ASAP7_75t_R _22038_ (.A(_15280_),
    .B(_00962_),
    .Y(_16217_));
 OA211x2_ASAP7_75t_R _22039_ (.A1(_14844_),
    .A2(_16155_),
    .B(_16217_),
    .C(_14850_),
    .Y(_16218_));
 OR3x1_ASAP7_75t_R _22040_ (.A(_14853_),
    .B(_16216_),
    .C(_16218_),
    .Y(_16219_));
 OA211x2_ASAP7_75t_R _22041_ (.A1(_14740_),
    .A2(_16214_),
    .B(_16219_),
    .C(_14863_),
    .Y(_16220_));
 NAND2x1_ASAP7_75t_R _22042_ (.A(_13952_),
    .B(_00959_),
    .Y(_16221_));
 OA211x2_ASAP7_75t_R _22043_ (.A1(_14987_),
    .A2(_16162_),
    .B(_16221_),
    .C(_15129_),
    .Y(_16222_));
 NAND2x1_ASAP7_75t_R _22044_ (.A(_13956_),
    .B(_00958_),
    .Y(_16223_));
 OA211x2_ASAP7_75t_R _22045_ (.A1(_15126_),
    .A2(_16165_),
    .B(_16223_),
    .C(_15134_),
    .Y(_16224_));
 OR3x1_ASAP7_75t_R _22046_ (.A(_14985_),
    .B(_16222_),
    .C(_16224_),
    .Y(_16225_));
 NAND2x1_ASAP7_75t_R _22047_ (.A(_13956_),
    .B(_00967_),
    .Y(_16226_));
 OA211x2_ASAP7_75t_R _22048_ (.A1(_14987_),
    .A2(_16169_),
    .B(_16226_),
    .C(_15129_),
    .Y(_16227_));
 NAND2x1_ASAP7_75t_R _22049_ (.A(_13956_),
    .B(_00966_),
    .Y(_16228_));
 OA211x2_ASAP7_75t_R _22050_ (.A1(_15126_),
    .A2(_16172_),
    .B(_16228_),
    .C(_15134_),
    .Y(_16229_));
 OR3x1_ASAP7_75t_R _22051_ (.A(_15125_),
    .B(_16227_),
    .C(_16229_),
    .Y(_16230_));
 AND3x1_ASAP7_75t_R _22052_ (.A(_15289_),
    .B(_16225_),
    .C(_16230_),
    .Y(_16231_));
 OR3x4_ASAP7_75t_R _22053_ (.A(_14814_),
    .B(_16220_),
    .C(_16231_),
    .Y(_16232_));
 NAND2x1_ASAP7_75t_R _22054_ (.A(_13952_),
    .B(_00975_),
    .Y(_16233_));
 OA211x2_ASAP7_75t_R _22055_ (.A1(_14987_),
    .A2(_16178_),
    .B(_16233_),
    .C(_15129_),
    .Y(_16234_));
 NAND2x1_ASAP7_75t_R _22056_ (.A(_13956_),
    .B(_00974_),
    .Y(_16235_));
 OA211x2_ASAP7_75t_R _22057_ (.A1(_15126_),
    .A2(_16181_),
    .B(_16235_),
    .C(_15134_),
    .Y(_16236_));
 OR3x1_ASAP7_75t_R _22058_ (.A(_14985_),
    .B(_16234_),
    .C(_16236_),
    .Y(_16237_));
 NAND2x1_ASAP7_75t_R _22059_ (.A(_13956_),
    .B(_00983_),
    .Y(_16238_));
 OA211x2_ASAP7_75t_R _22060_ (.A1(_14987_),
    .A2(_16185_),
    .B(_16238_),
    .C(_15129_),
    .Y(_16239_));
 NAND2x1_ASAP7_75t_R _22061_ (.A(_13956_),
    .B(_00982_),
    .Y(_16240_));
 OA211x2_ASAP7_75t_R _22062_ (.A1(_15126_),
    .A2(_16188_),
    .B(_16240_),
    .C(_15134_),
    .Y(_16241_));
 OR3x1_ASAP7_75t_R _22063_ (.A(_15125_),
    .B(_16239_),
    .C(_16241_),
    .Y(_16242_));
 AND3x1_ASAP7_75t_R _22064_ (.A(_15289_),
    .B(_16237_),
    .C(_16242_),
    .Y(_16243_));
 NOR2x1_ASAP7_75t_R _22065_ (.A(_14831_),
    .B(_00980_),
    .Y(_16244_));
 AO21x1_ASAP7_75t_R _22066_ (.A1(_15013_),
    .A2(_16193_),
    .B(_16244_),
    .Y(_16245_));
 NAND2x1_ASAP7_75t_R _22067_ (.A(_14764_),
    .B(_00979_),
    .Y(_16246_));
 OA211x2_ASAP7_75t_R _22068_ (.A1(_13865_),
    .A2(_16196_),
    .B(_16246_),
    .C(_13932_),
    .Y(_16247_));
 AO21x1_ASAP7_75t_R _22069_ (.A1(_13716_),
    .A2(_16245_),
    .B(_16247_),
    .Y(_16248_));
 NAND2x1_ASAP7_75t_R _22070_ (.A(_13756_),
    .B(_00971_),
    .Y(_16249_));
 OA211x2_ASAP7_75t_R _22071_ (.A1(_14854_),
    .A2(_16200_),
    .B(_16249_),
    .C(_14846_),
    .Y(_16250_));
 NAND2x1_ASAP7_75t_R _22072_ (.A(_14858_),
    .B(_00970_),
    .Y(_16251_));
 OA211x2_ASAP7_75t_R _22073_ (.A1(_14857_),
    .A2(_16203_),
    .B(_16251_),
    .C(_14850_),
    .Y(_16252_));
 OR3x1_ASAP7_75t_R _22074_ (.A(_13676_),
    .B(_16250_),
    .C(_16252_),
    .Y(_16253_));
 OA211x2_ASAP7_75t_R _22075_ (.A1(_15318_),
    .A2(_16248_),
    .B(_16253_),
    .C(_14863_),
    .Y(_16254_));
 OR3x4_ASAP7_75t_R _22076_ (.A(_14842_),
    .B(_16243_),
    .C(_16254_),
    .Y(_16255_));
 INVx1_ASAP7_75t_R _22077_ (.A(_00052_),
    .Y(_16256_));
 OA211x2_ASAP7_75t_R _22078_ (.A1(_13647_),
    .A2(_13658_),
    .B(_16256_),
    .C(_15334_),
    .Y(_16257_));
 AO31x2_ASAP7_75t_R _22079_ (.A1(_13947_),
    .A2(_16232_),
    .A3(_16255_),
    .B(_16257_),
    .Y(_16258_));
 INVx1_ASAP7_75t_R _22080_ (.A(_01535_),
    .Y(_16259_));
 AO32x1_ASAP7_75t_R _22081_ (.A1(_13771_),
    .A2(_13772_),
    .A3(_16258_),
    .B1(_13642_),
    .B2(_16259_),
    .Y(_16260_));
 BUFx4f_ASAP7_75t_R _22082_ (.A(_16260_),
    .Y(_18692_));
 INVx4_ASAP7_75t_R _22083_ (.A(_18692_),
    .Y(_18694_));
 OR4x1_ASAP7_75t_R _22084_ (.A(_15469_),
    .B(net1976),
    .C(net1986),
    .D(_00888_),
    .Y(_16261_));
 OA22x2_ASAP7_75t_R _22085_ (.A1(_00889_),
    .A2(_00888_),
    .B1(_16012_),
    .B2(_16261_),
    .Y(_16262_));
 AND5x1_ASAP7_75t_R _22086_ (.A(_00922_),
    .B(_00955_),
    .C(_00988_),
    .D(_16016_),
    .E(_16262_),
    .Y(_16263_));
 OR3x1_ASAP7_75t_R _22087_ (.A(_16009_),
    .B(_15478_),
    .C(_16010_),
    .Y(_16264_));
 OR4x1_ASAP7_75t_R _22088_ (.A(_15472_),
    .B(_15243_),
    .C(_16009_),
    .D(_16010_),
    .Y(_16265_));
 AO21x1_ASAP7_75t_R _22089_ (.A1(_00921_),
    .A2(_00955_),
    .B(_00954_),
    .Y(_16266_));
 AO32x2_ASAP7_75t_R _22090_ (.A1(_16263_),
    .A2(_16265_),
    .A3(_16264_),
    .B1(_16266_),
    .B2(_00988_),
    .Y(_16267_));
 XOR2x2_ASAP7_75t_R _22091_ (.A(_00987_),
    .B(_16267_),
    .Y(\alu_adder_result_ex[17] ));
 AND4x2_ASAP7_75t_R _22092_ (.A(_14898_),
    .B(_14909_),
    .C(_14914_),
    .D(_14925_),
    .Y(_16268_));
 AO21x1_ASAP7_75t_R _22093_ (.A1(_14920_),
    .A2(_14919_),
    .B(_15403_),
    .Y(_16269_));
 INVx1_ASAP7_75t_R _22094_ (.A(_00954_),
    .Y(_16270_));
 OA21x2_ASAP7_75t_R _22095_ (.A1(net1977),
    .A2(_15740_),
    .B(_00856_),
    .Y(_16271_));
 OR3x1_ASAP7_75t_R _22096_ (.A(net1985),
    .B(_16009_),
    .C(net2029),
    .Y(_16272_));
 OR5x1_ASAP7_75t_R _22097_ (.A(_16009_),
    .B(net2029),
    .C(_15405_),
    .D(_15473_),
    .E(_16010_),
    .Y(_16273_));
 OA21x2_ASAP7_75t_R _22098_ (.A1(_00922_),
    .A2(_00921_),
    .B(_00955_),
    .Y(_16274_));
 OR3x1_ASAP7_75t_R _22099_ (.A(_00889_),
    .B(_16009_),
    .C(net2029),
    .Y(_16275_));
 AND3x1_ASAP7_75t_R _22100_ (.A(_16273_),
    .B(_16274_),
    .C(_16275_),
    .Y(_16276_));
 OA21x2_ASAP7_75t_R _22101_ (.A1(_16271_),
    .A2(_16272_),
    .B(_16276_),
    .Y(_16277_));
 AND3x1_ASAP7_75t_R _22102_ (.A(_16270_),
    .B(_15408_),
    .C(_16277_),
    .Y(_16278_));
 OA21x2_ASAP7_75t_R _22103_ (.A1(_16268_),
    .A2(_16269_),
    .B(_16278_),
    .Y(_16279_));
 OR5x2_ASAP7_75t_R _22104_ (.A(_16009_),
    .B(net2029),
    .C(_15401_),
    .D(_15473_),
    .E(_16010_),
    .Y(_16280_));
 OAI21x1_ASAP7_75t_R _22105_ (.A1(_15408_),
    .A2(_16280_),
    .B(_16277_),
    .Y(_16281_));
 OA211x2_ASAP7_75t_R _22106_ (.A1(_16271_),
    .A2(_16272_),
    .B(_16276_),
    .C(_16280_),
    .Y(_16282_));
 AND2x2_ASAP7_75t_R _22107_ (.A(_16270_),
    .B(_16282_),
    .Y(_16283_));
 AO21x1_ASAP7_75t_R _22108_ (.A1(_00954_),
    .A2(_16281_),
    .B(_16283_),
    .Y(_16284_));
 OR3x1_ASAP7_75t_R _22109_ (.A(_15252_),
    .B(_15250_),
    .C(_15248_),
    .Y(_16285_));
 AND3x4_ASAP7_75t_R _22110_ (.A(_13602_),
    .B(_13587_),
    .C(_13606_),
    .Y(_16286_));
 AOI21x1_ASAP7_75t_R _22111_ (.A1(_14920_),
    .A2(_14919_),
    .B(_15403_),
    .Y(_16287_));
 NOR2x1_ASAP7_75t_R _22112_ (.A(_16270_),
    .B(_16280_),
    .Y(_16288_));
 OA211x2_ASAP7_75t_R _22113_ (.A1(_16285_),
    .A2(_16286_),
    .B(_16287_),
    .C(_16288_),
    .Y(_16289_));
 OR3x1_ASAP7_75t_R _22114_ (.A(_16279_),
    .B(_16284_),
    .C(_16289_),
    .Y(_16290_));
 BUFx6f_ASAP7_75t_R _22115_ (.A(_16290_),
    .Y(\alu_adder_result_ex[16] ));
 AND2x2_ASAP7_75t_R _22116_ (.A(_15767_),
    .B(_01805_),
    .Y(_16291_));
 AO21x1_ASAP7_75t_R _22117_ (.A1(_15871_),
    .A2(_00990_),
    .B(_16291_),
    .Y(_16292_));
 OAI22x1_ASAP7_75t_R _22118_ (.A1(_00989_),
    .A2(_15500_),
    .B1(_16292_),
    .B2(_15569_),
    .Y(_16293_));
 INVx1_ASAP7_75t_R _22119_ (.A(_00998_),
    .Y(_16294_));
 NAND2x1_ASAP7_75t_R _22120_ (.A(_15532_),
    .B(_00996_),
    .Y(_16295_));
 OA211x2_ASAP7_75t_R _22121_ (.A1(_16079_),
    .A2(_16294_),
    .B(_16295_),
    .C(_16082_),
    .Y(_16296_));
 INVx1_ASAP7_75t_R _22122_ (.A(_00997_),
    .Y(_16297_));
 NAND2x1_ASAP7_75t_R _22123_ (.A(_15891_),
    .B(_00995_),
    .Y(_16298_));
 OA211x2_ASAP7_75t_R _22124_ (.A1(_16079_),
    .A2(_16297_),
    .B(_16298_),
    .C(_15918_),
    .Y(_16299_));
 OR3x1_ASAP7_75t_R _22125_ (.A(_15567_),
    .B(_16296_),
    .C(_16299_),
    .Y(_16300_));
 OA211x2_ASAP7_75t_R _22126_ (.A1(_15870_),
    .A2(_16293_),
    .B(_16300_),
    .C(_16159_),
    .Y(_16301_));
 INVx1_ASAP7_75t_R _22127_ (.A(_00994_),
    .Y(_16302_));
 BUFx6f_ASAP7_75t_R _22128_ (.A(_15515_),
    .Y(_16303_));
 NAND2x1_ASAP7_75t_R _22129_ (.A(_16303_),
    .B(_00992_),
    .Y(_16304_));
 BUFx3_ASAP7_75t_R _22130_ (.A(_15537_),
    .Y(_16305_));
 OA211x2_ASAP7_75t_R _22131_ (.A1(_15573_),
    .A2(_16302_),
    .B(_16304_),
    .C(_16305_),
    .Y(_16306_));
 INVx1_ASAP7_75t_R _22132_ (.A(_00993_),
    .Y(_16307_));
 NAND2x1_ASAP7_75t_R _22133_ (.A(_16303_),
    .B(_00991_),
    .Y(_16308_));
 BUFx4f_ASAP7_75t_R _22134_ (.A(_13479_),
    .Y(_16309_));
 OA211x2_ASAP7_75t_R _22135_ (.A1(_15573_),
    .A2(_16307_),
    .B(_16308_),
    .C(_16309_),
    .Y(_16310_));
 OR3x1_ASAP7_75t_R _22136_ (.A(_15498_),
    .B(_16306_),
    .C(_16310_),
    .Y(_16311_));
 INVx1_ASAP7_75t_R _22137_ (.A(_01002_),
    .Y(_16312_));
 NAND2x1_ASAP7_75t_R _22138_ (.A(_16303_),
    .B(_01000_),
    .Y(_16313_));
 OA211x2_ASAP7_75t_R _22139_ (.A1(_15573_),
    .A2(_16312_),
    .B(_16313_),
    .C(_16305_),
    .Y(_16314_));
 INVx1_ASAP7_75t_R _22140_ (.A(_01001_),
    .Y(_16315_));
 NAND2x1_ASAP7_75t_R _22141_ (.A(_16303_),
    .B(_00999_),
    .Y(_16316_));
 OA211x2_ASAP7_75t_R _22142_ (.A1(_15573_),
    .A2(_16315_),
    .B(_16316_),
    .C(_16309_),
    .Y(_16317_));
 OR3x1_ASAP7_75t_R _22143_ (.A(_15512_),
    .B(_16314_),
    .C(_16317_),
    .Y(_16318_));
 AND3x1_ASAP7_75t_R _22144_ (.A(_15607_),
    .B(_16311_),
    .C(_16318_),
    .Y(_16319_));
 OR3x2_ASAP7_75t_R _22145_ (.A(_15497_),
    .B(_16319_),
    .C(_16301_),
    .Y(_16320_));
 BUFx10_ASAP7_75t_R clone5 (.A(net15),
    .Y(net5));
 INVx1_ASAP7_75t_R _22147_ (.A(_01010_),
    .Y(_16322_));
 NAND2x1_ASAP7_75t_R _22148_ (.A(_15872_),
    .B(_01008_),
    .Y(_16323_));
 OA211x2_ASAP7_75t_R _22149_ (.A1(_15586_),
    .A2(_16322_),
    .B(_16305_),
    .C(_16323_),
    .Y(_16324_));
 INVx1_ASAP7_75t_R _22150_ (.A(_01009_),
    .Y(_16325_));
 NAND2x1_ASAP7_75t_R _22151_ (.A(_16303_),
    .B(_01007_),
    .Y(_16326_));
 OA211x2_ASAP7_75t_R _22152_ (.A1(_15573_),
    .A2(_16325_),
    .B(_16326_),
    .C(_16309_),
    .Y(_16327_));
 OR3x1_ASAP7_75t_R _22153_ (.A(_15608_),
    .B(_16327_),
    .C(_16324_),
    .Y(_16328_));
 INVx1_ASAP7_75t_R _22154_ (.A(_01018_),
    .Y(_16329_));
 NAND2x1_ASAP7_75t_R _22155_ (.A(_16303_),
    .B(_01016_),
    .Y(_16330_));
 OA211x2_ASAP7_75t_R _22156_ (.A1(_15573_),
    .A2(_16329_),
    .B(_16305_),
    .C(_16330_),
    .Y(_16331_));
 INVx1_ASAP7_75t_R _22157_ (.A(_01017_),
    .Y(_16332_));
 NAND2x1_ASAP7_75t_R _22158_ (.A(_16303_),
    .B(_01015_),
    .Y(_16333_));
 OA211x2_ASAP7_75t_R _22159_ (.A1(_15573_),
    .A2(_16332_),
    .B(_16333_),
    .C(_16309_),
    .Y(_16334_));
 OR3x1_ASAP7_75t_R _22160_ (.A(_15512_),
    .B(_16334_),
    .C(_16331_),
    .Y(_16335_));
 AND3x1_ASAP7_75t_R _22161_ (.A(_15607_),
    .B(_16335_),
    .C(_16328_),
    .Y(_16336_));
 INVx2_ASAP7_75t_R _22162_ (.A(_01011_),
    .Y(_16337_));
 NOR2x1_ASAP7_75t_R _22163_ (.A(_15505_),
    .B(_01013_),
    .Y(_16338_));
 AO21x1_ASAP7_75t_R _22164_ (.A1(_15602_),
    .A2(_16337_),
    .B(_16338_),
    .Y(_16339_));
 INVx1_ASAP7_75t_R _22165_ (.A(_01014_),
    .Y(_16340_));
 NAND2x1_ASAP7_75t_R _22166_ (.A(_15570_),
    .B(_01012_),
    .Y(_16341_));
 BUFx3_ASAP7_75t_R _22167_ (.A(_15537_),
    .Y(_16342_));
 OA211x2_ASAP7_75t_R _22168_ (.A1(_15749_),
    .A2(_16340_),
    .B(_16342_),
    .C(_16341_),
    .Y(_16343_));
 AO21x1_ASAP7_75t_R _22169_ (.A1(_15649_),
    .A2(_16339_),
    .B(_16343_),
    .Y(_16344_));
 INVx1_ASAP7_75t_R _22170_ (.A(_01006_),
    .Y(_16345_));
 NAND2x1_ASAP7_75t_R _22171_ (.A(_15891_),
    .B(_01004_),
    .Y(_16346_));
 OA211x2_ASAP7_75t_R _22172_ (.A1(_15889_),
    .A2(_16345_),
    .B(_16346_),
    .C(_15893_),
    .Y(_16347_));
 INVx1_ASAP7_75t_R _22173_ (.A(_01005_),
    .Y(_16348_));
 NAND2x1_ASAP7_75t_R _22174_ (.A(_15609_),
    .B(_01003_),
    .Y(_16349_));
 OA211x2_ASAP7_75t_R _22175_ (.A1(_15895_),
    .A2(_16348_),
    .B(_16349_),
    .C(_15899_),
    .Y(_16350_));
 OR3x1_ASAP7_75t_R _22176_ (.A(_15888_),
    .B(_16347_),
    .C(_16350_),
    .Y(_16351_));
 OA211x2_ASAP7_75t_R _22177_ (.A1(_15929_),
    .A2(_16344_),
    .B(_16351_),
    .C(_16159_),
    .Y(_16352_));
 OR3x4_ASAP7_75t_R _22178_ (.A(_15912_),
    .B(_16352_),
    .C(_16336_),
    .Y(_16353_));
 AND2x4_ASAP7_75t_R _22179_ (.A(_16353_),
    .B(_16320_),
    .Y(_16354_));
 AO21x1_ASAP7_75t_R _22180_ (.A1(_13857_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_16355_));
 AND2x2_ASAP7_75t_R _22181_ (.A(_15491_),
    .B(_16355_),
    .Y(_16356_));
 AO21x2_ASAP7_75t_R _22182_ (.A1(_15496_),
    .A2(_16354_),
    .B(_16356_),
    .Y(_18698_));
 AND2x2_ASAP7_75t_R _22183_ (.A(_13763_),
    .B(_01805_),
    .Y(_16357_));
 AO21x1_ASAP7_75t_R _22184_ (.A1(_13709_),
    .A2(_00990_),
    .B(_16357_),
    .Y(_16358_));
 OAI22x1_ASAP7_75t_R _22185_ (.A1(_00989_),
    .A2(_13948_),
    .B1(_16358_),
    .B2(_13716_),
    .Y(_16359_));
 NAND2x1_ASAP7_75t_R _22186_ (.A(_14822_),
    .B(_00996_),
    .Y(_16360_));
 OA211x2_ASAP7_75t_R _22187_ (.A1(_14778_),
    .A2(_16294_),
    .B(_16360_),
    .C(_13724_),
    .Y(_16361_));
 NAND2x1_ASAP7_75t_R _22188_ (.A(_14822_),
    .B(_00995_),
    .Y(_16362_));
 OA211x2_ASAP7_75t_R _22189_ (.A1(_13866_),
    .A2(_16297_),
    .B(_16362_),
    .C(_13744_),
    .Y(_16363_));
 OR3x1_ASAP7_75t_R _22190_ (.A(_13696_),
    .B(_16361_),
    .C(_16363_),
    .Y(_16364_));
 OA211x2_ASAP7_75t_R _22191_ (.A1(_14815_),
    .A2(_16359_),
    .B(_16364_),
    .C(_13961_),
    .Y(_16365_));
 NAND2x1_ASAP7_75t_R _22192_ (.A(_13682_),
    .B(_00992_),
    .Y(_16366_));
 OA211x2_ASAP7_75t_R _22193_ (.A1(_14945_),
    .A2(_16302_),
    .B(_16366_),
    .C(_14940_),
    .Y(_16367_));
 NAND2x1_ASAP7_75t_R _22194_ (.A(_13701_),
    .B(_00991_),
    .Y(_16368_));
 OA211x2_ASAP7_75t_R _22195_ (.A1(_13904_),
    .A2(_16307_),
    .B(_16368_),
    .C(_14867_),
    .Y(_16369_));
 OR3x1_ASAP7_75t_R _22196_ (.A(_13676_),
    .B(_16367_),
    .C(_16369_),
    .Y(_16370_));
 NAND2x1_ASAP7_75t_R _22197_ (.A(_13690_),
    .B(_01000_),
    .Y(_16371_));
 OA211x2_ASAP7_75t_R _22198_ (.A1(_14945_),
    .A2(_16312_),
    .B(_16371_),
    .C(_14940_),
    .Y(_16372_));
 NAND2x1_ASAP7_75t_R _22199_ (.A(_13742_),
    .B(_00999_),
    .Y(_16373_));
 OA211x2_ASAP7_75t_R _22200_ (.A1(_13882_),
    .A2(_16315_),
    .B(_16373_),
    .C(_13693_),
    .Y(_16374_));
 OR3x1_ASAP7_75t_R _22201_ (.A(_13696_),
    .B(_16372_),
    .C(_16374_),
    .Y(_16375_));
 AND3x1_ASAP7_75t_R _22202_ (.A(_13674_),
    .B(_16370_),
    .C(_16375_),
    .Y(_16376_));
 OR3x4_ASAP7_75t_R _22203_ (.A(_13670_),
    .B(_16365_),
    .C(_16376_),
    .Y(_16377_));
 NAND2x1_ASAP7_75t_R _22204_ (.A(_13682_),
    .B(_01008_),
    .Y(_16378_));
 OA211x2_ASAP7_75t_R _22205_ (.A1(_15019_),
    .A2(_16322_),
    .B(_16378_),
    .C(_14940_),
    .Y(_16379_));
 NAND2x1_ASAP7_75t_R _22206_ (.A(_13690_),
    .B(_01007_),
    .Y(_16380_));
 OA211x2_ASAP7_75t_R _22207_ (.A1(_14945_),
    .A2(_16325_),
    .B(_16380_),
    .C(_14867_),
    .Y(_16381_));
 OR3x1_ASAP7_75t_R _22208_ (.A(_13676_),
    .B(_16379_),
    .C(_16381_),
    .Y(_16382_));
 NAND2x1_ASAP7_75t_R _22209_ (.A(_13682_),
    .B(_01016_),
    .Y(_16383_));
 OA211x2_ASAP7_75t_R _22210_ (.A1(_14938_),
    .A2(_16329_),
    .B(_16383_),
    .C(_14940_),
    .Y(_16384_));
 NAND2x1_ASAP7_75t_R _22211_ (.A(_13690_),
    .B(_01015_),
    .Y(_16385_));
 OA211x2_ASAP7_75t_R _22212_ (.A1(_13904_),
    .A2(_16332_),
    .B(_16385_),
    .C(_14867_),
    .Y(_16386_));
 OR3x1_ASAP7_75t_R _22213_ (.A(_14853_),
    .B(_16384_),
    .C(_16386_),
    .Y(_16387_));
 AND3x1_ASAP7_75t_R _22214_ (.A(_14843_),
    .B(_16382_),
    .C(_16387_),
    .Y(_16388_));
 NOR2x1_ASAP7_75t_R _22215_ (.A(_14993_),
    .B(_01013_),
    .Y(_16389_));
 AO21x1_ASAP7_75t_R _22216_ (.A1(_13930_),
    .A2(_16337_),
    .B(_16389_),
    .Y(_16390_));
 NAND2x1_ASAP7_75t_R _22217_ (.A(_13756_),
    .B(_01012_),
    .Y(_16391_));
 OA211x2_ASAP7_75t_R _22218_ (.A1(_14844_),
    .A2(_16340_),
    .B(_16391_),
    .C(_14846_),
    .Y(_16392_));
 AO21x1_ASAP7_75t_R _22219_ (.A1(_13749_),
    .A2(_16390_),
    .B(_16392_),
    .Y(_16393_));
 NAND2x1_ASAP7_75t_R _22220_ (.A(_14822_),
    .B(_01004_),
    .Y(_16394_));
 OA211x2_ASAP7_75t_R _22221_ (.A1(_13866_),
    .A2(_16345_),
    .B(_16394_),
    .C(_13724_),
    .Y(_16395_));
 NAND2x1_ASAP7_75t_R _22222_ (.A(_13722_),
    .B(_01003_),
    .Y(_16396_));
 OA211x2_ASAP7_75t_R _22223_ (.A1(_13872_),
    .A2(_16348_),
    .B(_16396_),
    .C(_13728_),
    .Y(_16397_));
 OR3x1_ASAP7_75t_R _22224_ (.A(_13706_),
    .B(_16395_),
    .C(_16397_),
    .Y(_16398_));
 OA211x2_ASAP7_75t_R _22225_ (.A1(_13748_),
    .A2(_16393_),
    .B(_16398_),
    .C(_13961_),
    .Y(_16399_));
 OR3x4_ASAP7_75t_R _22226_ (.A(_14842_),
    .B(_16388_),
    .C(_16399_),
    .Y(_16400_));
 INVx1_ASAP7_75t_R _22227_ (.A(_00053_),
    .Y(_16401_));
 OA211x2_ASAP7_75t_R _22228_ (.A1(_13647_),
    .A2(_13658_),
    .B(_16401_),
    .C(_13366_),
    .Y(_16402_));
 AO31x2_ASAP7_75t_R _22229_ (.A1(_13947_),
    .A2(_16377_),
    .A3(_16400_),
    .B(_16402_),
    .Y(_16403_));
 INVx1_ASAP7_75t_R _22230_ (.A(_01534_),
    .Y(_16404_));
 AO32x1_ASAP7_75t_R _22231_ (.A1(_13771_),
    .A2(_13772_),
    .A3(_16403_),
    .B1(_13642_),
    .B2(_16404_),
    .Y(_16405_));
 BUFx6f_ASAP7_75t_R _22232_ (.A(_16405_),
    .Y(_18697_));
 INVx3_ASAP7_75t_R _22233_ (.A(_18697_),
    .Y(_18699_));
 AND2x2_ASAP7_75t_R _22234_ (.A(_16046_),
    .B(_01804_),
    .Y(_16406_));
 AO21x1_ASAP7_75t_R _22235_ (.A1(_15502_),
    .A2(_01023_),
    .B(_16406_),
    .Y(_16407_));
 OAI22x1_ASAP7_75t_R _22236_ (.A1(_01022_),
    .A2(_15500_),
    .B1(_16407_),
    .B2(_15569_),
    .Y(_16408_));
 INVx1_ASAP7_75t_R _22237_ (.A(_01031_),
    .Y(_16409_));
 NAND2x1_ASAP7_75t_R _22238_ (.A(_15576_),
    .B(_01029_),
    .Y(_16410_));
 OA211x2_ASAP7_75t_R _22239_ (.A1(_16161_),
    .A2(_16409_),
    .B(_16410_),
    .C(_15807_),
    .Y(_16411_));
 INVx1_ASAP7_75t_R _22240_ (.A(_01030_),
    .Y(_16412_));
 NAND2x1_ASAP7_75t_R _22241_ (.A(_15936_),
    .B(_01028_),
    .Y(_16413_));
 OA211x2_ASAP7_75t_R _22242_ (.A1(_15505_),
    .A2(_16412_),
    .B(_16413_),
    .C(_15811_),
    .Y(_16414_));
 OR3x1_ASAP7_75t_R _22243_ (.A(_15567_),
    .B(_16411_),
    .C(_16414_),
    .Y(_16415_));
 OA211x2_ASAP7_75t_R _22244_ (.A1(_15499_),
    .A2(_16408_),
    .B(_16415_),
    .C(_16159_),
    .Y(_16416_));
 INVx1_ASAP7_75t_R _22245_ (.A(_01027_),
    .Y(_16417_));
 NAND2x1_ASAP7_75t_R _22246_ (.A(_15570_),
    .B(_01025_),
    .Y(_16418_));
 OA211x2_ASAP7_75t_R _22247_ (.A1(_15749_),
    .A2(_16417_),
    .B(_16418_),
    .C(net22),
    .Y(_16419_));
 BUFx4f_ASAP7_75t_R _22248_ (.A(_15748_),
    .Y(_16420_));
 INVx1_ASAP7_75t_R _22249_ (.A(_01026_),
    .Y(_16421_));
 BUFx6f_ASAP7_75t_R _22250_ (.A(_15534_),
    .Y(_16422_));
 NAND2x1_ASAP7_75t_R _22251_ (.A(_16422_),
    .B(_01024_),
    .Y(_16423_));
 OA211x2_ASAP7_75t_R _22252_ (.A1(_16420_),
    .A2(_16421_),
    .B(_16423_),
    .C(_15619_),
    .Y(_16424_));
 OR3x1_ASAP7_75t_R _22253_ (.A(_15608_),
    .B(_16419_),
    .C(_16424_),
    .Y(_16425_));
 INVx1_ASAP7_75t_R _22254_ (.A(_01035_),
    .Y(_16426_));
 NAND2x1_ASAP7_75t_R _22255_ (.A(_15570_),
    .B(_01033_),
    .Y(_16427_));
 OA211x2_ASAP7_75t_R _22256_ (.A1(_15749_),
    .A2(_16426_),
    .B(_16427_),
    .C(net22),
    .Y(_16428_));
 INVx1_ASAP7_75t_R _22257_ (.A(_01034_),
    .Y(_16429_));
 NAND2x1_ASAP7_75t_R _22258_ (.A(_16422_),
    .B(_01032_),
    .Y(_16430_));
 OA211x2_ASAP7_75t_R _22259_ (.A1(_16420_),
    .A2(_16429_),
    .B(_16430_),
    .C(_15619_),
    .Y(_16431_));
 OR3x1_ASAP7_75t_R _22260_ (.A(_15547_),
    .B(_16428_),
    .C(_16431_),
    .Y(_16432_));
 AND3x1_ASAP7_75t_R _22261_ (.A(_15607_),
    .B(_16432_),
    .C(_16425_),
    .Y(_16433_));
 OR3x2_ASAP7_75t_R _22262_ (.A(_15497_),
    .B(_16433_),
    .C(_16416_),
    .Y(_16434_));
 INVx1_ASAP7_75t_R _22263_ (.A(_01043_),
    .Y(_16435_));
 NAND2x1_ASAP7_75t_R _22264_ (.A(_15570_),
    .B(_01041_),
    .Y(_16436_));
 OA211x2_ASAP7_75t_R _22265_ (.A1(_15749_),
    .A2(_16435_),
    .B(_16436_),
    .C(_16342_),
    .Y(_16437_));
 INVx2_ASAP7_75t_R _22266_ (.A(_01042_),
    .Y(_16438_));
 NAND2x1_ASAP7_75t_R _22267_ (.A(_15570_),
    .B(_01040_),
    .Y(_16439_));
 OA211x2_ASAP7_75t_R _22268_ (.A1(_15749_),
    .A2(_16438_),
    .B(_16439_),
    .C(_15619_),
    .Y(_16440_));
 OR3x1_ASAP7_75t_R _22269_ (.A(_15608_),
    .B(_16437_),
    .C(_16440_),
    .Y(_16441_));
 INVx2_ASAP7_75t_R _22270_ (.A(_01051_),
    .Y(_16442_));
 NAND2x1_ASAP7_75t_R _22271_ (.A(_15570_),
    .B(_01049_),
    .Y(_16443_));
 OA211x2_ASAP7_75t_R _22272_ (.A1(_15749_),
    .A2(_16442_),
    .B(_16443_),
    .C(_16342_),
    .Y(_16444_));
 INVx2_ASAP7_75t_R _22273_ (.A(_01050_),
    .Y(_16445_));
 NAND2x1_ASAP7_75t_R _22274_ (.A(_16422_),
    .B(_01048_),
    .Y(_16446_));
 OA211x2_ASAP7_75t_R _22275_ (.A1(_16420_),
    .A2(_16445_),
    .B(_16446_),
    .C(_15619_),
    .Y(_16447_));
 OR3x1_ASAP7_75t_R _22276_ (.A(_15547_),
    .B(_16444_),
    .C(_16447_),
    .Y(_16448_));
 AND3x1_ASAP7_75t_R _22277_ (.A(_15607_),
    .B(_16441_),
    .C(_16448_),
    .Y(_16449_));
 INVx1_ASAP7_75t_R _22278_ (.A(_01044_),
    .Y(_16450_));
 NOR2x1_ASAP7_75t_R _22279_ (.A(net5),
    .B(_01046_),
    .Y(_16451_));
 AO21x1_ASAP7_75t_R _22280_ (.A1(_15602_),
    .A2(_16450_),
    .B(_16451_),
    .Y(_16452_));
 INVx1_ASAP7_75t_R _22281_ (.A(_01047_),
    .Y(_16453_));
 NAND2x1_ASAP7_75t_R _22282_ (.A(_15627_),
    .B(_01045_),
    .Y(_16454_));
 OA211x2_ASAP7_75t_R _22283_ (.A1(_15625_),
    .A2(_16453_),
    .B(_16454_),
    .C(_15614_),
    .Y(_16455_));
 AO21x1_ASAP7_75t_R _22284_ (.A1(_15649_),
    .A2(_16452_),
    .B(_16455_),
    .Y(_16456_));
 INVx1_ASAP7_75t_R _22285_ (.A(_01039_),
    .Y(_16457_));
 NAND2x1_ASAP7_75t_R _22286_ (.A(_15936_),
    .B(_01037_),
    .Y(_16458_));
 OA211x2_ASAP7_75t_R _22287_ (.A1(_15594_),
    .A2(_16457_),
    .B(_16458_),
    .C(_16082_),
    .Y(_16459_));
 INVx2_ASAP7_75t_R _22288_ (.A(_01038_),
    .Y(_16460_));
 NAND2x1_ASAP7_75t_R _22289_ (.A(_15532_),
    .B(_01036_),
    .Y(_16461_));
 OA211x2_ASAP7_75t_R _22290_ (.A1(_15594_),
    .A2(_16460_),
    .B(_16461_),
    .C(_15918_),
    .Y(_16462_));
 OR3x1_ASAP7_75t_R _22291_ (.A(_15888_),
    .B(_16459_),
    .C(_16462_),
    .Y(_16463_));
 OA211x2_ASAP7_75t_R _22292_ (.A1(_15568_),
    .A2(_16456_),
    .B(_16463_),
    .C(_16159_),
    .Y(_16464_));
 OR3x2_ASAP7_75t_R _22293_ (.A(_15555_),
    .B(_16464_),
    .C(_16449_),
    .Y(_16465_));
 AND2x4_ASAP7_75t_R _22294_ (.A(_16465_),
    .B(_16434_),
    .Y(_16466_));
 AO21x1_ASAP7_75t_R _22295_ (.A1(_14733_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_16467_));
 AND2x2_ASAP7_75t_R _22296_ (.A(_15491_),
    .B(_16467_),
    .Y(_16468_));
 AO21x2_ASAP7_75t_R _22297_ (.A1(_15496_),
    .A2(_16466_),
    .B(_16468_),
    .Y(_18703_));
 AND2x2_ASAP7_75t_R _22298_ (.A(_15061_),
    .B(_01804_),
    .Y(_16469_));
 AO21x1_ASAP7_75t_R _22299_ (.A1(_13859_),
    .A2(_01023_),
    .B(_16469_),
    .Y(_16470_));
 OAI22x1_ASAP7_75t_R _22300_ (.A1(_01022_),
    .A2(_14741_),
    .B1(_16470_),
    .B2(_13863_),
    .Y(_16471_));
 NAND2x1_ASAP7_75t_R _22301_ (.A(_14764_),
    .B(_01029_),
    .Y(_16472_));
 OA211x2_ASAP7_75t_R _22302_ (.A1(_13865_),
    .A2(_16409_),
    .B(_16472_),
    .C(_13932_),
    .Y(_16473_));
 NAND2x1_ASAP7_75t_R _22303_ (.A(_15067_),
    .B(_01028_),
    .Y(_16474_));
 OA211x2_ASAP7_75t_R _22304_ (.A1(_13930_),
    .A2(_16412_),
    .B(_16474_),
    .C(_13937_),
    .Y(_16475_));
 OR3x2_ASAP7_75t_R _22305_ (.A(_14768_),
    .B(_16473_),
    .C(_16475_),
    .Y(_16476_));
 OA211x2_ASAP7_75t_R _22306_ (.A1(_14986_),
    .A2(_16471_),
    .B(_16476_),
    .C(_13877_),
    .Y(_16477_));
 NAND2x1_ASAP7_75t_R _22307_ (.A(_13888_),
    .B(_01025_),
    .Y(_16478_));
 OA211x2_ASAP7_75t_R _22308_ (.A1(_13887_),
    .A2(_16417_),
    .B(_16478_),
    .C(_13884_),
    .Y(_16479_));
 NAND2x1_ASAP7_75t_R _22309_ (.A(_13755_),
    .B(_01024_),
    .Y(_16480_));
 OA211x2_ASAP7_75t_R _22310_ (.A1(_13895_),
    .A2(_16421_),
    .B(_16480_),
    .C(_13897_),
    .Y(_16481_));
 OR3x1_ASAP7_75t_R _22311_ (.A(_15039_),
    .B(_16479_),
    .C(_16481_),
    .Y(_16482_));
 NAND2x1_ASAP7_75t_R _22312_ (.A(_13888_),
    .B(_01033_),
    .Y(_16483_));
 OA211x2_ASAP7_75t_R _22313_ (.A1(_13887_),
    .A2(_16426_),
    .B(_16483_),
    .C(_13884_),
    .Y(_16484_));
 NAND2x1_ASAP7_75t_R _22314_ (.A(_15075_),
    .B(_01032_),
    .Y(_16485_));
 OA211x2_ASAP7_75t_R _22315_ (.A1(_15074_),
    .A2(_16429_),
    .B(_16485_),
    .C(_13897_),
    .Y(_16486_));
 OR3x1_ASAP7_75t_R _22316_ (.A(_15012_),
    .B(_16484_),
    .C(_16486_),
    .Y(_16487_));
 AND3x2_ASAP7_75t_R _22317_ (.A(_13879_),
    .B(_16482_),
    .C(_16487_),
    .Y(_16488_));
 OR3x4_ASAP7_75t_R _22318_ (.A(_14738_),
    .B(_16477_),
    .C(_16488_),
    .Y(_16489_));
 NAND2x1_ASAP7_75t_R _22319_ (.A(_13882_),
    .B(_01041_),
    .Y(_16490_));
 OA211x2_ASAP7_75t_R _22320_ (.A1(_13881_),
    .A2(_16435_),
    .B(_16490_),
    .C(_13884_),
    .Y(_16491_));
 NAND2x1_ASAP7_75t_R _22321_ (.A(_13888_),
    .B(_01040_),
    .Y(_16492_));
 OA211x2_ASAP7_75t_R _22322_ (.A1(_13887_),
    .A2(_16438_),
    .B(_16492_),
    .C(_13890_),
    .Y(_16493_));
 OR3x1_ASAP7_75t_R _22323_ (.A(_15039_),
    .B(_16491_),
    .C(_16493_),
    .Y(_16494_));
 NAND2x1_ASAP7_75t_R _22324_ (.A(_13882_),
    .B(_01049_),
    .Y(_16495_));
 OA211x2_ASAP7_75t_R _22325_ (.A1(_13881_),
    .A2(_16442_),
    .B(_16495_),
    .C(_13884_),
    .Y(_16496_));
 NAND2x1_ASAP7_75t_R _22326_ (.A(_13755_),
    .B(_01048_),
    .Y(_16497_));
 OA211x2_ASAP7_75t_R _22327_ (.A1(_13895_),
    .A2(_16445_),
    .B(_16497_),
    .C(_13890_),
    .Y(_16498_));
 OR3x1_ASAP7_75t_R _22328_ (.A(_15012_),
    .B(_16496_),
    .C(_16498_),
    .Y(_16499_));
 AND3x1_ASAP7_75t_R _22329_ (.A(_13879_),
    .B(_16494_),
    .C(_16499_),
    .Y(_16500_));
 NOR2x1_ASAP7_75t_R _22330_ (.A(_15718_),
    .B(_01046_),
    .Y(_16501_));
 AO21x1_ASAP7_75t_R _22331_ (.A1(_13920_),
    .A2(_16450_),
    .B(_16501_),
    .Y(_16502_));
 NAND2x1_ASAP7_75t_R _22332_ (.A(_14872_),
    .B(_01045_),
    .Y(_16503_));
 OA211x2_ASAP7_75t_R _22333_ (.A1(_15013_),
    .A2(_16453_),
    .B(_16503_),
    .C(_13927_),
    .Y(_16504_));
 AO21x1_ASAP7_75t_R _22334_ (.A1(_13918_),
    .A2(_16502_),
    .B(_16504_),
    .Y(_16505_));
 NAND2x1_ASAP7_75t_R _22335_ (.A(_15067_),
    .B(_01037_),
    .Y(_16506_));
 OA211x2_ASAP7_75t_R _22336_ (.A1(_13930_),
    .A2(_16457_),
    .B(_16506_),
    .C(_15305_),
    .Y(_16507_));
 NAND2x1_ASAP7_75t_R _22337_ (.A(_14816_),
    .B(_01036_),
    .Y(_16508_));
 OA211x2_ASAP7_75t_R _22338_ (.A1(_15307_),
    .A2(_16460_),
    .B(_16508_),
    .C(_15309_),
    .Y(_16509_));
 OR3x1_ASAP7_75t_R _22339_ (.A(_14760_),
    .B(_16507_),
    .C(_16509_),
    .Y(_16510_));
 OA211x2_ASAP7_75t_R _22340_ (.A1(_15318_),
    .A2(_16505_),
    .B(_16510_),
    .C(_13877_),
    .Y(_16511_));
 OR3x4_ASAP7_75t_R _22341_ (.A(_14776_),
    .B(_16500_),
    .C(_16511_),
    .Y(_16512_));
 INVx1_ASAP7_75t_R _22342_ (.A(_00054_),
    .Y(_16513_));
 OA211x2_ASAP7_75t_R _22343_ (.A1(_15114_),
    .A2(_15115_),
    .B(_16513_),
    .C(_14807_),
    .Y(_16514_));
 AO31x2_ASAP7_75t_R _22344_ (.A1(_13660_),
    .A2(_16489_),
    .A3(_16512_),
    .B(_16514_),
    .Y(_16515_));
 INVx1_ASAP7_75t_R _22345_ (.A(_01533_),
    .Y(_16516_));
 AO32x1_ASAP7_75t_R _22346_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_16515_),
    .B1(_15119_),
    .B2(_16516_),
    .Y(_16517_));
 BUFx6f_ASAP7_75t_R _22347_ (.A(_16517_),
    .Y(_18702_));
 INVx2_ASAP7_75t_R _22348_ (.A(_18702_),
    .Y(_18704_));
 BUFx3_ASAP7_75t_R _22349_ (.A(_01020_),
    .Y(_16518_));
 OA21x2_ASAP7_75t_R _22350_ (.A1(_00987_),
    .A2(_16267_),
    .B(_01021_),
    .Y(_16519_));
 OA21x2_ASAP7_75t_R _22351_ (.A1(_16518_),
    .A2(_16519_),
    .B(_01054_),
    .Y(_16520_));
 XOR2x2_ASAP7_75t_R _22352_ (.A(_01053_),
    .B(_16520_),
    .Y(\alu_adder_result_ex[19] ));
 OR2x2_ASAP7_75t_R _22353_ (.A(_00954_),
    .B(_00987_),
    .Y(_16521_));
 OR3x1_ASAP7_75t_R _22354_ (.A(_16009_),
    .B(net2028),
    .C(_16521_),
    .Y(_16522_));
 OR3x1_ASAP7_75t_R _22355_ (.A(_15471_),
    .B(_16010_),
    .C(_16522_),
    .Y(_16523_));
 NOR2x1_ASAP7_75t_R _22356_ (.A(_15266_),
    .B(_16523_),
    .Y(_16524_));
 OA31x2_ASAP7_75t_R _22357_ (.A1(net1975),
    .A2(_15262_),
    .A3(_15258_),
    .B1(_16524_),
    .Y(_16525_));
 OA21x2_ASAP7_75t_R _22358_ (.A1(_00988_),
    .A2(_00987_),
    .B(_01021_),
    .Y(_16526_));
 OA21x2_ASAP7_75t_R _22359_ (.A1(_16274_),
    .A2(_16521_),
    .B(_16526_),
    .Y(_16527_));
 AO21x2_ASAP7_75t_R _22360_ (.A1(_16021_),
    .A2(_16024_),
    .B(_16522_),
    .Y(_16528_));
 NAND2x1_ASAP7_75t_R _22361_ (.A(_16527_),
    .B(_16528_),
    .Y(_16529_));
 AO21x1_ASAP7_75t_R _22362_ (.A1(_15260_),
    .A2(_16525_),
    .B(_16529_),
    .Y(_16530_));
 XOR2x2_ASAP7_75t_R _22363_ (.A(_16518_),
    .B(_16530_),
    .Y(_16531_));
 INVx4_ASAP7_75t_R _22364_ (.A(_16531_),
    .Y(\alu_adder_result_ex[18] ));
 BUFx6f_ASAP7_75t_R _22365_ (.A(_15496_),
    .Y(_16532_));
 AND2x2_ASAP7_75t_R _22366_ (.A(_15586_),
    .B(_01802_),
    .Y(_16533_));
 AO21x1_ASAP7_75t_R _22367_ (.A1(_15502_),
    .A2(_01056_),
    .B(_16533_),
    .Y(_16534_));
 OAI22x1_ASAP7_75t_R _22368_ (.A1(_01055_),
    .A2(_15500_),
    .B1(_16534_),
    .B2(_15510_),
    .Y(_16535_));
 INVx1_ASAP7_75t_R _22369_ (.A(_01064_),
    .Y(_16536_));
 NAND2x1_ASAP7_75t_R _22370_ (.A(_16046_),
    .B(_01062_),
    .Y(_16537_));
 OA211x2_ASAP7_75t_R _22371_ (.A1(_15602_),
    .A2(_16536_),
    .B(_16537_),
    .C(_15758_),
    .Y(_16538_));
 INVx1_ASAP7_75t_R _22372_ (.A(_01063_),
    .Y(_16539_));
 BUFx6f_ASAP7_75t_R _22373_ (.A(_15541_),
    .Y(_16540_));
 NAND2x1_ASAP7_75t_R _22374_ (.A(_16540_),
    .B(_01061_),
    .Y(_16541_));
 OA211x2_ASAP7_75t_R _22375_ (.A1(_15602_),
    .A2(_16539_),
    .B(_16541_),
    .C(_15509_),
    .Y(_16542_));
 OR3x1_ASAP7_75t_R _22376_ (.A(_15753_),
    .B(_16538_),
    .C(_16542_),
    .Y(_16543_));
 OA21x2_ASAP7_75t_R _22377_ (.A1(_15499_),
    .A2(_16535_),
    .B(_16543_),
    .Y(_16544_));
 INVx1_ASAP7_75t_R _22378_ (.A(_01060_),
    .Y(_16545_));
 NAND2x1_ASAP7_75t_R _22379_ (.A(_16149_),
    .B(_01058_),
    .Y(_16546_));
 OA211x2_ASAP7_75t_R _22380_ (.A1(_15577_),
    .A2(_16545_),
    .B(_16546_),
    .C(_15581_),
    .Y(_16547_));
 INVx1_ASAP7_75t_R _22381_ (.A(_01059_),
    .Y(_16548_));
 NAND2x1_ASAP7_75t_R _22382_ (.A(_15656_),
    .B(_01057_),
    .Y(_16549_));
 OA211x2_ASAP7_75t_R _22383_ (.A1(_15533_),
    .A2(_16548_),
    .B(_16549_),
    .C(_15648_),
    .Y(_16550_));
 OR3x1_ASAP7_75t_R _22384_ (.A(_15531_),
    .B(_16547_),
    .C(_16550_),
    .Y(_16551_));
 INVx1_ASAP7_75t_R _22385_ (.A(_01068_),
    .Y(_16552_));
 NAND2x1_ASAP7_75t_R _22386_ (.A(_15656_),
    .B(_01066_),
    .Y(_16553_));
 OA211x2_ASAP7_75t_R _22387_ (.A1(_15577_),
    .A2(_16552_),
    .B(_16553_),
    .C(_15538_),
    .Y(_16554_));
 INVx1_ASAP7_75t_R _22388_ (.A(_01067_),
    .Y(_16555_));
 NAND2x1_ASAP7_75t_R _22389_ (.A(_15656_),
    .B(_01065_),
    .Y(_16556_));
 OA211x2_ASAP7_75t_R _22390_ (.A1(_15533_),
    .A2(_16555_),
    .B(_16556_),
    .C(_15648_),
    .Y(_16557_));
 OR3x1_ASAP7_75t_R _22391_ (.A(_15753_),
    .B(_16554_),
    .C(_16557_),
    .Y(_16558_));
 AND3x1_ASAP7_75t_R _22392_ (.A(_15529_),
    .B(_16551_),
    .C(_16558_),
    .Y(_16559_));
 AO21x1_ASAP7_75t_R _22393_ (.A1(_15747_),
    .A2(_16544_),
    .B(_16559_),
    .Y(_16560_));
 INVx1_ASAP7_75t_R _22394_ (.A(_01076_),
    .Y(_16561_));
 NAND2x1_ASAP7_75t_R _22395_ (.A(_16422_),
    .B(_01074_),
    .Y(_16562_));
 OA211x2_ASAP7_75t_R _22396_ (.A1(_16420_),
    .A2(_16561_),
    .B(_16562_),
    .C(_16342_),
    .Y(_16563_));
 INVx1_ASAP7_75t_R _22397_ (.A(_01075_),
    .Y(_16564_));
 NAND2x1_ASAP7_75t_R _22398_ (.A(_15872_),
    .B(_01073_),
    .Y(_16565_));
 OA211x2_ASAP7_75t_R _22399_ (.A1(_15586_),
    .A2(_16564_),
    .B(_16565_),
    .C(_16309_),
    .Y(_16566_));
 OR3x1_ASAP7_75t_R _22400_ (.A(_15608_),
    .B(_16563_),
    .C(_16566_),
    .Y(_16567_));
 INVx1_ASAP7_75t_R _22401_ (.A(_01084_),
    .Y(_16568_));
 NAND2x1_ASAP7_75t_R _22402_ (.A(_16422_),
    .B(_01082_),
    .Y(_16569_));
 OA211x2_ASAP7_75t_R _22403_ (.A1(_16420_),
    .A2(_16568_),
    .B(_16569_),
    .C(_16342_),
    .Y(_16570_));
 INVx1_ASAP7_75t_R _22404_ (.A(_01083_),
    .Y(_16571_));
 NAND2x1_ASAP7_75t_R _22405_ (.A(_15872_),
    .B(_01081_),
    .Y(_16572_));
 OA211x2_ASAP7_75t_R _22406_ (.A1(_15586_),
    .A2(_16571_),
    .B(_16572_),
    .C(_16309_),
    .Y(_16573_));
 OR3x1_ASAP7_75t_R _22407_ (.A(_15512_),
    .B(_16570_),
    .C(_16573_),
    .Y(_16574_));
 AND3x1_ASAP7_75t_R _22408_ (.A(_15607_),
    .B(_16567_),
    .C(_16574_),
    .Y(_16575_));
 INVx1_ASAP7_75t_R _22409_ (.A(_01077_),
    .Y(_16576_));
 NOR2x1_ASAP7_75t_R _22410_ (.A(_16161_),
    .B(_01079_),
    .Y(_16577_));
 AO21x1_ASAP7_75t_R _22411_ (.A1(_15602_),
    .A2(_16576_),
    .B(_16577_),
    .Y(_16578_));
 INVx1_ASAP7_75t_R _22412_ (.A(_01080_),
    .Y(_16579_));
 NAND2x1_ASAP7_75t_R _22413_ (.A(_16036_),
    .B(_01078_),
    .Y(_16580_));
 OA211x2_ASAP7_75t_R _22414_ (.A1(_15749_),
    .A2(_16579_),
    .B(_16580_),
    .C(_15614_),
    .Y(_16581_));
 AO21x1_ASAP7_75t_R _22415_ (.A1(_15649_),
    .A2(_16578_),
    .B(_16581_),
    .Y(_16582_));
 INVx1_ASAP7_75t_R _22416_ (.A(_01072_),
    .Y(_16583_));
 NAND2x1_ASAP7_75t_R _22417_ (.A(_15532_),
    .B(_01070_),
    .Y(_16584_));
 OA211x2_ASAP7_75t_R _22418_ (.A1(_16079_),
    .A2(_16583_),
    .B(_16584_),
    .C(_16082_),
    .Y(_16585_));
 INVx1_ASAP7_75t_R _22419_ (.A(_01071_),
    .Y(_16586_));
 NAND2x1_ASAP7_75t_R _22420_ (.A(_15532_),
    .B(_01069_),
    .Y(_16587_));
 OA211x2_ASAP7_75t_R _22421_ (.A1(_16079_),
    .A2(_16586_),
    .B(_16587_),
    .C(_15918_),
    .Y(_16588_));
 OR3x1_ASAP7_75t_R _22422_ (.A(_15888_),
    .B(_16585_),
    .C(_16588_),
    .Y(_16589_));
 OA211x2_ASAP7_75t_R _22423_ (.A1(_15568_),
    .A2(_16582_),
    .B(_16589_),
    .C(_16159_),
    .Y(_16590_));
 OR3x1_ASAP7_75t_R _22424_ (.A(_15555_),
    .B(_16575_),
    .C(_16590_),
    .Y(_16591_));
 OAI21x1_ASAP7_75t_R _22425_ (.A1(_15745_),
    .A2(_16560_),
    .B(_16591_),
    .Y(_16592_));
 NAND2x2_ASAP7_75t_R _22426_ (.A(_14309_),
    .B(_13435_),
    .Y(_16593_));
 BUFx4f_ASAP7_75t_R _22427_ (.A(_16593_),
    .Y(_16594_));
 AO21x1_ASAP7_75t_R _22428_ (.A1(_14312_),
    .A2(_14313_),
    .B(_13576_),
    .Y(_16595_));
 BUFx3_ASAP7_75t_R _22429_ (.A(_16595_),
    .Y(_16596_));
 OA211x2_ASAP7_75t_R _22430_ (.A1(_15510_),
    .A2(_16594_),
    .B(_15491_),
    .C(_16596_),
    .Y(_16597_));
 AOI21x1_ASAP7_75t_R _22431_ (.A1(_16532_),
    .A2(_16592_),
    .B(_16597_),
    .Y(_18708_));
 AND2x2_ASAP7_75t_R _22432_ (.A(_14945_),
    .B(_01802_),
    .Y(_16598_));
 AO21x1_ASAP7_75t_R _22433_ (.A1(_14742_),
    .A2(_01056_),
    .B(_16598_),
    .Y(_16599_));
 OAI22x1_ASAP7_75t_R _22434_ (.A1(_01055_),
    .A2(_14741_),
    .B1(_16599_),
    .B2(_14746_),
    .Y(_16600_));
 NAND2x1_ASAP7_75t_R _22435_ (.A(_13711_),
    .B(_01062_),
    .Y(_16601_));
 OA211x2_ASAP7_75t_R _22436_ (.A1(_14831_),
    .A2(_16536_),
    .B(_16601_),
    .C(_14751_),
    .Y(_16602_));
 NAND2x1_ASAP7_75t_R _22437_ (.A(_15424_),
    .B(_01061_),
    .Y(_16603_));
 OA211x2_ASAP7_75t_R _22438_ (.A1(_14831_),
    .A2(_16539_),
    .B(_16603_),
    .C(_14754_),
    .Y(_16604_));
 OR3x1_ASAP7_75t_R _22439_ (.A(_14748_),
    .B(_16602_),
    .C(_16604_),
    .Y(_16605_));
 OA211x2_ASAP7_75t_R _22440_ (.A1(_14740_),
    .A2(_16600_),
    .B(_16605_),
    .C(_14757_),
    .Y(_16606_));
 NAND2x1_ASAP7_75t_R _22441_ (.A(_14764_),
    .B(_01058_),
    .Y(_16607_));
 OA211x2_ASAP7_75t_R _22442_ (.A1(_13871_),
    .A2(_16545_),
    .B(_16607_),
    .C(_13932_),
    .Y(_16608_));
 NAND2x1_ASAP7_75t_R _22443_ (.A(_15067_),
    .B(_01057_),
    .Y(_16609_));
 OA211x2_ASAP7_75t_R _22444_ (.A1(_13930_),
    .A2(_16548_),
    .B(_16609_),
    .C(_13937_),
    .Y(_16610_));
 OR3x1_ASAP7_75t_R _22445_ (.A(_14760_),
    .B(_16608_),
    .C(_16610_),
    .Y(_16611_));
 NAND2x1_ASAP7_75t_R _22446_ (.A(_13872_),
    .B(_01066_),
    .Y(_16612_));
 OA211x2_ASAP7_75t_R _22447_ (.A1(_13871_),
    .A2(_16552_),
    .B(_16612_),
    .C(_13932_),
    .Y(_16613_));
 NAND2x1_ASAP7_75t_R _22448_ (.A(_15067_),
    .B(_01065_),
    .Y(_16614_));
 OA211x2_ASAP7_75t_R _22449_ (.A1(_13934_),
    .A2(_16555_),
    .B(_16614_),
    .C(_13937_),
    .Y(_16615_));
 OR3x1_ASAP7_75t_R _22450_ (.A(_14768_),
    .B(_16613_),
    .C(_16615_),
    .Y(_16616_));
 AND3x1_ASAP7_75t_R _22451_ (.A(_15289_),
    .B(_16611_),
    .C(_16616_),
    .Y(_16617_));
 OR3x4_ASAP7_75t_R _22452_ (.A(_14814_),
    .B(_16606_),
    .C(_16617_),
    .Y(_16618_));
 NAND2x1_ASAP7_75t_R _22453_ (.A(_14764_),
    .B(_01074_),
    .Y(_16619_));
 OA211x2_ASAP7_75t_R _22454_ (.A1(_13865_),
    .A2(_16561_),
    .B(_16619_),
    .C(_13869_),
    .Y(_16620_));
 NAND2x1_ASAP7_75t_R _22455_ (.A(_13872_),
    .B(_01073_),
    .Y(_16621_));
 OA211x2_ASAP7_75t_R _22456_ (.A1(_13871_),
    .A2(_16564_),
    .B(_16621_),
    .C(_13874_),
    .Y(_16622_));
 OR3x1_ASAP7_75t_R _22457_ (.A(_14760_),
    .B(_16620_),
    .C(_16622_),
    .Y(_16623_));
 NAND2x1_ASAP7_75t_R _22458_ (.A(_14764_),
    .B(_01082_),
    .Y(_16624_));
 OA211x2_ASAP7_75t_R _22459_ (.A1(_13865_),
    .A2(_16568_),
    .B(_16624_),
    .C(_13932_),
    .Y(_16625_));
 NAND2x1_ASAP7_75t_R _22460_ (.A(_15067_),
    .B(_01081_),
    .Y(_16626_));
 OA211x2_ASAP7_75t_R _22461_ (.A1(_13930_),
    .A2(_16571_),
    .B(_16626_),
    .C(_13937_),
    .Y(_16627_));
 OR3x1_ASAP7_75t_R _22462_ (.A(_14768_),
    .B(_16625_),
    .C(_16627_),
    .Y(_16628_));
 AND3x1_ASAP7_75t_R _22463_ (.A(_15289_),
    .B(_16623_),
    .C(_16628_),
    .Y(_16629_));
 NOR2x1_ASAP7_75t_R _22464_ (.A(_15967_),
    .B(_01079_),
    .Y(_16630_));
 AO21x1_ASAP7_75t_R _22465_ (.A1(_15712_),
    .A2(_16576_),
    .B(_16630_),
    .Y(_16631_));
 NAND2x1_ASAP7_75t_R _22466_ (.A(_13751_),
    .B(_01078_),
    .Y(_16632_));
 OA211x2_ASAP7_75t_R _22467_ (.A1(_13921_),
    .A2(_16579_),
    .B(_16632_),
    .C(_14780_),
    .Y(_16633_));
 AO21x1_ASAP7_75t_R _22468_ (.A1(_13716_),
    .A2(_16631_),
    .B(_16633_),
    .Y(_16634_));
 NAND2x1_ASAP7_75t_R _22469_ (.A(_15424_),
    .B(_01070_),
    .Y(_16635_));
 OA211x2_ASAP7_75t_R _22470_ (.A1(_15423_),
    .A2(_16583_),
    .B(_16635_),
    .C(_15282_),
    .Y(_16636_));
 NAND2x1_ASAP7_75t_R _22471_ (.A(_15280_),
    .B(_01069_),
    .Y(_16637_));
 OA211x2_ASAP7_75t_R _22472_ (.A1(_15423_),
    .A2(_16586_),
    .B(_16637_),
    .C(_14850_),
    .Y(_16638_));
 OR3x1_ASAP7_75t_R _22473_ (.A(_14739_),
    .B(_16636_),
    .C(_16638_),
    .Y(_16639_));
 OA211x2_ASAP7_75t_R _22474_ (.A1(_15318_),
    .A2(_16634_),
    .B(_16639_),
    .C(_14863_),
    .Y(_16640_));
 OR3x4_ASAP7_75t_R _22475_ (.A(_14776_),
    .B(_16629_),
    .C(_16640_),
    .Y(_16641_));
 INVx1_ASAP7_75t_R _22476_ (.A(_00055_),
    .Y(_16642_));
 OA211x2_ASAP7_75t_R _22477_ (.A1(_14804_),
    .A2(_14805_),
    .B(_16642_),
    .C(_15334_),
    .Y(_16643_));
 AO31x2_ASAP7_75t_R _22478_ (.A1(_14737_),
    .A2(_16618_),
    .A3(_16641_),
    .B(_16643_),
    .Y(_16644_));
 INVx1_ASAP7_75t_R _22479_ (.A(_01531_),
    .Y(_16645_));
 AO32x1_ASAP7_75t_R _22480_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_16644_),
    .B1(_15337_),
    .B2(_16645_),
    .Y(_16646_));
 BUFx6f_ASAP7_75t_R _22481_ (.A(_16646_),
    .Y(_18707_));
 INVx1_ASAP7_75t_R _22482_ (.A(_18707_),
    .Y(_18709_));
 AND2x2_ASAP7_75t_R _22483_ (.A(_15571_),
    .B(_01801_),
    .Y(_16647_));
 AO21x1_ASAP7_75t_R _22484_ (.A1(_15502_),
    .A2(_01089_),
    .B(_16647_),
    .Y(_16648_));
 OAI22x1_ASAP7_75t_R _22485_ (.A1(_01088_),
    .A2(_15500_),
    .B1(_16648_),
    .B2(_15510_),
    .Y(_16649_));
 BUFx10_ASAP7_75t_R _22486_ (.A(_15579_),
    .Y(_16650_));
 INVx1_ASAP7_75t_R _22487_ (.A(_01097_),
    .Y(_16651_));
 NAND2x1_ASAP7_75t_R _22488_ (.A(_15625_),
    .B(_01095_),
    .Y(_16652_));
 OA211x2_ASAP7_75t_R _22489_ (.A1(_16650_),
    .A2(_16651_),
    .B(_16652_),
    .C(net19),
    .Y(_16653_));
 INVx1_ASAP7_75t_R _22490_ (.A(_01096_),
    .Y(_16654_));
 NAND2x1_ASAP7_75t_R _22491_ (.A(_15625_),
    .B(_01094_),
    .Y(_16655_));
 OA211x2_ASAP7_75t_R _22492_ (.A1(_16650_),
    .A2(_16654_),
    .B(_16655_),
    .C(_15509_),
    .Y(_16656_));
 OR3x1_ASAP7_75t_R _22493_ (.A(_15929_),
    .B(_16653_),
    .C(_16656_),
    .Y(_16657_));
 OA21x2_ASAP7_75t_R _22494_ (.A1(_15499_),
    .A2(_16649_),
    .B(_16657_),
    .Y(_16658_));
 INVx1_ASAP7_75t_R _22495_ (.A(_01093_),
    .Y(_16659_));
 NAND2x1_ASAP7_75t_R _22496_ (.A(_15586_),
    .B(_01091_),
    .Y(_16660_));
 OA211x2_ASAP7_75t_R _22497_ (.A1(_16650_),
    .A2(_16659_),
    .B(_16660_),
    .C(net19),
    .Y(_16661_));
 INVx1_ASAP7_75t_R _22498_ (.A(_01092_),
    .Y(_16662_));
 NAND2x1_ASAP7_75t_R _22499_ (.A(_15586_),
    .B(_01090_),
    .Y(_16663_));
 OA211x2_ASAP7_75t_R _22500_ (.A1(_16650_),
    .A2(_16662_),
    .B(_16663_),
    .C(_15509_),
    .Y(_16664_));
 OR3x1_ASAP7_75t_R _22501_ (.A(_15870_),
    .B(_16661_),
    .C(_16664_),
    .Y(_16665_));
 INVx1_ASAP7_75t_R _22502_ (.A(_01101_),
    .Y(_16666_));
 NAND2x1_ASAP7_75t_R _22503_ (.A(_15586_),
    .B(_01099_),
    .Y(_16667_));
 OA211x2_ASAP7_75t_R _22504_ (.A1(_16650_),
    .A2(_16666_),
    .B(_16667_),
    .C(_15758_),
    .Y(_16668_));
 INVx1_ASAP7_75t_R _22505_ (.A(_01100_),
    .Y(_16669_));
 NAND2x1_ASAP7_75t_R _22506_ (.A(_15586_),
    .B(_01098_),
    .Y(_16670_));
 OA211x2_ASAP7_75t_R _22507_ (.A1(_16650_),
    .A2(_16669_),
    .B(_16670_),
    .C(_15509_),
    .Y(_16671_));
 OR3x1_ASAP7_75t_R _22508_ (.A(_15929_),
    .B(_16668_),
    .C(_16671_),
    .Y(_16672_));
 AND3x1_ASAP7_75t_R _22509_ (.A(_15529_),
    .B(_16665_),
    .C(_16672_),
    .Y(_16673_));
 AO21x1_ASAP7_75t_R _22510_ (.A1(_15747_),
    .A2(_16658_),
    .B(_16673_),
    .Y(_16674_));
 INVx1_ASAP7_75t_R _22511_ (.A(_01109_),
    .Y(_16675_));
 NAND2x1_ASAP7_75t_R _22512_ (.A(net5),
    .B(_01107_),
    .Y(_16676_));
 OA211x2_ASAP7_75t_R _22513_ (.A1(_15571_),
    .A2(_16675_),
    .B(_16676_),
    .C(_15758_),
    .Y(_16677_));
 INVx1_ASAP7_75t_R _22514_ (.A(_01108_),
    .Y(_16678_));
 NAND2x1_ASAP7_75t_R _22515_ (.A(_16161_),
    .B(_01106_),
    .Y(_16679_));
 OA211x2_ASAP7_75t_R _22516_ (.A1(_15571_),
    .A2(_16678_),
    .B(_16679_),
    .C(_15509_),
    .Y(_16680_));
 OR3x1_ASAP7_75t_R _22517_ (.A(_15531_),
    .B(_16677_),
    .C(_16680_),
    .Y(_16681_));
 INVx1_ASAP7_75t_R _22518_ (.A(_01117_),
    .Y(_16682_));
 NAND2x1_ASAP7_75t_R _22519_ (.A(_16161_),
    .B(_01115_),
    .Y(_16683_));
 OA211x2_ASAP7_75t_R _22520_ (.A1(_15571_),
    .A2(_16682_),
    .B(_16683_),
    .C(_15758_),
    .Y(_16684_));
 INVx1_ASAP7_75t_R _22521_ (.A(_01116_),
    .Y(_16685_));
 NAND2x1_ASAP7_75t_R _22522_ (.A(_16161_),
    .B(_01114_),
    .Y(_16686_));
 OA211x2_ASAP7_75t_R _22523_ (.A1(_15571_),
    .A2(_16685_),
    .B(_16686_),
    .C(_15509_),
    .Y(_16687_));
 OR3x1_ASAP7_75t_R _22524_ (.A(_15929_),
    .B(_16684_),
    .C(_16687_),
    .Y(_16688_));
 AND3x1_ASAP7_75t_R _22525_ (.A(_15529_),
    .B(_16681_),
    .C(_16688_),
    .Y(_16689_));
 INVx2_ASAP7_75t_R _22526_ (.A(_01110_),
    .Y(_16690_));
 NOR2x1_ASAP7_75t_R _22527_ (.A(_15765_),
    .B(_01112_),
    .Y(_16691_));
 AO21x1_ASAP7_75t_R _22528_ (.A1(_16650_),
    .A2(_16690_),
    .B(_16691_),
    .Y(_16692_));
 INVx1_ASAP7_75t_R _22529_ (.A(_01113_),
    .Y(_16693_));
 NAND2x1_ASAP7_75t_R _22530_ (.A(_15513_),
    .B(_01111_),
    .Y(_16694_));
 OA211x2_ASAP7_75t_R _22531_ (.A1(_15571_),
    .A2(_16693_),
    .B(_16694_),
    .C(_15758_),
    .Y(_16695_));
 AO21x1_ASAP7_75t_R _22532_ (.A1(_15510_),
    .A2(_16692_),
    .B(_16695_),
    .Y(_16696_));
 INVx1_ASAP7_75t_R _22533_ (.A(_01105_),
    .Y(_16697_));
 NAND2x1_ASAP7_75t_R _22534_ (.A(_16149_),
    .B(_01103_),
    .Y(_16698_));
 OA211x2_ASAP7_75t_R _22535_ (.A1(_15577_),
    .A2(_16697_),
    .B(_16698_),
    .C(_15581_),
    .Y(_16699_));
 INVx2_ASAP7_75t_R _22536_ (.A(_01104_),
    .Y(_16700_));
 NAND2x1_ASAP7_75t_R _22537_ (.A(_16149_),
    .B(_01102_),
    .Y(_16701_));
 OA211x2_ASAP7_75t_R _22538_ (.A1(_15577_),
    .A2(_16700_),
    .B(_16701_),
    .C(_15648_),
    .Y(_16702_));
 OR3x1_ASAP7_75t_R _22539_ (.A(_15531_),
    .B(_16699_),
    .C(_16702_),
    .Y(_16703_));
 OA211x2_ASAP7_75t_R _22540_ (.A1(_15568_),
    .A2(_16696_),
    .B(_16703_),
    .C(_15526_),
    .Y(_16704_));
 OR3x1_ASAP7_75t_R _22541_ (.A(_15555_),
    .B(_16689_),
    .C(_16704_),
    .Y(_16705_));
 OAI21x1_ASAP7_75t_R _22542_ (.A1(_15745_),
    .A2(_16674_),
    .B(_16705_),
    .Y(_16706_));
 OA211x2_ASAP7_75t_R _22543_ (.A1(_16650_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_16707_));
 AOI21x1_ASAP7_75t_R _22544_ (.A1(_16532_),
    .A2(_16706_),
    .B(_16707_),
    .Y(_18714_));
 AND2x2_ASAP7_75t_R _22545_ (.A(_15278_),
    .B(_01801_),
    .Y(_16708_));
 AO21x1_ASAP7_75t_R _22546_ (.A1(_14742_),
    .A2(_01089_),
    .B(_16708_),
    .Y(_16709_));
 OAI22x1_ASAP7_75t_R _22547_ (.A1(_01088_),
    .A2(_14741_),
    .B1(_16709_),
    .B2(_13863_),
    .Y(_16710_));
 NAND2x1_ASAP7_75t_R _22548_ (.A(_13880_),
    .B(_01095_),
    .Y(_16711_));
 OA211x2_ASAP7_75t_R _22549_ (.A1(_15061_),
    .A2(_16651_),
    .B(_16711_),
    .C(_14751_),
    .Y(_16712_));
 NAND2x1_ASAP7_75t_R _22550_ (.A(_13886_),
    .B(_01094_),
    .Y(_16713_));
 OA211x2_ASAP7_75t_R _22551_ (.A1(_15967_),
    .A2(_16654_),
    .B(_16713_),
    .C(_14754_),
    .Y(_16714_));
 OR3x1_ASAP7_75t_R _22552_ (.A(_14748_),
    .B(_16712_),
    .C(_16714_),
    .Y(_16715_));
 OA211x2_ASAP7_75t_R _22553_ (.A1(_14740_),
    .A2(_16710_),
    .B(_16715_),
    .C(_14757_),
    .Y(_16716_));
 NAND2x1_ASAP7_75t_R _22554_ (.A(_14820_),
    .B(_01091_),
    .Y(_16717_));
 OA211x2_ASAP7_75t_R _22555_ (.A1(_15677_),
    .A2(_16659_),
    .B(_16717_),
    .C(_14995_),
    .Y(_16718_));
 NAND2x1_ASAP7_75t_R _22556_ (.A(_14993_),
    .B(_01090_),
    .Y(_16719_));
 OA211x2_ASAP7_75t_R _22557_ (.A1(_14992_),
    .A2(_16662_),
    .B(_16719_),
    .C(_15681_),
    .Y(_16720_));
 OR3x1_ASAP7_75t_R _22558_ (.A(_14777_),
    .B(_16718_),
    .C(_16720_),
    .Y(_16721_));
 NAND2x1_ASAP7_75t_R _22559_ (.A(_14993_),
    .B(_01099_),
    .Y(_16722_));
 OA211x2_ASAP7_75t_R _22560_ (.A1(_15677_),
    .A2(_16666_),
    .B(_16722_),
    .C(_14995_),
    .Y(_16723_));
 NAND2x1_ASAP7_75t_R _22561_ (.A(_13751_),
    .B(_01098_),
    .Y(_16724_));
 OA211x2_ASAP7_75t_R _22562_ (.A1(_14992_),
    .A2(_16669_),
    .B(_16724_),
    .C(_15681_),
    .Y(_16725_));
 OR3x1_ASAP7_75t_R _22563_ (.A(_13902_),
    .B(_16723_),
    .C(_16725_),
    .Y(_16726_));
 AND3x1_ASAP7_75t_R _22564_ (.A(_14759_),
    .B(_16721_),
    .C(_16726_),
    .Y(_16727_));
 OR3x4_ASAP7_75t_R _22565_ (.A(_14738_),
    .B(_16716_),
    .C(_16727_),
    .Y(_16728_));
 NAND2x1_ASAP7_75t_R _22566_ (.A(_14820_),
    .B(_01107_),
    .Y(_16729_));
 OA211x2_ASAP7_75t_R _22567_ (.A1(_15677_),
    .A2(_16675_),
    .B(_16729_),
    .C(_14995_),
    .Y(_16730_));
 NAND2x1_ASAP7_75t_R _22568_ (.A(_14993_),
    .B(_01106_),
    .Y(_16731_));
 OA211x2_ASAP7_75t_R _22569_ (.A1(_14992_),
    .A2(_16678_),
    .B(_16731_),
    .C(_15681_),
    .Y(_16732_));
 OR3x1_ASAP7_75t_R _22570_ (.A(_14777_),
    .B(_16730_),
    .C(_16732_),
    .Y(_16733_));
 NAND2x1_ASAP7_75t_R _22571_ (.A(_14820_),
    .B(_01115_),
    .Y(_16734_));
 OA211x2_ASAP7_75t_R _22572_ (.A1(_15677_),
    .A2(_16682_),
    .B(_16734_),
    .C(_14995_),
    .Y(_16735_));
 NAND2x1_ASAP7_75t_R _22573_ (.A(_13751_),
    .B(_01114_),
    .Y(_16736_));
 OA211x2_ASAP7_75t_R _22574_ (.A1(_14992_),
    .A2(_16685_),
    .B(_16736_),
    .C(_15681_),
    .Y(_16737_));
 OR3x1_ASAP7_75t_R _22575_ (.A(_13902_),
    .B(_16735_),
    .C(_16737_),
    .Y(_16738_));
 AND3x1_ASAP7_75t_R _22576_ (.A(_14759_),
    .B(_16733_),
    .C(_16738_),
    .Y(_16739_));
 NOR2x1_ASAP7_75t_R _22577_ (.A(_13860_),
    .B(_01112_),
    .Y(_16740_));
 AO21x1_ASAP7_75t_R _22578_ (.A1(_15712_),
    .A2(_16690_),
    .B(_16740_),
    .Y(_16741_));
 NAND2x1_ASAP7_75t_R _22579_ (.A(_13919_),
    .B(_01111_),
    .Y(_16742_));
 OA211x2_ASAP7_75t_R _22580_ (.A1(_15143_),
    .A2(_16693_),
    .B(_16742_),
    .C(_15141_),
    .Y(_16743_));
 AO21x1_ASAP7_75t_R _22581_ (.A1(_13918_),
    .A2(_16741_),
    .B(_16743_),
    .Y(_16744_));
 NAND2x1_ASAP7_75t_R _22582_ (.A(_13886_),
    .B(_01103_),
    .Y(_16745_));
 OA211x2_ASAP7_75t_R _22583_ (.A1(_15967_),
    .A2(_16697_),
    .B(_16745_),
    .C(_14751_),
    .Y(_16746_));
 NAND2x1_ASAP7_75t_R _22584_ (.A(_13886_),
    .B(_01102_),
    .Y(_16747_));
 OA211x2_ASAP7_75t_R _22585_ (.A1(_14749_),
    .A2(_16700_),
    .B(_16747_),
    .C(_14754_),
    .Y(_16748_));
 OR3x1_ASAP7_75t_R _22586_ (.A(_14739_),
    .B(_16746_),
    .C(_16748_),
    .Y(_16749_));
 OA211x2_ASAP7_75t_R _22587_ (.A1(_15318_),
    .A2(_16744_),
    .B(_16749_),
    .C(_14757_),
    .Y(_16750_));
 OR3x4_ASAP7_75t_R _22588_ (.A(_14776_),
    .B(_16739_),
    .C(_16750_),
    .Y(_16751_));
 INVx2_ASAP7_75t_R _22589_ (.A(_00056_),
    .Y(_16752_));
 OA211x2_ASAP7_75t_R _22590_ (.A1(_14804_),
    .A2(_14805_),
    .B(_16752_),
    .C(_15334_),
    .Y(_16753_));
 AO31x2_ASAP7_75t_R _22591_ (.A1(_13947_),
    .A2(_16728_),
    .A3(_16751_),
    .B(_16753_),
    .Y(_16754_));
 INVx1_ASAP7_75t_R _22592_ (.A(_01530_),
    .Y(_16755_));
 AO32x1_ASAP7_75t_R _22593_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_16754_),
    .B1(_15337_),
    .B2(_16755_),
    .Y(_16756_));
 BUFx6f_ASAP7_75t_R _22594_ (.A(_16756_),
    .Y(_18715_));
 INVx1_ASAP7_75t_R _22595_ (.A(_18715_),
    .Y(_18713_));
 BUFx3_ASAP7_75t_R _22596_ (.A(_01119_),
    .Y(_16757_));
 OA211x2_ASAP7_75t_R _22597_ (.A1(_01087_),
    .A2(_01086_),
    .B(_01120_),
    .C(_01054_),
    .Y(_16758_));
 OA21x2_ASAP7_75t_R _22598_ (.A1(_01021_),
    .A2(_16518_),
    .B(_16758_),
    .Y(_16759_));
 AO21x1_ASAP7_75t_R _22599_ (.A1(_00987_),
    .A2(_01021_),
    .B(_16518_),
    .Y(_16760_));
 AO21x1_ASAP7_75t_R _22600_ (.A1(_01054_),
    .A2(_16760_),
    .B(_01053_),
    .Y(_16761_));
 AND2x2_ASAP7_75t_R _22601_ (.A(_01087_),
    .B(_01120_),
    .Y(_16762_));
 AO22x1_ASAP7_75t_R _22602_ (.A1(_01086_),
    .A2(_01120_),
    .B1(_16761_),
    .B2(_16762_),
    .Y(_16763_));
 AO21x1_ASAP7_75t_R _22603_ (.A1(_16267_),
    .A2(_16759_),
    .B(_16763_),
    .Y(_16764_));
 XOR2x2_ASAP7_75t_R _22604_ (.A(_16757_),
    .B(_16764_),
    .Y(\alu_adder_result_ex[21] ));
 OA21x2_ASAP7_75t_R _22605_ (.A1(_14925_),
    .A2(_15403_),
    .B(_15408_),
    .Y(_16765_));
 OA21x2_ASAP7_75t_R _22606_ (.A1(_14922_),
    .A2(_15403_),
    .B(_16765_),
    .Y(_16766_));
 INVx1_ASAP7_75t_R _22607_ (.A(_01086_),
    .Y(_16767_));
 OR3x4_ASAP7_75t_R _22608_ (.A(_16518_),
    .B(_01053_),
    .C(_16521_),
    .Y(_16768_));
 OR3x1_ASAP7_75t_R _22609_ (.A(_16767_),
    .B(_16280_),
    .C(_16768_),
    .Y(_16769_));
 OA21x2_ASAP7_75t_R _22610_ (.A1(_16518_),
    .A2(_16526_),
    .B(_01054_),
    .Y(_16770_));
 OA21x2_ASAP7_75t_R _22611_ (.A1(_01053_),
    .A2(_16770_),
    .B(_01087_),
    .Y(_16771_));
 OAI21x1_ASAP7_75t_R _22612_ (.A1(_16277_),
    .A2(_16768_),
    .B(_16771_),
    .Y(_16772_));
 OA211x2_ASAP7_75t_R _22613_ (.A1(_16282_),
    .A2(_16768_),
    .B(_16771_),
    .C(_16767_),
    .Y(_16773_));
 AOI21x1_ASAP7_75t_R _22614_ (.A1(_01086_),
    .A2(_16772_),
    .B(_16773_),
    .Y(_16774_));
 AND4x1_ASAP7_75t_R _22615_ (.A(_16767_),
    .B(_16277_),
    .C(_16765_),
    .D(_16771_),
    .Y(_16775_));
 OAI21x1_ASAP7_75t_R _22616_ (.A1(net2003),
    .A2(_15403_),
    .B(_16775_),
    .Y(_16776_));
 OA211x2_ASAP7_75t_R _22617_ (.A1(_16766_),
    .A2(_16769_),
    .B(_16774_),
    .C(_16776_),
    .Y(_16777_));
 INVx4_ASAP7_75t_R _22618_ (.A(_16777_),
    .Y(\alu_adder_result_ex[20] ));
 AND2x2_ASAP7_75t_R _22619_ (.A(_15535_),
    .B(_01800_),
    .Y(_16778_));
 AO21x1_ASAP7_75t_R _22620_ (.A1(_15871_),
    .A2(_01122_),
    .B(_16778_),
    .Y(_16779_));
 OAI22x1_ASAP7_75t_R _22621_ (.A1(_01121_),
    .A2(_15500_),
    .B1(_16779_),
    .B2(_15569_),
    .Y(_16780_));
 INVx1_ASAP7_75t_R _22622_ (.A(_01130_),
    .Y(_16781_));
 NAND2x1_ASAP7_75t_R _22623_ (.A(_15665_),
    .B(_01128_),
    .Y(_16782_));
 OA211x2_ASAP7_75t_R _22624_ (.A1(net5),
    .A2(_16781_),
    .B(_16782_),
    .C(_15807_),
    .Y(_16783_));
 INVx2_ASAP7_75t_R _22625_ (.A(_01129_),
    .Y(_16784_));
 NAND2x1_ASAP7_75t_R _22626_ (.A(_15665_),
    .B(_01127_),
    .Y(_16785_));
 OA211x2_ASAP7_75t_R _22627_ (.A1(_16161_),
    .A2(_16784_),
    .B(_16785_),
    .C(_15811_),
    .Y(_16786_));
 OR3x1_ASAP7_75t_R _22628_ (.A(_15567_),
    .B(_16783_),
    .C(_16786_),
    .Y(_16787_));
 OA21x2_ASAP7_75t_R _22629_ (.A1(_15870_),
    .A2(_16780_),
    .B(_16787_),
    .Y(_16788_));
 INVx1_ASAP7_75t_R _22630_ (.A(_01126_),
    .Y(_16789_));
 NAND2x1_ASAP7_75t_R _22631_ (.A(_15532_),
    .B(_01124_),
    .Y(_16790_));
 OA211x2_ASAP7_75t_R _22632_ (.A1(_16079_),
    .A2(_16789_),
    .B(_16790_),
    .C(_16082_),
    .Y(_16791_));
 INVx1_ASAP7_75t_R _22633_ (.A(_01125_),
    .Y(_16792_));
 NAND2x1_ASAP7_75t_R _22634_ (.A(_15891_),
    .B(_01123_),
    .Y(_16793_));
 OA211x2_ASAP7_75t_R _22635_ (.A1(_15889_),
    .A2(_16792_),
    .B(_16793_),
    .C(_15918_),
    .Y(_16794_));
 OR3x1_ASAP7_75t_R _22636_ (.A(_15888_),
    .B(_16791_),
    .C(_16794_),
    .Y(_16795_));
 INVx1_ASAP7_75t_R _22637_ (.A(_01134_),
    .Y(_16796_));
 NAND2x1_ASAP7_75t_R _22638_ (.A(_15532_),
    .B(_01132_),
    .Y(_16797_));
 OA211x2_ASAP7_75t_R _22639_ (.A1(_16079_),
    .A2(_16796_),
    .B(_16797_),
    .C(_16082_),
    .Y(_16798_));
 INVx1_ASAP7_75t_R _22640_ (.A(_01133_),
    .Y(_16799_));
 NAND2x1_ASAP7_75t_R _22641_ (.A(_15891_),
    .B(_01131_),
    .Y(_16800_));
 OA211x2_ASAP7_75t_R _22642_ (.A1(_15889_),
    .A2(_16799_),
    .B(_16800_),
    .C(_15918_),
    .Y(_16801_));
 OR3x1_ASAP7_75t_R _22643_ (.A(_15902_),
    .B(_16798_),
    .C(_16801_),
    .Y(_16802_));
 AND3x1_ASAP7_75t_R _22644_ (.A(_15887_),
    .B(_16795_),
    .C(_16802_),
    .Y(_16803_));
 AO21x1_ASAP7_75t_R _22645_ (.A1(_15747_),
    .A2(_16788_),
    .B(_16803_),
    .Y(_16804_));
 INVx1_ASAP7_75t_R _22646_ (.A(_01142_),
    .Y(_16805_));
 NAND2x1_ASAP7_75t_R _22647_ (.A(_16151_),
    .B(_01140_),
    .Y(_16806_));
 OA211x2_ASAP7_75t_R _22648_ (.A1(_16149_),
    .A2(_16805_),
    .B(_16806_),
    .C(_16153_),
    .Y(_16807_));
 INVx1_ASAP7_75t_R _22649_ (.A(_01141_),
    .Y(_16808_));
 NAND2x1_ASAP7_75t_R _22650_ (.A(_16151_),
    .B(_01139_),
    .Y(_16809_));
 OA211x2_ASAP7_75t_R _22651_ (.A1(_15656_),
    .A2(_16808_),
    .B(_16809_),
    .C(_15883_),
    .Y(_16810_));
 OR3x1_ASAP7_75t_R _22652_ (.A(_15869_),
    .B(_16807_),
    .C(_16810_),
    .Y(_16811_));
 INVx1_ASAP7_75t_R _22653_ (.A(_01150_),
    .Y(_16812_));
 NAND2x1_ASAP7_75t_R _22654_ (.A(_16151_),
    .B(_01148_),
    .Y(_16813_));
 OA211x2_ASAP7_75t_R _22655_ (.A1(_16149_),
    .A2(_16812_),
    .B(_16813_),
    .C(_16153_),
    .Y(_16814_));
 INVx1_ASAP7_75t_R _22656_ (.A(_01149_),
    .Y(_16815_));
 NAND2x1_ASAP7_75t_R _22657_ (.A(_15572_),
    .B(_01147_),
    .Y(_16816_));
 OA211x2_ASAP7_75t_R _22658_ (.A1(_15656_),
    .A2(_16815_),
    .B(_16816_),
    .C(_15883_),
    .Y(_16817_));
 OR3x1_ASAP7_75t_R _22659_ (.A(_15876_),
    .B(_16814_),
    .C(_16817_),
    .Y(_16818_));
 AND3x1_ASAP7_75t_R _22660_ (.A(_15528_),
    .B(_16811_),
    .C(_16818_),
    .Y(_16819_));
 INVx1_ASAP7_75t_R _22661_ (.A(_01143_),
    .Y(_16820_));
 NOR2x1_ASAP7_75t_R _22662_ (.A(_15872_),
    .B(_01145_),
    .Y(_16821_));
 AO21x1_ASAP7_75t_R _22663_ (.A1(_15513_),
    .A2(_16820_),
    .B(_16821_),
    .Y(_16822_));
 INVx2_ASAP7_75t_R _22664_ (.A(_01146_),
    .Y(_16823_));
 NAND2x1_ASAP7_75t_R _22665_ (.A(_15748_),
    .B(_01144_),
    .Y(_16824_));
 OA211x2_ASAP7_75t_R _22666_ (.A1(_16540_),
    .A2(_16823_),
    .B(_16824_),
    .C(_16044_),
    .Y(_16825_));
 AO21x1_ASAP7_75t_R _22667_ (.A1(_15931_),
    .A2(_16822_),
    .B(_16825_),
    .Y(_16826_));
 INVx1_ASAP7_75t_R _22668_ (.A(_01138_),
    .Y(_16827_));
 NAND2x1_ASAP7_75t_R _22669_ (.A(net5),
    .B(_01136_),
    .Y(_16828_));
 OA211x2_ASAP7_75t_R _22670_ (.A1(_16029_),
    .A2(_16827_),
    .B(_16828_),
    .C(net18),
    .Y(_16829_));
 INVx2_ASAP7_75t_R _22671_ (.A(_01137_),
    .Y(_16830_));
 NAND2x1_ASAP7_75t_R _22672_ (.A(_15541_),
    .B(_01135_),
    .Y(_16831_));
 OA211x2_ASAP7_75t_R _22673_ (.A1(_15516_),
    .A2(_16830_),
    .B(_16831_),
    .C(_15945_),
    .Y(_16832_));
 OR3x1_ASAP7_75t_R _22674_ (.A(_15530_),
    .B(_16829_),
    .C(_16832_),
    .Y(_16833_));
 OA211x2_ASAP7_75t_R _22675_ (.A1(_15753_),
    .A2(_16826_),
    .B(_16833_),
    .C(_15746_),
    .Y(_16834_));
 OR3x1_ASAP7_75t_R _22676_ (.A(_15912_),
    .B(_16819_),
    .C(_16834_),
    .Y(_16835_));
 OAI21x1_ASAP7_75t_R _22677_ (.A1(_15745_),
    .A2(_16804_),
    .B(_16835_),
    .Y(_16836_));
 OA211x2_ASAP7_75t_R _22678_ (.A1(_15747_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_16837_));
 AOI21x1_ASAP7_75t_R _22679_ (.A1(_16532_),
    .A2(_16836_),
    .B(_16837_),
    .Y(_18718_));
 AND2x2_ASAP7_75t_R _22680_ (.A(_14854_),
    .B(_01800_),
    .Y(_16838_));
 AO21x1_ASAP7_75t_R _22681_ (.A1(_14742_),
    .A2(_01122_),
    .B(_16838_),
    .Y(_16839_));
 OAI22x1_ASAP7_75t_R _22682_ (.A1(_01121_),
    .A2(_14741_),
    .B1(_16839_),
    .B2(_14746_),
    .Y(_16840_));
 NAND2x1_ASAP7_75t_R _22683_ (.A(_13886_),
    .B(_01128_),
    .Y(_16841_));
 OA211x2_ASAP7_75t_R _22684_ (.A1(_15967_),
    .A2(_16781_),
    .B(_16841_),
    .C(_14751_),
    .Y(_16842_));
 NAND2x1_ASAP7_75t_R _22685_ (.A(_13886_),
    .B(_01127_),
    .Y(_16843_));
 OA211x2_ASAP7_75t_R _22686_ (.A1(_14749_),
    .A2(_16784_),
    .B(_16843_),
    .C(_14754_),
    .Y(_16844_));
 OR3x1_ASAP7_75t_R _22687_ (.A(_14748_),
    .B(_16842_),
    .C(_16844_),
    .Y(_16845_));
 OA211x2_ASAP7_75t_R _22688_ (.A1(_14740_),
    .A2(_16840_),
    .B(_16845_),
    .C(_14757_),
    .Y(_16846_));
 NAND2x1_ASAP7_75t_R _22689_ (.A(_15190_),
    .B(_01124_),
    .Y(_16847_));
 OA211x2_ASAP7_75t_R _22690_ (.A1(_13921_),
    .A2(_16789_),
    .B(_16847_),
    .C(_14780_),
    .Y(_16848_));
 NAND2x1_ASAP7_75t_R _22691_ (.A(_15190_),
    .B(_01123_),
    .Y(_16849_));
 OA211x2_ASAP7_75t_R _22692_ (.A1(_15718_),
    .A2(_16792_),
    .B(_16849_),
    .C(_13715_),
    .Y(_16850_));
 OR3x1_ASAP7_75t_R _22693_ (.A(_14777_),
    .B(_16848_),
    .C(_16850_),
    .Y(_16851_));
 NAND2x1_ASAP7_75t_R _22694_ (.A(_15190_),
    .B(_01132_),
    .Y(_16852_));
 OA211x2_ASAP7_75t_R _22695_ (.A1(_15718_),
    .A2(_16796_),
    .B(_16852_),
    .C(_14780_),
    .Y(_16853_));
 NAND2x1_ASAP7_75t_R _22696_ (.A(_14778_),
    .B(_01131_),
    .Y(_16854_));
 OA211x2_ASAP7_75t_R _22697_ (.A1(_15718_),
    .A2(_16799_),
    .B(_16854_),
    .C(_13874_),
    .Y(_16855_));
 OR3x1_ASAP7_75t_R _22698_ (.A(_13902_),
    .B(_16853_),
    .C(_16855_),
    .Y(_16856_));
 AND3x1_ASAP7_75t_R _22699_ (.A(_14759_),
    .B(_16851_),
    .C(_16856_),
    .Y(_16857_));
 OR3x4_ASAP7_75t_R _22700_ (.A(_14738_),
    .B(_16846_),
    .C(_16857_),
    .Y(_16858_));
 NAND2x1_ASAP7_75t_R _22701_ (.A(_13751_),
    .B(_01140_),
    .Y(_16859_));
 OA211x2_ASAP7_75t_R _22702_ (.A1(_13921_),
    .A2(_16805_),
    .B(_16859_),
    .C(_14780_),
    .Y(_16860_));
 NAND2x1_ASAP7_75t_R _22703_ (.A(_15190_),
    .B(_01139_),
    .Y(_16861_));
 OA211x2_ASAP7_75t_R _22704_ (.A1(_15718_),
    .A2(_16808_),
    .B(_16861_),
    .C(_13715_),
    .Y(_16862_));
 OR3x1_ASAP7_75t_R _22705_ (.A(_14777_),
    .B(_16860_),
    .C(_16862_),
    .Y(_16863_));
 NAND2x1_ASAP7_75t_R _22706_ (.A(_15190_),
    .B(_01148_),
    .Y(_16864_));
 OA211x2_ASAP7_75t_R _22707_ (.A1(_15718_),
    .A2(_16812_),
    .B(_16864_),
    .C(_14780_),
    .Y(_16865_));
 NAND2x1_ASAP7_75t_R _22708_ (.A(_14778_),
    .B(_01147_),
    .Y(_16866_));
 OA211x2_ASAP7_75t_R _22709_ (.A1(_15718_),
    .A2(_16815_),
    .B(_16866_),
    .C(_13715_),
    .Y(_16867_));
 OR3x1_ASAP7_75t_R _22710_ (.A(_13902_),
    .B(_16865_),
    .C(_16867_),
    .Y(_16868_));
 AND3x1_ASAP7_75t_R _22711_ (.A(_14759_),
    .B(_16863_),
    .C(_16868_),
    .Y(_16869_));
 NOR2x1_ASAP7_75t_R _22712_ (.A(_15061_),
    .B(_01145_),
    .Y(_16870_));
 AO21x1_ASAP7_75t_R _22713_ (.A1(_15712_),
    .A2(_16820_),
    .B(_16870_),
    .Y(_16871_));
 BUFx10_ASAP7_75t_R _22714_ (.A(_13699_),
    .Y(_16872_));
 NAND2x1_ASAP7_75t_R _22715_ (.A(_16872_),
    .B(_01144_),
    .Y(_16873_));
 OA211x2_ASAP7_75t_R _22716_ (.A1(_15954_),
    .A2(_16823_),
    .B(_16873_),
    .C(_14995_),
    .Y(_16874_));
 AO21x1_ASAP7_75t_R _22717_ (.A1(_13918_),
    .A2(_16871_),
    .B(_16874_),
    .Y(_16875_));
 NAND2x1_ASAP7_75t_R _22718_ (.A(_13711_),
    .B(_01136_),
    .Y(_16876_));
 OA211x2_ASAP7_75t_R _22719_ (.A1(_14749_),
    .A2(_16827_),
    .B(_16876_),
    .C(_14751_),
    .Y(_16877_));
 NAND2x1_ASAP7_75t_R _22720_ (.A(_13711_),
    .B(_01135_),
    .Y(_16878_));
 OA211x2_ASAP7_75t_R _22721_ (.A1(_14749_),
    .A2(_16830_),
    .B(_16878_),
    .C(_14754_),
    .Y(_16879_));
 OR3x1_ASAP7_75t_R _22722_ (.A(_14739_),
    .B(_16877_),
    .C(_16879_),
    .Y(_16880_));
 OA211x2_ASAP7_75t_R _22723_ (.A1(_15318_),
    .A2(_16875_),
    .B(_16880_),
    .C(_14757_),
    .Y(_16881_));
 OR3x4_ASAP7_75t_R _22724_ (.A(_14776_),
    .B(_16869_),
    .C(_16881_),
    .Y(_16882_));
 INVx2_ASAP7_75t_R _22725_ (.A(_00057_),
    .Y(_16883_));
 OA211x2_ASAP7_75t_R _22726_ (.A1(_13647_),
    .A2(_13658_),
    .B(_16883_),
    .C(_15334_),
    .Y(_16884_));
 AO31x2_ASAP7_75t_R _22727_ (.A1(_13947_),
    .A2(_16858_),
    .A3(_16882_),
    .B(_16884_),
    .Y(_16885_));
 INVx1_ASAP7_75t_R _22728_ (.A(_01529_),
    .Y(_16886_));
 AO32x1_ASAP7_75t_R _22729_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_16885_),
    .B1(_15337_),
    .B2(_16886_),
    .Y(_16887_));
 BUFx6f_ASAP7_75t_R _22730_ (.A(_16887_),
    .Y(_18717_));
 INVx3_ASAP7_75t_R _22731_ (.A(_18717_),
    .Y(_18719_));
 AND2x2_ASAP7_75t_R _22732_ (.A(_15872_),
    .B(_01799_),
    .Y(_16888_));
 AO21x1_ASAP7_75t_R _22733_ (.A1(_15871_),
    .A2(_01155_),
    .B(_16888_),
    .Y(_16889_));
 OAI22x1_ASAP7_75t_R _22734_ (.A1(_01154_),
    .A2(_15500_),
    .B1(_16889_),
    .B2(_15649_),
    .Y(_16890_));
 INVx1_ASAP7_75t_R _22735_ (.A(_01163_),
    .Y(_16891_));
 NAND2x1_ASAP7_75t_R _22736_ (.A(_15586_),
    .B(_01161_),
    .Y(_16892_));
 OA211x2_ASAP7_75t_R _22737_ (.A1(_15617_),
    .A2(_16891_),
    .B(_16892_),
    .C(_15879_),
    .Y(_16893_));
 INVx2_ASAP7_75t_R _22738_ (.A(_01162_),
    .Y(_16894_));
 NAND2x1_ASAP7_75t_R _22739_ (.A(_15586_),
    .B(_01160_),
    .Y(_16895_));
 OA211x2_ASAP7_75t_R _22740_ (.A1(_15627_),
    .A2(_16894_),
    .B(_16895_),
    .C(_15883_),
    .Y(_16896_));
 OR3x1_ASAP7_75t_R _22741_ (.A(_15876_),
    .B(_16893_),
    .C(_16896_),
    .Y(_16897_));
 OA211x2_ASAP7_75t_R _22742_ (.A1(_15870_),
    .A2(_16890_),
    .B(_16897_),
    .C(_15746_),
    .Y(_16898_));
 INVx1_ASAP7_75t_R _22743_ (.A(_01159_),
    .Y(_16899_));
 NAND2x1_ASAP7_75t_R _22744_ (.A(_15609_),
    .B(_01157_),
    .Y(_16900_));
 OA211x2_ASAP7_75t_R _22745_ (.A1(_15889_),
    .A2(_16899_),
    .B(_16900_),
    .C(_15893_),
    .Y(_16901_));
 INVx2_ASAP7_75t_R _22746_ (.A(_01158_),
    .Y(_16902_));
 NAND2x1_ASAP7_75t_R _22747_ (.A(_15897_),
    .B(_01156_),
    .Y(_16903_));
 OA211x2_ASAP7_75t_R _22748_ (.A1(_15895_),
    .A2(_16902_),
    .B(_16903_),
    .C(_15899_),
    .Y(_16904_));
 OR3x1_ASAP7_75t_R _22749_ (.A(_15888_),
    .B(_16901_),
    .C(_16904_),
    .Y(_16905_));
 INVx1_ASAP7_75t_R _22750_ (.A(_01167_),
    .Y(_16906_));
 NAND2x1_ASAP7_75t_R _22751_ (.A(_15609_),
    .B(_01165_),
    .Y(_16907_));
 OA211x2_ASAP7_75t_R _22752_ (.A1(_15895_),
    .A2(_16906_),
    .B(_16907_),
    .C(_15893_),
    .Y(_16908_));
 INVx1_ASAP7_75t_R _22753_ (.A(_01166_),
    .Y(_16909_));
 NAND2x1_ASAP7_75t_R _22754_ (.A(_15897_),
    .B(_01164_),
    .Y(_16910_));
 OA211x2_ASAP7_75t_R _22755_ (.A1(_15756_),
    .A2(_16909_),
    .B(_16910_),
    .C(_15899_),
    .Y(_16911_));
 OR3x1_ASAP7_75t_R _22756_ (.A(_15902_),
    .B(_16908_),
    .C(_16911_),
    .Y(_16912_));
 AND3x1_ASAP7_75t_R _22757_ (.A(_15528_),
    .B(_16905_),
    .C(_16912_),
    .Y(_16913_));
 OR3x4_ASAP7_75t_R _22758_ (.A(_15497_),
    .B(_16898_),
    .C(_16913_),
    .Y(_16914_));
 INVx1_ASAP7_75t_R _22759_ (.A(_01175_),
    .Y(_16915_));
 NAND2x1_ASAP7_75t_R _22760_ (.A(_15891_),
    .B(_01173_),
    .Y(_16916_));
 OA211x2_ASAP7_75t_R _22761_ (.A1(_15889_),
    .A2(_16915_),
    .B(_16916_),
    .C(_15893_),
    .Y(_16917_));
 INVx1_ASAP7_75t_R _22762_ (.A(_01174_),
    .Y(_16918_));
 NAND2x1_ASAP7_75t_R _22763_ (.A(_15609_),
    .B(_01172_),
    .Y(_16919_));
 OA211x2_ASAP7_75t_R _22764_ (.A1(_15895_),
    .A2(_16918_),
    .B(_16919_),
    .C(_15899_),
    .Y(_16920_));
 OR3x1_ASAP7_75t_R _22765_ (.A(_15888_),
    .B(_16917_),
    .C(_16920_),
    .Y(_16921_));
 INVx1_ASAP7_75t_R _22766_ (.A(_01183_),
    .Y(_16922_));
 NAND2x1_ASAP7_75t_R _22767_ (.A(_15609_),
    .B(_01181_),
    .Y(_16923_));
 OA211x2_ASAP7_75t_R _22768_ (.A1(_15889_),
    .A2(_16922_),
    .B(_16923_),
    .C(_15893_),
    .Y(_16924_));
 INVx1_ASAP7_75t_R _22769_ (.A(_01182_),
    .Y(_16925_));
 NAND2x1_ASAP7_75t_R _22770_ (.A(_15897_),
    .B(_01180_),
    .Y(_16926_));
 OA211x2_ASAP7_75t_R _22771_ (.A1(_15895_),
    .A2(_16925_),
    .B(_16926_),
    .C(_15899_),
    .Y(_16927_));
 OR3x1_ASAP7_75t_R _22772_ (.A(_15902_),
    .B(_16924_),
    .C(_16927_),
    .Y(_16928_));
 AND3x1_ASAP7_75t_R _22773_ (.A(_15887_),
    .B(_16921_),
    .C(_16928_),
    .Y(_16929_));
 INVx2_ASAP7_75t_R _22774_ (.A(_01176_),
    .Y(_16930_));
 NOR2x1_ASAP7_75t_R _22775_ (.A(_15535_),
    .B(_01178_),
    .Y(_16931_));
 AO21x1_ASAP7_75t_R _22776_ (.A1(_15625_),
    .A2(_16930_),
    .B(_16931_),
    .Y(_16932_));
 INVx1_ASAP7_75t_R _22777_ (.A(_01179_),
    .Y(_16933_));
 NAND2x1_ASAP7_75t_R _22778_ (.A(_15936_),
    .B(_01177_),
    .Y(_16934_));
 OA211x2_ASAP7_75t_R _22779_ (.A1(_15594_),
    .A2(_16933_),
    .B(_16934_),
    .C(_16082_),
    .Y(_16935_));
 AO21x1_ASAP7_75t_R _22780_ (.A1(_15931_),
    .A2(_16932_),
    .B(_16935_),
    .Y(_16936_));
 INVx1_ASAP7_75t_R _22781_ (.A(_01171_),
    .Y(_16937_));
 NAND2x1_ASAP7_75t_R _22782_ (.A(_15586_),
    .B(_01169_),
    .Y(_16938_));
 OA211x2_ASAP7_75t_R _22783_ (.A1(_15627_),
    .A2(_16937_),
    .B(_16938_),
    .C(_15879_),
    .Y(_16939_));
 INVx1_ASAP7_75t_R _22784_ (.A(_01170_),
    .Y(_16940_));
 NAND2x1_ASAP7_75t_R _22785_ (.A(_15651_),
    .B(_01168_),
    .Y(_16941_));
 OA211x2_ASAP7_75t_R _22786_ (.A1(_16036_),
    .A2(_16940_),
    .B(_16941_),
    .C(_15945_),
    .Y(_16942_));
 OR3x1_ASAP7_75t_R _22787_ (.A(_15530_),
    .B(_16939_),
    .C(_16942_),
    .Y(_16943_));
 OA211x2_ASAP7_75t_R _22788_ (.A1(_15929_),
    .A2(_16936_),
    .B(_16943_),
    .C(_15746_),
    .Y(_16944_));
 OR3x4_ASAP7_75t_R _22789_ (.A(_15912_),
    .B(_16929_),
    .C(_16944_),
    .Y(_16945_));
 AND2x4_ASAP7_75t_R _22790_ (.A(_16914_),
    .B(_16945_),
    .Y(_16946_));
 INVx1_ASAP7_75t_R _22791_ (.A(_16946_),
    .Y(_16947_));
 OA211x2_ASAP7_75t_R _22792_ (.A1(_15568_),
    .A2(_16594_),
    .B(_15491_),
    .C(_16596_),
    .Y(_16948_));
 AOI21x1_ASAP7_75t_R _22793_ (.A1(_16532_),
    .A2(_16947_),
    .B(_16948_),
    .Y(_18724_));
 AND2x2_ASAP7_75t_R _22794_ (.A(_14831_),
    .B(_01799_),
    .Y(_16949_));
 AO21x1_ASAP7_75t_R _22795_ (.A1(_13859_),
    .A2(_01155_),
    .B(_16949_),
    .Y(_16950_));
 OAI22x1_ASAP7_75t_R _22796_ (.A1(_01154_),
    .A2(_14741_),
    .B1(_16950_),
    .B2(_13863_),
    .Y(_16951_));
 NAND2x1_ASAP7_75t_R _22797_ (.A(_13880_),
    .B(_01161_),
    .Y(_16952_));
 OA211x2_ASAP7_75t_R _22798_ (.A1(_13860_),
    .A2(_16891_),
    .B(_16952_),
    .C(_14751_),
    .Y(_16953_));
 NAND2x1_ASAP7_75t_R _22799_ (.A(_13880_),
    .B(_01160_),
    .Y(_16954_));
 OA211x2_ASAP7_75t_R _22800_ (.A1(_15061_),
    .A2(_16894_),
    .B(_16954_),
    .C(_15355_),
    .Y(_16955_));
 OR3x1_ASAP7_75t_R _22801_ (.A(_14748_),
    .B(_16953_),
    .C(_16955_),
    .Y(_16956_));
 OA211x2_ASAP7_75t_R _22802_ (.A1(_14986_),
    .A2(_16951_),
    .B(_16956_),
    .C(_14757_),
    .Y(_16957_));
 NAND2x1_ASAP7_75t_R _22803_ (.A(_16872_),
    .B(_01157_),
    .Y(_16958_));
 OA211x2_ASAP7_75t_R _22804_ (.A1(_15954_),
    .A2(_16899_),
    .B(_16958_),
    .C(_15141_),
    .Y(_16959_));
 NAND2x1_ASAP7_75t_R _22805_ (.A(_16872_),
    .B(_01156_),
    .Y(_16960_));
 OA211x2_ASAP7_75t_R _22806_ (.A1(_15954_),
    .A2(_16902_),
    .B(_16960_),
    .C(_15681_),
    .Y(_16961_));
 OR3x1_ASAP7_75t_R _22807_ (.A(_14777_),
    .B(_16959_),
    .C(_16961_),
    .Y(_16962_));
 NAND2x1_ASAP7_75t_R _22808_ (.A(_16872_),
    .B(_01165_),
    .Y(_16963_));
 OA211x2_ASAP7_75t_R _22809_ (.A1(_15954_),
    .A2(_16906_),
    .B(_16963_),
    .C(_15141_),
    .Y(_16964_));
 NAND2x1_ASAP7_75t_R _22810_ (.A(_14820_),
    .B(_01164_),
    .Y(_16965_));
 OA211x2_ASAP7_75t_R _22811_ (.A1(_15677_),
    .A2(_16909_),
    .B(_16965_),
    .C(_15681_),
    .Y(_16966_));
 OR3x1_ASAP7_75t_R _22812_ (.A(_15079_),
    .B(_16964_),
    .C(_16966_),
    .Y(_16967_));
 AND3x2_ASAP7_75t_R _22813_ (.A(_14759_),
    .B(_16962_),
    .C(_16967_),
    .Y(_16968_));
 OR3x4_ASAP7_75t_R _22814_ (.A(_14738_),
    .B(_16957_),
    .C(_16968_),
    .Y(_16969_));
 NAND2x1_ASAP7_75t_R _22815_ (.A(_16872_),
    .B(_01173_),
    .Y(_16970_));
 OA211x2_ASAP7_75t_R _22816_ (.A1(_15143_),
    .A2(_16915_),
    .B(_16970_),
    .C(_15141_),
    .Y(_16971_));
 NAND2x1_ASAP7_75t_R _22817_ (.A(_16872_),
    .B(_01172_),
    .Y(_16972_));
 OA211x2_ASAP7_75t_R _22818_ (.A1(_15954_),
    .A2(_16918_),
    .B(_16972_),
    .C(_15109_),
    .Y(_16973_));
 OR3x1_ASAP7_75t_R _22819_ (.A(_13856_),
    .B(_16971_),
    .C(_16973_),
    .Y(_16974_));
 NAND2x1_ASAP7_75t_R _22820_ (.A(_16872_),
    .B(_01181_),
    .Y(_16975_));
 OA211x2_ASAP7_75t_R _22821_ (.A1(_15954_),
    .A2(_16922_),
    .B(_16975_),
    .C(_15141_),
    .Y(_16976_));
 NAND2x1_ASAP7_75t_R _22822_ (.A(_16872_),
    .B(_01180_),
    .Y(_16977_));
 OA211x2_ASAP7_75t_R _22823_ (.A1(_15954_),
    .A2(_16925_),
    .B(_16977_),
    .C(_15681_),
    .Y(_16978_));
 OR3x1_ASAP7_75t_R _22824_ (.A(_15079_),
    .B(_16976_),
    .C(_16978_),
    .Y(_16979_));
 AND3x1_ASAP7_75t_R _22825_ (.A(_14759_),
    .B(_16974_),
    .C(_16979_),
    .Y(_16980_));
 NOR2x1_ASAP7_75t_R _22826_ (.A(_15126_),
    .B(_01178_),
    .Y(_16981_));
 AO21x1_ASAP7_75t_R _22827_ (.A1(_15964_),
    .A2(_16930_),
    .B(_16981_),
    .Y(_16982_));
 NAND2x1_ASAP7_75t_R _22828_ (.A(_13689_),
    .B(_01177_),
    .Y(_16983_));
 OA211x2_ASAP7_75t_R _22829_ (.A1(_15138_),
    .A2(_16933_),
    .B(_16983_),
    .C(_15081_),
    .Y(_16984_));
 AO21x1_ASAP7_75t_R _22830_ (.A1(_13918_),
    .A2(_16982_),
    .B(_16984_),
    .Y(_16985_));
 NAND2x1_ASAP7_75t_R _22831_ (.A(_13880_),
    .B(_01169_),
    .Y(_16986_));
 OA211x2_ASAP7_75t_R _22832_ (.A1(_15061_),
    .A2(_16937_),
    .B(_16986_),
    .C(_14751_),
    .Y(_16987_));
 NAND2x1_ASAP7_75t_R _22833_ (.A(_13880_),
    .B(_01168_),
    .Y(_16988_));
 OA211x2_ASAP7_75t_R _22834_ (.A1(_15061_),
    .A2(_16940_),
    .B(_16988_),
    .C(_15355_),
    .Y(_16989_));
 OR3x1_ASAP7_75t_R _22835_ (.A(_14739_),
    .B(_16987_),
    .C(_16989_),
    .Y(_16990_));
 OA211x2_ASAP7_75t_R _22836_ (.A1(_15318_),
    .A2(_16985_),
    .B(_16990_),
    .C(_14757_),
    .Y(_16991_));
 OR3x4_ASAP7_75t_R _22837_ (.A(_14776_),
    .B(_16980_),
    .C(_16991_),
    .Y(_16992_));
 INVx1_ASAP7_75t_R _22838_ (.A(_00058_),
    .Y(_16993_));
 OA211x2_ASAP7_75t_R _22839_ (.A1(_14804_),
    .A2(_14805_),
    .B(_16993_),
    .C(_15334_),
    .Y(_16994_));
 AO31x2_ASAP7_75t_R _22840_ (.A1(_14737_),
    .A2(_16969_),
    .A3(_16992_),
    .B(_16994_),
    .Y(_16995_));
 INVx1_ASAP7_75t_R _22841_ (.A(_01528_),
    .Y(_16996_));
 AO32x1_ASAP7_75t_R _22842_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_16995_),
    .B1(_15337_),
    .B2(_16996_),
    .Y(_16997_));
 BUFx6f_ASAP7_75t_R _22843_ (.A(_16997_),
    .Y(_18725_));
 INVx1_ASAP7_75t_R _22844_ (.A(_18725_),
    .Y(_18723_));
 BUFx3_ASAP7_75t_R _22845_ (.A(_01185_),
    .Y(_16998_));
 OR2x2_ASAP7_75t_R _22846_ (.A(_16757_),
    .B(_01152_),
    .Y(_16999_));
 OA21x2_ASAP7_75t_R _22847_ (.A1(_01153_),
    .A2(_01152_),
    .B(_01186_),
    .Y(_17000_));
 OA21x2_ASAP7_75t_R _22848_ (.A1(_16764_),
    .A2(_16999_),
    .B(_17000_),
    .Y(_17001_));
 XNOR2x2_ASAP7_75t_R _22849_ (.A(_16998_),
    .B(_17001_),
    .Y(_17002_));
 CKINVDCx8_ASAP7_75t_R _22850_ (.A(_17002_),
    .Y(\alu_adder_result_ex[23] ));
 INVx2_ASAP7_75t_R _22851_ (.A(_01152_),
    .Y(_17003_));
 OA21x2_ASAP7_75t_R _22852_ (.A1(_16518_),
    .A2(_16527_),
    .B(_01054_),
    .Y(_17004_));
 OA21x2_ASAP7_75t_R _22853_ (.A1(_01053_),
    .A2(_17004_),
    .B(_01087_),
    .Y(_17005_));
 OA21x2_ASAP7_75t_R _22854_ (.A1(_01086_),
    .A2(_17005_),
    .B(_01120_),
    .Y(_17006_));
 OR4x2_ASAP7_75t_R _22855_ (.A(_16518_),
    .B(_01053_),
    .C(_01086_),
    .D(_16757_),
    .Y(_17007_));
 OR2x2_ASAP7_75t_R _22856_ (.A(_16528_),
    .B(_17007_),
    .Y(_17008_));
 OA211x2_ASAP7_75t_R _22857_ (.A1(_16757_),
    .A2(_17006_),
    .B(_17008_),
    .C(_01153_),
    .Y(_17009_));
 NAND2x1_ASAP7_75t_R _22858_ (.A(_17003_),
    .B(_17007_),
    .Y(_17010_));
 OAI21x1_ASAP7_75t_R _22859_ (.A1(_16757_),
    .A2(_17006_),
    .B(_01153_),
    .Y(_17011_));
 OAI22x1_ASAP7_75t_R _22860_ (.A1(_17003_),
    .A2(_17009_),
    .B1(_17010_),
    .B2(_17011_),
    .Y(_17012_));
 NAND2x1_ASAP7_75t_R _22861_ (.A(_17003_),
    .B(_16528_),
    .Y(_17013_));
 AOI211x1_ASAP7_75t_R _22862_ (.A1(_15260_),
    .A2(_16525_),
    .B(_17011_),
    .C(_17013_),
    .Y(_17014_));
 INVx1_ASAP7_75t_R _22863_ (.A(_17007_),
    .Y(_17015_));
 AND4x2_ASAP7_75t_R _22864_ (.A(_01152_),
    .B(_15260_),
    .C(_16525_),
    .D(_17015_),
    .Y(_17016_));
 NOR3x2_ASAP7_75t_R _22865_ (.B(_17014_),
    .C(_17016_),
    .Y(_17017_),
    .A(_17012_));
 INVx4_ASAP7_75t_R _22866_ (.A(_17017_),
    .Y(\alu_adder_result_ex[22] ));
 AND2x2_ASAP7_75t_R _22867_ (.A(_16036_),
    .B(_01798_),
    .Y(_17018_));
 AO21x1_ASAP7_75t_R _22868_ (.A1(_15871_),
    .A2(_01188_),
    .B(_17018_),
    .Y(_17019_));
 OAI22x1_ASAP7_75t_R _22869_ (.A1(_01187_),
    .A2(_15500_),
    .B1(_17019_),
    .B2(_15649_),
    .Y(_17020_));
 INVx1_ASAP7_75t_R _22870_ (.A(_01196_),
    .Y(_17021_));
 NAND2x1_ASAP7_75t_R _22871_ (.A(_15532_),
    .B(_01194_),
    .Y(_17022_));
 OA211x2_ASAP7_75t_R _22872_ (.A1(_16079_),
    .A2(_17021_),
    .B(_17022_),
    .C(_16082_),
    .Y(_17023_));
 INVx1_ASAP7_75t_R _22873_ (.A(_01195_),
    .Y(_17024_));
 NAND2x1_ASAP7_75t_R _22874_ (.A(_15891_),
    .B(_01193_),
    .Y(_17025_));
 OA211x2_ASAP7_75t_R _22875_ (.A1(_16079_),
    .A2(_17024_),
    .B(_17025_),
    .C(_15918_),
    .Y(_17026_));
 OR3x1_ASAP7_75t_R _22876_ (.A(_15567_),
    .B(_17023_),
    .C(_17026_),
    .Y(_17027_));
 OA21x2_ASAP7_75t_R _22877_ (.A1(_15870_),
    .A2(_17020_),
    .B(_17027_),
    .Y(_17028_));
 INVx1_ASAP7_75t_R _22878_ (.A(_01192_),
    .Y(_17029_));
 NAND2x1_ASAP7_75t_R _22879_ (.A(_16048_),
    .B(_01190_),
    .Y(_17030_));
 OA211x2_ASAP7_75t_R _22880_ (.A1(_16540_),
    .A2(_17029_),
    .B(_17030_),
    .C(_16044_),
    .Y(_17031_));
 INVx1_ASAP7_75t_R _22881_ (.A(_01191_),
    .Y(_17032_));
 NAND2x1_ASAP7_75t_R _22882_ (.A(_15748_),
    .B(_01189_),
    .Y(_17033_));
 OA211x2_ASAP7_75t_R _22883_ (.A1(_16540_),
    .A2(_17032_),
    .B(_17033_),
    .C(_15930_),
    .Y(_17034_));
 OR3x1_ASAP7_75t_R _22884_ (.A(_15869_),
    .B(_17031_),
    .C(_17034_),
    .Y(_17035_));
 INVx1_ASAP7_75t_R _22885_ (.A(_01200_),
    .Y(_17036_));
 NAND2x1_ASAP7_75t_R _22886_ (.A(_16048_),
    .B(_01198_),
    .Y(_17037_));
 OA211x2_ASAP7_75t_R _22887_ (.A1(_16540_),
    .A2(_17036_),
    .B(_17037_),
    .C(_16044_),
    .Y(_17038_));
 INVx1_ASAP7_75t_R _22888_ (.A(_01199_),
    .Y(_17039_));
 NAND2x1_ASAP7_75t_R _22889_ (.A(_15748_),
    .B(_01197_),
    .Y(_17040_));
 OA211x2_ASAP7_75t_R _22890_ (.A1(_16540_),
    .A2(_17039_),
    .B(_17040_),
    .C(_15930_),
    .Y(_17041_));
 OR3x1_ASAP7_75t_R _22891_ (.A(_15902_),
    .B(_17038_),
    .C(_17041_),
    .Y(_17042_));
 AND3x1_ASAP7_75t_R _22892_ (.A(_15528_),
    .B(_17035_),
    .C(_17042_),
    .Y(_17043_));
 AO21x1_ASAP7_75t_R _22893_ (.A1(_15747_),
    .A2(_17028_),
    .B(_17043_),
    .Y(_17044_));
 INVx1_ASAP7_75t_R _22894_ (.A(_01208_),
    .Y(_17045_));
 NAND2x1_ASAP7_75t_R _22895_ (.A(_15572_),
    .B(_01206_),
    .Y(_17046_));
 OA211x2_ASAP7_75t_R _22896_ (.A1(_15542_),
    .A2(_17045_),
    .B(_17046_),
    .C(_16153_),
    .Y(_17047_));
 INVx1_ASAP7_75t_R _22897_ (.A(_01207_),
    .Y(_17048_));
 NAND2x1_ASAP7_75t_R _22898_ (.A(_15586_),
    .B(_01205_),
    .Y(_17049_));
 OA211x2_ASAP7_75t_R _22899_ (.A1(_15617_),
    .A2(_17048_),
    .B(_17049_),
    .C(_15883_),
    .Y(_17050_));
 OR3x1_ASAP7_75t_R _22900_ (.A(_15530_),
    .B(_17047_),
    .C(_17050_),
    .Y(_17051_));
 INVx1_ASAP7_75t_R _22901_ (.A(_01216_),
    .Y(_17052_));
 NAND2x1_ASAP7_75t_R _22902_ (.A(_15572_),
    .B(_01214_),
    .Y(_17053_));
 OA211x2_ASAP7_75t_R _22903_ (.A1(_15612_),
    .A2(_17052_),
    .B(_17053_),
    .C(_15879_),
    .Y(_17054_));
 INVx1_ASAP7_75t_R _22904_ (.A(_01215_),
    .Y(_17055_));
 NAND2x1_ASAP7_75t_R _22905_ (.A(_15586_),
    .B(_01213_),
    .Y(_17056_));
 OA211x2_ASAP7_75t_R _22906_ (.A1(_15617_),
    .A2(_17055_),
    .B(_17056_),
    .C(_15883_),
    .Y(_17057_));
 OR3x1_ASAP7_75t_R _22907_ (.A(_15876_),
    .B(_17054_),
    .C(_17057_),
    .Y(_17058_));
 AND3x1_ASAP7_75t_R _22908_ (.A(_15528_),
    .B(_17051_),
    .C(_17058_),
    .Y(_17059_));
 INVx1_ASAP7_75t_R _22909_ (.A(_01209_),
    .Y(_17060_));
 NOR2x1_ASAP7_75t_R _22910_ (.A(_16029_),
    .B(_01211_),
    .Y(_17061_));
 AO21x1_ASAP7_75t_R _22911_ (.A1(net5),
    .A2(_17060_),
    .B(_17061_),
    .Y(_17062_));
 INVx1_ASAP7_75t_R _22912_ (.A(_01212_),
    .Y(_17063_));
 NAND2x1_ASAP7_75t_R _22913_ (.A(_15572_),
    .B(_01210_),
    .Y(_17064_));
 OA211x2_ASAP7_75t_R _22914_ (.A1(_15656_),
    .A2(_17063_),
    .B(_17064_),
    .C(_16153_),
    .Y(_17065_));
 AO21x1_ASAP7_75t_R _22915_ (.A1(_15931_),
    .A2(_17062_),
    .B(_17065_),
    .Y(_17066_));
 INVx1_ASAP7_75t_R _22916_ (.A(_01204_),
    .Y(_17067_));
 NAND2x1_ASAP7_75t_R _22917_ (.A(_15541_),
    .B(_01202_),
    .Y(_17068_));
 OA211x2_ASAP7_75t_R _22918_ (.A1(_15602_),
    .A2(_17067_),
    .B(_17068_),
    .C(net18),
    .Y(_17069_));
 INVx1_ASAP7_75t_R _22919_ (.A(_01203_),
    .Y(_17070_));
 NAND2x1_ASAP7_75t_R _22920_ (.A(_15541_),
    .B(_01201_),
    .Y(_17071_));
 OA211x2_ASAP7_75t_R _22921_ (.A1(_15602_),
    .A2(_17070_),
    .B(_17071_),
    .C(_15945_),
    .Y(_17072_));
 OR3x1_ASAP7_75t_R _22922_ (.A(_15530_),
    .B(_17069_),
    .C(_17072_),
    .Y(_17073_));
 OA211x2_ASAP7_75t_R _22923_ (.A1(_15753_),
    .A2(_17066_),
    .B(_17073_),
    .C(_15746_),
    .Y(_17074_));
 OR3x1_ASAP7_75t_R _22924_ (.A(_15912_),
    .B(_17059_),
    .C(_17074_),
    .Y(_17075_));
 OAI21x1_ASAP7_75t_R _22925_ (.A1(_15745_),
    .A2(_17044_),
    .B(_17075_),
    .Y(_17076_));
 OA211x2_ASAP7_75t_R _22926_ (.A1(_15555_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_17077_));
 AOI21x1_ASAP7_75t_R _22927_ (.A1(_16532_),
    .A2(_17076_),
    .B(_17077_),
    .Y(_18729_));
 AND2x2_ASAP7_75t_R _22928_ (.A(_15131_),
    .B(_01798_),
    .Y(_17078_));
 AO21x1_ASAP7_75t_R _22929_ (.A1(_13859_),
    .A2(_01188_),
    .B(_17078_),
    .Y(_17079_));
 OAI22x1_ASAP7_75t_R _22930_ (.A1(_01187_),
    .A2(_13858_),
    .B1(_17079_),
    .B2(_14990_),
    .Y(_17080_));
 NAND2x1_ASAP7_75t_R _22931_ (.A(_15190_),
    .B(_01194_),
    .Y(_17081_));
 OA211x2_ASAP7_75t_R _22932_ (.A1(_13921_),
    .A2(_17021_),
    .B(_17081_),
    .C(_14780_),
    .Y(_17082_));
 NAND2x1_ASAP7_75t_R _22933_ (.A(_15190_),
    .B(_01193_),
    .Y(_17083_));
 OA211x2_ASAP7_75t_R _22934_ (.A1(_15718_),
    .A2(_17024_),
    .B(_17083_),
    .C(_13715_),
    .Y(_17084_));
 OR3x2_ASAP7_75t_R _22935_ (.A(_13902_),
    .B(_17082_),
    .C(_17084_),
    .Y(_17085_));
 OA211x2_ASAP7_75t_R _22936_ (.A1(_14986_),
    .A2(_17080_),
    .B(_17085_),
    .C(_13877_),
    .Y(_17086_));
 NAND2x1_ASAP7_75t_R _22937_ (.A(_14743_),
    .B(_01190_),
    .Y(_17087_));
 OA211x2_ASAP7_75t_R _22938_ (.A1(_15017_),
    .A2(_17029_),
    .B(_17087_),
    .C(_13906_),
    .Y(_17088_));
 NAND2x1_ASAP7_75t_R _22939_ (.A(_14938_),
    .B(_01189_),
    .Y(_17089_));
 OA211x2_ASAP7_75t_R _22940_ (.A1(_15042_),
    .A2(_17032_),
    .B(_17089_),
    .C(_13917_),
    .Y(_17090_));
 OR3x1_ASAP7_75t_R _22941_ (.A(_15039_),
    .B(_17088_),
    .C(_17090_),
    .Y(_17091_));
 NAND2x1_ASAP7_75t_R _22942_ (.A(_15019_),
    .B(_01198_),
    .Y(_17092_));
 OA211x2_ASAP7_75t_R _22943_ (.A1(_15017_),
    .A2(_17036_),
    .B(_17092_),
    .C(_13906_),
    .Y(_17093_));
 NAND2x1_ASAP7_75t_R _22944_ (.A(_14945_),
    .B(_01197_),
    .Y(_17094_));
 OA211x2_ASAP7_75t_R _22945_ (.A1(_15042_),
    .A2(_17039_),
    .B(_17094_),
    .C(_13890_),
    .Y(_17095_));
 OR3x1_ASAP7_75t_R _22946_ (.A(_15012_),
    .B(_17093_),
    .C(_17095_),
    .Y(_17096_));
 AND3x2_ASAP7_75t_R _22947_ (.A(_13879_),
    .B(_17091_),
    .C(_17096_),
    .Y(_17097_));
 OR3x4_ASAP7_75t_R _22948_ (.A(_14738_),
    .B(_17086_),
    .C(_17097_),
    .Y(_17098_));
 NAND2x1_ASAP7_75t_R _22949_ (.A(_14743_),
    .B(_01206_),
    .Y(_17099_));
 OA211x2_ASAP7_75t_R _22950_ (.A1(_15006_),
    .A2(_17045_),
    .B(_17099_),
    .C(_13906_),
    .Y(_17100_));
 NAND2x1_ASAP7_75t_R _22951_ (.A(_14938_),
    .B(_01205_),
    .Y(_17101_));
 OA211x2_ASAP7_75t_R _22952_ (.A1(_15042_),
    .A2(_17048_),
    .B(_17101_),
    .C(_13917_),
    .Y(_17102_));
 OR3x1_ASAP7_75t_R _22953_ (.A(_15039_),
    .B(_17100_),
    .C(_17102_),
    .Y(_17103_));
 NAND2x1_ASAP7_75t_R _22954_ (.A(_15019_),
    .B(_01214_),
    .Y(_17104_));
 OA211x2_ASAP7_75t_R _22955_ (.A1(_15017_),
    .A2(_17052_),
    .B(_17104_),
    .C(_13906_),
    .Y(_17105_));
 NAND2x1_ASAP7_75t_R _22956_ (.A(_14945_),
    .B(_01213_),
    .Y(_17106_));
 OA211x2_ASAP7_75t_R _22957_ (.A1(_15042_),
    .A2(_17055_),
    .B(_17106_),
    .C(_13890_),
    .Y(_17107_));
 OR3x1_ASAP7_75t_R _22958_ (.A(_15012_),
    .B(_17105_),
    .C(_17107_),
    .Y(_17108_));
 AND3x1_ASAP7_75t_R _22959_ (.A(_13879_),
    .B(_17103_),
    .C(_17108_),
    .Y(_17109_));
 NOR2x1_ASAP7_75t_R _22960_ (.A(_15677_),
    .B(_01211_),
    .Y(_17110_));
 AO21x1_ASAP7_75t_R _22961_ (.A1(_14011_),
    .A2(_17060_),
    .B(_17110_),
    .Y(_17111_));
 NAND2x1_ASAP7_75t_R _22962_ (.A(_15278_),
    .B(_01210_),
    .Y(_17112_));
 OA211x2_ASAP7_75t_R _22963_ (.A1(_15712_),
    .A2(_17063_),
    .B(_17112_),
    .C(_15686_),
    .Y(_17113_));
 AO21x1_ASAP7_75t_R _22964_ (.A1(_14746_),
    .A2(_17111_),
    .B(_17113_),
    .Y(_17114_));
 NAND2x1_ASAP7_75t_R _22965_ (.A(_14778_),
    .B(_01202_),
    .Y(_17115_));
 OA211x2_ASAP7_75t_R _22966_ (.A1(_14761_),
    .A2(_17067_),
    .B(_17115_),
    .C(_13869_),
    .Y(_17116_));
 NAND2x1_ASAP7_75t_R _22967_ (.A(_14764_),
    .B(_01201_),
    .Y(_17117_));
 OA211x2_ASAP7_75t_R _22968_ (.A1(_13865_),
    .A2(_17070_),
    .B(_17117_),
    .C(_13874_),
    .Y(_17118_));
 OR3x1_ASAP7_75t_R _22969_ (.A(_14777_),
    .B(_17116_),
    .C(_17118_),
    .Y(_17119_));
 OA211x2_ASAP7_75t_R _22970_ (.A1(_13903_),
    .A2(_17114_),
    .B(_17119_),
    .C(_13877_),
    .Y(_17120_));
 OR3x4_ASAP7_75t_R _22971_ (.A(_14776_),
    .B(_17109_),
    .C(_17120_),
    .Y(_17121_));
 INVx2_ASAP7_75t_R _22972_ (.A(_00059_),
    .Y(_17122_));
 OA211x2_ASAP7_75t_R _22973_ (.A1(_14804_),
    .A2(_14805_),
    .B(_17122_),
    .C(_14807_),
    .Y(_17123_));
 AO31x2_ASAP7_75t_R _22974_ (.A1(_14737_),
    .A2(_17098_),
    .A3(_17121_),
    .B(_17123_),
    .Y(_17124_));
 INVx1_ASAP7_75t_R _22975_ (.A(_01527_),
    .Y(_17125_));
 AO32x1_ASAP7_75t_R _22976_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_17124_),
    .B1(_15119_),
    .B2(_17125_),
    .Y(_17126_));
 BUFx6f_ASAP7_75t_R _22977_ (.A(_17126_),
    .Y(_18730_));
 INVx1_ASAP7_75t_R _22978_ (.A(_18730_),
    .Y(_18728_));
 AND2x2_ASAP7_75t_R _22979_ (.A(_15872_),
    .B(_01797_),
    .Y(_17127_));
 AO21x1_ASAP7_75t_R _22980_ (.A1(_15871_),
    .A2(_01221_),
    .B(_17127_),
    .Y(_17128_));
 OAI22x1_ASAP7_75t_R _22981_ (.A1(_01220_),
    .A2(_15500_),
    .B1(_17128_),
    .B2(_15649_),
    .Y(_17129_));
 INVx1_ASAP7_75t_R _22982_ (.A(_01229_),
    .Y(_17130_));
 NAND2x1_ASAP7_75t_R _22983_ (.A(_16048_),
    .B(_01227_),
    .Y(_17131_));
 OA211x2_ASAP7_75t_R _22984_ (.A1(_16046_),
    .A2(_17130_),
    .B(_17131_),
    .C(_16044_),
    .Y(_17132_));
 INVx1_ASAP7_75t_R _22985_ (.A(_01228_),
    .Y(_17133_));
 NAND2x1_ASAP7_75t_R _22986_ (.A(_16048_),
    .B(_01226_),
    .Y(_17134_));
 OA211x2_ASAP7_75t_R _22987_ (.A1(_16046_),
    .A2(_17133_),
    .B(_17134_),
    .C(_15930_),
    .Y(_17135_));
 OR3x1_ASAP7_75t_R _22988_ (.A(_15902_),
    .B(_17132_),
    .C(_17135_),
    .Y(_17136_));
 OA21x2_ASAP7_75t_R _22989_ (.A1(_15870_),
    .A2(_17129_),
    .B(_17136_),
    .Y(_17137_));
 INVx1_ASAP7_75t_R _22990_ (.A(_01225_),
    .Y(_17138_));
 NAND2x1_ASAP7_75t_R _22991_ (.A(_16151_),
    .B(_01223_),
    .Y(_17139_));
 OA211x2_ASAP7_75t_R _22992_ (.A1(_15579_),
    .A2(_17138_),
    .B(_17139_),
    .C(_16153_),
    .Y(_17140_));
 INVx1_ASAP7_75t_R _22993_ (.A(_01224_),
    .Y(_17141_));
 NAND2x1_ASAP7_75t_R _22994_ (.A(_16151_),
    .B(_01222_),
    .Y(_17142_));
 OA211x2_ASAP7_75t_R _22995_ (.A1(_16149_),
    .A2(_17141_),
    .B(_17142_),
    .C(_15883_),
    .Y(_17143_));
 OR3x1_ASAP7_75t_R _22996_ (.A(_15869_),
    .B(_17140_),
    .C(_17143_),
    .Y(_17144_));
 INVx1_ASAP7_75t_R _22997_ (.A(_01233_),
    .Y(_17145_));
 NAND2x1_ASAP7_75t_R _22998_ (.A(_16151_),
    .B(_01231_),
    .Y(_17146_));
 OA211x2_ASAP7_75t_R _22999_ (.A1(_16149_),
    .A2(_17145_),
    .B(_17146_),
    .C(_16153_),
    .Y(_17147_));
 INVx1_ASAP7_75t_R _23000_ (.A(_01232_),
    .Y(_17148_));
 NAND2x1_ASAP7_75t_R _23001_ (.A(_16151_),
    .B(_01230_),
    .Y(_17149_));
 OA211x2_ASAP7_75t_R _23002_ (.A1(_15656_),
    .A2(_17148_),
    .B(_17149_),
    .C(_15883_),
    .Y(_17150_));
 OR3x1_ASAP7_75t_R _23003_ (.A(_15876_),
    .B(_17147_),
    .C(_17150_),
    .Y(_17151_));
 AND3x1_ASAP7_75t_R _23004_ (.A(_15528_),
    .B(_17144_),
    .C(_17151_),
    .Y(_17152_));
 AO21x1_ASAP7_75t_R _23005_ (.A1(_15747_),
    .A2(_17137_),
    .B(_17152_),
    .Y(_17153_));
 INVx1_ASAP7_75t_R _23006_ (.A(_01241_),
    .Y(_17154_));
 NAND2x1_ASAP7_75t_R _23007_ (.A(_15651_),
    .B(_01239_),
    .Y(_17155_));
 OA211x2_ASAP7_75t_R _23008_ (.A1(_16036_),
    .A2(_17154_),
    .B(_17155_),
    .C(_15879_),
    .Y(_17156_));
 INVx2_ASAP7_75t_R _23009_ (.A(_01240_),
    .Y(_17157_));
 NAND2x1_ASAP7_75t_R _23010_ (.A(_15651_),
    .B(_01238_),
    .Y(_17158_));
 OA211x2_ASAP7_75t_R _23011_ (.A1(_16036_),
    .A2(_17157_),
    .B(_17158_),
    .C(_15945_),
    .Y(_17159_));
 OR3x1_ASAP7_75t_R _23012_ (.A(_15530_),
    .B(_17156_),
    .C(_17159_),
    .Y(_17160_));
 INVx1_ASAP7_75t_R _23013_ (.A(_01249_),
    .Y(_17161_));
 NAND2x1_ASAP7_75t_R _23014_ (.A(_15651_),
    .B(_01247_),
    .Y(_17162_));
 OA211x2_ASAP7_75t_R _23015_ (.A1(_16036_),
    .A2(_17161_),
    .B(_17162_),
    .C(_15879_),
    .Y(_17163_));
 INVx1_ASAP7_75t_R _23016_ (.A(_01248_),
    .Y(_17164_));
 NAND2x1_ASAP7_75t_R _23017_ (.A(_15651_),
    .B(_01246_),
    .Y(_17165_));
 OA211x2_ASAP7_75t_R _23018_ (.A1(_16036_),
    .A2(_17164_),
    .B(_17165_),
    .C(_15945_),
    .Y(_17166_));
 OR3x1_ASAP7_75t_R _23019_ (.A(_15876_),
    .B(_17163_),
    .C(_17166_),
    .Y(_17167_));
 AND3x1_ASAP7_75t_R _23020_ (.A(_15528_),
    .B(_17160_),
    .C(_17167_),
    .Y(_17168_));
 INVx2_ASAP7_75t_R _23021_ (.A(_01242_),
    .Y(_17169_));
 NOR2x1_ASAP7_75t_R _23022_ (.A(_15602_),
    .B(_01244_),
    .Y(_17170_));
 AO21x1_ASAP7_75t_R _23023_ (.A1(_15505_),
    .A2(_17169_),
    .B(_17170_),
    .Y(_17171_));
 INVx1_ASAP7_75t_R _23024_ (.A(_01245_),
    .Y(_17172_));
 NAND2x1_ASAP7_75t_R _23025_ (.A(_15572_),
    .B(_01243_),
    .Y(_17173_));
 OA211x2_ASAP7_75t_R _23026_ (.A1(_15612_),
    .A2(_17172_),
    .B(_17173_),
    .C(_15879_),
    .Y(_17174_));
 AO21x1_ASAP7_75t_R _23027_ (.A1(_15509_),
    .A2(_17171_),
    .B(_17174_),
    .Y(_17175_));
 INVx1_ASAP7_75t_R _23028_ (.A(_01237_),
    .Y(_17176_));
 NAND2x1_ASAP7_75t_R _23029_ (.A(_15541_),
    .B(_01235_),
    .Y(_17177_));
 OA211x2_ASAP7_75t_R _23030_ (.A1(_15665_),
    .A2(_17176_),
    .B(_17177_),
    .C(net18),
    .Y(_17178_));
 INVx2_ASAP7_75t_R _23031_ (.A(_01236_),
    .Y(_17179_));
 NAND2x1_ASAP7_75t_R _23032_ (.A(_15541_),
    .B(_01234_),
    .Y(_17180_));
 OA211x2_ASAP7_75t_R _23033_ (.A1(_15576_),
    .A2(_17179_),
    .B(_17180_),
    .C(_15945_),
    .Y(_17181_));
 OR3x1_ASAP7_75t_R _23034_ (.A(_15530_),
    .B(_17178_),
    .C(_17181_),
    .Y(_17182_));
 OA211x2_ASAP7_75t_R _23035_ (.A1(_15753_),
    .A2(_17175_),
    .B(_17182_),
    .C(_13512_),
    .Y(_17183_));
 OR3x1_ASAP7_75t_R _23036_ (.A(_13518_),
    .B(_17168_),
    .C(_17183_),
    .Y(_17184_));
 OAI21x1_ASAP7_75t_R _23037_ (.A1(_15745_),
    .A2(_17153_),
    .B(_17184_),
    .Y(_17185_));
 OA211x2_ASAP7_75t_R _23038_ (.A1(_13601_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_17186_));
 AOI21x1_ASAP7_75t_R _23039_ (.A1(_16532_),
    .A2(_17185_),
    .B(_17186_),
    .Y(_18733_));
 AND2x2_ASAP7_75t_R _23040_ (.A(_14987_),
    .B(_01797_),
    .Y(_17187_));
 AO21x1_ASAP7_75t_R _23041_ (.A1(_13859_),
    .A2(_01221_),
    .B(_17187_),
    .Y(_17188_));
 OAI22x1_ASAP7_75t_R _23042_ (.A1(_01220_),
    .A2(_13858_),
    .B1(_17188_),
    .B2(_14990_),
    .Y(_17189_));
 NAND2x1_ASAP7_75t_R _23043_ (.A(_14820_),
    .B(_01227_),
    .Y(_17190_));
 OA211x2_ASAP7_75t_R _23044_ (.A1(_15677_),
    .A2(_17130_),
    .B(_17190_),
    .C(_14995_),
    .Y(_17191_));
 NAND2x1_ASAP7_75t_R _23045_ (.A(_13751_),
    .B(_01226_),
    .Y(_17192_));
 OA211x2_ASAP7_75t_R _23046_ (.A1(_14992_),
    .A2(_17133_),
    .B(_17192_),
    .C(_15681_),
    .Y(_17193_));
 OR3x2_ASAP7_75t_R _23047_ (.A(_13902_),
    .B(_17191_),
    .C(_17193_),
    .Y(_17194_));
 OA211x2_ASAP7_75t_R _23048_ (.A1(_14986_),
    .A2(_17189_),
    .B(_17194_),
    .C(_14791_),
    .Y(_17195_));
 NAND2x1_ASAP7_75t_R _23049_ (.A(_14848_),
    .B(_01223_),
    .Y(_17196_));
 OA211x2_ASAP7_75t_R _23050_ (.A1(_15207_),
    .A2(_17138_),
    .B(_17196_),
    .C(_15004_),
    .Y(_17197_));
 NAND2x1_ASAP7_75t_R _23051_ (.A(_13925_),
    .B(_01222_),
    .Y(_17198_));
 OA211x2_ASAP7_75t_R _23052_ (.A1(_15013_),
    .A2(_17141_),
    .B(_17198_),
    .C(_15009_),
    .Y(_17199_));
 OR3x1_ASAP7_75t_R _23053_ (.A(_13707_),
    .B(_17197_),
    .C(_17199_),
    .Y(_17200_));
 NAND2x1_ASAP7_75t_R _23054_ (.A(_14857_),
    .B(_01231_),
    .Y(_17201_));
 OA211x2_ASAP7_75t_R _23055_ (.A1(_13924_),
    .A2(_17145_),
    .B(_17201_),
    .C(_15004_),
    .Y(_17202_));
 NAND2x1_ASAP7_75t_R _23056_ (.A(_14872_),
    .B(_01230_),
    .Y(_17203_));
 OA211x2_ASAP7_75t_R _23057_ (.A1(_15006_),
    .A2(_17148_),
    .B(_17203_),
    .C(_15009_),
    .Y(_17204_));
 OR3x1_ASAP7_75t_R _23058_ (.A(_15031_),
    .B(_17202_),
    .C(_17204_),
    .Y(_17205_));
 AND3x2_ASAP7_75t_R _23059_ (.A(_15002_),
    .B(_17200_),
    .C(_17205_),
    .Y(_17206_));
 OR3x4_ASAP7_75t_R _23060_ (.A(_14733_),
    .B(_17195_),
    .C(_17206_),
    .Y(_17207_));
 NAND2x1_ASAP7_75t_R _23061_ (.A(_14854_),
    .B(_01239_),
    .Y(_17208_));
 OA211x2_ASAP7_75t_R _23062_ (.A1(_15207_),
    .A2(_17154_),
    .B(_17208_),
    .C(_15004_),
    .Y(_17209_));
 NAND2x1_ASAP7_75t_R _23063_ (.A(_13925_),
    .B(_01238_),
    .Y(_17210_));
 OA211x2_ASAP7_75t_R _23064_ (.A1(_13924_),
    .A2(_17157_),
    .B(_17210_),
    .C(_15689_),
    .Y(_17211_));
 OR3x1_ASAP7_75t_R _23065_ (.A(_13707_),
    .B(_17209_),
    .C(_17211_),
    .Y(_17212_));
 NAND2x1_ASAP7_75t_R _23066_ (.A(_14848_),
    .B(_01247_),
    .Y(_17213_));
 OA211x2_ASAP7_75t_R _23067_ (.A1(_15207_),
    .A2(_17161_),
    .B(_17213_),
    .C(_15004_),
    .Y(_17214_));
 NAND2x1_ASAP7_75t_R _23068_ (.A(_14872_),
    .B(_01246_),
    .Y(_17215_));
 OA211x2_ASAP7_75t_R _23069_ (.A1(_15013_),
    .A2(_17164_),
    .B(_17215_),
    .C(_15009_),
    .Y(_17216_));
 OR3x1_ASAP7_75t_R _23070_ (.A(_15031_),
    .B(_17214_),
    .C(_17216_),
    .Y(_17217_));
 AND3x1_ASAP7_75t_R _23071_ (.A(_15002_),
    .B(_17212_),
    .C(_17217_),
    .Y(_17218_));
 NOR2x1_ASAP7_75t_R _23072_ (.A(_15954_),
    .B(_01244_),
    .Y(_17219_));
 AO21x1_ASAP7_75t_R _23073_ (.A1(_14011_),
    .A2(_17169_),
    .B(_17219_),
    .Y(_17220_));
 NAND2x1_ASAP7_75t_R _23074_ (.A(_15423_),
    .B(_01243_),
    .Y(_17221_));
 OA211x2_ASAP7_75t_R _23075_ (.A1(_15712_),
    .A2(_17172_),
    .B(_17221_),
    .C(_15686_),
    .Y(_17222_));
 AO21x1_ASAP7_75t_R _23076_ (.A1(_14746_),
    .A2(_17220_),
    .B(_17222_),
    .Y(_17223_));
 NAND2x1_ASAP7_75t_R _23077_ (.A(_15190_),
    .B(_01235_),
    .Y(_17224_));
 OA211x2_ASAP7_75t_R _23078_ (.A1(_13921_),
    .A2(_17176_),
    .B(_17224_),
    .C(_14780_),
    .Y(_17225_));
 NAND2x1_ASAP7_75t_R _23079_ (.A(_14778_),
    .B(_01234_),
    .Y(_17226_));
 OA211x2_ASAP7_75t_R _23080_ (.A1(_15718_),
    .A2(_17179_),
    .B(_17226_),
    .C(_13715_),
    .Y(_17227_));
 OR3x1_ASAP7_75t_R _23081_ (.A(_14777_),
    .B(_17225_),
    .C(_17227_),
    .Y(_17228_));
 OA211x2_ASAP7_75t_R _23082_ (.A1(_13903_),
    .A2(_17223_),
    .B(_17228_),
    .C(_13877_),
    .Y(_17229_));
 OR3x4_ASAP7_75t_R _23083_ (.A(_15025_),
    .B(_17218_),
    .C(_17229_),
    .Y(_17230_));
 INVx1_ASAP7_75t_R _23084_ (.A(_00060_),
    .Y(_17231_));
 OA211x2_ASAP7_75t_R _23085_ (.A1(_15114_),
    .A2(_15115_),
    .B(_17231_),
    .C(_14807_),
    .Y(_17232_));
 AO31x2_ASAP7_75t_R _23086_ (.A1(_14737_),
    .A2(_17207_),
    .A3(_17230_),
    .B(_17232_),
    .Y(_17233_));
 INVx1_ASAP7_75t_R _23087_ (.A(_01526_),
    .Y(_17234_));
 AO32x1_ASAP7_75t_R _23088_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_17233_),
    .B1(_15119_),
    .B2(_17234_),
    .Y(_17235_));
 BUFx6f_ASAP7_75t_R _23089_ (.A(_17235_),
    .Y(_18732_));
 INVx1_ASAP7_75t_R _23090_ (.A(_18732_),
    .Y(_18734_));
 OAI21x1_ASAP7_75t_R _23091_ (.A1(_16998_),
    .A2(_17001_),
    .B(_01219_),
    .Y(_17236_));
 BUFx3_ASAP7_75t_R _23092_ (.A(_01218_),
    .Y(_17237_));
 INVx1_ASAP7_75t_R _23093_ (.A(_01251_),
    .Y(_17238_));
 NOR2x1_ASAP7_75t_R _23094_ (.A(_17237_),
    .B(_17238_),
    .Y(_17239_));
 AND2x2_ASAP7_75t_R _23095_ (.A(_01252_),
    .B(_17238_),
    .Y(_17240_));
 OA211x2_ASAP7_75t_R _23096_ (.A1(_16998_),
    .A2(_17001_),
    .B(_17240_),
    .C(_01219_),
    .Y(_17241_));
 INVx1_ASAP7_75t_R _23097_ (.A(_01252_),
    .Y(_17242_));
 AND3x1_ASAP7_75t_R _23098_ (.A(_17237_),
    .B(_01252_),
    .C(_17238_),
    .Y(_17243_));
 AO21x1_ASAP7_75t_R _23099_ (.A1(_17242_),
    .A2(_01251_),
    .B(_17243_),
    .Y(_17244_));
 AO211x2_ASAP7_75t_R _23100_ (.A1(_17236_),
    .A2(_17239_),
    .B(_17241_),
    .C(_17244_),
    .Y(_17245_));
 BUFx10_ASAP7_75t_R _23101_ (.A(_17245_),
    .Y(\alu_adder_result_ex[25] ));
 OA21x2_ASAP7_75t_R _23102_ (.A1(_01120_),
    .A2(_16757_),
    .B(_01153_),
    .Y(_17246_));
 OA211x2_ASAP7_75t_R _23103_ (.A1(_01152_),
    .A2(_17246_),
    .B(_01219_),
    .C(_01186_),
    .Y(_17247_));
 OR3x1_ASAP7_75t_R _23104_ (.A(_01086_),
    .B(_16757_),
    .C(_01152_),
    .Y(_17248_));
 AO22x1_ASAP7_75t_R _23105_ (.A1(_16998_),
    .A2(_01219_),
    .B1(_17247_),
    .B2(_17248_),
    .Y(_17249_));
 OR2x2_ASAP7_75t_R _23106_ (.A(_16280_),
    .B(_16768_),
    .Y(_17250_));
 OR3x1_ASAP7_75t_R _23107_ (.A(_15408_),
    .B(_16280_),
    .C(_16768_),
    .Y(_17251_));
 AND2x2_ASAP7_75t_R _23108_ (.A(_16771_),
    .B(_17247_),
    .Y(_17252_));
 OA211x2_ASAP7_75t_R _23109_ (.A1(_16277_),
    .A2(_16768_),
    .B(_17251_),
    .C(_17252_),
    .Y(_17253_));
 OA31x2_ASAP7_75t_R _23110_ (.A1(_16268_),
    .A2(_16269_),
    .A3(_17250_),
    .B1(_17253_),
    .Y(_17254_));
 OAI21x1_ASAP7_75t_R _23111_ (.A1(_17249_),
    .A2(_17254_),
    .B(_17237_),
    .Y(_17255_));
 OR3x2_ASAP7_75t_R _23112_ (.A(_17237_),
    .B(_17249_),
    .C(_17254_),
    .Y(_17256_));
 NAND2x2_ASAP7_75t_R _23113_ (.A(_17255_),
    .B(_17256_),
    .Y(_17257_));
 INVx3_ASAP7_75t_R _23114_ (.A(_17257_),
    .Y(\alu_adder_result_ex[24] ));
 AND2x2_ASAP7_75t_R _23115_ (.A(_15767_),
    .B(_01796_),
    .Y(_17258_));
 AO21x1_ASAP7_75t_R _23116_ (.A1(_15871_),
    .A2(_01254_),
    .B(_17258_),
    .Y(_17259_));
 OAI22x1_ASAP7_75t_R _23117_ (.A1(_01253_),
    .A2(_15500_),
    .B1(_17259_),
    .B2(_15569_),
    .Y(_17260_));
 INVx1_ASAP7_75t_R _23118_ (.A(_01262_),
    .Y(_17261_));
 NAND2x1_ASAP7_75t_R _23119_ (.A(_15891_),
    .B(_01260_),
    .Y(_17262_));
 OA211x2_ASAP7_75t_R _23120_ (.A1(_16079_),
    .A2(_17261_),
    .B(_17262_),
    .C(_16082_),
    .Y(_17263_));
 INVx2_ASAP7_75t_R _23121_ (.A(_01261_),
    .Y(_17264_));
 NAND2x1_ASAP7_75t_R _23122_ (.A(_15609_),
    .B(_01259_),
    .Y(_17265_));
 OA211x2_ASAP7_75t_R _23123_ (.A1(_15889_),
    .A2(_17264_),
    .B(_17265_),
    .C(_15918_),
    .Y(_17266_));
 OR3x1_ASAP7_75t_R _23124_ (.A(_15902_),
    .B(_17263_),
    .C(_17266_),
    .Y(_17267_));
 OA211x2_ASAP7_75t_R _23125_ (.A1(_15870_),
    .A2(_17260_),
    .B(_17267_),
    .C(_16159_),
    .Y(_17268_));
 INVx1_ASAP7_75t_R _23126_ (.A(_01258_),
    .Y(_17269_));
 NAND2x1_ASAP7_75t_R _23127_ (.A(_16303_),
    .B(_01256_),
    .Y(_17270_));
 OA211x2_ASAP7_75t_R _23128_ (.A1(_15573_),
    .A2(_17269_),
    .B(_17270_),
    .C(net21),
    .Y(_17271_));
 INVx1_ASAP7_75t_R _23129_ (.A(_01257_),
    .Y(_17272_));
 NAND2x1_ASAP7_75t_R _23130_ (.A(_16029_),
    .B(_01255_),
    .Y(_17273_));
 OA211x2_ASAP7_75t_R _23131_ (.A1(_15652_),
    .A2(_17272_),
    .B(_17273_),
    .C(_16309_),
    .Y(_17274_));
 OR3x1_ASAP7_75t_R _23132_ (.A(_15498_),
    .B(_17271_),
    .C(_17274_),
    .Y(_17275_));
 INVx1_ASAP7_75t_R _23133_ (.A(_01266_),
    .Y(_17276_));
 NAND2x1_ASAP7_75t_R _23134_ (.A(_16029_),
    .B(_01264_),
    .Y(_17277_));
 OA211x2_ASAP7_75t_R _23135_ (.A1(_15652_),
    .A2(_17276_),
    .B(_17277_),
    .C(net21),
    .Y(_17278_));
 INVx1_ASAP7_75t_R _23136_ (.A(_01265_),
    .Y(_17279_));
 NAND2x1_ASAP7_75t_R _23137_ (.A(_16029_),
    .B(_01263_),
    .Y(_17280_));
 OA211x2_ASAP7_75t_R _23138_ (.A1(_15652_),
    .A2(_17279_),
    .B(_17280_),
    .C(_15523_),
    .Y(_17281_));
 OR3x1_ASAP7_75t_R _23139_ (.A(_15512_),
    .B(_17278_),
    .C(_17281_),
    .Y(_17282_));
 AND3x1_ASAP7_75t_R _23140_ (.A(_15887_),
    .B(_17275_),
    .C(_17282_),
    .Y(_17283_));
 OR3x4_ASAP7_75t_R _23141_ (.A(_15497_),
    .B(_17268_),
    .C(_17283_),
    .Y(_17284_));
 INVx1_ASAP7_75t_R _23142_ (.A(_01274_),
    .Y(_17285_));
 NAND2x1_ASAP7_75t_R _23143_ (.A(_16029_),
    .B(_01272_),
    .Y(_17286_));
 OA211x2_ASAP7_75t_R _23144_ (.A1(_15652_),
    .A2(_17285_),
    .B(_17286_),
    .C(net21),
    .Y(_17287_));
 INVx2_ASAP7_75t_R _23145_ (.A(_01273_),
    .Y(_17288_));
 NAND2x1_ASAP7_75t_R _23146_ (.A(_16029_),
    .B(_01271_),
    .Y(_17289_));
 OA211x2_ASAP7_75t_R _23147_ (.A1(_15652_),
    .A2(_17288_),
    .B(_17289_),
    .C(_15523_),
    .Y(_17290_));
 OR3x1_ASAP7_75t_R _23148_ (.A(_15498_),
    .B(_17287_),
    .C(_17290_),
    .Y(_17291_));
 INVx1_ASAP7_75t_R _23149_ (.A(_01282_),
    .Y(_17292_));
 NAND2x1_ASAP7_75t_R _23150_ (.A(_16029_),
    .B(_01280_),
    .Y(_17293_));
 OA211x2_ASAP7_75t_R _23151_ (.A1(_15652_),
    .A2(_17292_),
    .B(_17293_),
    .C(net21),
    .Y(_17294_));
 INVx2_ASAP7_75t_R _23152_ (.A(_01281_),
    .Y(_17295_));
 NAND2x1_ASAP7_75t_R _23153_ (.A(_16029_),
    .B(_01279_),
    .Y(_17296_));
 OA211x2_ASAP7_75t_R _23154_ (.A1(_15652_),
    .A2(_17295_),
    .B(_17296_),
    .C(_15523_),
    .Y(_17297_));
 OR3x1_ASAP7_75t_R _23155_ (.A(_15512_),
    .B(_17294_),
    .C(_17297_),
    .Y(_17298_));
 AND3x1_ASAP7_75t_R _23156_ (.A(_15887_),
    .B(_17291_),
    .C(_17298_),
    .Y(_17299_));
 INVx2_ASAP7_75t_R _23157_ (.A(_01275_),
    .Y(_17300_));
 NOR2x1_ASAP7_75t_R _23158_ (.A(_15594_),
    .B(_01277_),
    .Y(_17301_));
 AO21x1_ASAP7_75t_R _23159_ (.A1(_15602_),
    .A2(_17300_),
    .B(_17301_),
    .Y(_17302_));
 INVx2_ASAP7_75t_R _23160_ (.A(_01278_),
    .Y(_17303_));
 NAND2x1_ASAP7_75t_R _23161_ (.A(_16422_),
    .B(_01276_),
    .Y(_17304_));
 OA211x2_ASAP7_75t_R _23162_ (.A1(_16420_),
    .A2(_17303_),
    .B(_17304_),
    .C(_16305_),
    .Y(_17305_));
 AO21x1_ASAP7_75t_R _23163_ (.A1(_15931_),
    .A2(_17302_),
    .B(_17305_),
    .Y(_17306_));
 INVx1_ASAP7_75t_R _23164_ (.A(_01270_),
    .Y(_17307_));
 NAND2x1_ASAP7_75t_R _23165_ (.A(_15897_),
    .B(_01268_),
    .Y(_17308_));
 OA211x2_ASAP7_75t_R _23166_ (.A1(_15756_),
    .A2(_17307_),
    .B(_17308_),
    .C(_16044_),
    .Y(_17309_));
 INVx2_ASAP7_75t_R _23167_ (.A(_01269_),
    .Y(_17310_));
 NAND2x1_ASAP7_75t_R _23168_ (.A(_16048_),
    .B(_01267_),
    .Y(_17311_));
 OA211x2_ASAP7_75t_R _23169_ (.A1(_16046_),
    .A2(_17310_),
    .B(_17311_),
    .C(_15930_),
    .Y(_17312_));
 OR3x1_ASAP7_75t_R _23170_ (.A(_15869_),
    .B(_17309_),
    .C(_17312_),
    .Y(_17313_));
 OA211x2_ASAP7_75t_R _23171_ (.A1(_15929_),
    .A2(_17306_),
    .B(_17313_),
    .C(_16159_),
    .Y(_17314_));
 OR3x4_ASAP7_75t_R _23172_ (.A(_15912_),
    .B(_17299_),
    .C(_17314_),
    .Y(_17315_));
 NAND2x2_ASAP7_75t_R _23173_ (.A(_17284_),
    .B(_17315_),
    .Y(_17316_));
 OA211x2_ASAP7_75t_R _23174_ (.A1(_13589_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_17317_));
 AOI21x1_ASAP7_75t_R _23175_ (.A1(_16532_),
    .A2(_17316_),
    .B(_17317_),
    .Y(_18739_));
 AND2x2_ASAP7_75t_R _23176_ (.A(_13689_),
    .B(_01796_),
    .Y(_17318_));
 AO21x1_ASAP7_75t_R _23177_ (.A1(_14742_),
    .A2(_01254_),
    .B(_17318_),
    .Y(_17319_));
 OAI22x1_ASAP7_75t_R _23178_ (.A1(_01253_),
    .A2(_13948_),
    .B1(_17319_),
    .B2(_13918_),
    .Y(_17320_));
 NAND2x1_ASAP7_75t_R _23179_ (.A(_14858_),
    .B(_01260_),
    .Y(_17321_));
 OA211x2_ASAP7_75t_R _23180_ (.A1(_14857_),
    .A2(_17261_),
    .B(_17321_),
    .C(_14846_),
    .Y(_17322_));
 NAND2x1_ASAP7_75t_R _23181_ (.A(_13682_),
    .B(_01259_),
    .Y(_17323_));
 OA211x2_ASAP7_75t_R _23182_ (.A1(_14872_),
    .A2(_17264_),
    .B(_17323_),
    .C(_14867_),
    .Y(_17324_));
 OR3x1_ASAP7_75t_R _23183_ (.A(_14853_),
    .B(_17322_),
    .C(_17324_),
    .Y(_17325_));
 OA211x2_ASAP7_75t_R _23184_ (.A1(_14740_),
    .A2(_17320_),
    .B(_17325_),
    .C(_13961_),
    .Y(_17326_));
 NAND2x1_ASAP7_75t_R _23185_ (.A(_13726_),
    .B(_01256_),
    .Y(_17327_));
 OA211x2_ASAP7_75t_R _23186_ (.A1(_15358_),
    .A2(_17269_),
    .B(_17327_),
    .C(_15352_),
    .Y(_17328_));
 NAND2x1_ASAP7_75t_R _23187_ (.A(_13763_),
    .B(_01255_),
    .Y(_17329_));
 OA211x2_ASAP7_75t_R _23188_ (.A1(_13750_),
    .A2(_17272_),
    .B(_17329_),
    .C(_15355_),
    .Y(_17330_));
 OR3x1_ASAP7_75t_R _23189_ (.A(_14985_),
    .B(_17328_),
    .C(_17330_),
    .Y(_17331_));
 NAND2x1_ASAP7_75t_R _23190_ (.A(_13763_),
    .B(_01264_),
    .Y(_17332_));
 OA211x2_ASAP7_75t_R _23191_ (.A1(_13750_),
    .A2(_17276_),
    .B(_17332_),
    .C(_15352_),
    .Y(_17333_));
 NAND2x1_ASAP7_75t_R _23192_ (.A(_13880_),
    .B(_01263_),
    .Y(_17334_));
 OA211x2_ASAP7_75t_R _23193_ (.A1(_13860_),
    .A2(_17279_),
    .B(_17334_),
    .C(_15355_),
    .Y(_17335_));
 OR3x1_ASAP7_75t_R _23194_ (.A(_14748_),
    .B(_17333_),
    .C(_17335_),
    .Y(_17336_));
 AND3x1_ASAP7_75t_R _23195_ (.A(_14843_),
    .B(_17331_),
    .C(_17336_),
    .Y(_17337_));
 OR3x4_ASAP7_75t_R _23196_ (.A(_14814_),
    .B(_17326_),
    .C(_17337_),
    .Y(_17338_));
 NAND2x1_ASAP7_75t_R _23197_ (.A(_13721_),
    .B(_01272_),
    .Y(_17339_));
 OA211x2_ASAP7_75t_R _23198_ (.A1(_15126_),
    .A2(_17285_),
    .B(_17339_),
    .C(_15352_),
    .Y(_17340_));
 NAND2x1_ASAP7_75t_R _23199_ (.A(_13726_),
    .B(_01271_),
    .Y(_17341_));
 OA211x2_ASAP7_75t_R _23200_ (.A1(_15358_),
    .A2(_17288_),
    .B(_17341_),
    .C(_15134_),
    .Y(_17342_));
 OR3x1_ASAP7_75t_R _23201_ (.A(_14985_),
    .B(_17340_),
    .C(_17342_),
    .Y(_04261_));
 NAND2x1_ASAP7_75t_R _23202_ (.A(_13721_),
    .B(_01280_),
    .Y(_04262_));
 OA211x2_ASAP7_75t_R _23203_ (.A1(_15131_),
    .A2(_17292_),
    .B(_04262_),
    .C(_15352_),
    .Y(_04263_));
 NAND2x1_ASAP7_75t_R _23204_ (.A(_13726_),
    .B(_01279_),
    .Y(_04264_));
 OA211x2_ASAP7_75t_R _23205_ (.A1(_15358_),
    .A2(_17295_),
    .B(_04264_),
    .C(_15355_),
    .Y(_04265_));
 OR3x1_ASAP7_75t_R _23206_ (.A(_15125_),
    .B(_04263_),
    .C(_04265_),
    .Y(_04266_));
 AND3x1_ASAP7_75t_R _23207_ (.A(_14843_),
    .B(_04261_),
    .C(_04266_),
    .Y(_04267_));
 NOR2x1_ASAP7_75t_R _23208_ (.A(_15278_),
    .B(_01277_),
    .Y(_04268_));
 AO21x1_ASAP7_75t_R _23209_ (.A1(_15042_),
    .A2(_17300_),
    .B(_04268_),
    .Y(_04269_));
 NAND2x1_ASAP7_75t_R _23210_ (.A(_13935_),
    .B(_01276_),
    .Y(_04270_));
 OA211x2_ASAP7_75t_R _23211_ (.A1(_15307_),
    .A2(_17303_),
    .B(_04270_),
    .C(_15305_),
    .Y(_04271_));
 AO21x1_ASAP7_75t_R _23212_ (.A1(_13716_),
    .A2(_04269_),
    .B(_04271_),
    .Y(_04272_));
 NAND2x1_ASAP7_75t_R _23213_ (.A(_13682_),
    .B(_01268_),
    .Y(_04273_));
 OA211x2_ASAP7_75t_R _23214_ (.A1(_14743_),
    .A2(_17307_),
    .B(_04273_),
    .C(_14846_),
    .Y(_04274_));
 NAND2x1_ASAP7_75t_R _23215_ (.A(_13682_),
    .B(_01267_),
    .Y(_04275_));
 OA211x2_ASAP7_75t_R _23216_ (.A1(_14938_),
    .A2(_17310_),
    .B(_04275_),
    .C(_14867_),
    .Y(_04276_));
 OR3x1_ASAP7_75t_R _23217_ (.A(_13676_),
    .B(_04274_),
    .C(_04276_),
    .Y(_04277_));
 OA211x2_ASAP7_75t_R _23218_ (.A1(_15318_),
    .A2(_04272_),
    .B(_04277_),
    .C(_13961_),
    .Y(_04278_));
 OR3x4_ASAP7_75t_R _23219_ (.A(_14842_),
    .B(_04267_),
    .C(_04278_),
    .Y(_04279_));
 INVx1_ASAP7_75t_R _23220_ (.A(_00061_),
    .Y(_04280_));
 OA211x2_ASAP7_75t_R _23221_ (.A1(_14804_),
    .A2(_14805_),
    .B(_04280_),
    .C(_15334_),
    .Y(_04281_));
 AO31x2_ASAP7_75t_R _23222_ (.A1(_13947_),
    .A2(_17338_),
    .A3(_04279_),
    .B(_04281_),
    .Y(_04282_));
 INVx1_ASAP7_75t_R _23223_ (.A(_01525_),
    .Y(_04283_));
 AO32x1_ASAP7_75t_R _23224_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_04282_),
    .B1(_15337_),
    .B2(_04283_),
    .Y(_04284_));
 BUFx4f_ASAP7_75t_R _23225_ (.A(_04284_),
    .Y(_18740_));
 INVx3_ASAP7_75t_R _23226_ (.A(_18740_),
    .Y(_18738_));
 AND2x2_ASAP7_75t_R _23227_ (.A(_15505_),
    .B(_01795_),
    .Y(_04285_));
 AO21x1_ASAP7_75t_R _23228_ (.A1(_15502_),
    .A2(_01287_),
    .B(_04285_),
    .Y(_04286_));
 OAI22x1_ASAP7_75t_R _23229_ (.A1(_01286_),
    .A2(_15500_),
    .B1(_04286_),
    .B2(_15569_),
    .Y(_04287_));
 INVx1_ASAP7_75t_R _23230_ (.A(_01295_),
    .Y(_04288_));
 NAND2x1_ASAP7_75t_R _23231_ (.A(_15516_),
    .B(_01293_),
    .Y(_04289_));
 OA211x2_ASAP7_75t_R _23232_ (.A1(_15513_),
    .A2(_04288_),
    .B(_04289_),
    .C(_15519_),
    .Y(_04290_));
 INVx1_ASAP7_75t_R _23233_ (.A(_01294_),
    .Y(_04291_));
 NAND2x1_ASAP7_75t_R _23234_ (.A(_15516_),
    .B(_01292_),
    .Y(_04292_));
 OA211x2_ASAP7_75t_R _23235_ (.A1(_15513_),
    .A2(_04291_),
    .B(_04292_),
    .C(_15523_),
    .Y(_04293_));
 OR3x1_ASAP7_75t_R _23236_ (.A(_15512_),
    .B(_04290_),
    .C(_04293_),
    .Y(_04294_));
 OA211x2_ASAP7_75t_R _23237_ (.A1(_15499_),
    .A2(_04287_),
    .B(_04294_),
    .C(_15526_),
    .Y(_04295_));
 INVx1_ASAP7_75t_R _23238_ (.A(_01291_),
    .Y(_04296_));
 NAND2x1_ASAP7_75t_R _23239_ (.A(_15535_),
    .B(_01289_),
    .Y(_04297_));
 OA211x2_ASAP7_75t_R _23240_ (.A1(_15533_),
    .A2(_04296_),
    .B(_04297_),
    .C(_15538_),
    .Y(_04298_));
 INVx1_ASAP7_75t_R _23241_ (.A(_01290_),
    .Y(_04299_));
 NAND2x1_ASAP7_75t_R _23242_ (.A(_15542_),
    .B(_01288_),
    .Y(_04300_));
 OA211x2_ASAP7_75t_R _23243_ (.A1(_15540_),
    .A2(_04299_),
    .B(_04300_),
    .C(_15544_),
    .Y(_04301_));
 OR3x1_ASAP7_75t_R _23244_ (.A(_15531_),
    .B(_04298_),
    .C(_04301_),
    .Y(_04302_));
 INVx1_ASAP7_75t_R _23245_ (.A(_01299_),
    .Y(_04303_));
 NAND2x1_ASAP7_75t_R _23246_ (.A(_15542_),
    .B(_01297_),
    .Y(_04304_));
 OA211x2_ASAP7_75t_R _23247_ (.A1(_15540_),
    .A2(_04303_),
    .B(_04304_),
    .C(_15538_),
    .Y(_04305_));
 INVx1_ASAP7_75t_R _23248_ (.A(_01298_),
    .Y(_04306_));
 NAND2x1_ASAP7_75t_R _23249_ (.A(_15612_),
    .B(_01296_),
    .Y(_04307_));
 OA211x2_ASAP7_75t_R _23250_ (.A1(_15540_),
    .A2(_04306_),
    .B(_04307_),
    .C(_15544_),
    .Y(_04308_));
 OR3x1_ASAP7_75t_R _23251_ (.A(_15547_),
    .B(_04305_),
    .C(_04308_),
    .Y(_04309_));
 AND3x1_ASAP7_75t_R _23252_ (.A(_15529_),
    .B(_04302_),
    .C(_04309_),
    .Y(_04310_));
 OR3x4_ASAP7_75t_R _23253_ (.A(_15497_),
    .B(_04295_),
    .C(_04310_),
    .Y(_04311_));
 INVx2_ASAP7_75t_R _23254_ (.A(_01307_),
    .Y(_04312_));
 NAND2x1_ASAP7_75t_R _23255_ (.A(_15542_),
    .B(_01305_),
    .Y(_04313_));
 OA211x2_ASAP7_75t_R _23256_ (.A1(_15540_),
    .A2(_04312_),
    .B(_04313_),
    .C(_15538_),
    .Y(_04314_));
 INVx2_ASAP7_75t_R _23257_ (.A(_01306_),
    .Y(_04315_));
 NAND2x1_ASAP7_75t_R _23258_ (.A(_15612_),
    .B(_01304_),
    .Y(_04316_));
 OA211x2_ASAP7_75t_R _23259_ (.A1(_15540_),
    .A2(_04315_),
    .B(_04316_),
    .C(_15544_),
    .Y(_04317_));
 OR3x1_ASAP7_75t_R _23260_ (.A(_15608_),
    .B(_04314_),
    .C(_04317_),
    .Y(_04318_));
 INVx2_ASAP7_75t_R _23261_ (.A(_01315_),
    .Y(_04319_));
 NAND2x1_ASAP7_75t_R _23262_ (.A(_15542_),
    .B(_01313_),
    .Y(_04320_));
 OA211x2_ASAP7_75t_R _23263_ (.A1(_15540_),
    .A2(_04319_),
    .B(_04320_),
    .C(net145),
    .Y(_04321_));
 INVx1_ASAP7_75t_R _23264_ (.A(_01314_),
    .Y(_04322_));
 NAND2x1_ASAP7_75t_R _23265_ (.A(_15612_),
    .B(_01312_),
    .Y(_04323_));
 OA211x2_ASAP7_75t_R _23266_ (.A1(_15610_),
    .A2(_04322_),
    .B(_04323_),
    .C(_15544_),
    .Y(_04324_));
 OR3x1_ASAP7_75t_R _23267_ (.A(_15547_),
    .B(_04321_),
    .C(_04324_),
    .Y(_04325_));
 AND3x1_ASAP7_75t_R _23268_ (.A(_15607_),
    .B(_04318_),
    .C(_04325_),
    .Y(_04326_));
 INVx1_ASAP7_75t_R _23269_ (.A(_01308_),
    .Y(_04327_));
 NOR2x1_ASAP7_75t_R _23270_ (.A(_15652_),
    .B(_01310_),
    .Y(_04328_));
 AO21x1_ASAP7_75t_R _23271_ (.A1(_15571_),
    .A2(_04327_),
    .B(_04328_),
    .Y(_04329_));
 INVx2_ASAP7_75t_R _23272_ (.A(_01311_),
    .Y(_04330_));
 NAND2x1_ASAP7_75t_R _23273_ (.A(_16149_),
    .B(_01309_),
    .Y(_04331_));
 OA211x2_ASAP7_75t_R _23274_ (.A1(_15577_),
    .A2(_04330_),
    .B(_04331_),
    .C(_15581_),
    .Y(_04332_));
 AO21x1_ASAP7_75t_R _23275_ (.A1(_15569_),
    .A2(_04329_),
    .B(_04332_),
    .Y(_04333_));
 INVx1_ASAP7_75t_R _23276_ (.A(_01303_),
    .Y(_04334_));
 NAND2x1_ASAP7_75t_R _23277_ (.A(_15602_),
    .B(_01301_),
    .Y(_04335_));
 OA211x2_ASAP7_75t_R _23278_ (.A1(_15587_),
    .A2(_04334_),
    .B(_04335_),
    .C(_15519_),
    .Y(_04336_));
 INVx2_ASAP7_75t_R _23279_ (.A(_01302_),
    .Y(_04337_));
 NAND2x1_ASAP7_75t_R _23280_ (.A(_15602_),
    .B(_01300_),
    .Y(_04338_));
 OA211x2_ASAP7_75t_R _23281_ (.A1(_15587_),
    .A2(_04337_),
    .B(_04338_),
    .C(_15523_),
    .Y(_04339_));
 OR3x1_ASAP7_75t_R _23282_ (.A(_15498_),
    .B(_04336_),
    .C(_04339_),
    .Y(_04340_));
 OA211x2_ASAP7_75t_R _23283_ (.A1(_15568_),
    .A2(_04333_),
    .B(_04340_),
    .C(_15526_),
    .Y(_04341_));
 OR3x4_ASAP7_75t_R _23284_ (.A(_15555_),
    .B(_04326_),
    .C(_04341_),
    .Y(_04342_));
 NAND2x2_ASAP7_75t_R _23285_ (.A(_04311_),
    .B(_04342_),
    .Y(_04343_));
 OA211x2_ASAP7_75t_R _23286_ (.A1(_13579_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_04344_));
 AOI21x1_ASAP7_75t_R _23287_ (.A1(_16532_),
    .A2(_04343_),
    .B(_04344_),
    .Y(_18743_));
 AND2x2_ASAP7_75t_R _23288_ (.A(_15061_),
    .B(_01795_),
    .Y(_04345_));
 AO21x1_ASAP7_75t_R _23289_ (.A1(_13859_),
    .A2(_01287_),
    .B(_04345_),
    .Y(_04346_));
 OAI22x1_ASAP7_75t_R _23290_ (.A1(_01286_),
    .A2(_14741_),
    .B1(_04346_),
    .B2(_13863_),
    .Y(_04347_));
 NAND2x1_ASAP7_75t_R _23291_ (.A(_13872_),
    .B(_01293_),
    .Y(_04348_));
 OA211x2_ASAP7_75t_R _23292_ (.A1(_13871_),
    .A2(_04288_),
    .B(_04348_),
    .C(_13932_),
    .Y(_04349_));
 NAND2x1_ASAP7_75t_R _23293_ (.A(_13935_),
    .B(_01292_),
    .Y(_04350_));
 OA211x2_ASAP7_75t_R _23294_ (.A1(_13934_),
    .A2(_04291_),
    .B(_04350_),
    .C(_13937_),
    .Y(_04351_));
 OR3x2_ASAP7_75t_R _23295_ (.A(_14768_),
    .B(_04349_),
    .C(_04351_),
    .Y(_04352_));
 OA211x2_ASAP7_75t_R _23296_ (.A1(_14986_),
    .A2(_04347_),
    .B(_04352_),
    .C(_13877_),
    .Y(_04353_));
 NAND2x1_ASAP7_75t_R _23297_ (.A(_13755_),
    .B(_01289_),
    .Y(_04354_));
 OA211x2_ASAP7_75t_R _23298_ (.A1(_13887_),
    .A2(_04296_),
    .B(_04354_),
    .C(_15081_),
    .Y(_04355_));
 NAND2x1_ASAP7_75t_R _23299_ (.A(_15075_),
    .B(_01288_),
    .Y(_04356_));
 OA211x2_ASAP7_75t_R _23300_ (.A1(_15074_),
    .A2(_04299_),
    .B(_04356_),
    .C(_13897_),
    .Y(_04357_));
 OR3x1_ASAP7_75t_R _23301_ (.A(_13856_),
    .B(_04355_),
    .C(_04357_),
    .Y(_04358_));
 NAND2x1_ASAP7_75t_R _23302_ (.A(_15075_),
    .B(_01297_),
    .Y(_04359_));
 OA211x2_ASAP7_75t_R _23303_ (.A1(_13895_),
    .A2(_04303_),
    .B(_04359_),
    .C(_15081_),
    .Y(_04360_));
 NAND2x1_ASAP7_75t_R _23304_ (.A(_13680_),
    .B(_01296_),
    .Y(_04361_));
 OA211x2_ASAP7_75t_R _23305_ (.A1(_15074_),
    .A2(_04306_),
    .B(_04361_),
    .C(_15109_),
    .Y(_04362_));
 OR3x1_ASAP7_75t_R _23306_ (.A(_15079_),
    .B(_04360_),
    .C(_04362_),
    .Y(_04363_));
 AND3x2_ASAP7_75t_R _23307_ (.A(_13879_),
    .B(_04358_),
    .C(_04363_),
    .Y(_04364_));
 OR3x4_ASAP7_75t_R _23308_ (.A(_14738_),
    .B(_04353_),
    .C(_04364_),
    .Y(_04365_));
 NAND2x1_ASAP7_75t_R _23309_ (.A(_13755_),
    .B(_01305_),
    .Y(_04366_));
 OA211x2_ASAP7_75t_R _23310_ (.A1(_13887_),
    .A2(_04312_),
    .B(_04366_),
    .C(_15081_),
    .Y(_04367_));
 NAND2x1_ASAP7_75t_R _23311_ (.A(_15075_),
    .B(_01304_),
    .Y(_04368_));
 OA211x2_ASAP7_75t_R _23312_ (.A1(_15074_),
    .A2(_04315_),
    .B(_04368_),
    .C(_13897_),
    .Y(_04369_));
 OR3x1_ASAP7_75t_R _23313_ (.A(_13856_),
    .B(_04367_),
    .C(_04369_),
    .Y(_04370_));
 NAND2x1_ASAP7_75t_R _23314_ (.A(_13755_),
    .B(_01313_),
    .Y(_04371_));
 OA211x2_ASAP7_75t_R _23315_ (.A1(_13895_),
    .A2(_04319_),
    .B(_04371_),
    .C(_15081_),
    .Y(_04372_));
 NAND2x1_ASAP7_75t_R _23316_ (.A(_13680_),
    .B(_01312_),
    .Y(_04373_));
 OA211x2_ASAP7_75t_R _23317_ (.A1(_15074_),
    .A2(_04322_),
    .B(_04373_),
    .C(_13897_),
    .Y(_04374_));
 OR3x1_ASAP7_75t_R _23318_ (.A(_15079_),
    .B(_04372_),
    .C(_04374_),
    .Y(_04375_));
 AND3x1_ASAP7_75t_R _23319_ (.A(_13879_),
    .B(_04370_),
    .C(_04375_),
    .Y(_04376_));
 NOR2x1_ASAP7_75t_R _23320_ (.A(_14761_),
    .B(_01310_),
    .Y(_04377_));
 AO21x1_ASAP7_75t_R _23321_ (.A1(_13920_),
    .A2(_04327_),
    .B(_04377_),
    .Y(_04378_));
 NAND2x1_ASAP7_75t_R _23322_ (.A(_15019_),
    .B(_01309_),
    .Y(_04379_));
 OA211x2_ASAP7_75t_R _23323_ (.A1(_15017_),
    .A2(_04330_),
    .B(_04379_),
    .C(_13906_),
    .Y(_04380_));
 AO21x1_ASAP7_75t_R _23324_ (.A1(_13918_),
    .A2(_04378_),
    .B(_04380_),
    .Y(_04381_));
 NAND2x1_ASAP7_75t_R _23325_ (.A(_14816_),
    .B(_01301_),
    .Y(_04382_));
 OA211x2_ASAP7_75t_R _23326_ (.A1(_15307_),
    .A2(_04334_),
    .B(_04382_),
    .C(_15129_),
    .Y(_04383_));
 NAND2x1_ASAP7_75t_R _23327_ (.A(_13952_),
    .B(_01300_),
    .Y(_04384_));
 OA211x2_ASAP7_75t_R _23328_ (.A1(_14987_),
    .A2(_04337_),
    .B(_04384_),
    .C(_15309_),
    .Y(_04385_));
 OR3x1_ASAP7_75t_R _23329_ (.A(_14985_),
    .B(_04383_),
    .C(_04385_),
    .Y(_04386_));
 OA211x2_ASAP7_75t_R _23330_ (.A1(_15318_),
    .A2(_04381_),
    .B(_04386_),
    .C(_14757_),
    .Y(_04387_));
 OR3x4_ASAP7_75t_R _23331_ (.A(_14776_),
    .B(_04376_),
    .C(_04387_),
    .Y(_04388_));
 INVx2_ASAP7_75t_R _23332_ (.A(_00062_),
    .Y(_04389_));
 OA211x2_ASAP7_75t_R _23333_ (.A1(_14804_),
    .A2(_14805_),
    .B(_04389_),
    .C(_14807_),
    .Y(_04390_));
 AO31x2_ASAP7_75t_R _23334_ (.A1(_14737_),
    .A2(_04365_),
    .A3(_04388_),
    .B(_04390_),
    .Y(_04391_));
 INVx1_ASAP7_75t_R _23335_ (.A(_01524_),
    .Y(_04392_));
 AO32x1_ASAP7_75t_R _23336_ (.A1(_15273_),
    .A2(_15274_),
    .A3(_04391_),
    .B1(_15337_),
    .B2(_04392_),
    .Y(_04393_));
 BUFx6f_ASAP7_75t_R _23337_ (.A(_04393_),
    .Y(_18742_));
 INVx1_ASAP7_75t_R _23338_ (.A(_18742_),
    .Y(_18744_));
 OR5x1_ASAP7_75t_R _23339_ (.A(_16998_),
    .B(_17237_),
    .C(_01251_),
    .D(_16763_),
    .E(_16999_),
    .Y(_04394_));
 AO21x1_ASAP7_75t_R _23340_ (.A1(_16759_),
    .A2(_16267_),
    .B(_04394_),
    .Y(_04395_));
 OA21x2_ASAP7_75t_R _23341_ (.A1(_01219_),
    .A2(_17237_),
    .B(_01252_),
    .Y(_04396_));
 OR4x1_ASAP7_75t_R _23342_ (.A(_16998_),
    .B(_17237_),
    .C(_01251_),
    .D(_17000_),
    .Y(_04397_));
 OA211x2_ASAP7_75t_R _23343_ (.A1(_01251_),
    .A2(_04396_),
    .B(_04397_),
    .C(_01285_),
    .Y(_04398_));
 AND2x2_ASAP7_75t_R _23344_ (.A(_01318_),
    .B(_04398_),
    .Y(_04399_));
 AO22x1_ASAP7_75t_R _23345_ (.A1(_01284_),
    .A2(_01318_),
    .B1(_04395_),
    .B2(_04399_),
    .Y(_04400_));
 XOR2x2_ASAP7_75t_R _23346_ (.A(_01317_),
    .B(_04400_),
    .Y(\alu_adder_result_ex[27] ));
 OR2x2_ASAP7_75t_R _23347_ (.A(_15266_),
    .B(_16523_),
    .Y(_04401_));
 AO31x2_ASAP7_75t_R _23348_ (.A1(_14920_),
    .A2(_14919_),
    .A3(_15484_),
    .B(_04401_),
    .Y(_04402_));
 OA21x2_ASAP7_75t_R _23349_ (.A1(_01186_),
    .A2(_16998_),
    .B(_01219_),
    .Y(_04403_));
 OA21x2_ASAP7_75t_R _23350_ (.A1(_17237_),
    .A2(_04403_),
    .B(_01252_),
    .Y(_04404_));
 OA21x2_ASAP7_75t_R _23351_ (.A1(_01251_),
    .A2(_04404_),
    .B(_01285_),
    .Y(_04405_));
 AND2x2_ASAP7_75t_R _23352_ (.A(_16528_),
    .B(_04405_),
    .Y(_04406_));
 OA211x2_ASAP7_75t_R _23353_ (.A1(_16757_),
    .A2(_17006_),
    .B(_04406_),
    .C(_01153_),
    .Y(_04407_));
 OA21x2_ASAP7_75t_R _23354_ (.A1(_15485_),
    .A2(_04402_),
    .B(_04407_),
    .Y(_04408_));
 OA211x2_ASAP7_75t_R _23355_ (.A1(_16757_),
    .A2(_17006_),
    .B(_17007_),
    .C(_01153_),
    .Y(_04409_));
 OR4x1_ASAP7_75t_R _23356_ (.A(_01152_),
    .B(_16998_),
    .C(_17237_),
    .D(_01251_),
    .Y(_04410_));
 OA21x2_ASAP7_75t_R _23357_ (.A1(_04409_),
    .A2(_04410_),
    .B(_04405_),
    .Y(_04411_));
 OAI21x1_ASAP7_75t_R _23358_ (.A1(_04408_),
    .A2(_04411_),
    .B(_01284_),
    .Y(_04412_));
 OR3x2_ASAP7_75t_R _23359_ (.A(_01284_),
    .B(_04408_),
    .C(_04411_),
    .Y(_04413_));
 NAND2x2_ASAP7_75t_R _23360_ (.A(_04412_),
    .B(_04413_),
    .Y(_04414_));
 INVx3_ASAP7_75t_R _23361_ (.A(_04414_),
    .Y(\alu_adder_result_ex[26] ));
 AND2x2_ASAP7_75t_R _23362_ (.A(_16161_),
    .B(_01794_),
    .Y(_04415_));
 AO21x1_ASAP7_75t_R _23363_ (.A1(_15502_),
    .A2(_01320_),
    .B(_04415_),
    .Y(_04416_));
 OAI22x1_ASAP7_75t_R _23364_ (.A1(_01319_),
    .A2(_15500_),
    .B1(_04416_),
    .B2(_15510_),
    .Y(_04417_));
 INVx2_ASAP7_75t_R _23365_ (.A(_01328_),
    .Y(_04418_));
 NAND2x1_ASAP7_75t_R _23366_ (.A(_15612_),
    .B(_01326_),
    .Y(_04419_));
 OA211x2_ASAP7_75t_R _23367_ (.A1(_15610_),
    .A2(_04418_),
    .B(_04419_),
    .C(_15614_),
    .Y(_04420_));
 INVx1_ASAP7_75t_R _23368_ (.A(_01327_),
    .Y(_04421_));
 NAND2x1_ASAP7_75t_R _23369_ (.A(_15617_),
    .B(_01325_),
    .Y(_04422_));
 OA211x2_ASAP7_75t_R _23370_ (.A1(_15610_),
    .A2(_04421_),
    .B(_04422_),
    .C(_15544_),
    .Y(_04423_));
 OR3x1_ASAP7_75t_R _23371_ (.A(_15547_),
    .B(_04420_),
    .C(_04423_),
    .Y(_04424_));
 OA21x2_ASAP7_75t_R _23372_ (.A1(_15499_),
    .A2(_04417_),
    .B(_04424_),
    .Y(_04425_));
 INVx1_ASAP7_75t_R _23373_ (.A(_01324_),
    .Y(_04426_));
 NAND2x1_ASAP7_75t_R _23374_ (.A(_15570_),
    .B(_01322_),
    .Y(_04427_));
 OA211x2_ASAP7_75t_R _23375_ (.A1(_15749_),
    .A2(_04426_),
    .B(_04427_),
    .C(net22),
    .Y(_04428_));
 INVx1_ASAP7_75t_R _23376_ (.A(_01323_),
    .Y(_04429_));
 NAND2x1_ASAP7_75t_R _23377_ (.A(_16422_),
    .B(_01321_),
    .Y(_04430_));
 OA211x2_ASAP7_75t_R _23378_ (.A1(_16420_),
    .A2(_04429_),
    .B(_04430_),
    .C(_15619_),
    .Y(_04431_));
 OR3x1_ASAP7_75t_R _23379_ (.A(_15608_),
    .B(_04428_),
    .C(_04431_),
    .Y(_04432_));
 INVx2_ASAP7_75t_R _23380_ (.A(_01332_),
    .Y(_04433_));
 NAND2x1_ASAP7_75t_R _23381_ (.A(_16422_),
    .B(_01330_),
    .Y(_04434_));
 OA211x2_ASAP7_75t_R _23382_ (.A1(_16420_),
    .A2(_04433_),
    .B(_04434_),
    .C(net22),
    .Y(_04435_));
 INVx1_ASAP7_75t_R _23383_ (.A(_01331_),
    .Y(_04436_));
 NAND2x1_ASAP7_75t_R _23384_ (.A(_16422_),
    .B(_01329_),
    .Y(_04437_));
 OA211x2_ASAP7_75t_R _23385_ (.A1(_16420_),
    .A2(_04436_),
    .B(_04437_),
    .C(_16309_),
    .Y(_04438_));
 OR3x1_ASAP7_75t_R _23386_ (.A(_15512_),
    .B(_04435_),
    .C(_04438_),
    .Y(_04439_));
 AND3x1_ASAP7_75t_R _23387_ (.A(_15607_),
    .B(_04432_),
    .C(_04439_),
    .Y(_04440_));
 AO21x1_ASAP7_75t_R _23388_ (.A1(_15747_),
    .A2(_04425_),
    .B(_04440_),
    .Y(_04441_));
 INVx1_ASAP7_75t_R _23389_ (.A(_01340_),
    .Y(_04442_));
 NAND2x1_ASAP7_75t_R _23390_ (.A(_15665_),
    .B(_01338_),
    .Y(_04443_));
 OA211x2_ASAP7_75t_R _23391_ (.A1(_15587_),
    .A2(_04442_),
    .B(_04443_),
    .C(_15519_),
    .Y(_04444_));
 INVx1_ASAP7_75t_R _23392_ (.A(_01339_),
    .Y(_04445_));
 NAND2x1_ASAP7_75t_R _23393_ (.A(_15665_),
    .B(_01337_),
    .Y(_04446_));
 OA211x2_ASAP7_75t_R _23394_ (.A1(net5),
    .A2(_04445_),
    .B(_04446_),
    .C(_15811_),
    .Y(_04447_));
 OR3x1_ASAP7_75t_R _23395_ (.A(_15498_),
    .B(_04444_),
    .C(_04447_),
    .Y(_04448_));
 INVx2_ASAP7_75t_R _23396_ (.A(_01348_),
    .Y(_04449_));
 NAND2x1_ASAP7_75t_R _23397_ (.A(_15665_),
    .B(_01346_),
    .Y(_04450_));
 OA211x2_ASAP7_75t_R _23398_ (.A1(net5),
    .A2(_04449_),
    .B(_04450_),
    .C(_15807_),
    .Y(_04451_));
 INVx2_ASAP7_75t_R _23399_ (.A(_01347_),
    .Y(_04452_));
 NAND2x1_ASAP7_75t_R _23400_ (.A(_15665_),
    .B(_01345_),
    .Y(_04453_));
 OA211x2_ASAP7_75t_R _23401_ (.A1(net5),
    .A2(_04452_),
    .B(_04453_),
    .C(_15811_),
    .Y(_04454_));
 OR3x1_ASAP7_75t_R _23402_ (.A(_15567_),
    .B(_04451_),
    .C(_04454_),
    .Y(_04455_));
 AND3x1_ASAP7_75t_R _23403_ (.A(_15887_),
    .B(_04448_),
    .C(_04455_),
    .Y(_04456_));
 INVx1_ASAP7_75t_R _23404_ (.A(_01341_),
    .Y(_04457_));
 NOR2x1_ASAP7_75t_R _23405_ (.A(_16046_),
    .B(_01343_),
    .Y(_04458_));
 AO21x1_ASAP7_75t_R _23406_ (.A1(_15577_),
    .A2(_04457_),
    .B(_04458_),
    .Y(_04459_));
 INVx2_ASAP7_75t_R _23407_ (.A(_01344_),
    .Y(_04460_));
 NAND2x1_ASAP7_75t_R _23408_ (.A(_15516_),
    .B(_01342_),
    .Y(_04461_));
 OA211x2_ASAP7_75t_R _23409_ (.A1(_15513_),
    .A2(_04460_),
    .B(_04461_),
    .C(_15519_),
    .Y(_04462_));
 AO21x1_ASAP7_75t_R _23410_ (.A1(_15931_),
    .A2(_04459_),
    .B(_04462_),
    .Y(_04463_));
 INVx1_ASAP7_75t_R _23411_ (.A(_01336_),
    .Y(_04464_));
 NAND2x1_ASAP7_75t_R _23412_ (.A(_15748_),
    .B(_01334_),
    .Y(_04465_));
 OA211x2_ASAP7_75t_R _23413_ (.A1(_15579_),
    .A2(_04464_),
    .B(_04465_),
    .C(_16153_),
    .Y(_04466_));
 INVx2_ASAP7_75t_R _23414_ (.A(_01335_),
    .Y(_04467_));
 NAND2x1_ASAP7_75t_R _23415_ (.A(_16151_),
    .B(_01333_),
    .Y(_04468_));
 OA211x2_ASAP7_75t_R _23416_ (.A1(_16149_),
    .A2(_04467_),
    .B(_04468_),
    .C(_15930_),
    .Y(_04469_));
 OR3x1_ASAP7_75t_R _23417_ (.A(_15869_),
    .B(_04466_),
    .C(_04469_),
    .Y(_04470_));
 OA211x2_ASAP7_75t_R _23418_ (.A1(_15929_),
    .A2(_04463_),
    .B(_04470_),
    .C(_16159_),
    .Y(_04471_));
 OR3x1_ASAP7_75t_R _23419_ (.A(_15912_),
    .B(_04456_),
    .C(_04471_),
    .Y(_04472_));
 OAI21x1_ASAP7_75t_R _23420_ (.A1(_15745_),
    .A2(_04441_),
    .B(_04472_),
    .Y(_04473_));
 OA211x2_ASAP7_75t_R _23421_ (.A1(_13578_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_04474_));
 AOI21x1_ASAP7_75t_R _23422_ (.A1(_16532_),
    .A2(_04473_),
    .B(_04474_),
    .Y(_18748_));
 AND2x2_ASAP7_75t_R _23423_ (.A(_15138_),
    .B(_01794_),
    .Y(_04475_));
 AO21x1_ASAP7_75t_R _23424_ (.A1(_13777_),
    .A2(_01320_),
    .B(_04475_),
    .Y(_04476_));
 OAI22x1_ASAP7_75t_R _23425_ (.A1(_01319_),
    .A2(_13858_),
    .B1(_04476_),
    .B2(_14990_),
    .Y(_04477_));
 NAND2x1_ASAP7_75t_R _23426_ (.A(_13925_),
    .B(_01326_),
    .Y(_04478_));
 OA211x2_ASAP7_75t_R _23427_ (.A1(_13924_),
    .A2(_04418_),
    .B(_04478_),
    .C(_13927_),
    .Y(_04479_));
 NAND2x1_ASAP7_75t_R _23428_ (.A(_14743_),
    .B(_01325_),
    .Y(_04480_));
 OA211x2_ASAP7_75t_R _23429_ (.A1(_15006_),
    .A2(_04421_),
    .B(_04480_),
    .C(_15009_),
    .Y(_04481_));
 OR3x1_ASAP7_75t_R _23430_ (.A(_15031_),
    .B(_04479_),
    .C(_04481_),
    .Y(_04482_));
 OA211x2_ASAP7_75t_R _23431_ (.A1(_13857_),
    .A2(_04477_),
    .B(_04482_),
    .C(_15038_),
    .Y(_04483_));
 NAND2x1_ASAP7_75t_R _23432_ (.A(_15358_),
    .B(_01322_),
    .Y(_04484_));
 OA211x2_ASAP7_75t_R _23433_ (.A1(_15992_),
    .A2(_04426_),
    .B(_04484_),
    .C(_15854_),
    .Y(_04485_));
 NAND2x1_ASAP7_75t_R _23434_ (.A(_13860_),
    .B(_01321_),
    .Y(_04486_));
 OA211x2_ASAP7_75t_R _23435_ (.A1(_15992_),
    .A2(_04429_),
    .B(_04486_),
    .C(_15969_),
    .Y(_04487_));
 OR3x1_ASAP7_75t_R _23436_ (.A(_14815_),
    .B(_04485_),
    .C(_04487_),
    .Y(_04488_));
 NAND2x1_ASAP7_75t_R _23437_ (.A(_13750_),
    .B(_01330_),
    .Y(_04489_));
 OA211x2_ASAP7_75t_R _23438_ (.A1(_15992_),
    .A2(_04433_),
    .B(_04489_),
    .C(_15854_),
    .Y(_04490_));
 NAND2x1_ASAP7_75t_R _23439_ (.A(_13860_),
    .B(_01329_),
    .Y(_04491_));
 OA211x2_ASAP7_75t_R _23440_ (.A1(_15964_),
    .A2(_04436_),
    .B(_04491_),
    .C(_15969_),
    .Y(_04492_));
 OR3x1_ASAP7_75t_R _23441_ (.A(_13748_),
    .B(_04490_),
    .C(_04492_),
    .Y(_04493_));
 AND3x2_ASAP7_75t_R _23442_ (.A(_14732_),
    .B(_04488_),
    .C(_04493_),
    .Y(_04494_));
 OR3x4_ASAP7_75t_R _23443_ (.A(_14733_),
    .B(_04483_),
    .C(_04494_),
    .Y(_04495_));
 NAND2x1_ASAP7_75t_R _23444_ (.A(_15358_),
    .B(_01338_),
    .Y(_04496_));
 OA211x2_ASAP7_75t_R _23445_ (.A1(_15992_),
    .A2(_04442_),
    .B(_04496_),
    .C(_15854_),
    .Y(_04497_));
 NAND2x1_ASAP7_75t_R _23446_ (.A(_13750_),
    .B(_01337_),
    .Y(_04498_));
 OA211x2_ASAP7_75t_R _23447_ (.A1(_15992_),
    .A2(_04445_),
    .B(_04498_),
    .C(_15969_),
    .Y(_04499_));
 OR3x1_ASAP7_75t_R _23448_ (.A(_14815_),
    .B(_04497_),
    .C(_04499_),
    .Y(_04500_));
 NAND2x1_ASAP7_75t_R _23449_ (.A(_13750_),
    .B(_01346_),
    .Y(_04501_));
 OA211x2_ASAP7_75t_R _23450_ (.A1(_15992_),
    .A2(_04449_),
    .B(_04501_),
    .C(_15854_),
    .Y(_04502_));
 NAND2x1_ASAP7_75t_R _23451_ (.A(_13860_),
    .B(_01345_),
    .Y(_04503_));
 OA211x2_ASAP7_75t_R _23452_ (.A1(_15992_),
    .A2(_04452_),
    .B(_04503_),
    .C(_15969_),
    .Y(_04504_));
 OR3x1_ASAP7_75t_R _23453_ (.A(_13748_),
    .B(_04502_),
    .C(_04504_),
    .Y(_04505_));
 AND3x1_ASAP7_75t_R _23454_ (.A(_14732_),
    .B(_04500_),
    .C(_04505_),
    .Y(_04506_));
 NOR2x1_ASAP7_75t_R _23455_ (.A(_15712_),
    .B(_01343_),
    .Y(_04507_));
 AO21x1_ASAP7_75t_R _23456_ (.A1(_14011_),
    .A2(_04457_),
    .B(_04507_),
    .Y(_04508_));
 NAND2x1_ASAP7_75t_R _23457_ (.A(_15290_),
    .B(_01342_),
    .Y(_04509_));
 OA211x2_ASAP7_75t_R _23458_ (.A1(_13920_),
    .A2(_04460_),
    .B(_04509_),
    .C(_13945_),
    .Y(_04510_));
 AO21x1_ASAP7_75t_R _23459_ (.A1(_13863_),
    .A2(_04508_),
    .B(_04510_),
    .Y(_04511_));
 NAND2x1_ASAP7_75t_R _23460_ (.A(_14938_),
    .B(_01334_),
    .Y(_04512_));
 OA211x2_ASAP7_75t_R _23461_ (.A1(_15042_),
    .A2(_04464_),
    .B(_04512_),
    .C(_13906_),
    .Y(_04513_));
 NAND2x1_ASAP7_75t_R _23462_ (.A(_14945_),
    .B(_01333_),
    .Y(_04514_));
 OA211x2_ASAP7_75t_R _23463_ (.A1(_13881_),
    .A2(_04467_),
    .B(_04514_),
    .C(_13890_),
    .Y(_04515_));
 OR3x1_ASAP7_75t_R _23464_ (.A(_15039_),
    .B(_04513_),
    .C(_04515_),
    .Y(_04516_));
 OA211x2_ASAP7_75t_R _23465_ (.A1(_13903_),
    .A2(_04511_),
    .B(_04516_),
    .C(_15038_),
    .Y(_04517_));
 OR3x4_ASAP7_75t_R _23466_ (.A(_15025_),
    .B(_04506_),
    .C(_04517_),
    .Y(_04518_));
 INVx2_ASAP7_75t_R _23467_ (.A(_00063_),
    .Y(_04519_));
 OA211x2_ASAP7_75t_R _23468_ (.A1(_15114_),
    .A2(_15115_),
    .B(_04519_),
    .C(_13367_),
    .Y(_04520_));
 AO31x2_ASAP7_75t_R _23469_ (.A1(_13660_),
    .A2(_04495_),
    .A3(_04518_),
    .B(_04520_),
    .Y(_04521_));
 BUFx3_ASAP7_75t_R _23470_ (.A(_13642_),
    .Y(_04522_));
 INVx1_ASAP7_75t_R _23471_ (.A(_01523_),
    .Y(_04523_));
 AO32x1_ASAP7_75t_R _23472_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_04521_),
    .B1(_04522_),
    .B2(_04523_),
    .Y(_04524_));
 BUFx4f_ASAP7_75t_R _23473_ (.A(_04524_),
    .Y(_18747_));
 INVx1_ASAP7_75t_R _23474_ (.A(_18747_),
    .Y(_18749_));
 AND2x2_ASAP7_75t_R _23475_ (.A(_15587_),
    .B(_01793_),
    .Y(_04525_));
 AO21x1_ASAP7_75t_R _23476_ (.A1(_15502_),
    .A2(_01353_),
    .B(_04525_),
    .Y(_04526_));
 OAI22x1_ASAP7_75t_R _23477_ (.A1(_01352_),
    .A2(_15500_),
    .B1(_04526_),
    .B2(_15510_),
    .Y(_04527_));
 INVx1_ASAP7_75t_R _23478_ (.A(_01361_),
    .Y(_04528_));
 NAND2x1_ASAP7_75t_R _23479_ (.A(_15872_),
    .B(_01359_),
    .Y(_04529_));
 OA211x2_ASAP7_75t_R _23480_ (.A1(_15586_),
    .A2(_04528_),
    .B(_04529_),
    .C(net21),
    .Y(_04530_));
 INVx1_ASAP7_75t_R _23481_ (.A(_01360_),
    .Y(_04531_));
 NAND2x1_ASAP7_75t_R _23482_ (.A(_15872_),
    .B(_01358_),
    .Y(_04532_));
 OA211x2_ASAP7_75t_R _23483_ (.A1(_15573_),
    .A2(_04531_),
    .B(_04532_),
    .C(_16309_),
    .Y(_04533_));
 OR3x1_ASAP7_75t_R _23484_ (.A(_15512_),
    .B(_04530_),
    .C(_04533_),
    .Y(_04534_));
 OA211x2_ASAP7_75t_R _23485_ (.A1(_15499_),
    .A2(_04527_),
    .B(_04534_),
    .C(_15526_),
    .Y(_04535_));
 INVx1_ASAP7_75t_R _23486_ (.A(_01357_),
    .Y(_04536_));
 NAND2x1_ASAP7_75t_R _23487_ (.A(_15767_),
    .B(_01355_),
    .Y(_04537_));
 OA211x2_ASAP7_75t_R _23488_ (.A1(_15765_),
    .A2(_04536_),
    .B(_04537_),
    .C(_15581_),
    .Y(_04538_));
 INVx1_ASAP7_75t_R _23489_ (.A(_01356_),
    .Y(_04539_));
 NAND2x1_ASAP7_75t_R _23490_ (.A(_15579_),
    .B(_01354_),
    .Y(_04540_));
 OA211x2_ASAP7_75t_R _23491_ (.A1(_15765_),
    .A2(_04539_),
    .B(_04540_),
    .C(_15648_),
    .Y(_04541_));
 OR3x1_ASAP7_75t_R _23492_ (.A(_15531_),
    .B(_04538_),
    .C(_04541_),
    .Y(_04542_));
 INVx1_ASAP7_75t_R _23493_ (.A(_01365_),
    .Y(_04543_));
 NAND2x1_ASAP7_75t_R _23494_ (.A(_15767_),
    .B(_01363_),
    .Y(_04544_));
 OA211x2_ASAP7_75t_R _23495_ (.A1(_15765_),
    .A2(_04543_),
    .B(_04544_),
    .C(_15581_),
    .Y(_04545_));
 INVx1_ASAP7_75t_R _23496_ (.A(_01364_),
    .Y(_04546_));
 NAND2x1_ASAP7_75t_R _23497_ (.A(_15579_),
    .B(_01362_),
    .Y(_04547_));
 OA211x2_ASAP7_75t_R _23498_ (.A1(_15577_),
    .A2(_04546_),
    .B(_04547_),
    .C(_15648_),
    .Y(_04548_));
 OR3x1_ASAP7_75t_R _23499_ (.A(_15753_),
    .B(_04545_),
    .C(_04548_),
    .Y(_04549_));
 AND3x1_ASAP7_75t_R _23500_ (.A(_15529_),
    .B(_04542_),
    .C(_04549_),
    .Y(_04550_));
 OR3x4_ASAP7_75t_R _23501_ (.A(_15745_),
    .B(_04535_),
    .C(_04550_),
    .Y(_04551_));
 INVx1_ASAP7_75t_R _23502_ (.A(_01373_),
    .Y(_04552_));
 NAND2x1_ASAP7_75t_R _23503_ (.A(_16540_),
    .B(_01371_),
    .Y(_04553_));
 OA211x2_ASAP7_75t_R _23504_ (.A1(_15602_),
    .A2(_04552_),
    .B(_04553_),
    .C(_15581_),
    .Y(_04554_));
 INVx1_ASAP7_75t_R _23505_ (.A(_01372_),
    .Y(_04555_));
 NAND2x1_ASAP7_75t_R _23506_ (.A(_16540_),
    .B(_01370_),
    .Y(_04556_));
 OA211x2_ASAP7_75t_R _23507_ (.A1(_15765_),
    .A2(_04555_),
    .B(_04556_),
    .C(_15648_),
    .Y(_04557_));
 OR3x1_ASAP7_75t_R _23508_ (.A(_15531_),
    .B(_04554_),
    .C(_04557_),
    .Y(_04558_));
 INVx1_ASAP7_75t_R _23509_ (.A(_01381_),
    .Y(_04559_));
 NAND2x1_ASAP7_75t_R _23510_ (.A(_16540_),
    .B(_01379_),
    .Y(_04560_));
 OA211x2_ASAP7_75t_R _23511_ (.A1(_15765_),
    .A2(_04559_),
    .B(_04560_),
    .C(_15581_),
    .Y(_04561_));
 INVx2_ASAP7_75t_R _23512_ (.A(_01380_),
    .Y(_04562_));
 NAND2x1_ASAP7_75t_R _23513_ (.A(_16540_),
    .B(_01378_),
    .Y(_04563_));
 OA211x2_ASAP7_75t_R _23514_ (.A1(_15765_),
    .A2(_04562_),
    .B(_04563_),
    .C(_15648_),
    .Y(_04564_));
 OR3x1_ASAP7_75t_R _23515_ (.A(_15753_),
    .B(_04561_),
    .C(_04564_),
    .Y(_04565_));
 AND3x1_ASAP7_75t_R _23516_ (.A(_15529_),
    .B(_04558_),
    .C(_04565_),
    .Y(_04566_));
 INVx1_ASAP7_75t_R _23517_ (.A(_01374_),
    .Y(_04567_));
 NOR2x1_ASAP7_75t_R _23518_ (.A(_15625_),
    .B(_01376_),
    .Y(_04568_));
 AO21x1_ASAP7_75t_R _23519_ (.A1(_16650_),
    .A2(_04567_),
    .B(_04568_),
    .Y(_04569_));
 INVx1_ASAP7_75t_R _23520_ (.A(_01377_),
    .Y(_04570_));
 NAND2x1_ASAP7_75t_R _23521_ (.A(_15756_),
    .B(_01375_),
    .Y(_04571_));
 OA211x2_ASAP7_75t_R _23522_ (.A1(_15602_),
    .A2(_04570_),
    .B(_04571_),
    .C(net19),
    .Y(_04572_));
 AO21x1_ASAP7_75t_R _23523_ (.A1(_15569_),
    .A2(_04569_),
    .B(_04572_),
    .Y(_04573_));
 INVx1_ASAP7_75t_R _23524_ (.A(_01369_),
    .Y(_04574_));
 NAND2x1_ASAP7_75t_R _23525_ (.A(_16422_),
    .B(_01367_),
    .Y(_04575_));
 OA211x2_ASAP7_75t_R _23526_ (.A1(_16420_),
    .A2(_04574_),
    .B(_04575_),
    .C(net22),
    .Y(_04576_));
 INVx2_ASAP7_75t_R _23527_ (.A(_01368_),
    .Y(_04577_));
 NAND2x1_ASAP7_75t_R _23528_ (.A(_15872_),
    .B(_01366_),
    .Y(_04578_));
 OA211x2_ASAP7_75t_R _23529_ (.A1(_15586_),
    .A2(_04577_),
    .B(_04578_),
    .C(_16309_),
    .Y(_04579_));
 OR3x1_ASAP7_75t_R _23530_ (.A(_15608_),
    .B(_04576_),
    .C(_04579_),
    .Y(_04580_));
 OA211x2_ASAP7_75t_R _23531_ (.A1(_15568_),
    .A2(_04573_),
    .B(_04580_),
    .C(_15526_),
    .Y(_04581_));
 OR3x4_ASAP7_75t_R _23532_ (.A(_15555_),
    .B(_04566_),
    .C(_04581_),
    .Y(_04582_));
 NAND2x2_ASAP7_75t_R _23533_ (.A(_04551_),
    .B(_04582_),
    .Y(_04583_));
 OA211x2_ASAP7_75t_R _23534_ (.A1(_13577_),
    .A2(_16594_),
    .B(_15490_),
    .C(_16596_),
    .Y(_04584_));
 AOI21x1_ASAP7_75t_R _23535_ (.A1(_16532_),
    .A2(_04583_),
    .B(_04584_),
    .Y(_18753_));
 AND2x2_ASAP7_75t_R _23536_ (.A(_15138_),
    .B(_01793_),
    .Y(_04585_));
 AO21x1_ASAP7_75t_R _23537_ (.A1(_13777_),
    .A2(_01353_),
    .B(_04585_),
    .Y(_04586_));
 OAI22x1_ASAP7_75t_R _23538_ (.A1(_01352_),
    .A2(_13858_),
    .B1(_04586_),
    .B2(_14990_),
    .Y(_04587_));
 NAND2x1_ASAP7_75t_R _23539_ (.A(_14854_),
    .B(_01359_),
    .Y(_04588_));
 OA211x2_ASAP7_75t_R _23540_ (.A1(_15319_),
    .A2(_04528_),
    .B(_04588_),
    .C(_15686_),
    .Y(_04589_));
 NAND2x1_ASAP7_75t_R _23541_ (.A(_14848_),
    .B(_01358_),
    .Y(_04590_));
 OA211x2_ASAP7_75t_R _23542_ (.A1(_15207_),
    .A2(_04531_),
    .B(_04590_),
    .C(_15689_),
    .Y(_04591_));
 OR3x1_ASAP7_75t_R _23543_ (.A(_15031_),
    .B(_04589_),
    .C(_04591_),
    .Y(_04592_));
 OA211x2_ASAP7_75t_R _23544_ (.A1(_13857_),
    .A2(_04587_),
    .B(_04592_),
    .C(_15038_),
    .Y(_04593_));
 NAND2x1_ASAP7_75t_R _23545_ (.A(_15126_),
    .B(_01355_),
    .Y(_04594_));
 OA211x2_ASAP7_75t_R _23546_ (.A1(_13920_),
    .A2(_04536_),
    .B(_04594_),
    .C(_13945_),
    .Y(_04595_));
 NAND2x1_ASAP7_75t_R _23547_ (.A(_15131_),
    .B(_01354_),
    .Y(_04596_));
 OA211x2_ASAP7_75t_R _23548_ (.A1(_13920_),
    .A2(_04539_),
    .B(_04596_),
    .C(_13749_),
    .Y(_04597_));
 OR3x1_ASAP7_75t_R _23549_ (.A(_14815_),
    .B(_04595_),
    .C(_04597_),
    .Y(_04598_));
 NAND2x1_ASAP7_75t_R _23550_ (.A(_15131_),
    .B(_01363_),
    .Y(_04599_));
 OA211x2_ASAP7_75t_R _23551_ (.A1(_13920_),
    .A2(_04543_),
    .B(_04599_),
    .C(_13945_),
    .Y(_04600_));
 NAND2x1_ASAP7_75t_R _23552_ (.A(_15358_),
    .B(_01362_),
    .Y(_04601_));
 OA211x2_ASAP7_75t_R _23553_ (.A1(_15992_),
    .A2(_04546_),
    .B(_04601_),
    .C(_15969_),
    .Y(_04602_));
 OR3x1_ASAP7_75t_R _23554_ (.A(_13748_),
    .B(_04600_),
    .C(_04602_),
    .Y(_04603_));
 AND3x2_ASAP7_75t_R _23555_ (.A(_14732_),
    .B(_04598_),
    .C(_04603_),
    .Y(_04604_));
 OR3x4_ASAP7_75t_R _23556_ (.A(_14733_),
    .B(_04593_),
    .C(_04604_),
    .Y(_04605_));
 NAND2x1_ASAP7_75t_R _23557_ (.A(_15126_),
    .B(_01371_),
    .Y(_04606_));
 OA211x2_ASAP7_75t_R _23558_ (.A1(_13920_),
    .A2(_04552_),
    .B(_04606_),
    .C(_13945_),
    .Y(_04607_));
 NAND2x1_ASAP7_75t_R _23559_ (.A(_15131_),
    .B(_01370_),
    .Y(_04608_));
 OA211x2_ASAP7_75t_R _23560_ (.A1(_13920_),
    .A2(_04555_),
    .B(_04608_),
    .C(_13749_),
    .Y(_04609_));
 OR3x1_ASAP7_75t_R _23561_ (.A(_14815_),
    .B(_04607_),
    .C(_04609_),
    .Y(_04610_));
 NAND2x1_ASAP7_75t_R _23562_ (.A(_15131_),
    .B(_01379_),
    .Y(_04611_));
 OA211x2_ASAP7_75t_R _23563_ (.A1(_13920_),
    .A2(_04559_),
    .B(_04611_),
    .C(_13945_),
    .Y(_04612_));
 NAND2x1_ASAP7_75t_R _23564_ (.A(_15358_),
    .B(_01378_),
    .Y(_04613_));
 OA211x2_ASAP7_75t_R _23565_ (.A1(_15992_),
    .A2(_04562_),
    .B(_04613_),
    .C(_15969_),
    .Y(_04614_));
 OR3x1_ASAP7_75t_R _23566_ (.A(_13748_),
    .B(_04612_),
    .C(_04614_),
    .Y(_04615_));
 AND3x1_ASAP7_75t_R _23567_ (.A(_14732_),
    .B(_04610_),
    .C(_04615_),
    .Y(_04616_));
 NOR2x1_ASAP7_75t_R _23568_ (.A(_15712_),
    .B(_01376_),
    .Y(_04617_));
 AO21x1_ASAP7_75t_R _23569_ (.A1(_14011_),
    .A2(_04567_),
    .B(_04617_),
    .Y(_04618_));
 NAND2x1_ASAP7_75t_R _23570_ (.A(_13934_),
    .B(_01375_),
    .Y(_04619_));
 OA211x2_ASAP7_75t_R _23571_ (.A1(_14011_),
    .A2(_04570_),
    .B(_04619_),
    .C(_13945_),
    .Y(_04620_));
 AO21x1_ASAP7_75t_R _23572_ (.A1(_13863_),
    .A2(_04618_),
    .B(_04620_),
    .Y(_04621_));
 NAND2x1_ASAP7_75t_R _23573_ (.A(_14872_),
    .B(_01367_),
    .Y(_04622_));
 OA211x2_ASAP7_75t_R _23574_ (.A1(_15013_),
    .A2(_04574_),
    .B(_04622_),
    .C(_13927_),
    .Y(_04623_));
 NAND2x1_ASAP7_75t_R _23575_ (.A(_15019_),
    .B(_01366_),
    .Y(_04624_));
 OA211x2_ASAP7_75t_R _23576_ (.A1(_15017_),
    .A2(_04577_),
    .B(_04624_),
    .C(_13917_),
    .Y(_04625_));
 OR3x1_ASAP7_75t_R _23577_ (.A(_15039_),
    .B(_04623_),
    .C(_04625_),
    .Y(_04626_));
 OA211x2_ASAP7_75t_R _23578_ (.A1(_13903_),
    .A2(_04621_),
    .B(_04626_),
    .C(_15038_),
    .Y(_04627_));
 OR3x4_ASAP7_75t_R _23579_ (.A(_15025_),
    .B(_04616_),
    .C(_04627_),
    .Y(_04628_));
 INVx1_ASAP7_75t_R _23580_ (.A(_00064_),
    .Y(_04629_));
 OA211x2_ASAP7_75t_R _23581_ (.A1(_15114_),
    .A2(_15115_),
    .B(_04629_),
    .C(_13367_),
    .Y(_04630_));
 AO31x2_ASAP7_75t_R _23582_ (.A1(_13660_),
    .A2(_04605_),
    .A3(_04628_),
    .B(_04630_),
    .Y(_04631_));
 INVx1_ASAP7_75t_R _23583_ (.A(_01522_),
    .Y(_04632_));
 AO32x1_ASAP7_75t_R _23584_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_04631_),
    .B1(_04522_),
    .B2(_04632_),
    .Y(_04633_));
 BUFx6f_ASAP7_75t_R _23585_ (.A(_04633_),
    .Y(_18752_));
 INVx1_ASAP7_75t_R _23586_ (.A(_18752_),
    .Y(_18754_));
 OA21x2_ASAP7_75t_R _23587_ (.A1(_01317_),
    .A2(_04400_),
    .B(_01351_),
    .Y(_04634_));
 OA21x2_ASAP7_75t_R _23588_ (.A1(_01350_),
    .A2(_04634_),
    .B(_01384_),
    .Y(_04635_));
 XOR2x2_ASAP7_75t_R _23589_ (.A(_01383_),
    .B(_04635_),
    .Y(\alu_adder_result_ex[29] ));
 OA31x2_ASAP7_75t_R _23590_ (.A1(_01284_),
    .A2(_04408_),
    .A3(_04411_),
    .B1(_01318_),
    .Y(_04636_));
 OA21x2_ASAP7_75t_R _23591_ (.A1(_01317_),
    .A2(_04636_),
    .B(_01351_),
    .Y(_04637_));
 XOR2x2_ASAP7_75t_R _23592_ (.A(_01350_),
    .B(_04637_),
    .Y(_04638_));
 BUFx12_ASAP7_75t_R _23593_ (.A(_04638_),
    .Y(\alu_adder_result_ex[28] ));
 AND2x2_ASAP7_75t_R _23594_ (.A(_15579_),
    .B(_01791_),
    .Y(_04639_));
 AO21x1_ASAP7_75t_R _23595_ (.A1(_15871_),
    .A2(_01386_),
    .B(_04639_),
    .Y(_04640_));
 OAI22x1_ASAP7_75t_R _23596_ (.A1(_01385_),
    .A2(_15500_),
    .B1(_04640_),
    .B2(_15569_),
    .Y(_04641_));
 INVx1_ASAP7_75t_R _23597_ (.A(_01394_),
    .Y(_04642_));
 NAND2x1_ASAP7_75t_R _23598_ (.A(_15516_),
    .B(_01392_),
    .Y(_04643_));
 OA211x2_ASAP7_75t_R _23599_ (.A1(_15587_),
    .A2(_04642_),
    .B(_04643_),
    .C(_15519_),
    .Y(_04644_));
 INVx1_ASAP7_75t_R _23600_ (.A(_01393_),
    .Y(_04645_));
 NAND2x1_ASAP7_75t_R _23601_ (.A(_15602_),
    .B(_01391_),
    .Y(_04646_));
 OA211x2_ASAP7_75t_R _23602_ (.A1(_15587_),
    .A2(_04645_),
    .B(_04646_),
    .C(_15523_),
    .Y(_04647_));
 OR3x1_ASAP7_75t_R _23603_ (.A(_15567_),
    .B(_04644_),
    .C(_04647_),
    .Y(_04648_));
 OA21x2_ASAP7_75t_R _23604_ (.A1(_15870_),
    .A2(_04641_),
    .B(_04648_),
    .Y(_04649_));
 INVx2_ASAP7_75t_R _23605_ (.A(_01390_),
    .Y(_04650_));
 NAND2x1_ASAP7_75t_R _23606_ (.A(_15936_),
    .B(_01388_),
    .Y(_04651_));
 OA211x2_ASAP7_75t_R _23607_ (.A1(_15505_),
    .A2(_04650_),
    .B(_04651_),
    .C(_15807_),
    .Y(_04652_));
 INVx1_ASAP7_75t_R _23608_ (.A(_01389_),
    .Y(_04653_));
 NAND2x1_ASAP7_75t_R _23609_ (.A(_15936_),
    .B(_01387_),
    .Y(_04654_));
 OA211x2_ASAP7_75t_R _23610_ (.A1(_15594_),
    .A2(_04653_),
    .B(_04654_),
    .C(_15918_),
    .Y(_04655_));
 OR3x1_ASAP7_75t_R _23611_ (.A(_15888_),
    .B(_04652_),
    .C(_04655_),
    .Y(_04656_));
 INVx2_ASAP7_75t_R _23612_ (.A(_01398_),
    .Y(_04657_));
 NAND2x1_ASAP7_75t_R _23613_ (.A(_15936_),
    .B(_01396_),
    .Y(_04658_));
 OA211x2_ASAP7_75t_R _23614_ (.A1(_15594_),
    .A2(_04657_),
    .B(_04658_),
    .C(_16082_),
    .Y(_04659_));
 INVx1_ASAP7_75t_R _23615_ (.A(_01397_),
    .Y(_04660_));
 NAND2x1_ASAP7_75t_R _23616_ (.A(_15936_),
    .B(_01395_),
    .Y(_04661_));
 OA211x2_ASAP7_75t_R _23617_ (.A1(_15594_),
    .A2(_04660_),
    .B(_04661_),
    .C(_15918_),
    .Y(_04662_));
 OR3x1_ASAP7_75t_R _23618_ (.A(_15567_),
    .B(_04659_),
    .C(_04662_),
    .Y(_04663_));
 AND3x1_ASAP7_75t_R _23619_ (.A(_15887_),
    .B(_04656_),
    .C(_04663_),
    .Y(_04664_));
 AO21x1_ASAP7_75t_R _23620_ (.A1(_15747_),
    .A2(_04649_),
    .B(_04664_),
    .Y(_04665_));
 INVx1_ASAP7_75t_R _23621_ (.A(_01406_),
    .Y(_04666_));
 NAND2x1_ASAP7_75t_R _23622_ (.A(_15748_),
    .B(_01404_),
    .Y(_04667_));
 OA211x2_ASAP7_75t_R _23623_ (.A1(_15767_),
    .A2(_04666_),
    .B(_04667_),
    .C(_16044_),
    .Y(_04668_));
 INVx1_ASAP7_75t_R _23624_ (.A(_01405_),
    .Y(_04669_));
 NAND2x1_ASAP7_75t_R _23625_ (.A(_15748_),
    .B(_01403_),
    .Y(_04670_));
 OA211x2_ASAP7_75t_R _23626_ (.A1(_15767_),
    .A2(_04669_),
    .B(_04670_),
    .C(_15930_),
    .Y(_04671_));
 OR3x1_ASAP7_75t_R _23627_ (.A(_15869_),
    .B(_04668_),
    .C(_04671_),
    .Y(_04672_));
 INVx2_ASAP7_75t_R _23628_ (.A(_01414_),
    .Y(_04673_));
 NAND2x1_ASAP7_75t_R _23629_ (.A(_15748_),
    .B(_01412_),
    .Y(_04674_));
 OA211x2_ASAP7_75t_R _23630_ (.A1(_15767_),
    .A2(_04673_),
    .B(_04674_),
    .C(_16153_),
    .Y(_04675_));
 INVx1_ASAP7_75t_R _23631_ (.A(_01413_),
    .Y(_04676_));
 NAND2x1_ASAP7_75t_R _23632_ (.A(_15748_),
    .B(_01411_),
    .Y(_04677_));
 OA211x2_ASAP7_75t_R _23633_ (.A1(_15579_),
    .A2(_04676_),
    .B(_04677_),
    .C(_15930_),
    .Y(_04678_));
 OR3x1_ASAP7_75t_R _23634_ (.A(_15876_),
    .B(_04675_),
    .C(_04678_),
    .Y(_04679_));
 AND3x1_ASAP7_75t_R _23635_ (.A(_15528_),
    .B(_04672_),
    .C(_04679_),
    .Y(_04680_));
 INVx1_ASAP7_75t_R _23636_ (.A(_01407_),
    .Y(_04681_));
 NOR2x1_ASAP7_75t_R _23637_ (.A(_15570_),
    .B(_01409_),
    .Y(_04682_));
 AO21x1_ASAP7_75t_R _23638_ (.A1(_15652_),
    .A2(_04681_),
    .B(_04682_),
    .Y(_04683_));
 INVx2_ASAP7_75t_R _23639_ (.A(_01410_),
    .Y(_04684_));
 NAND2x1_ASAP7_75t_R _23640_ (.A(_16048_),
    .B(_01408_),
    .Y(_04685_));
 OA211x2_ASAP7_75t_R _23641_ (.A1(_16046_),
    .A2(_04684_),
    .B(_04685_),
    .C(_16044_),
    .Y(_04686_));
 AO21x1_ASAP7_75t_R _23642_ (.A1(_15931_),
    .A2(_04683_),
    .B(_04686_),
    .Y(_04687_));
 INVx2_ASAP7_75t_R _23643_ (.A(_01402_),
    .Y(_04688_));
 NAND2x1_ASAP7_75t_R _23644_ (.A(net5),
    .B(_01400_),
    .Y(_04689_));
 OA211x2_ASAP7_75t_R _23645_ (.A1(_16303_),
    .A2(_04688_),
    .B(_04689_),
    .C(net18),
    .Y(_04690_));
 INVx2_ASAP7_75t_R _23646_ (.A(_01401_),
    .Y(_04691_));
 NAND2x1_ASAP7_75t_R _23647_ (.A(net5),
    .B(_01399_),
    .Y(_04692_));
 OA211x2_ASAP7_75t_R _23648_ (.A1(_16303_),
    .A2(_04691_),
    .B(_04692_),
    .C(_15945_),
    .Y(_04693_));
 OR3x1_ASAP7_75t_R _23649_ (.A(_15530_),
    .B(_04690_),
    .C(_04693_),
    .Y(_04694_));
 OA211x2_ASAP7_75t_R _23650_ (.A1(_15753_),
    .A2(_04687_),
    .B(_04694_),
    .C(_15746_),
    .Y(_04695_));
 OR3x1_ASAP7_75t_R _23651_ (.A(_15912_),
    .B(_04680_),
    .C(_04695_),
    .Y(_04696_));
 OAI21x1_ASAP7_75t_R _23652_ (.A1(_15745_),
    .A2(_04665_),
    .B(_04696_),
    .Y(_04697_));
 OA211x2_ASAP7_75t_R _23653_ (.A1(_13575_),
    .A2(_16593_),
    .B(_15490_),
    .C(_16595_),
    .Y(_04698_));
 AOI21x1_ASAP7_75t_R _23654_ (.A1(_15496_),
    .A2(_04697_),
    .B(_04698_),
    .Y(_18759_));
 AND2x2_ASAP7_75t_R _23655_ (.A(_13866_),
    .B(_01791_),
    .Y(_04699_));
 AO21x1_ASAP7_75t_R _23656_ (.A1(_13709_),
    .A2(_01386_),
    .B(_04699_),
    .Y(_04700_));
 OAI22x1_ASAP7_75t_R _23657_ (.A1(_01385_),
    .A2(_13948_),
    .B1(_04700_),
    .B2(_13918_),
    .Y(_04701_));
 NAND2x1_ASAP7_75t_R _23658_ (.A(_13964_),
    .B(_01392_),
    .Y(_04702_));
 OA211x2_ASAP7_75t_R _23659_ (.A1(_13919_),
    .A2(_04642_),
    .B(_04702_),
    .C(_13724_),
    .Y(_04703_));
 NAND2x1_ASAP7_75t_R _23660_ (.A(_13964_),
    .B(_01391_),
    .Y(_04704_));
 OA211x2_ASAP7_75t_R _23661_ (.A1(_13919_),
    .A2(_04645_),
    .B(_04704_),
    .C(_13744_),
    .Y(_04705_));
 OR3x1_ASAP7_75t_R _23662_ (.A(_13696_),
    .B(_04703_),
    .C(_04705_),
    .Y(_04706_));
 OA211x2_ASAP7_75t_R _23663_ (.A1(_14815_),
    .A2(_04701_),
    .B(_04706_),
    .C(_13961_),
    .Y(_04707_));
 NAND2x1_ASAP7_75t_R _23664_ (.A(_15424_),
    .B(_01388_),
    .Y(_04708_));
 OA211x2_ASAP7_75t_R _23665_ (.A1(_14831_),
    .A2(_04650_),
    .B(_04708_),
    .C(_15282_),
    .Y(_04709_));
 NAND2x1_ASAP7_75t_R _23666_ (.A(_15424_),
    .B(_01387_),
    .Y(_04710_));
 OA211x2_ASAP7_75t_R _23667_ (.A1(_15423_),
    .A2(_04653_),
    .B(_04710_),
    .C(_14754_),
    .Y(_04711_));
 OR3x1_ASAP7_75t_R _23668_ (.A(_14739_),
    .B(_04709_),
    .C(_04711_),
    .Y(_04712_));
 NAND2x1_ASAP7_75t_R _23669_ (.A(_15424_),
    .B(_01396_),
    .Y(_04713_));
 OA211x2_ASAP7_75t_R _23670_ (.A1(_15423_),
    .A2(_04657_),
    .B(_04713_),
    .C(_15282_),
    .Y(_04714_));
 NAND2x1_ASAP7_75t_R _23671_ (.A(_15280_),
    .B(_01395_),
    .Y(_04715_));
 OA211x2_ASAP7_75t_R _23672_ (.A1(_15278_),
    .A2(_04660_),
    .B(_04715_),
    .C(_14850_),
    .Y(_04716_));
 OR3x1_ASAP7_75t_R _23673_ (.A(_14853_),
    .B(_04714_),
    .C(_04716_),
    .Y(_04717_));
 AND3x1_ASAP7_75t_R _23674_ (.A(_14843_),
    .B(_04712_),
    .C(_04717_),
    .Y(_04718_));
 OR3x4_ASAP7_75t_R _23675_ (.A(_14814_),
    .B(_04707_),
    .C(_04718_),
    .Y(_04719_));
 NAND2x1_ASAP7_75t_R _23676_ (.A(_15424_),
    .B(_01404_),
    .Y(_04720_));
 OA211x2_ASAP7_75t_R _23677_ (.A1(_14831_),
    .A2(_04666_),
    .B(_04720_),
    .C(_15282_),
    .Y(_04721_));
 NAND2x1_ASAP7_75t_R _23678_ (.A(_15424_),
    .B(_01403_),
    .Y(_04722_));
 OA211x2_ASAP7_75t_R _23679_ (.A1(_15423_),
    .A2(_04669_),
    .B(_04722_),
    .C(_14754_),
    .Y(_04723_));
 OR3x1_ASAP7_75t_R _23680_ (.A(_14739_),
    .B(_04721_),
    .C(_04723_),
    .Y(_04724_));
 NAND2x1_ASAP7_75t_R _23681_ (.A(_15424_),
    .B(_01412_),
    .Y(_04725_));
 OA211x2_ASAP7_75t_R _23682_ (.A1(_15423_),
    .A2(_04673_),
    .B(_04725_),
    .C(_15282_),
    .Y(_04726_));
 NAND2x1_ASAP7_75t_R _23683_ (.A(_15280_),
    .B(_01411_),
    .Y(_04727_));
 OA211x2_ASAP7_75t_R _23684_ (.A1(_15423_),
    .A2(_04676_),
    .B(_04727_),
    .C(_14754_),
    .Y(_04728_));
 OR3x1_ASAP7_75t_R _23685_ (.A(_14748_),
    .B(_04726_),
    .C(_04728_),
    .Y(_04729_));
 AND3x1_ASAP7_75t_R _23686_ (.A(_14843_),
    .B(_04724_),
    .C(_04729_),
    .Y(_04730_));
 NOR2x1_ASAP7_75t_R _23687_ (.A(_13680_),
    .B(_01409_),
    .Y(_04731_));
 AO21x1_ASAP7_75t_R _23688_ (.A1(_15954_),
    .A2(_04681_),
    .B(_04731_),
    .Y(_04732_));
 NAND2x1_ASAP7_75t_R _23689_ (.A(_13711_),
    .B(_01408_),
    .Y(_04733_));
 OA211x2_ASAP7_75t_R _23690_ (.A1(_14749_),
    .A2(_04684_),
    .B(_04733_),
    .C(_14751_),
    .Y(_04734_));
 AO21x1_ASAP7_75t_R _23691_ (.A1(_13749_),
    .A2(_04732_),
    .B(_04734_),
    .Y(_04735_));
 NAND2x1_ASAP7_75t_R _23692_ (.A(_13964_),
    .B(_01400_),
    .Y(_04736_));
 OA211x2_ASAP7_75t_R _23693_ (.A1(_16872_),
    .A2(_04688_),
    .B(_04736_),
    .C(_13724_),
    .Y(_04737_));
 NAND2x1_ASAP7_75t_R _23694_ (.A(_13964_),
    .B(_01399_),
    .Y(_04738_));
 OA211x2_ASAP7_75t_R _23695_ (.A1(_16872_),
    .A2(_04691_),
    .B(_04738_),
    .C(_13744_),
    .Y(_04739_));
 OR3x1_ASAP7_75t_R _23696_ (.A(_13706_),
    .B(_04737_),
    .C(_04739_),
    .Y(_04740_));
 OA211x2_ASAP7_75t_R _23697_ (.A1(_13748_),
    .A2(_04735_),
    .B(_04740_),
    .C(_13961_),
    .Y(_04741_));
 OR3x4_ASAP7_75t_R _23698_ (.A(_14842_),
    .B(_04730_),
    .C(_04741_),
    .Y(_04742_));
 INVx1_ASAP7_75t_R _23699_ (.A(_00065_),
    .Y(_04743_));
 OA211x2_ASAP7_75t_R _23700_ (.A1(_13647_),
    .A2(_13658_),
    .B(_04743_),
    .C(_13366_),
    .Y(_04744_));
 AO31x2_ASAP7_75t_R _23701_ (.A1(_13947_),
    .A2(_04719_),
    .A3(_04742_),
    .B(_04744_),
    .Y(_04745_));
 INVx1_ASAP7_75t_R _23702_ (.A(_01520_),
    .Y(_04746_));
 AO32x1_ASAP7_75t_R _23703_ (.A1(_13771_),
    .A2(_13772_),
    .A3(_04745_),
    .B1(_13642_),
    .B2(_04746_),
    .Y(_04747_));
 BUFx6f_ASAP7_75t_R _23704_ (.A(_04747_),
    .Y(_18760_));
 INVx2_ASAP7_75t_R _23705_ (.A(_18760_),
    .Y(_18758_));
 AO32x1_ASAP7_75t_R _23706_ (.A1(_13435_),
    .A2(_13406_),
    .A3(_13412_),
    .B1(_13421_),
    .B2(_13428_),
    .Y(_04748_));
 AO21x2_ASAP7_75t_R _23707_ (.A1(_14058_),
    .A2(_04748_),
    .B(_13788_),
    .Y(_04749_));
 AND2x2_ASAP7_75t_R _23708_ (.A(net20),
    .B(_01790_),
    .Y(_04750_));
 AO21x1_ASAP7_75t_R _23709_ (.A1(_13390_),
    .A2(_01419_),
    .B(_04750_),
    .Y(_04751_));
 OAI22x1_ASAP7_75t_R _23710_ (.A1(_01418_),
    .A2(_13497_),
    .B1(_04751_),
    .B2(_13492_),
    .Y(_04752_));
 INVx1_ASAP7_75t_R _23711_ (.A(_01435_),
    .Y(_04753_));
 NAND2x1_ASAP7_75t_R _23712_ (.A(_13462_),
    .B(_01433_),
    .Y(_04754_));
 OA211x2_ASAP7_75t_R _23713_ (.A1(_13457_),
    .A2(_04753_),
    .B(_04754_),
    .C(_14117_),
    .Y(_04755_));
 INVx1_ASAP7_75t_R _23714_ (.A(_01434_),
    .Y(_04756_));
 NAND2x1_ASAP7_75t_R _23715_ (.A(_13462_),
    .B(_01432_),
    .Y(_04757_));
 OA211x2_ASAP7_75t_R _23716_ (.A1(_13457_),
    .A2(_04756_),
    .B(_04757_),
    .C(_13491_),
    .Y(_04758_));
 OR3x1_ASAP7_75t_R _23717_ (.A(_13517_),
    .B(_04755_),
    .C(_04758_),
    .Y(_04759_));
 OA211x2_ASAP7_75t_R _23718_ (.A1(_13447_),
    .A2(_04752_),
    .B(_04759_),
    .C(_13483_),
    .Y(_04760_));
 INVx1_ASAP7_75t_R _23719_ (.A(_01427_),
    .Y(_04761_));
 NAND2x1_ASAP7_75t_R _23720_ (.A(_14495_),
    .B(_01425_),
    .Y(_04762_));
 OA211x2_ASAP7_75t_R _23721_ (.A1(_13801_),
    .A2(_04761_),
    .B(_04762_),
    .C(net11),
    .Y(_04763_));
 INVx1_ASAP7_75t_R _23722_ (.A(_01426_),
    .Y(_04764_));
 NAND2x1_ASAP7_75t_R _23723_ (.A(_14495_),
    .B(_01424_),
    .Y(_04765_));
 OA211x2_ASAP7_75t_R _23724_ (.A1(net20),
    .A2(_04764_),
    .B(_04765_),
    .C(_13491_),
    .Y(_04766_));
 OR3x1_ASAP7_75t_R _23725_ (.A(_13446_),
    .B(_04763_),
    .C(_04766_),
    .Y(_04767_));
 INVx1_ASAP7_75t_R _23726_ (.A(_01443_),
    .Y(_04768_));
 NAND2x1_ASAP7_75t_R _23727_ (.A(_14495_),
    .B(_01441_),
    .Y(_04769_));
 OA211x2_ASAP7_75t_R _23728_ (.A1(net20),
    .A2(_04768_),
    .B(_04769_),
    .C(net11),
    .Y(_04770_));
 INVx1_ASAP7_75t_R _23729_ (.A(_01442_),
    .Y(_04771_));
 NAND2x1_ASAP7_75t_R _23730_ (.A(_14262_),
    .B(_01440_),
    .Y(_04772_));
 OA211x2_ASAP7_75t_R _23731_ (.A1(net20),
    .A2(_04771_),
    .B(_04772_),
    .C(_13491_),
    .Y(_04773_));
 OR3x1_ASAP7_75t_R _23732_ (.A(_13517_),
    .B(_04770_),
    .C(_04773_),
    .Y(_04774_));
 AND3x1_ASAP7_75t_R _23733_ (.A(_13453_),
    .B(_04767_),
    .C(_04774_),
    .Y(_04775_));
 INVx1_ASAP7_75t_R _23734_ (.A(_01439_),
    .Y(_04776_));
 NAND2x1_ASAP7_75t_R _23735_ (.A(_13472_),
    .B(_01437_),
    .Y(_04777_));
 OA211x2_ASAP7_75t_R _23736_ (.A1(_13502_),
    .A2(_04776_),
    .B(_04777_),
    .C(_13795_),
    .Y(_04778_));
 INVx1_ASAP7_75t_R _23737_ (.A(_01438_),
    .Y(_04779_));
 NAND2x1_ASAP7_75t_R _23738_ (.A(_13463_),
    .B(_01436_),
    .Y(_04780_));
 OA211x2_ASAP7_75t_R _23739_ (.A1(net12),
    .A2(_04779_),
    .B(_04780_),
    .C(_13478_),
    .Y(_04781_));
 OA21x2_ASAP7_75t_R _23740_ (.A1(_04778_),
    .A2(_04781_),
    .B(_14205_),
    .Y(_04782_));
 OR5x2_ASAP7_75t_R _23741_ (.A(_13451_),
    .B(_14373_),
    .C(_04760_),
    .D(_04775_),
    .E(_04782_),
    .Y(_04783_));
 INVx1_ASAP7_75t_R _23742_ (.A(_01431_),
    .Y(_04784_));
 NAND2x1_ASAP7_75t_R _23743_ (.A(_14110_),
    .B(_01429_),
    .Y(_04785_));
 OA211x2_ASAP7_75t_R _23744_ (.A1(_13801_),
    .A2(_04784_),
    .B(_04785_),
    .C(net11),
    .Y(_04786_));
 INVx1_ASAP7_75t_R _23745_ (.A(_01430_),
    .Y(_04787_));
 NAND2x1_ASAP7_75t_R _23746_ (.A(_14110_),
    .B(_01428_),
    .Y(_04788_));
 OA211x2_ASAP7_75t_R _23747_ (.A1(_13801_),
    .A2(_04787_),
    .B(_04788_),
    .C(_14036_),
    .Y(_04789_));
 OR3x1_ASAP7_75t_R _23748_ (.A(_13447_),
    .B(_04786_),
    .C(_04789_),
    .Y(_04790_));
 INVx1_ASAP7_75t_R _23749_ (.A(_01447_),
    .Y(_04791_));
 NAND2x1_ASAP7_75t_R _23750_ (.A(_14495_),
    .B(_01445_),
    .Y(_04792_));
 OA211x2_ASAP7_75t_R _23751_ (.A1(_13801_),
    .A2(_04791_),
    .B(_04792_),
    .C(_13469_),
    .Y(_04793_));
 INVx1_ASAP7_75t_R _23752_ (.A(_01446_),
    .Y(_04794_));
 NAND2x1_ASAP7_75t_R _23753_ (.A(_14495_),
    .B(_01444_),
    .Y(_04795_));
 OA211x2_ASAP7_75t_R _23754_ (.A1(_13801_),
    .A2(_04794_),
    .B(_04795_),
    .C(_14036_),
    .Y(_04796_));
 OR3x1_ASAP7_75t_R _23755_ (.A(_13517_),
    .B(_04793_),
    .C(_04796_),
    .Y(_04797_));
 AND2x2_ASAP7_75t_R _23756_ (.A(_13483_),
    .B(_13517_),
    .Y(_04798_));
 INVx1_ASAP7_75t_R _23757_ (.A(_01420_),
    .Y(_04799_));
 NOR2x1_ASAP7_75t_R _23758_ (.A(_13801_),
    .B(_01422_),
    .Y(_04800_));
 AO21x1_ASAP7_75t_R _23759_ (.A1(_13472_),
    .A2(_04799_),
    .B(_04800_),
    .Y(_04801_));
 INVx1_ASAP7_75t_R _23760_ (.A(_01423_),
    .Y(_04802_));
 NAND2x1_ASAP7_75t_R _23761_ (.A(net20),
    .B(_01421_),
    .Y(_04803_));
 OA211x2_ASAP7_75t_R _23762_ (.A1(_13463_),
    .A2(_04802_),
    .B(_04803_),
    .C(net11),
    .Y(_04804_));
 AO21x1_ASAP7_75t_R _23763_ (.A1(_13492_),
    .A2(_04801_),
    .B(_04804_),
    .Y(_04805_));
 AO32x1_ASAP7_75t_R _23764_ (.A1(_13453_),
    .A2(_04790_),
    .A3(_04797_),
    .B1(_04798_),
    .B2(_04805_),
    .Y(_04806_));
 OR4x2_ASAP7_75t_R _23765_ (.A(_13512_),
    .B(_14373_),
    .C(_04782_),
    .D(_04806_),
    .Y(_04807_));
 NAND3x2_ASAP7_75t_R _23766_ (.B(_04783_),
    .C(_04807_),
    .Y(_18844_),
    .A(_04749_));
 INVx3_ASAP7_75t_R _23767_ (.A(_18844_),
    .Y(_18846_));
 NAND2x1_ASAP7_75t_R _23768_ (.A(_13671_),
    .B(_01426_),
    .Y(_04808_));
 OA211x2_ASAP7_75t_R _23769_ (.A1(_13980_),
    .A2(_04787_),
    .B(_04808_),
    .C(_13708_),
    .Y(_04809_));
 INVx1_ASAP7_75t_R _23770_ (.A(_01428_),
    .Y(_04810_));
 NAND2x1_ASAP7_75t_R _23771_ (.A(_13671_),
    .B(_01424_),
    .Y(_04811_));
 OA211x2_ASAP7_75t_R _23772_ (.A1(_13980_),
    .A2(_04810_),
    .B(_04811_),
    .C(_13719_),
    .Y(_04812_));
 OA21x2_ASAP7_75t_R _23773_ (.A1(_04809_),
    .A2(_04812_),
    .B(_13714_),
    .Y(_04813_));
 NAND2x1_ASAP7_75t_R _23774_ (.A(_13671_),
    .B(_01427_),
    .Y(_04814_));
 OA211x2_ASAP7_75t_R _23775_ (.A1(_13980_),
    .A2(_04784_),
    .B(_04814_),
    .C(_13708_),
    .Y(_04815_));
 INVx1_ASAP7_75t_R _23776_ (.A(_01429_),
    .Y(_04816_));
 NAND2x1_ASAP7_75t_R _23777_ (.A(_13671_),
    .B(_01425_),
    .Y(_04817_));
 OA211x2_ASAP7_75t_R _23778_ (.A1(_13980_),
    .A2(_04816_),
    .B(_04817_),
    .C(_13719_),
    .Y(_04818_));
 OA21x2_ASAP7_75t_R _23779_ (.A1(_04815_),
    .A2(_04818_),
    .B(_13868_),
    .Y(_04819_));
 OR4x1_ASAP7_75t_R _23780_ (.A(_00410_),
    .B(_13669_),
    .C(_04813_),
    .D(_04819_),
    .Y(_04820_));
 NAND2x1_ASAP7_75t_R _23781_ (.A(_13719_),
    .B(_01444_),
    .Y(_04821_));
 OA211x2_ASAP7_75t_R _23782_ (.A1(_13678_),
    .A2(_04794_),
    .B(_04821_),
    .C(_00413_),
    .Y(_04822_));
 NAND2x1_ASAP7_75t_R _23783_ (.A(_13719_),
    .B(_01445_),
    .Y(_04823_));
 OA211x2_ASAP7_75t_R _23784_ (.A1(_13678_),
    .A2(_04791_),
    .B(_04823_),
    .C(_13684_),
    .Y(_04824_));
 OA21x2_ASAP7_75t_R _23785_ (.A1(_04822_),
    .A2(_04824_),
    .B(_13673_),
    .Y(_04825_));
 INVx1_ASAP7_75t_R _23786_ (.A(_01441_),
    .Y(_04826_));
 NOR2x1_ASAP7_75t_R _23787_ (.A(_13719_),
    .B(_01443_),
    .Y(_04827_));
 AO21x1_ASAP7_75t_R _23788_ (.A1(_13678_),
    .A2(_04826_),
    .B(_04827_),
    .Y(_04828_));
 AND3x1_ASAP7_75t_R _23789_ (.A(_13685_),
    .B(_13672_),
    .C(_04828_),
    .Y(_04829_));
 INVx1_ASAP7_75t_R _23790_ (.A(_01440_),
    .Y(_04830_));
 NOR2x1_ASAP7_75t_R _23791_ (.A(_13719_),
    .B(_01442_),
    .Y(_04831_));
 AO21x1_ASAP7_75t_R _23792_ (.A1(_13678_),
    .A2(_04830_),
    .B(_04831_),
    .Y(_04832_));
 AND3x1_ASAP7_75t_R _23793_ (.A(_13692_),
    .B(_13672_),
    .C(_04832_),
    .Y(_04833_));
 OR5x1_ASAP7_75t_R _23794_ (.A(_00410_),
    .B(_13668_),
    .C(_04825_),
    .D(_04829_),
    .E(_04833_),
    .Y(_04834_));
 INVx1_ASAP7_75t_R _23795_ (.A(_01419_),
    .Y(_04835_));
 NAND2x1_ASAP7_75t_R _23796_ (.A(_13720_),
    .B(_01790_),
    .Y(_04836_));
 OA211x2_ASAP7_75t_R _23797_ (.A1(_13754_),
    .A2(_04835_),
    .B(_04836_),
    .C(_13868_),
    .Y(_04837_));
 AND3x1_ASAP7_75t_R _23798_ (.A(_13672_),
    .B(_00410_),
    .C(_13668_),
    .Y(_04838_));
 OAI21x1_ASAP7_75t_R _23799_ (.A1(_01418_),
    .A2(_13710_),
    .B(_04838_),
    .Y(_04839_));
 NAND2x1_ASAP7_75t_R _23800_ (.A(_13671_),
    .B(_01435_),
    .Y(_04840_));
 OA211x2_ASAP7_75t_R _23801_ (.A1(_13980_),
    .A2(_04776_),
    .B(_04840_),
    .C(_13708_),
    .Y(_04841_));
 INVx1_ASAP7_75t_R _23802_ (.A(_01437_),
    .Y(_04842_));
 NAND2x1_ASAP7_75t_R _23803_ (.A(_13671_),
    .B(_01433_),
    .Y(_04843_));
 OA211x2_ASAP7_75t_R _23804_ (.A1(_13980_),
    .A2(_04842_),
    .B(_04843_),
    .C(_13719_),
    .Y(_04844_));
 OR5x1_ASAP7_75t_R _23805_ (.A(_13714_),
    .B(_13675_),
    .C(_13668_),
    .D(_04841_),
    .E(_04844_),
    .Y(_04845_));
 OA21x2_ASAP7_75t_R _23806_ (.A1(_04837_),
    .A2(_04839_),
    .B(_04845_),
    .Y(_04846_));
 INVx1_ASAP7_75t_R _23807_ (.A(_01422_),
    .Y(_04847_));
 NAND2x1_ASAP7_75t_R _23808_ (.A(_13719_),
    .B(_01420_),
    .Y(_04848_));
 OA211x2_ASAP7_75t_R _23809_ (.A1(_13678_),
    .A2(_04847_),
    .B(_04848_),
    .C(_00413_),
    .Y(_04849_));
 NAND2x1_ASAP7_75t_R _23810_ (.A(_13719_),
    .B(_01421_),
    .Y(_04850_));
 OA211x2_ASAP7_75t_R _23811_ (.A1(_13678_),
    .A2(_04802_),
    .B(_04850_),
    .C(_13685_),
    .Y(_04851_));
 OR4x1_ASAP7_75t_R _23812_ (.A(_13672_),
    .B(_13669_),
    .C(_04849_),
    .D(_04851_),
    .Y(_04852_));
 INVx1_ASAP7_75t_R _23813_ (.A(_01436_),
    .Y(_04853_));
 NAND2x1_ASAP7_75t_R _23814_ (.A(_13980_),
    .B(_01432_),
    .Y(_04854_));
 OA211x2_ASAP7_75t_R _23815_ (.A1(_13980_),
    .A2(_04853_),
    .B(_04854_),
    .C(_13678_),
    .Y(_04855_));
 NAND2x1_ASAP7_75t_R _23816_ (.A(_13671_),
    .B(_01434_),
    .Y(_04856_));
 OA211x2_ASAP7_75t_R _23817_ (.A1(_13980_),
    .A2(_04779_),
    .B(_04856_),
    .C(_13708_),
    .Y(_04857_));
 OR4x1_ASAP7_75t_R _23818_ (.A(_13868_),
    .B(_13668_),
    .C(_04855_),
    .D(_04857_),
    .Y(_04858_));
 AO21x1_ASAP7_75t_R _23819_ (.A1(_04852_),
    .A2(_04858_),
    .B(_13675_),
    .Y(_04859_));
 AND4x2_ASAP7_75t_R _23820_ (.A(_04820_),
    .B(_04834_),
    .C(_04846_),
    .D(_04859_),
    .Y(_04860_));
 BUFx6f_ASAP7_75t_R _23821_ (.A(_04860_),
    .Y(_04861_));
 NAND3x2_ASAP7_75t_R _23822_ (.B(_13667_),
    .C(_04861_),
    .Y(_04862_),
    .A(_13659_));
 INVx1_ASAP7_75t_R _23823_ (.A(_01519_),
    .Y(_04863_));
 INVx2_ASAP7_75t_R _23824_ (.A(_00066_),
    .Y(_04864_));
 AND3x1_ASAP7_75t_R _23825_ (.A(_04864_),
    .B(_13664_),
    .C(_13665_),
    .Y(_04865_));
 AOI22x1_ASAP7_75t_R _23826_ (.A1(_04863_),
    .A2(_13414_),
    .B1(_13770_),
    .B2(_04865_),
    .Y(_04866_));
 AND2x6_ASAP7_75t_R _23827_ (.A(_04862_),
    .B(_04866_),
    .Y(_18845_));
 BUFx6f_ASAP7_75t_R _23828_ (.A(_14925_),
    .Y(_04867_));
 BUFx4f_ASAP7_75t_R _23829_ (.A(_01448_),
    .Y(_04868_));
 INVx3_ASAP7_75t_R _23830_ (.A(_04868_),
    .Y(_04869_));
 NAND2x2_ASAP7_75t_R _23831_ (.A(_01816_),
    .B(_02217_),
    .Y(_04870_));
 INVx3_ASAP7_75t_R _23832_ (.A(_00408_),
    .Y(_04871_));
 AOI22x1_ASAP7_75t_R _23833_ (.A1(_04871_),
    .A2(_04868_),
    .B1(_01751_),
    .B2(_04870_),
    .Y(_04872_));
 OAI21x1_ASAP7_75t_R _23834_ (.A1(_00407_),
    .A2(_04861_),
    .B(_04872_),
    .Y(_04873_));
 AND3x1_ASAP7_75t_R _23835_ (.A(_04869_),
    .B(_04870_),
    .C(_04873_),
    .Y(_04874_));
 OR3x4_ASAP7_75t_R _23836_ (.A(_13451_),
    .B(_04760_),
    .C(_04775_),
    .Y(_04875_));
 OR3x4_ASAP7_75t_R _23837_ (.A(_13512_),
    .B(_04782_),
    .C(_04806_),
    .Y(_04876_));
 INVx1_ASAP7_75t_R _23838_ (.A(_00407_),
    .Y(_04877_));
 OR3x1_ASAP7_75t_R _23839_ (.A(_04871_),
    .B(_04877_),
    .C(_04870_),
    .Y(_04878_));
 BUFx4f_ASAP7_75t_R _23840_ (.A(_04878_),
    .Y(_04879_));
 AOI21x1_ASAP7_75t_R _23841_ (.A1(_04875_),
    .A2(_04876_),
    .B(_04879_),
    .Y(_04880_));
 AOI211x1_ASAP7_75t_R _23842_ (.A1(_04869_),
    .A2(_04870_),
    .B(_04873_),
    .C(_04880_),
    .Y(_04881_));
 OR3x1_ASAP7_75t_R _23843_ (.A(_04867_),
    .B(_04874_),
    .C(_04881_),
    .Y(_04882_));
 AND3x2_ASAP7_75t_R _23844_ (.A(_13659_),
    .B(_13666_),
    .C(_04861_),
    .Y(_04883_));
 AO32x2_ASAP7_75t_R _23845_ (.A1(_04864_),
    .A2(_13770_),
    .A3(_13666_),
    .B1(_04863_),
    .B2(_13414_),
    .Y(_04884_));
 OR3x2_ASAP7_75t_R _23846_ (.A(_18844_),
    .B(_04883_),
    .C(_04884_),
    .Y(_04885_));
 AO21x1_ASAP7_75t_R _23847_ (.A1(_04862_),
    .A2(_04866_),
    .B(_18846_),
    .Y(_04886_));
 AO21x2_ASAP7_75t_R _23848_ (.A1(_04885_),
    .A2(_04886_),
    .B(_17344_),
    .Y(_04887_));
 AND3x1_ASAP7_75t_R _23849_ (.A(_18846_),
    .B(_04862_),
    .C(_04866_),
    .Y(_04888_));
 OA21x2_ASAP7_75t_R _23850_ (.A1(_04883_),
    .A2(_04884_),
    .B(_18844_),
    .Y(_04889_));
 OR4x2_ASAP7_75t_R _23851_ (.A(_14922_),
    .B(_16286_),
    .C(_04888_),
    .D(_04889_),
    .Y(_04890_));
 OA21x2_ASAP7_75t_R _23852_ (.A1(_01318_),
    .A2(_01317_),
    .B(_01351_),
    .Y(_04891_));
 OA21x2_ASAP7_75t_R _23853_ (.A1(_01350_),
    .A2(_04891_),
    .B(_01384_),
    .Y(_04892_));
 OA21x2_ASAP7_75t_R _23854_ (.A1(_01383_),
    .A2(_04892_),
    .B(_01417_),
    .Y(_04893_));
 OR4x1_ASAP7_75t_R _23855_ (.A(_01284_),
    .B(_01317_),
    .C(_01350_),
    .D(_01383_),
    .Y(_04894_));
 AND2x2_ASAP7_75t_R _23856_ (.A(_01449_),
    .B(_04894_),
    .Y(_04895_));
 AND4x1_ASAP7_75t_R _23857_ (.A(_01449_),
    .B(_04395_),
    .C(_04398_),
    .D(_04893_),
    .Y(_04896_));
 AOI221x1_ASAP7_75t_R _23858_ (.A1(_01416_),
    .A2(_01449_),
    .B1(_04893_),
    .B2(_04895_),
    .C(_04896_),
    .Y(_04897_));
 AO31x2_ASAP7_75t_R _23859_ (.A1(_04882_),
    .A2(_04887_),
    .A3(_04890_),
    .B(_04897_),
    .Y(_04898_));
 AO221x2_ASAP7_75t_R _23860_ (.A1(_01416_),
    .A2(_01449_),
    .B1(_04893_),
    .B2(_04895_),
    .C(_04896_),
    .Y(_04899_));
 AOI21x1_ASAP7_75t_R _23861_ (.A1(_04885_),
    .A2(_04886_),
    .B(_17344_),
    .Y(_04900_));
 OA21x2_ASAP7_75t_R _23862_ (.A1(net1973),
    .A2(_15262_),
    .B(_16285_),
    .Y(_04901_));
 AND4x2_ASAP7_75t_R _23863_ (.A(_04901_),
    .B(_04867_),
    .C(_04885_),
    .D(_04886_),
    .Y(_04902_));
 AO21x2_ASAP7_75t_R _23864_ (.A1(_01816_),
    .A2(_02217_),
    .B(_04868_),
    .Y(_04903_));
 AND2x2_ASAP7_75t_R _23865_ (.A(_16286_),
    .B(_04903_),
    .Y(_04904_));
 OAI21x1_ASAP7_75t_R _23866_ (.A1(_04873_),
    .A2(_04880_),
    .B(_04904_),
    .Y(_04905_));
 OR4x2_ASAP7_75t_R _23867_ (.A(_14925_),
    .B(_04873_),
    .C(_04880_),
    .D(_04903_),
    .Y(_04906_));
 NAND2x1_ASAP7_75t_R _23868_ (.A(_04905_),
    .B(_04906_),
    .Y(_04907_));
 OR4x2_ASAP7_75t_R _23869_ (.A(_04899_),
    .B(_04900_),
    .C(_04902_),
    .D(_04907_),
    .Y(_04908_));
 NAND2x2_ASAP7_75t_R _23870_ (.A(_04898_),
    .B(_04908_),
    .Y(\alu_adder_result_ex[31] ));
 OR3x1_ASAP7_75t_R _23871_ (.A(_15485_),
    .B(_04402_),
    .C(_17007_),
    .Y(_04909_));
 OR2x2_ASAP7_75t_R _23872_ (.A(_04410_),
    .B(_04894_),
    .Y(_04910_));
 OA21x2_ASAP7_75t_R _23873_ (.A1(_01284_),
    .A2(_04405_),
    .B(_01318_),
    .Y(_04911_));
 OA21x2_ASAP7_75t_R _23874_ (.A1(_01317_),
    .A2(_04911_),
    .B(_01351_),
    .Y(_04912_));
 OA21x2_ASAP7_75t_R _23875_ (.A1(_01350_),
    .A2(_04912_),
    .B(_01384_),
    .Y(_04913_));
 OA21x2_ASAP7_75t_R _23876_ (.A1(_01383_),
    .A2(_04913_),
    .B(_01417_),
    .Y(_04914_));
 OR2x2_ASAP7_75t_R _23877_ (.A(_17009_),
    .B(_04910_),
    .Y(_04915_));
 OA211x2_ASAP7_75t_R _23878_ (.A1(_04909_),
    .A2(_04910_),
    .B(_04914_),
    .C(_04915_),
    .Y(_04916_));
 XNOR2x2_ASAP7_75t_R _23879_ (.A(_01416_),
    .B(_04916_),
    .Y(_04917_));
 INVx4_ASAP7_75t_R _23880_ (.A(_04917_),
    .Y(\alu_adder_result_ex[30] ));
 INVx1_ASAP7_75t_R _23881_ (.A(_18845_),
    .Y(_18847_));
 BUFx4f_ASAP7_75t_R _23882_ (.A(_01454_),
    .Y(_04918_));
 BUFx4f_ASAP7_75t_R _23883_ (.A(_04918_),
    .Y(_04919_));
 INVx2_ASAP7_75t_R _23884_ (.A(net47),
    .Y(_04920_));
 NAND2x2_ASAP7_75t_R _23885_ (.A(_04920_),
    .B(_01508_),
    .Y(_04921_));
 AND3x2_ASAP7_75t_R _23886_ (.A(_00399_),
    .B(_13359_),
    .C(_13357_),
    .Y(_04922_));
 AND2x4_ASAP7_75t_R _23887_ (.A(net104),
    .B(_04922_),
    .Y(_04923_));
 AND3x1_ASAP7_75t_R _23888_ (.A(_04919_),
    .B(_04921_),
    .C(_04923_),
    .Y(\id_stage_i.controller_i.load_err_d ));
 INVx1_ASAP7_75t_R _23889_ (.A(_01454_),
    .Y(_04924_));
 AND3x1_ASAP7_75t_R _23890_ (.A(_04924_),
    .B(_04921_),
    .C(_04923_),
    .Y(\id_stage_i.controller_i.store_err_d ));
 AND3x4_ASAP7_75t_R _23891_ (.A(_14022_),
    .B(_14034_),
    .C(_14068_),
    .Y(_04925_));
 OR3x4_ASAP7_75t_R _23892_ (.A(_13631_),
    .B(_13632_),
    .C(_13774_),
    .Y(_04926_));
 AND2x2_ASAP7_75t_R _23893_ (.A(_04925_),
    .B(_04926_),
    .Y(_04927_));
 BUFx6f_ASAP7_75t_R _23894_ (.A(_04927_),
    .Y(_04928_));
 BUFx6f_ASAP7_75t_R _23895_ (.A(_14668_),
    .Y(_18658_));
 AND2x2_ASAP7_75t_R _23896_ (.A(_18658_),
    .B(_18663_),
    .Y(_04929_));
 BUFx4f_ASAP7_75t_R _23897_ (.A(_01555_),
    .Y(_04930_));
 BUFx4f_ASAP7_75t_R _23898_ (.A(_01782_),
    .Y(_04931_));
 BUFx4f_ASAP7_75t_R _23899_ (.A(_01779_),
    .Y(_04932_));
 INVx3_ASAP7_75t_R _23900_ (.A(_04932_),
    .Y(_04933_));
 BUFx3_ASAP7_75t_R _23901_ (.A(_01780_),
    .Y(_04934_));
 BUFx4f_ASAP7_75t_R _23902_ (.A(_01781_),
    .Y(_04935_));
 INVx3_ASAP7_75t_R _23903_ (.A(_04935_),
    .Y(_04936_));
 OR3x4_ASAP7_75t_R _23904_ (.A(_04933_),
    .B(_04934_),
    .C(_04936_),
    .Y(_04937_));
 NOR2x2_ASAP7_75t_R _23905_ (.A(_04931_),
    .B(_04937_),
    .Y(_04938_));
 AND3x1_ASAP7_75t_R _23906_ (.A(_13407_),
    .B(_04930_),
    .C(_04938_),
    .Y(_04939_));
 BUFx6f_ASAP7_75t_R _23907_ (.A(_04939_),
    .Y(_04940_));
 AND3x1_ASAP7_75t_R _23908_ (.A(_02310_),
    .B(_04929_),
    .C(_04940_),
    .Y(_04941_));
 INVx1_ASAP7_75t_R _23909_ (.A(_02302_),
    .Y(_04942_));
 OA21x2_ASAP7_75t_R _23910_ (.A1(_04942_),
    .A2(_02301_),
    .B(_02300_),
    .Y(_04943_));
 NOR2x1_ASAP7_75t_R _23911_ (.A(_01452_),
    .B(_02301_),
    .Y(_04944_));
 BUFx6f_ASAP7_75t_R _23912_ (.A(_01455_),
    .Y(_04945_));
 BUFx4f_ASAP7_75t_R _23913_ (.A(_00571_),
    .Y(_04946_));
 NAND2x2_ASAP7_75t_R _23914_ (.A(_00479_),
    .B(_04946_),
    .Y(_04947_));
 BUFx4f_ASAP7_75t_R _23915_ (.A(_00572_),
    .Y(_04948_));
 NAND2x2_ASAP7_75t_R _23916_ (.A(_04948_),
    .B(_14299_),
    .Y(_04949_));
 OR2x4_ASAP7_75t_R _23917_ (.A(_04947_),
    .B(_04949_),
    .Y(_04950_));
 NAND2x1_ASAP7_75t_R _23918_ (.A(_04945_),
    .B(_04950_),
    .Y(_04951_));
 NAND2x2_ASAP7_75t_R _23919_ (.A(_14298_),
    .B(_14668_),
    .Y(_04952_));
 OR3x4_ASAP7_75t_R _23920_ (.A(_14059_),
    .B(_13579_),
    .C(_14314_),
    .Y(_04953_));
 AND4x1_ASAP7_75t_R _23921_ (.A(_13511_),
    .B(_13447_),
    .C(_14384_),
    .D(_14440_),
    .Y(_04954_));
 AND4x1_ASAP7_75t_R _23922_ (.A(_13511_),
    .B(_13518_),
    .C(_14377_),
    .D(_14433_),
    .Y(_04955_));
 AND2x2_ASAP7_75t_R _23923_ (.A(_13450_),
    .B(_13518_),
    .Y(_04956_));
 OA211x2_ASAP7_75t_R _23924_ (.A1(_14449_),
    .A2(_14452_),
    .B(_14391_),
    .C(_14393_),
    .Y(_04957_));
 OA211x2_ASAP7_75t_R _23925_ (.A1(_14443_),
    .A2(_14446_),
    .B(_14387_),
    .C(_14389_),
    .Y(_04958_));
 NOR2x1_ASAP7_75t_R _23926_ (.A(_13511_),
    .B(_13518_),
    .Y(_04959_));
 AO22x1_ASAP7_75t_R _23927_ (.A1(_04956_),
    .A2(_04957_),
    .B1(_04958_),
    .B2(_04959_),
    .Y(_04960_));
 OA31x2_ASAP7_75t_R _23928_ (.A1(_04954_),
    .A2(_04955_),
    .A3(_04960_),
    .B1(_13484_),
    .Y(_04961_));
 AND5x2_ASAP7_75t_R _23929_ (.A(_13518_),
    .B(_14417_),
    .C(_14424_),
    .D(_14461_),
    .E(_14468_),
    .Y(_04962_));
 AOI221x1_ASAP7_75t_R _23930_ (.A1(_14402_),
    .A2(_14409_),
    .B1(_14477_),
    .B2(_14484_),
    .C(_13518_),
    .Y(_04963_));
 OA21x2_ASAP7_75t_R _23931_ (.A1(_04962_),
    .A2(_04963_),
    .B(_13454_),
    .Y(_04964_));
 OAI21x1_ASAP7_75t_R _23932_ (.A1(_04961_),
    .A2(_04964_),
    .B(_13788_),
    .Y(_04965_));
 NAND2x2_ASAP7_75t_R _23933_ (.A(_13775_),
    .B(_04925_),
    .Y(_04966_));
 AO211x2_ASAP7_75t_R _23934_ (.A1(_04953_),
    .A2(_04965_),
    .B(_04966_),
    .C(_18634_),
    .Y(_04967_));
 OA21x2_ASAP7_75t_R _23935_ (.A1(_14545_),
    .A2(_14547_),
    .B(_14069_),
    .Y(_04968_));
 INVx2_ASAP7_75t_R _23936_ (.A(_04968_),
    .Y(_18851_));
 OR3x4_ASAP7_75t_R _23937_ (.A(_18654_),
    .B(_14729_),
    .C(_18851_),
    .Y(_04969_));
 OR5x1_ASAP7_75t_R _23938_ (.A(_14306_),
    .B(_04951_),
    .C(_04952_),
    .D(_04967_),
    .E(_04969_),
    .Y(_04970_));
 OA21x2_ASAP7_75t_R _23939_ (.A1(_04943_),
    .A2(_04944_),
    .B(_04970_),
    .Y(_04971_));
 NAND2x2_ASAP7_75t_R _23940_ (.A(_18627_),
    .B(_18634_),
    .Y(_04972_));
 NAND2x1_ASAP7_75t_R _23941_ (.A(_13365_),
    .B(_13551_),
    .Y(_04973_));
 OR4x2_ASAP7_75t_R _23942_ (.A(_14151_),
    .B(_14152_),
    .C(_14154_),
    .D(_04973_),
    .Y(_04974_));
 BUFx6f_ASAP7_75t_R _23943_ (.A(_04974_),
    .Y(_04975_));
 INVx3_ASAP7_75t_R _23944_ (.A(_14299_),
    .Y(_04976_));
 AND2x4_ASAP7_75t_R _23945_ (.A(_04976_),
    .B(_14069_),
    .Y(_04977_));
 NAND3x2_ASAP7_75t_R _23946_ (.B(_04975_),
    .C(_04977_),
    .Y(_04978_),
    .A(_14229_));
 OR3x2_ASAP7_75t_R _23947_ (.A(_18643_),
    .B(_04972_),
    .C(_04978_),
    .Y(_04979_));
 OAI21x1_ASAP7_75t_R _23948_ (.A1(_14151_),
    .A2(_14152_),
    .B(_13551_),
    .Y(_04980_));
 AOI21x1_ASAP7_75t_R _23949_ (.A1(_13387_),
    .A2(_14148_),
    .B(_14154_),
    .Y(_04981_));
 AND4x2_ASAP7_75t_R _23950_ (.A(_13367_),
    .B(_04980_),
    .C(_04981_),
    .D(_14229_),
    .Y(_04982_));
 NOR2x2_ASAP7_75t_R _23951_ (.A(_04947_),
    .B(_04949_),
    .Y(_04983_));
 BUFx3_ASAP7_75t_R _23952_ (.A(_04967_),
    .Y(_04984_));
 OR5x2_ASAP7_75t_R _23953_ (.A(_04966_),
    .B(_18627_),
    .C(_04982_),
    .D(_04983_),
    .E(_04984_),
    .Y(_04985_));
 OR4x2_ASAP7_75t_R _23954_ (.A(_18654_),
    .B(_14668_),
    .C(_14729_),
    .D(_18851_),
    .Y(_04986_));
 BUFx4f_ASAP7_75t_R _23955_ (.A(_04986_),
    .Y(_04987_));
 AOI21x1_ASAP7_75t_R _23956_ (.A1(_04979_),
    .A2(_04985_),
    .B(_04987_),
    .Y(_04988_));
 AND2x2_ASAP7_75t_R _23957_ (.A(_14069_),
    .B(_18632_),
    .Y(_04989_));
 AO33x2_ASAP7_75t_R _23958_ (.A1(_14395_),
    .A2(_14410_),
    .A3(_14425_),
    .B1(_14454_),
    .B2(_14469_),
    .B3(_14485_),
    .Y(_04990_));
 NAND2x1_ASAP7_75t_R _23959_ (.A(_13589_),
    .B(_13579_),
    .Y(_04991_));
 AO32x2_ASAP7_75t_R _23960_ (.A1(_13366_),
    .A2(_13387_),
    .A3(_04990_),
    .B1(_04991_),
    .B2(_14429_),
    .Y(_04992_));
 OR5x2_ASAP7_75t_R _23961_ (.A(_18654_),
    .B(_14668_),
    .C(_14729_),
    .D(_18851_),
    .E(_04992_),
    .Y(_04993_));
 INVx1_ASAP7_75t_R _23962_ (.A(_04993_),
    .Y(_04994_));
 INVx1_ASAP7_75t_R _23963_ (.A(_04948_),
    .Y(_04995_));
 AO21x2_ASAP7_75t_R _23964_ (.A1(_14149_),
    .A2(_14155_),
    .B(_14305_),
    .Y(_04996_));
 OR3x1_ASAP7_75t_R _23965_ (.A(_04995_),
    .B(_14298_),
    .C(_04996_),
    .Y(_04997_));
 AND4x1_ASAP7_75t_R _23966_ (.A(_04950_),
    .B(_04989_),
    .C(_04994_),
    .D(_04997_),
    .Y(_04998_));
 NAND2x2_ASAP7_75t_R _23967_ (.A(_14070_),
    .B(_04996_),
    .Y(_04999_));
 OR5x2_ASAP7_75t_R _23968_ (.A(_04966_),
    .B(_14298_),
    .C(_18632_),
    .D(_18640_),
    .E(_18643_),
    .Y(_05000_));
 NOR2x2_ASAP7_75t_R _23969_ (.A(_04986_),
    .B(_05000_),
    .Y(_05001_));
 NAND2x2_ASAP7_75t_R _23970_ (.A(_04953_),
    .B(_04965_),
    .Y(_05002_));
 NAND2x1_ASAP7_75t_R _23971_ (.A(_14297_),
    .B(_18658_),
    .Y(_05003_));
 AND4x1_ASAP7_75t_R _23972_ (.A(_04950_),
    .B(_05002_),
    .C(_04989_),
    .D(_05003_),
    .Y(_05004_));
 OR3x4_ASAP7_75t_R _23973_ (.A(_18654_),
    .B(_14729_),
    .C(_18851_),
    .Y(_05005_));
 NOR2x1_ASAP7_75t_R _23974_ (.A(_14306_),
    .B(_05005_),
    .Y(_05006_));
 AO32x1_ASAP7_75t_R _23975_ (.A1(_04999_),
    .A2(_04950_),
    .A3(_05001_),
    .B1(_05004_),
    .B2(_05006_),
    .Y(_05007_));
 OR3x1_ASAP7_75t_R _23976_ (.A(_14298_),
    .B(_18632_),
    .C(_04992_),
    .Y(_05008_));
 BUFx4f_ASAP7_75t_R _23977_ (.A(_05008_),
    .Y(_05009_));
 NOR2x1_ASAP7_75t_R _23978_ (.A(_04986_),
    .B(_05009_),
    .Y(_05010_));
 INVx1_ASAP7_75t_R _23979_ (.A(_04946_),
    .Y(_05011_));
 AND2x2_ASAP7_75t_R _23980_ (.A(_05011_),
    .B(_14069_),
    .Y(_05012_));
 NAND3x2_ASAP7_75t_R _23981_ (.B(_04975_),
    .C(_05012_),
    .Y(_05013_),
    .A(_18625_));
 OAI21x1_ASAP7_75t_R _23982_ (.A1(_14299_),
    .A2(_14306_),
    .B(_05013_),
    .Y(_05014_));
 OA21x2_ASAP7_75t_R _23983_ (.A1(_05011_),
    .A2(_04976_),
    .B(_14668_),
    .Y(_05015_));
 OA211x2_ASAP7_75t_R _23984_ (.A1(_14427_),
    .A2(_14428_),
    .B(_14059_),
    .C(_14487_),
    .Y(_05016_));
 AND3x1_ASAP7_75t_R _23985_ (.A(_13788_),
    .B(_14426_),
    .C(_14486_),
    .Y(_05017_));
 AO21x2_ASAP7_75t_R _23986_ (.A1(_14373_),
    .A2(_05016_),
    .B(_05017_),
    .Y(_05018_));
 AND5x1_ASAP7_75t_R _23987_ (.A(_18652_),
    .B(_18665_),
    .C(_04968_),
    .D(_05015_),
    .E(_05018_),
    .Y(_05019_));
 NOR2x1_ASAP7_75t_R _23988_ (.A(_04996_),
    .B(_04972_),
    .Y(_05020_));
 INVx1_ASAP7_75t_R _23989_ (.A(_04992_),
    .Y(_05021_));
 OA221x2_ASAP7_75t_R _23990_ (.A1(_13601_),
    .A2(_14314_),
    .B1(_14371_),
    .B2(_14373_),
    .C(_14069_),
    .Y(_05022_));
 AO32x2_ASAP7_75t_R _23991_ (.A1(_14604_),
    .A2(_14546_),
    .A3(_14429_),
    .B1(_14545_),
    .B2(_14603_),
    .Y(_05023_));
 AND5x1_ASAP7_75t_R _23992_ (.A(_14229_),
    .B(_14729_),
    .C(_04974_),
    .D(_04977_),
    .E(_05023_),
    .Y(_05024_));
 AND5x2_ASAP7_75t_R _23993_ (.A(_14298_),
    .B(_18658_),
    .C(_05021_),
    .D(_05022_),
    .E(_05024_),
    .Y(_05025_));
 AO221x1_ASAP7_75t_R _23994_ (.A1(_05010_),
    .A2(_05014_),
    .B1(_05019_),
    .B2(_05020_),
    .C(_05025_),
    .Y(_05026_));
 OR4x1_ASAP7_75t_R _23995_ (.A(_04988_),
    .B(_04998_),
    .C(_05007_),
    .D(_05026_),
    .Y(_05027_));
 AND2x2_ASAP7_75t_R _23996_ (.A(_18652_),
    .B(_04968_),
    .Y(_05028_));
 AND2x2_ASAP7_75t_R _23997_ (.A(_04953_),
    .B(_04965_),
    .Y(_05029_));
 AND2x2_ASAP7_75t_R _23998_ (.A(_14070_),
    .B(_04992_),
    .Y(_05030_));
 NAND2x2_ASAP7_75t_R _23999_ (.A(_05029_),
    .B(_05030_),
    .Y(_05031_));
 AND3x1_ASAP7_75t_R _24000_ (.A(_05028_),
    .B(_04971_),
    .C(_05031_),
    .Y(_05032_));
 AND4x1_ASAP7_75t_R _24001_ (.A(_14069_),
    .B(_14298_),
    .C(_18634_),
    .D(_04947_),
    .Y(_05033_));
 BUFx4f_ASAP7_75t_R _24002_ (.A(_00479_),
    .Y(_05034_));
 INVx1_ASAP7_75t_R _24003_ (.A(_05034_),
    .Y(_05035_));
 OR2x2_ASAP7_75t_R _24004_ (.A(_05035_),
    .B(_04949_),
    .Y(_05036_));
 AO32x1_ASAP7_75t_R _24005_ (.A1(_18619_),
    .A2(_18625_),
    .A3(_05033_),
    .B1(_05036_),
    .B2(_04966_),
    .Y(_05037_));
 AND4x1_ASAP7_75t_R _24006_ (.A(_18627_),
    .B(_04982_),
    .C(_18634_),
    .D(_05036_),
    .Y(_05038_));
 AND2x2_ASAP7_75t_R _24007_ (.A(_18660_),
    .B(_18663_),
    .Y(_05039_));
 OAI21x1_ASAP7_75t_R _24008_ (.A1(_05037_),
    .A2(_05038_),
    .B(_05039_),
    .Y(_05040_));
 NAND2x1_ASAP7_75t_R _24009_ (.A(_14230_),
    .B(_18627_),
    .Y(_05041_));
 OAI22x1_ASAP7_75t_R _24010_ (.A1(_18627_),
    .A2(_04975_),
    .B1(_05041_),
    .B2(_18617_),
    .Y(_05042_));
 AND3x1_ASAP7_75t_R _24011_ (.A(_04949_),
    .B(_05022_),
    .C(_05039_),
    .Y(_05043_));
 OR2x2_ASAP7_75t_R _24012_ (.A(_14373_),
    .B(_14148_),
    .Y(_05044_));
 OA211x2_ASAP7_75t_R _24013_ (.A1(_14230_),
    .A2(_05044_),
    .B(_04975_),
    .C(_04995_),
    .Y(_05045_));
 AND4x1_ASAP7_75t_R _24014_ (.A(_05034_),
    .B(_04946_),
    .C(_15334_),
    .D(_13551_),
    .Y(_05046_));
 INVx1_ASAP7_75t_R _24015_ (.A(_05046_),
    .Y(_05047_));
 OR3x1_ASAP7_75t_R _24016_ (.A(_14151_),
    .B(_14152_),
    .C(_14154_),
    .Y(_05048_));
 OA222x2_ASAP7_75t_R _24017_ (.A1(_04976_),
    .A2(_04947_),
    .B1(_04975_),
    .B2(_14230_),
    .C1(_05047_),
    .C2(_05048_),
    .Y(_05049_));
 OA211x2_ASAP7_75t_R _24018_ (.A1(_05045_),
    .A2(_05049_),
    .B(_05022_),
    .C(_05039_),
    .Y(_05050_));
 AOI21x1_ASAP7_75t_R _24019_ (.A1(_05042_),
    .A2(_05043_),
    .B(_05050_),
    .Y(_05051_));
 NAND2x1_ASAP7_75t_R _24020_ (.A(_05040_),
    .B(_05051_),
    .Y(_05052_));
 OA21x2_ASAP7_75t_R _24021_ (.A1(_04996_),
    .A2(_04972_),
    .B(_14070_),
    .Y(_05053_));
 NAND2x1_ASAP7_75t_R _24022_ (.A(_18627_),
    .B(_04982_),
    .Y(_05054_));
 NAND2x1_ASAP7_75t_R _24023_ (.A(_18632_),
    .B(_04977_),
    .Y(_05055_));
 OAI22x1_ASAP7_75t_R _24024_ (.A1(_04946_),
    .A2(_05053_),
    .B1(_05054_),
    .B2(_05055_),
    .Y(_05056_));
 AND3x1_ASAP7_75t_R _24025_ (.A(_04971_),
    .B(_04994_),
    .C(_05056_),
    .Y(_05057_));
 AOI221x1_ASAP7_75t_R _24026_ (.A1(_04971_),
    .A2(_05027_),
    .B1(_05032_),
    .B2(_05052_),
    .C(_05057_),
    .Y(_05058_));
 BUFx6f_ASAP7_75t_R _24027_ (.A(_05058_),
    .Y(_05059_));
 OAI21x1_ASAP7_75t_R _24028_ (.A1(_04941_),
    .A2(_05059_),
    .B(_14071_),
    .Y(_05060_));
 BUFx6f_ASAP7_75t_R _24029_ (.A(net2018),
    .Y(_05061_));
 BUFx4f_ASAP7_75t_R _24030_ (.A(_05061_),
    .Y(_05062_));
 AO21x1_ASAP7_75t_R _24031_ (.A1(_04928_),
    .A2(_05060_),
    .B(_05062_),
    .Y(_05063_));
 OR5x1_ASAP7_75t_R _24032_ (.A(_05061_),
    .B(_13403_),
    .C(_13623_),
    .D(_13648_),
    .E(_13650_),
    .Y(_05064_));
 BUFx3_ASAP7_75t_R _24033_ (.A(_05064_),
    .Y(_05065_));
 OR3x4_ASAP7_75t_R _24034_ (.A(_14057_),
    .B(_14062_),
    .C(_05065_),
    .Y(_05066_));
 INVx1_ASAP7_75t_R _24035_ (.A(_05066_),
    .Y(_05067_));
 BUFx4f_ASAP7_75t_R _24036_ (.A(_18850_),
    .Y(_05068_));
 NOR2x1_ASAP7_75t_R _24037_ (.A(_14065_),
    .B(_05065_),
    .Y(_05069_));
 INVx1_ASAP7_75t_R _24038_ (.A(_01855_),
    .Y(_05070_));
 AND4x2_ASAP7_75t_R _24039_ (.A(_13577_),
    .B(_14546_),
    .C(_14292_),
    .D(_14138_),
    .Y(_05071_));
 AO21x1_ASAP7_75t_R _24040_ (.A1(_05070_),
    .A2(_05071_),
    .B(_14039_),
    .Y(_05072_));
 OA211x2_ASAP7_75t_R _24041_ (.A1(_05068_),
    .A2(_14812_),
    .B(_05069_),
    .C(_05072_),
    .Y(_05073_));
 AOI21x1_ASAP7_75t_R _24042_ (.A1(_04945_),
    .A2(_05067_),
    .B(_05073_),
    .Y(_05074_));
 INVx2_ASAP7_75t_R _24043_ (.A(_01780_),
    .Y(_05075_));
 AND4x1_ASAP7_75t_R _24044_ (.A(_04932_),
    .B(_05075_),
    .C(_04936_),
    .D(_04931_),
    .Y(_05076_));
 BUFx4f_ASAP7_75t_R _24045_ (.A(_05076_),
    .Y(_05077_));
 AOI21x1_ASAP7_75t_R _24046_ (.A1(_05063_),
    .A2(_05074_),
    .B(_05077_),
    .Y(\id_stage_i.controller_i.illegal_insn_d ));
 BUFx4f_ASAP7_75t_R _24047_ (.A(_13776_),
    .Y(_05078_));
 INVx2_ASAP7_75t_R _24048_ (.A(_04930_),
    .Y(_05079_));
 AND2x2_ASAP7_75t_R _24049_ (.A(_13605_),
    .B(_14064_),
    .Y(_05080_));
 AND5x2_ASAP7_75t_R _24050_ (.A(net12),
    .B(_13511_),
    .C(_13482_),
    .D(_13577_),
    .E(_13578_),
    .Y(_05081_));
 AND2x2_ASAP7_75t_R _24051_ (.A(_13603_),
    .B(_05081_),
    .Y(_05082_));
 AND3x1_ASAP7_75t_R _24052_ (.A(_13774_),
    .B(_05080_),
    .C(_05082_),
    .Y(_05083_));
 NOR2x1_ASAP7_75t_R _24053_ (.A(_05079_),
    .B(_05083_),
    .Y(_05084_));
 AND3x4_ASAP7_75t_R _24054_ (.A(_02310_),
    .B(_14070_),
    .C(_04940_),
    .Y(_05085_));
 NAND2x1_ASAP7_75t_R _24055_ (.A(_04929_),
    .B(_05085_),
    .Y(_05086_));
 OA211x2_ASAP7_75t_R _24056_ (.A1(_05061_),
    .A2(_05084_),
    .B(_05086_),
    .C(_05074_),
    .Y(_05087_));
 NAND2x1_ASAP7_75t_R _24057_ (.A(_04928_),
    .B(_05087_),
    .Y(_05088_));
 AO21x1_ASAP7_75t_R _24058_ (.A1(_05078_),
    .A2(_05059_),
    .B(_05088_),
    .Y(_05089_));
 NOR2x1_ASAP7_75t_R _24059_ (.A(_05061_),
    .B(_05077_),
    .Y(_05090_));
 AND2x2_ASAP7_75t_R _24060_ (.A(_05089_),
    .B(_05090_),
    .Y(\id_stage_i.controller_i.exc_req_d ));
 INVx5_ASAP7_75t_R _24061_ (.A(_01816_),
    .Y(_05091_));
 BUFx3_ASAP7_75t_R _24062_ (.A(_05091_),
    .Y(_05092_));
 BUFx4f_ASAP7_75t_R _24063_ (.A(_01458_),
    .Y(_05093_));
 BUFx4f_ASAP7_75t_R _24064_ (.A(_00070_),
    .Y(_05094_));
 INVx2_ASAP7_75t_R _24065_ (.A(_05094_),
    .Y(_05095_));
 NOR2x2_ASAP7_75t_R _24066_ (.A(_13593_),
    .B(_04867_),
    .Y(_05096_));
 AND3x4_ASAP7_75t_R _24067_ (.A(_04925_),
    .B(_04926_),
    .C(_04940_),
    .Y(_05097_));
 NAND2x2_ASAP7_75t_R _24068_ (.A(_05096_),
    .B(_05097_),
    .Y(_05098_));
 BUFx6f_ASAP7_75t_R _24069_ (.A(_05098_),
    .Y(_05099_));
 BUFx4f_ASAP7_75t_R _24070_ (.A(_01457_),
    .Y(_05100_));
 BUFx6f_ASAP7_75t_R _24071_ (.A(_00069_),
    .Y(_05101_));
 NAND2x1_ASAP7_75t_R _24072_ (.A(_05100_),
    .B(_05101_),
    .Y(_05102_));
 BUFx3_ASAP7_75t_R _24073_ (.A(_05102_),
    .Y(_05103_));
 OR4x1_ASAP7_75t_R _24074_ (.A(_05093_),
    .B(_05095_),
    .C(_05099_),
    .D(_05103_),
    .Y(_05104_));
 INVx3_ASAP7_75t_R _24075_ (.A(_02212_),
    .Y(_05105_));
 AND3x2_ASAP7_75t_R _24076_ (.A(_04928_),
    .B(_04940_),
    .C(_05096_),
    .Y(_05106_));
 AND2x2_ASAP7_75t_R _24077_ (.A(_05105_),
    .B(_05106_),
    .Y(_05107_));
 BUFx4f_ASAP7_75t_R _24078_ (.A(_05107_),
    .Y(_05108_));
 AO21x1_ASAP7_75t_R _24079_ (.A1(_05092_),
    .A2(_05104_),
    .B(_05108_),
    .Y(_00005_));
 BUFx4f_ASAP7_75t_R _24080_ (.A(_04877_),
    .Y(_05109_));
 NOR3x1_ASAP7_75t_R _24081_ (.A(_04867_),
    .B(_04874_),
    .C(_04881_),
    .Y(_05110_));
 OA31x2_ASAP7_75t_R _24082_ (.A1(_05110_),
    .A2(_04900_),
    .A3(_04902_),
    .B1(_04899_),
    .Y(_05111_));
 AND4x1_ASAP7_75t_R _24083_ (.A(_04897_),
    .B(_04882_),
    .C(_04887_),
    .D(_04890_),
    .Y(_05112_));
 AO22x1_ASAP7_75t_R _24084_ (.A1(_17255_),
    .A2(_17256_),
    .B1(_04412_),
    .B2(_04413_),
    .Y(_05113_));
 OR5x2_ASAP7_75t_R _24085_ (.A(\alu_adder_result_ex[29] ),
    .B(_05111_),
    .C(_05112_),
    .D(\alu_adder_result_ex[30] ),
    .E(_05113_),
    .Y(_05114_));
 OR5x2_ASAP7_75t_R _24086_ (.A(\alu_adder_result_ex[10] ),
    .B(\alu_adder_result_ex[16] ),
    .C(\alu_adder_result_ex[20] ),
    .D(\alu_adder_result_ex[25] ),
    .E(\alu_adder_result_ex[27] ),
    .Y(_05115_));
 OA21x2_ASAP7_75t_R _24087_ (.A1(_15240_),
    .A2(_15241_),
    .B(_00800_),
    .Y(_05116_));
 OA21x2_ASAP7_75t_R _24088_ (.A1(_00799_),
    .A2(_05116_),
    .B(_00803_),
    .Y(_05117_));
 XOR2x2_ASAP7_75t_R _24089_ (.A(_00802_),
    .B(_05117_),
    .Y(\alu_adder_result_ex[5] ));
 OA21x2_ASAP7_75t_R _24090_ (.A1(_00415_),
    .A2(_02229_),
    .B(_00794_),
    .Y(_05118_));
 OA21x2_ASAP7_75t_R _24091_ (.A1(net1993),
    .A2(_05118_),
    .B(_00797_),
    .Y(_05119_));
 XOR2x2_ASAP7_75t_R _24092_ (.A(_00796_),
    .B(_05119_),
    .Y(\alu_adder_result_ex[3] ));
 OR4x1_ASAP7_75t_R _24093_ (.A(_18762_),
    .B(\alu_adder_result_ex[7] ),
    .C(\alu_adder_result_ex[5] ),
    .D(\alu_adder_result_ex[3] ),
    .Y(_05120_));
 OR4x1_ASAP7_75t_R _24094_ (.A(\alu_adder_result_ex[9] ),
    .B(\alu_adder_result_ex[11] ),
    .C(\alu_adder_result_ex[17] ),
    .D(_05120_),
    .Y(_05121_));
 OR5x1_ASAP7_75t_R _24095_ (.A(\alu_adder_result_ex[13] ),
    .B(\alu_adder_result_ex[15] ),
    .C(\alu_adder_result_ex[21] ),
    .D(\alu_adder_result_ex[23] ),
    .E(_05121_),
    .Y(_05122_));
 OR4x1_ASAP7_75t_R _24096_ (.A(\alu_adder_result_ex[12] ),
    .B(\alu_adder_result_ex[14] ),
    .C(\alu_adder_result_ex[19] ),
    .D(_05122_),
    .Y(_05123_));
 AO21x1_ASAP7_75t_R _24097_ (.A1(_14920_),
    .A2(_14919_),
    .B(_15263_),
    .Y(_05124_));
 OA21x2_ASAP7_75t_R _24098_ (.A1(_16268_),
    .A2(_05124_),
    .B(_15257_),
    .Y(_05125_));
 XNOR2x2_ASAP7_75t_R _24099_ (.A(net1994),
    .B(_05125_),
    .Y(_05126_));
 NAND2x1_ASAP7_75t_R _24100_ (.A(_15417_),
    .B(_05126_),
    .Y(_05127_));
 XNOR2x2_ASAP7_75t_R _24101_ (.A(_00799_),
    .B(_16766_),
    .Y(_05128_));
 CKINVDCx6p67_ASAP7_75t_R _24102_ (.A(_05128_),
    .Y(\alu_adder_result_ex[4] ));
 NAND2x1_ASAP7_75t_R _24103_ (.A(_16531_),
    .B(_17017_),
    .Y(_05129_));
 OR5x2_ASAP7_75t_R _24104_ (.A(\alu_adder_result_ex[6] ),
    .B(_05123_),
    .C(_05127_),
    .D(\alu_adder_result_ex[4] ),
    .E(_05129_),
    .Y(_05130_));
 OR3x4_ASAP7_75t_R _24105_ (.A(_05114_),
    .B(_05115_),
    .C(_05130_),
    .Y(_05131_));
 BUFx6f_ASAP7_75t_R _24106_ (.A(_05106_),
    .Y(_05132_));
 INVx2_ASAP7_75t_R _24107_ (.A(_02211_),
    .Y(_05133_));
 OA211x2_ASAP7_75t_R _24108_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_05131_),
    .B(_05132_),
    .C(_05133_),
    .Y(_05134_));
 AO21x1_ASAP7_75t_R _24109_ (.A1(_05109_),
    .A2(_05099_),
    .B(_05134_),
    .Y(_00004_));
 INVx3_ASAP7_75t_R _24110_ (.A(_04638_),
    .Y(_05135_));
 NOR3x2_ASAP7_75t_R _24111_ (.B(_05115_),
    .C(_05130_),
    .Y(_05136_),
    .A(_05114_));
 AND2x2_ASAP7_75t_R _24112_ (.A(_05135_),
    .B(_05136_),
    .Y(_05137_));
 BUFx4f_ASAP7_75t_R _24113_ (.A(_04871_),
    .Y(_05138_));
 BUFx4f_ASAP7_75t_R _24114_ (.A(_05138_),
    .Y(_05139_));
 AOI211x1_ASAP7_75t_R _24115_ (.A1(_05133_),
    .A2(_05137_),
    .B(_05099_),
    .C(_05139_),
    .Y(_05140_));
 AOI21x1_ASAP7_75t_R _24116_ (.A1(_02218_),
    .A2(_05099_),
    .B(_05140_),
    .Y(_00003_));
 BUFx6f_ASAP7_75t_R _24117_ (.A(_04867_),
    .Y(_05141_));
 BUFx6f_ASAP7_75t_R _24118_ (.A(_05141_),
    .Y(_05142_));
 NAND2x2_ASAP7_75t_R _24119_ (.A(_04928_),
    .B(_04940_),
    .Y(_05143_));
 OR3x4_ASAP7_75t_R _24120_ (.A(_13567_),
    .B(_05142_),
    .C(_05143_),
    .Y(_05144_));
 INVx3_ASAP7_75t_R _24121_ (.A(_05144_),
    .Y(_05145_));
 INVx1_ASAP7_75t_R _24122_ (.A(_13617_),
    .Y(_05146_));
 OA211x2_ASAP7_75t_R _24123_ (.A1(_13560_),
    .A2(_14059_),
    .B(_05146_),
    .C(_13585_),
    .Y(_05147_));
 NOR2x1_ASAP7_75t_R _24124_ (.A(_14925_),
    .B(_05147_),
    .Y(_05148_));
 OA21x2_ASAP7_75t_R _24125_ (.A1(_02213_),
    .A2(_05148_),
    .B(_01459_),
    .Y(_05149_));
 AND2x2_ASAP7_75t_R _24126_ (.A(_02216_),
    .B(_05144_),
    .Y(_05150_));
 AOI21x1_ASAP7_75t_R _24127_ (.A1(_05145_),
    .A2(_05149_),
    .B(_05150_),
    .Y(_00000_));
 OR3x1_ASAP7_75t_R _24128_ (.A(_02213_),
    .B(_04867_),
    .C(_05147_),
    .Y(_05151_));
 BUFx3_ASAP7_75t_R _24129_ (.A(_05151_),
    .Y(_05152_));
 BUFx6f_ASAP7_75t_R _24130_ (.A(_05152_),
    .Y(_05153_));
 BUFx10_ASAP7_75t_R _24131_ (.A(_01459_),
    .Y(_05154_));
 AND2x2_ASAP7_75t_R _24132_ (.A(_05154_),
    .B(_05144_),
    .Y(_05155_));
 AOI21x1_ASAP7_75t_R _24133_ (.A1(_05145_),
    .A2(_05153_),
    .B(_05155_),
    .Y(_00001_));
 BUFx4f_ASAP7_75t_R _24134_ (.A(_02217_),
    .Y(_05156_));
 BUFx4f_ASAP7_75t_R _24135_ (.A(_05156_),
    .Y(_05157_));
 BUFx4f_ASAP7_75t_R _24136_ (.A(_05132_),
    .Y(_05158_));
 BUFx4f_ASAP7_75t_R _24137_ (.A(_01816_),
    .Y(_05159_));
 BUFx6f_ASAP7_75t_R _24138_ (.A(_05159_),
    .Y(_05160_));
 OR5x1_ASAP7_75t_R _24139_ (.A(_05093_),
    .B(_05095_),
    .C(_05160_),
    .D(_05099_),
    .E(_05103_),
    .Y(_05161_));
 OAI21x1_ASAP7_75t_R _24140_ (.A1(_05157_),
    .A2(_05158_),
    .B(_05161_),
    .Y(_00002_));
 INVx1_ASAP7_75t_R _24141_ (.A(_00787_),
    .Y(\cs_registers_i.mhpmcounter[2][0] ));
 INVx1_ASAP7_75t_R _24142_ (.A(_00786_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[0] ));
 INVx6_ASAP7_75t_R _24143_ (.A(net52),
    .Y(\alu_adder_result_ex[0] ));
 INVx6_ASAP7_75t_R _24144_ (.A(_05126_),
    .Y(\alu_adder_result_ex[2] ));
 INVx1_ASAP7_75t_R _24145_ (.A(_18868_),
    .Y(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ));
 BUFx4f_ASAP7_75t_R _24146_ (.A(_18867_),
    .Y(_05162_));
 INVx4_ASAP7_75t_R _24147_ (.A(_05162_),
    .Y(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ));
 NAND2x2_ASAP7_75t_R _24148_ (.A(_05154_),
    .B(_02214_),
    .Y(_05163_));
 BUFx4f_ASAP7_75t_R _24149_ (.A(_05163_),
    .Y(_05164_));
 AND2x4_ASAP7_75t_R _24150_ (.A(_05154_),
    .B(_02214_),
    .Y(_05165_));
 AND3x1_ASAP7_75t_R _24151_ (.A(_13821_),
    .B(_13852_),
    .C(_05165_),
    .Y(_05166_));
 AO21x1_ASAP7_75t_R _24152_ (.A1(_16094_),
    .A2(_05164_),
    .B(_05166_),
    .Y(_05167_));
 BUFx6f_ASAP7_75t_R _24153_ (.A(_05167_),
    .Y(_05168_));
 AND2x4_ASAP7_75t_R _24154_ (.A(_16117_),
    .B(_16140_),
    .Y(_05169_));
 NAND2x2_ASAP7_75t_R _24155_ (.A(_05154_),
    .B(_02213_),
    .Y(_05170_));
 BUFx3_ASAP7_75t_R _24156_ (.A(_05170_),
    .Y(_05171_));
 AND2x4_ASAP7_75t_R _24157_ (.A(_05154_),
    .B(_02213_),
    .Y(_05172_));
 AND3x1_ASAP7_75t_R _24158_ (.A(_13901_),
    .B(_13941_),
    .C(_05172_),
    .Y(_05173_));
 AO21x2_ASAP7_75t_R _24159_ (.A1(_05169_),
    .A2(_05171_),
    .B(_05173_),
    .Y(_05174_));
 BUFx4f_ASAP7_75t_R _24160_ (.A(_05174_),
    .Y(_05175_));
 AND2x2_ASAP7_75t_R _24161_ (.A(_05168_),
    .B(_05175_),
    .Y(_18873_));
 BUFx6f_ASAP7_75t_R _24162_ (.A(_05152_),
    .Y(_05176_));
 BUFx4f_ASAP7_75t_R _24163_ (.A(_05165_),
    .Y(_05177_));
 OA21x2_ASAP7_75t_R _24164_ (.A1(_02213_),
    .A2(_05148_),
    .B(_05177_),
    .Y(_05178_));
 BUFx3_ASAP7_75t_R _24165_ (.A(_05178_),
    .Y(_05179_));
 BUFx4f_ASAP7_75t_R _24166_ (.A(_00953_),
    .Y(_05180_));
 OAI22x1_ASAP7_75t_R _24167_ (.A1(_00447_),
    .A2(_05176_),
    .B1(_05179_),
    .B2(_05180_),
    .Y(_18874_));
 AND3x1_ASAP7_75t_R _24168_ (.A(_13514_),
    .B(_13549_),
    .C(_05165_),
    .Y(_05181_));
 AO21x1_ASAP7_75t_R _24169_ (.A1(_16209_),
    .A2(_05164_),
    .B(_05181_),
    .Y(_05182_));
 BUFx4f_ASAP7_75t_R _24170_ (.A(_05182_),
    .Y(_05183_));
 BUFx6f_ASAP7_75t_R _24171_ (.A(_05183_),
    .Y(_05184_));
 NAND2x1_ASAP7_75t_R _24172_ (.A(_05175_),
    .B(_05184_),
    .Y(_17349_));
 BUFx4f_ASAP7_75t_R _24173_ (.A(_05165_),
    .Y(_05185_));
 AND2x2_ASAP7_75t_R _24174_ (.A(_14148_),
    .B(_05185_),
    .Y(_05186_));
 AO21x2_ASAP7_75t_R _24175_ (.A1(_05164_),
    .A2(_16354_),
    .B(_05186_),
    .Y(_05187_));
 BUFx3_ASAP7_75t_R _24176_ (.A(_05187_),
    .Y(_05188_));
 AND2x2_ASAP7_75t_R _24177_ (.A(_05175_),
    .B(_05188_),
    .Y(_18884_));
 AND2x2_ASAP7_75t_R _24178_ (.A(_16232_),
    .B(_16255_),
    .Y(_05189_));
 AND3x1_ASAP7_75t_R _24179_ (.A(_13733_),
    .B(_13768_),
    .C(_05172_),
    .Y(_05190_));
 AO21x2_ASAP7_75t_R _24180_ (.A1(_05189_),
    .A2(_05171_),
    .B(_05190_),
    .Y(_05191_));
 BUFx6f_ASAP7_75t_R _24181_ (.A(_05191_),
    .Y(_05192_));
 NAND2x1_ASAP7_75t_R _24182_ (.A(_05184_),
    .B(_05192_),
    .Y(_17351_));
 AND2x2_ASAP7_75t_R _24183_ (.A(_14225_),
    .B(_05185_),
    .Y(_05193_));
 AO21x2_ASAP7_75t_R _24184_ (.A1(_05164_),
    .A2(_16466_),
    .B(_05193_),
    .Y(_05194_));
 BUFx3_ASAP7_75t_R _24185_ (.A(_05194_),
    .Y(_05195_));
 AND2x2_ASAP7_75t_R _24186_ (.A(_05175_),
    .B(_05195_),
    .Y(_18887_));
 AND2x2_ASAP7_75t_R _24187_ (.A(_05188_),
    .B(_05192_),
    .Y(_18886_));
 AND2x6_ASAP7_75t_R _24188_ (.A(_14841_),
    .B(_14877_),
    .Y(_05196_));
 BUFx4f_ASAP7_75t_R _24189_ (.A(_05172_),
    .Y(_05197_));
 AND3x1_ASAP7_75t_R _24190_ (.A(_16377_),
    .B(_16400_),
    .C(_05170_),
    .Y(_05198_));
 AO21x2_ASAP7_75t_R _24191_ (.A1(_05196_),
    .A2(_05197_),
    .B(_05198_),
    .Y(_05199_));
 BUFx6f_ASAP7_75t_R _24192_ (.A(_05199_),
    .Y(_05200_));
 NAND2x1_ASAP7_75t_R _24193_ (.A(_05184_),
    .B(_05200_),
    .Y(_17353_));
 NOR2x1_ASAP7_75t_R _24194_ (.A(_05185_),
    .B(_16592_),
    .Y(_05201_));
 AO21x2_ASAP7_75t_R _24195_ (.A1(_14295_),
    .A2(_05177_),
    .B(_05201_),
    .Y(_05202_));
 BUFx4f_ASAP7_75t_R _24196_ (.A(_05202_),
    .Y(_05203_));
 AND2x2_ASAP7_75t_R _24197_ (.A(_05175_),
    .B(_05203_),
    .Y(_17357_));
 AND2x2_ASAP7_75t_R _24198_ (.A(_05192_),
    .B(_05195_),
    .Y(_17356_));
 AND2x2_ASAP7_75t_R _24199_ (.A(_05188_),
    .B(_05199_),
    .Y(_17358_));
 AND2x6_ASAP7_75t_R _24200_ (.A(_14953_),
    .B(_14977_),
    .Y(_05204_));
 AND3x1_ASAP7_75t_R _24201_ (.A(_16489_),
    .B(_16512_),
    .C(_05170_),
    .Y(_05205_));
 AO21x2_ASAP7_75t_R _24202_ (.A1(_05204_),
    .A2(_05197_),
    .B(_05205_),
    .Y(_05206_));
 BUFx6f_ASAP7_75t_R _24203_ (.A(_05206_),
    .Y(_05207_));
 NAND2x1_ASAP7_75t_R _24204_ (.A(_05184_),
    .B(_05207_),
    .Y(_17361_));
 OR2x2_ASAP7_75t_R _24205_ (.A(_14371_),
    .B(_05164_),
    .Y(_05208_));
 OAI21x1_ASAP7_75t_R _24206_ (.A1(_16706_),
    .A2(_05177_),
    .B(_05208_),
    .Y(_05209_));
 AND2x2_ASAP7_75t_R _24207_ (.A(_05175_),
    .B(_05209_),
    .Y(_18902_));
 AND2x2_ASAP7_75t_R _24208_ (.A(_05191_),
    .B(_05203_),
    .Y(_17373_));
 AND2x2_ASAP7_75t_R _24209_ (.A(_05195_),
    .B(_05199_),
    .Y(_17372_));
 AND2x2_ASAP7_75t_R _24210_ (.A(_05188_),
    .B(_05206_),
    .Y(_17374_));
 AND2x6_ASAP7_75t_R _24211_ (.A(_15024_),
    .B(_15052_),
    .Y(_05210_));
 AND3x1_ASAP7_75t_R _24212_ (.A(_16618_),
    .B(_16641_),
    .C(_05170_),
    .Y(_05211_));
 AO21x2_ASAP7_75t_R _24213_ (.A1(_05210_),
    .A2(_05197_),
    .B(_05211_),
    .Y(_05212_));
 BUFx6f_ASAP7_75t_R _24214_ (.A(_05212_),
    .Y(_05213_));
 NAND2x1_ASAP7_75t_R _24215_ (.A(_05184_),
    .B(_05213_),
    .Y(_17376_));
 NOR2x1_ASAP7_75t_R _24216_ (.A(_16836_),
    .B(_05185_),
    .Y(_05214_));
 AO21x1_ASAP7_75t_R _24217_ (.A1(_14426_),
    .A2(_05177_),
    .B(_05214_),
    .Y(_05215_));
 BUFx6f_ASAP7_75t_R _24218_ (.A(_05215_),
    .Y(_05216_));
 AND2x2_ASAP7_75t_R _24219_ (.A(_05175_),
    .B(_05216_),
    .Y(_18911_));
 AND2x2_ASAP7_75t_R _24220_ (.A(_05191_),
    .B(_05209_),
    .Y(_18912_));
 AND2x2_ASAP7_75t_R _24221_ (.A(_05199_),
    .B(_05203_),
    .Y(_17389_));
 AND2x2_ASAP7_75t_R _24222_ (.A(_05195_),
    .B(_05206_),
    .Y(_17388_));
 AND2x2_ASAP7_75t_R _24223_ (.A(_05188_),
    .B(_05212_),
    .Y(_17390_));
 AND2x4_ASAP7_75t_R _24224_ (.A(_16728_),
    .B(_16751_),
    .Y(_05217_));
 AND3x1_ASAP7_75t_R _24225_ (.A(_15087_),
    .B(_15113_),
    .C(_05197_),
    .Y(_05218_));
 AO21x2_ASAP7_75t_R _24226_ (.A1(_05217_),
    .A2(_05171_),
    .B(_05218_),
    .Y(_05219_));
 BUFx6f_ASAP7_75t_R _24227_ (.A(_05219_),
    .Y(_05220_));
 NAND2x1_ASAP7_75t_R _24228_ (.A(_05184_),
    .B(_05220_),
    .Y(_17394_));
 AND2x2_ASAP7_75t_R _24229_ (.A(_14486_),
    .B(_05165_),
    .Y(_05221_));
 AO21x1_ASAP7_75t_R _24230_ (.A1(_16946_),
    .A2(_05164_),
    .B(_05221_),
    .Y(_05222_));
 BUFx4f_ASAP7_75t_R _24231_ (.A(_05222_),
    .Y(_05223_));
 BUFx6f_ASAP7_75t_R _24232_ (.A(_05223_),
    .Y(_05224_));
 NAND2x1_ASAP7_75t_R _24233_ (.A(_05175_),
    .B(_05224_),
    .Y(_17401_));
 AND2x2_ASAP7_75t_R _24234_ (.A(_05203_),
    .B(_05206_),
    .Y(_17406_));
 AND2x2_ASAP7_75t_R _24235_ (.A(_05195_),
    .B(_05212_),
    .Y(_17405_));
 AND2x2_ASAP7_75t_R _24236_ (.A(_05188_),
    .B(_05219_),
    .Y(_17407_));
 AND2x4_ASAP7_75t_R _24237_ (.A(_16858_),
    .B(_16882_),
    .Y(_05225_));
 AND3x1_ASAP7_75t_R _24238_ (.A(_15154_),
    .B(_15179_),
    .C(_05197_),
    .Y(_05226_));
 AO21x2_ASAP7_75t_R _24239_ (.A1(_05225_),
    .A2(_05171_),
    .B(_05226_),
    .Y(_05227_));
 BUFx6f_ASAP7_75t_R _24240_ (.A(_05227_),
    .Y(_05228_));
 NAND2x1_ASAP7_75t_R _24241_ (.A(_05184_),
    .B(_05228_),
    .Y(_17414_));
 INVx1_ASAP7_75t_R _24242_ (.A(_02328_),
    .Y(_17385_));
 OR3x4_ASAP7_75t_R _24243_ (.A(_14500_),
    .B(_14515_),
    .C(_14544_),
    .Y(_05229_));
 BUFx4f_ASAP7_75t_R _24244_ (.A(_05229_),
    .Y(_05230_));
 NOR2x1_ASAP7_75t_R _24245_ (.A(_17076_),
    .B(_05185_),
    .Y(_05231_));
 AO21x1_ASAP7_75t_R _24246_ (.A1(_05230_),
    .A2(_05177_),
    .B(_05231_),
    .Y(_05232_));
 BUFx6f_ASAP7_75t_R _24247_ (.A(_05232_),
    .Y(_05233_));
 AND2x2_ASAP7_75t_R _24248_ (.A(_05175_),
    .B(_05233_),
    .Y(_18937_));
 NAND2x1_ASAP7_75t_R _24249_ (.A(_05192_),
    .B(_05224_),
    .Y(_17426_));
 AND2x2_ASAP7_75t_R _24250_ (.A(_05203_),
    .B(_05212_),
    .Y(_17430_));
 AND2x2_ASAP7_75t_R _24251_ (.A(_05195_),
    .B(_05219_),
    .Y(_17432_));
 AND2x2_ASAP7_75t_R _24252_ (.A(_05188_),
    .B(_05227_),
    .Y(_17431_));
 AND2x4_ASAP7_75t_R _24253_ (.A(_16969_),
    .B(_16992_),
    .Y(_05234_));
 AND3x1_ASAP7_75t_R _24254_ (.A(_15206_),
    .B(_15234_),
    .C(_05197_),
    .Y(_05235_));
 AO21x2_ASAP7_75t_R _24255_ (.A1(_05234_),
    .A2(_05171_),
    .B(_05235_),
    .Y(_05236_));
 BUFx6f_ASAP7_75t_R _24256_ (.A(_05236_),
    .Y(_05237_));
 NAND2x1_ASAP7_75t_R _24257_ (.A(_05184_),
    .B(_05237_),
    .Y(_17434_));
 NOR2x1_ASAP7_75t_R _24258_ (.A(_17185_),
    .B(_05185_),
    .Y(_05238_));
 AO21x1_ASAP7_75t_R _24259_ (.A1(_14603_),
    .A2(_05185_),
    .B(_05238_),
    .Y(_05239_));
 BUFx6f_ASAP7_75t_R _24260_ (.A(_05239_),
    .Y(_05240_));
 AND2x2_ASAP7_75t_R _24261_ (.A(_05174_),
    .B(_05240_),
    .Y(_18946_));
 AND2x2_ASAP7_75t_R _24262_ (.A(_05191_),
    .B(_05233_),
    .Y(_18945_));
 NAND2x1_ASAP7_75t_R _24263_ (.A(_05200_),
    .B(_05224_),
    .Y(_17450_));
 AND2x2_ASAP7_75t_R _24264_ (.A(_05203_),
    .B(_05219_),
    .Y(_17454_));
 AND2x2_ASAP7_75t_R _24265_ (.A(_05195_),
    .B(_05227_),
    .Y(_17453_));
 AND2x2_ASAP7_75t_R _24266_ (.A(_05188_),
    .B(_05236_),
    .Y(_17455_));
 AND2x4_ASAP7_75t_R _24267_ (.A(_17098_),
    .B(_17121_),
    .Y(_05241_));
 AND3x1_ASAP7_75t_R _24268_ (.A(_15303_),
    .B(_15332_),
    .C(_05197_),
    .Y(_05242_));
 AO21x2_ASAP7_75t_R _24269_ (.A1(_05241_),
    .A2(_05171_),
    .B(_05242_),
    .Y(_05243_));
 BUFx6f_ASAP7_75t_R _24270_ (.A(_05243_),
    .Y(_05244_));
 NAND2x1_ASAP7_75t_R _24271_ (.A(_05184_),
    .B(_05244_),
    .Y(_17459_));
 AND3x1_ASAP7_75t_R _24272_ (.A(_17284_),
    .B(_17315_),
    .C(_05163_),
    .Y(_05245_));
 AO21x2_ASAP7_75t_R _24273_ (.A1(_14666_),
    .A2(_05177_),
    .B(_05245_),
    .Y(_05246_));
 BUFx4f_ASAP7_75t_R _24274_ (.A(_05246_),
    .Y(_05247_));
 BUFx6f_ASAP7_75t_R _24275_ (.A(_05247_),
    .Y(_05248_));
 NAND2x1_ASAP7_75t_R _24276_ (.A(_05175_),
    .B(_05248_),
    .Y(_17477_));
 NAND2x1_ASAP7_75t_R _24277_ (.A(_05207_),
    .B(_05224_),
    .Y(_17480_));
 AND2x2_ASAP7_75t_R _24278_ (.A(_05203_),
    .B(_05227_),
    .Y(_17484_));
 AND2x2_ASAP7_75t_R _24279_ (.A(_05195_),
    .B(_05236_),
    .Y(_17483_));
 AND2x2_ASAP7_75t_R _24280_ (.A(_05188_),
    .B(_05243_),
    .Y(_17485_));
 AND2x4_ASAP7_75t_R _24281_ (.A(_17207_),
    .B(_17230_),
    .Y(_05249_));
 AND3x1_ASAP7_75t_R _24282_ (.A(_15365_),
    .B(_15390_),
    .C(_05197_),
    .Y(_05250_));
 AO21x2_ASAP7_75t_R _24283_ (.A1(_05249_),
    .A2(_05171_),
    .B(_05250_),
    .Y(_05251_));
 BUFx6f_ASAP7_75t_R _24284_ (.A(_05251_),
    .Y(_05252_));
 NAND2x1_ASAP7_75t_R _24285_ (.A(_05184_),
    .B(_05252_),
    .Y(_17490_));
 AND3x1_ASAP7_75t_R _24286_ (.A(_04311_),
    .B(_04342_),
    .C(_05164_),
    .Y(_05253_));
 AO21x2_ASAP7_75t_R _24287_ (.A1(_14723_),
    .A2(_05177_),
    .B(_05253_),
    .Y(_05254_));
 BUFx6f_ASAP7_75t_R _24288_ (.A(_05254_),
    .Y(_05255_));
 AND2x2_ASAP7_75t_R _24289_ (.A(_05174_),
    .B(_05255_),
    .Y(_18974_));
 NAND2x1_ASAP7_75t_R _24290_ (.A(_05192_),
    .B(_05248_),
    .Y(_17505_));
 NAND2x1_ASAP7_75t_R _24291_ (.A(_05213_),
    .B(_05224_),
    .Y(_17508_));
 AND2x2_ASAP7_75t_R _24292_ (.A(_05203_),
    .B(_05236_),
    .Y(_17512_));
 AND2x2_ASAP7_75t_R _24293_ (.A(_05195_),
    .B(_05243_),
    .Y(_17511_));
 AND2x2_ASAP7_75t_R _24294_ (.A(_05188_),
    .B(_05251_),
    .Y(_17513_));
 AND2x2_ASAP7_75t_R _24295_ (.A(_15440_),
    .B(_15463_),
    .Y(_05256_));
 AND3x1_ASAP7_75t_R _24296_ (.A(_17338_),
    .B(_04279_),
    .C(_05170_),
    .Y(_05257_));
 AO21x1_ASAP7_75t_R _24297_ (.A1(_05256_),
    .A2(_05197_),
    .B(_05257_),
    .Y(_05258_));
 BUFx4f_ASAP7_75t_R _24298_ (.A(_05258_),
    .Y(_05259_));
 BUFx6f_ASAP7_75t_R _24299_ (.A(_05259_),
    .Y(_05260_));
 NAND2x1_ASAP7_75t_R _24300_ (.A(_05183_),
    .B(_05260_),
    .Y(_17520_));
 AND2x4_ASAP7_75t_R _24301_ (.A(_15554_),
    .B(_15592_),
    .Y(_05261_));
 NOR2x1_ASAP7_75t_R _24302_ (.A(_04473_),
    .B(_05185_),
    .Y(_05262_));
 AO21x2_ASAP7_75t_R _24303_ (.A1(_05261_),
    .A2(_05177_),
    .B(_05262_),
    .Y(_05263_));
 BUFx6f_ASAP7_75t_R _24304_ (.A(_05263_),
    .Y(_05264_));
 AND2x2_ASAP7_75t_R _24305_ (.A(_05174_),
    .B(_05264_),
    .Y(_18989_));
 AND2x2_ASAP7_75t_R _24306_ (.A(_05191_),
    .B(_05255_),
    .Y(_18988_));
 NAND2x1_ASAP7_75t_R _24307_ (.A(_05200_),
    .B(_05248_),
    .Y(_17534_));
 NAND2x1_ASAP7_75t_R _24308_ (.A(_05220_),
    .B(_05224_),
    .Y(_17539_));
 AND2x2_ASAP7_75t_R _24309_ (.A(_05203_),
    .B(_05243_),
    .Y(_17543_));
 AND2x2_ASAP7_75t_R _24310_ (.A(_05195_),
    .B(_05251_),
    .Y(_17542_));
 AND2x2_ASAP7_75t_R _24311_ (.A(_05187_),
    .B(_05259_),
    .Y(_17544_));
 AND2x4_ASAP7_75t_R _24312_ (.A(_04365_),
    .B(_04388_),
    .Y(_05265_));
 AND3x1_ASAP7_75t_R _24313_ (.A(_14775_),
    .B(_14803_),
    .C(_05172_),
    .Y(_05266_));
 AO21x1_ASAP7_75t_R _24314_ (.A1(_05265_),
    .A2(_05171_),
    .B(_05266_),
    .Y(_05267_));
 BUFx4f_ASAP7_75t_R _24315_ (.A(_05267_),
    .Y(_05268_));
 BUFx6f_ASAP7_75t_R _24316_ (.A(_05268_),
    .Y(_05269_));
 NAND2x1_ASAP7_75t_R _24317_ (.A(_05183_),
    .B(_05269_),
    .Y(_17553_));
 AND3x1_ASAP7_75t_R _24318_ (.A(_04551_),
    .B(_04582_),
    .C(_05164_),
    .Y(_05270_));
 AO21x2_ASAP7_75t_R _24319_ (.A1(_15671_),
    .A2(_05177_),
    .B(_05270_),
    .Y(_05271_));
 BUFx6f_ASAP7_75t_R _24320_ (.A(_05271_),
    .Y(_05272_));
 AND2x2_ASAP7_75t_R _24321_ (.A(_05174_),
    .B(_05272_),
    .Y(_17567_));
 AND2x2_ASAP7_75t_R _24322_ (.A(_05191_),
    .B(_05264_),
    .Y(_17566_));
 AND2x2_ASAP7_75t_R _24323_ (.A(_05199_),
    .B(_05255_),
    .Y(_17568_));
 NAND2x1_ASAP7_75t_R _24324_ (.A(_05207_),
    .B(_05248_),
    .Y(_17572_));
 NAND2x1_ASAP7_75t_R _24325_ (.A(_05224_),
    .B(_05228_),
    .Y(_17577_));
 AND2x2_ASAP7_75t_R _24326_ (.A(_05202_),
    .B(_05251_),
    .Y(_17584_));
 AND2x2_ASAP7_75t_R _24327_ (.A(_05194_),
    .B(_05259_),
    .Y(_17583_));
 AND2x2_ASAP7_75t_R _24328_ (.A(_05187_),
    .B(_05268_),
    .Y(_17582_));
 AND2x4_ASAP7_75t_R _24329_ (.A(_04495_),
    .B(_04518_),
    .Y(_05273_));
 AND3x1_ASAP7_75t_R _24330_ (.A(_13979_),
    .B(_14013_),
    .C(_05172_),
    .Y(_05274_));
 AO21x1_ASAP7_75t_R _24331_ (.A1(_05273_),
    .A2(_05171_),
    .B(_05274_),
    .Y(_05275_));
 BUFx4f_ASAP7_75t_R _24332_ (.A(_05275_),
    .Y(_05276_));
 BUFx6f_ASAP7_75t_R _24333_ (.A(_05276_),
    .Y(_05277_));
 NAND2x1_ASAP7_75t_R _24334_ (.A(_05183_),
    .B(_05277_),
    .Y(_17592_));
 NOR2x1_ASAP7_75t_R _24335_ (.A(_04697_),
    .B(_05185_),
    .Y(_05278_));
 AO21x1_ASAP7_75t_R _24336_ (.A1(_15816_),
    .A2(_05177_),
    .B(_05278_),
    .Y(_05279_));
 BUFx6f_ASAP7_75t_R _24337_ (.A(_05279_),
    .Y(_05280_));
 AND2x2_ASAP7_75t_R _24338_ (.A(_05174_),
    .B(_05280_),
    .Y(_19020_));
 NAND2x1_ASAP7_75t_R _24339_ (.A(_05192_),
    .B(_05272_),
    .Y(_17609_));
 NAND2x1_ASAP7_75t_R _24340_ (.A(_05213_),
    .B(_05248_),
    .Y(_17612_));
 NAND2x1_ASAP7_75t_R _24341_ (.A(_05224_),
    .B(_05237_),
    .Y(_17619_));
 AND2x2_ASAP7_75t_R _24342_ (.A(_05202_),
    .B(_05259_),
    .Y(_17626_));
 AND2x2_ASAP7_75t_R _24343_ (.A(_05194_),
    .B(_05268_),
    .Y(_17625_));
 AND2x2_ASAP7_75t_R _24344_ (.A(_05187_),
    .B(_05276_),
    .Y(_17624_));
 AND2x4_ASAP7_75t_R _24345_ (.A(_04605_),
    .B(_04628_),
    .Y(_05281_));
 AND3x1_ASAP7_75t_R _24346_ (.A(_15698_),
    .B(_15723_),
    .C(_05172_),
    .Y(_05282_));
 AO21x1_ASAP7_75t_R _24347_ (.A1(_05281_),
    .A2(_05171_),
    .B(_05282_),
    .Y(_05283_));
 BUFx4f_ASAP7_75t_R _24348_ (.A(_05283_),
    .Y(_05284_));
 BUFx6f_ASAP7_75t_R _24349_ (.A(_05284_),
    .Y(_05285_));
 NAND2x1_ASAP7_75t_R _24350_ (.A(_05183_),
    .B(_05285_),
    .Y(_17633_));
 AO21x1_ASAP7_75t_R _24351_ (.A1(_04875_),
    .A2(_04876_),
    .B(_05185_),
    .Y(_05286_));
 OA21x2_ASAP7_75t_R _24352_ (.A1(_15950_),
    .A2(_05164_),
    .B(_05286_),
    .Y(_05287_));
 BUFx6f_ASAP7_75t_R _24353_ (.A(_05287_),
    .Y(_05288_));
 AND2x2_ASAP7_75t_R _24354_ (.A(_05174_),
    .B(_05288_),
    .Y(_19039_));
 AND2x2_ASAP7_75t_R _24355_ (.A(_05191_),
    .B(_05280_),
    .Y(_19038_));
 AND2x2_ASAP7_75t_R _24356_ (.A(_05199_),
    .B(_05272_),
    .Y(_17649_));
 AND2x2_ASAP7_75t_R _24357_ (.A(_05206_),
    .B(_05264_),
    .Y(_17648_));
 AND2x2_ASAP7_75t_R _24358_ (.A(_05212_),
    .B(_05255_),
    .Y(_17650_));
 NAND2x1_ASAP7_75t_R _24359_ (.A(_05220_),
    .B(_05248_),
    .Y(_17653_));
 NAND2x1_ASAP7_75t_R _24360_ (.A(_05224_),
    .B(_05244_),
    .Y(_17663_));
 AND2x2_ASAP7_75t_R _24361_ (.A(_05202_),
    .B(_05268_),
    .Y(_17667_));
 AND2x2_ASAP7_75t_R _24362_ (.A(_05194_),
    .B(_05276_),
    .Y(_17669_));
 AND2x2_ASAP7_75t_R _24363_ (.A(_05187_),
    .B(_05284_),
    .Y(_17668_));
 AND2x4_ASAP7_75t_R _24364_ (.A(_04719_),
    .B(_04742_),
    .Y(_05289_));
 AND3x1_ASAP7_75t_R _24365_ (.A(_15839_),
    .B(_15863_),
    .C(_05172_),
    .Y(_05290_));
 AO21x1_ASAP7_75t_R _24366_ (.A1(_05289_),
    .A2(_05170_),
    .B(_05290_),
    .Y(_05291_));
 BUFx4f_ASAP7_75t_R _24367_ (.A(_05291_),
    .Y(_05292_));
 BUFx6f_ASAP7_75t_R _24368_ (.A(_05292_),
    .Y(_05293_));
 NAND2x1_ASAP7_75t_R _24369_ (.A(_05183_),
    .B(_05293_),
    .Y(_17675_));
 AND2x2_ASAP7_75t_R _24370_ (.A(_13589_),
    .B(_13397_),
    .Y(_05294_));
 OA21x2_ASAP7_75t_R _24371_ (.A1(_13617_),
    .A2(_05294_),
    .B(_16286_),
    .Y(_05295_));
 AND3x4_ASAP7_75t_R _24372_ (.A(_04875_),
    .B(_04876_),
    .C(_05295_),
    .Y(_05296_));
 BUFx4f_ASAP7_75t_R _24373_ (.A(_05296_),
    .Y(_05297_));
 NAND2x2_ASAP7_75t_R _24374_ (.A(_05297_),
    .B(_05164_),
    .Y(_05298_));
 BUFx3_ASAP7_75t_R _24375_ (.A(_05298_),
    .Y(_05299_));
 INVx1_ASAP7_75t_R _24376_ (.A(_05299_),
    .Y(_17732_));
 OR2x2_ASAP7_75t_R _24377_ (.A(_05174_),
    .B(_05299_),
    .Y(_17692_));
 AND2x2_ASAP7_75t_R _24378_ (.A(_05206_),
    .B(_05272_),
    .Y(_17694_));
 AND2x2_ASAP7_75t_R _24379_ (.A(_05212_),
    .B(_05264_),
    .Y(_17696_));
 AND2x2_ASAP7_75t_R _24380_ (.A(_05219_),
    .B(_05255_),
    .Y(_17695_));
 NAND2x1_ASAP7_75t_R _24381_ (.A(_05228_),
    .B(_05248_),
    .Y(_17702_));
 NAND2x1_ASAP7_75t_R _24382_ (.A(_05224_),
    .B(_05252_),
    .Y(_17712_));
 AND2x2_ASAP7_75t_R _24383_ (.A(_05202_),
    .B(_05276_),
    .Y(_17716_));
 AND2x2_ASAP7_75t_R _24384_ (.A(_05194_),
    .B(_05284_),
    .Y(_17715_));
 AND2x2_ASAP7_75t_R _24385_ (.A(_05187_),
    .B(_05292_),
    .Y(_17717_));
 AND2x2_ASAP7_75t_R _24386_ (.A(_15978_),
    .B(_16002_),
    .Y(_05300_));
 AND2x2_ASAP7_75t_R _24387_ (.A(_04861_),
    .B(_05170_),
    .Y(_05301_));
 AO21x1_ASAP7_75t_R _24388_ (.A1(_05300_),
    .A2(_05197_),
    .B(_05301_),
    .Y(_05302_));
 BUFx4f_ASAP7_75t_R _24389_ (.A(_05302_),
    .Y(_05303_));
 AND2x2_ASAP7_75t_R _24390_ (.A(_05183_),
    .B(_05303_),
    .Y(_17728_));
 BUFx6f_ASAP7_75t_R _24391_ (.A(_16286_),
    .Y(_05304_));
 AO21x2_ASAP7_75t_R _24392_ (.A1(_13560_),
    .A2(_13396_),
    .B(_05294_),
    .Y(_05305_));
 AND2x2_ASAP7_75t_R _24393_ (.A(_05304_),
    .B(_05305_),
    .Y(_05306_));
 AND3x1_ASAP7_75t_R _24394_ (.A(_04861_),
    .B(_05306_),
    .C(_05170_),
    .Y(_05307_));
 BUFx10_ASAP7_75t_R _24395_ (.A(_05307_),
    .Y(_05308_));
 BUFx6f_ASAP7_75t_R _24396_ (.A(_05308_),
    .Y(_05309_));
 AND2x6_ASAP7_75t_R _24397_ (.A(_05168_),
    .B(_05309_),
    .Y(_17727_));
 OAI22x1_ASAP7_75t_R _24398_ (.A1(_05154_),
    .A2(_01747_),
    .B1(_05176_),
    .B2(_05180_),
    .Y(_17729_));
 OR2x2_ASAP7_75t_R _24399_ (.A(_05191_),
    .B(_05299_),
    .Y(_17743_));
 AND2x2_ASAP7_75t_R _24400_ (.A(_05212_),
    .B(_05271_),
    .Y(_17750_));
 AND2x2_ASAP7_75t_R _24401_ (.A(_05219_),
    .B(_05263_),
    .Y(_17749_));
 AND2x2_ASAP7_75t_R _24402_ (.A(_05227_),
    .B(_05254_),
    .Y(_17748_));
 NAND2x1_ASAP7_75t_R _24403_ (.A(_05237_),
    .B(_05248_),
    .Y(_17755_));
 NAND2x1_ASAP7_75t_R _24404_ (.A(_05223_),
    .B(_05260_),
    .Y(_17765_));
 AND2x2_ASAP7_75t_R _24405_ (.A(_05202_),
    .B(_05284_),
    .Y(_17772_));
 AND2x2_ASAP7_75t_R _24406_ (.A(_05194_),
    .B(_05292_),
    .Y(_17771_));
 AND2x2_ASAP7_75t_R _24407_ (.A(_05187_),
    .B(_05303_),
    .Y(_17770_));
 AND2x6_ASAP7_75t_R _24408_ (.A(_05183_),
    .B(_05309_),
    .Y(_17780_));
 OAI22x1_ASAP7_75t_R _24409_ (.A1(_05154_),
    .A2(_00232_),
    .B1(_05176_),
    .B2(_00986_),
    .Y(_17781_));
 OR2x2_ASAP7_75t_R _24410_ (.A(_05199_),
    .B(_05299_),
    .Y(_17793_));
 AND2x2_ASAP7_75t_R _24411_ (.A(_05219_),
    .B(_05271_),
    .Y(_17798_));
 AND2x2_ASAP7_75t_R _24412_ (.A(_05227_),
    .B(_05263_),
    .Y(_17797_));
 AND2x2_ASAP7_75t_R _24413_ (.A(_05236_),
    .B(_05254_),
    .Y(_17799_));
 NAND2x1_ASAP7_75t_R _24414_ (.A(_05244_),
    .B(_05248_),
    .Y(_17803_));
 NAND2x1_ASAP7_75t_R _24415_ (.A(_05223_),
    .B(_05269_),
    .Y(_17814_));
 AND2x2_ASAP7_75t_R _24416_ (.A(_05202_),
    .B(_05292_),
    .Y(_17819_));
 AND2x2_ASAP7_75t_R _24417_ (.A(_05194_),
    .B(_05303_),
    .Y(_17818_));
 NAND2x2_ASAP7_75t_R _24418_ (.A(_05309_),
    .B(_05187_),
    .Y(_17865_));
 INVx2_ASAP7_75t_R _24419_ (.A(_17865_),
    .Y(_17820_));
 NAND2x2_ASAP7_75t_R _24420_ (.A(_05304_),
    .B(_05305_),
    .Y(_05310_));
 OR3x1_ASAP7_75t_R _24421_ (.A(_05154_),
    .B(_00232_),
    .C(_05310_),
    .Y(_05311_));
 BUFx4f_ASAP7_75t_R _24422_ (.A(_05311_),
    .Y(_05312_));
 BUFx6f_ASAP7_75t_R _24423_ (.A(_05312_),
    .Y(_05313_));
 OAI21x1_ASAP7_75t_R _24424_ (.A1(_01019_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_17827_));
 OR2x2_ASAP7_75t_R _24425_ (.A(_05206_),
    .B(_05299_),
    .Y(_17838_));
 AND2x2_ASAP7_75t_R _24426_ (.A(_05227_),
    .B(_05271_),
    .Y(_17843_));
 AND2x2_ASAP7_75t_R _24427_ (.A(_05236_),
    .B(_05263_),
    .Y(_17842_));
 AND2x2_ASAP7_75t_R _24428_ (.A(_05243_),
    .B(_05254_),
    .Y(_17844_));
 NAND2x1_ASAP7_75t_R _24429_ (.A(_05248_),
    .B(_05252_),
    .Y(_17848_));
 NAND2x1_ASAP7_75t_R _24430_ (.A(_05223_),
    .B(_05277_),
    .Y(_17859_));
 BUFx6f_ASAP7_75t_R _24431_ (.A(_05303_),
    .Y(_05314_));
 NAND2x1_ASAP7_75t_R _24432_ (.A(_05203_),
    .B(_05314_),
    .Y(_17864_));
 NAND2x2_ASAP7_75t_R _24433_ (.A(_05308_),
    .B(_05194_),
    .Y(_17863_));
 INVx2_ASAP7_75t_R _24434_ (.A(_17863_),
    .Y(_17910_));
 OAI21x1_ASAP7_75t_R _24435_ (.A1(_01052_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_17873_));
 OR2x2_ASAP7_75t_R _24436_ (.A(_05212_),
    .B(_05299_),
    .Y(_17884_));
 AND2x2_ASAP7_75t_R _24437_ (.A(_05236_),
    .B(_05271_),
    .Y(_17891_));
 AND2x2_ASAP7_75t_R _24438_ (.A(_05243_),
    .B(_05263_),
    .Y(_17890_));
 AND2x2_ASAP7_75t_R _24439_ (.A(_05251_),
    .B(_05254_),
    .Y(_17889_));
 NAND2x1_ASAP7_75t_R _24440_ (.A(_05247_),
    .B(_05260_),
    .Y(_17896_));
 NAND2x1_ASAP7_75t_R _24441_ (.A(_05223_),
    .B(_05285_),
    .Y(_17905_));
 AND2x2_ASAP7_75t_R _24442_ (.A(_05202_),
    .B(_05309_),
    .Y(_17911_));
 BUFx4f_ASAP7_75t_R _24443_ (.A(_01085_),
    .Y(_05315_));
 OAI21x1_ASAP7_75t_R _24444_ (.A1(_05315_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_17920_));
 OR2x2_ASAP7_75t_R _24445_ (.A(_05219_),
    .B(_05299_),
    .Y(_17932_));
 AND2x2_ASAP7_75t_R _24446_ (.A(_05243_),
    .B(_05271_),
    .Y(_17936_));
 AND2x2_ASAP7_75t_R _24447_ (.A(_05251_),
    .B(_05263_),
    .Y(_17935_));
 AND2x2_ASAP7_75t_R _24448_ (.A(_05254_),
    .B(_05259_),
    .Y(_17937_));
 NAND2x1_ASAP7_75t_R _24449_ (.A(_05247_),
    .B(_05269_),
    .Y(_17942_));
 NAND2x1_ASAP7_75t_R _24450_ (.A(_05223_),
    .B(_05293_),
    .Y(_17953_));
 NAND2x2_ASAP7_75t_R _24451_ (.A(_05209_),
    .B(_05308_),
    .Y(_17951_));
 INVx1_ASAP7_75t_R _24452_ (.A(_17951_),
    .Y(_18033_));
 OAI21x1_ASAP7_75t_R _24453_ (.A1(_01118_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_17960_));
 OR2x2_ASAP7_75t_R _24454_ (.A(_05227_),
    .B(_05299_),
    .Y(_17972_));
 AND2x2_ASAP7_75t_R _24455_ (.A(_05251_),
    .B(_05271_),
    .Y(_17977_));
 AND2x2_ASAP7_75t_R _24456_ (.A(_05259_),
    .B(_05263_),
    .Y(_17976_));
 AND2x2_ASAP7_75t_R _24457_ (.A(_05254_),
    .B(_05268_),
    .Y(_17978_));
 NAND2x1_ASAP7_75t_R _24458_ (.A(_05247_),
    .B(_05277_),
    .Y(_17982_));
 NAND2x1_ASAP7_75t_R _24459_ (.A(_05223_),
    .B(_05314_),
    .Y(_17993_));
 NAND2x2_ASAP7_75t_R _24460_ (.A(_05216_),
    .B(_05308_),
    .Y(_17992_));
 INVx1_ASAP7_75t_R _24461_ (.A(_17992_),
    .Y(_18034_));
 BUFx6f_ASAP7_75t_R _24462_ (.A(_01151_),
    .Y(_05316_));
 OAI21x1_ASAP7_75t_R _24463_ (.A1(_05316_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_18001_));
 OR2x2_ASAP7_75t_R _24464_ (.A(_05236_),
    .B(_05299_),
    .Y(_18011_));
 NAND2x1_ASAP7_75t_R _24465_ (.A(_05260_),
    .B(_05272_),
    .Y(_18018_));
 NAND2x1_ASAP7_75t_R _24466_ (.A(_05247_),
    .B(_05285_),
    .Y(_18024_));
 AND2x2_ASAP7_75t_R _24467_ (.A(_05223_),
    .B(_05309_),
    .Y(_18035_));
 OAI21x1_ASAP7_75t_R _24468_ (.A1(_01184_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_18046_));
 OR2x2_ASAP7_75t_R _24469_ (.A(_05243_),
    .B(_05299_),
    .Y(_18058_));
 NAND2x1_ASAP7_75t_R _24470_ (.A(_05269_),
    .B(_05272_),
    .Y(_18062_));
 NAND2x1_ASAP7_75t_R _24471_ (.A(_05247_),
    .B(_05293_),
    .Y(_18069_));
 NAND2x2_ASAP7_75t_R _24472_ (.A(_05233_),
    .B(_05308_),
    .Y(_18070_));
 INVx1_ASAP7_75t_R _24473_ (.A(_18070_),
    .Y(_18141_));
 BUFx4f_ASAP7_75t_R _24474_ (.A(_01217_),
    .Y(_05317_));
 OAI21x1_ASAP7_75t_R _24475_ (.A1(_05317_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_18084_));
 OR2x2_ASAP7_75t_R _24476_ (.A(_05251_),
    .B(_05298_),
    .Y(_18095_));
 NAND2x1_ASAP7_75t_R _24477_ (.A(_05272_),
    .B(_05277_),
    .Y(_18100_));
 NAND2x1_ASAP7_75t_R _24478_ (.A(_05247_),
    .B(_05314_),
    .Y(_18106_));
 NAND2x1_ASAP7_75t_R _24479_ (.A(_05240_),
    .B(_05308_),
    .Y(_18107_));
 INVx1_ASAP7_75t_R _24480_ (.A(_18107_),
    .Y(_18142_));
 OAI21x1_ASAP7_75t_R _24481_ (.A1(_01250_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_18118_));
 OR2x2_ASAP7_75t_R _24482_ (.A(_05259_),
    .B(_05298_),
    .Y(_18130_));
 NAND2x1_ASAP7_75t_R _24483_ (.A(_05272_),
    .B(_05285_),
    .Y(_18135_));
 AND2x2_ASAP7_75t_R _24484_ (.A(_05247_),
    .B(_05309_),
    .Y(_18140_));
 BUFx6f_ASAP7_75t_R _24485_ (.A(_01283_),
    .Y(_05318_));
 OAI21x1_ASAP7_75t_R _24486_ (.A1(_05318_),
    .A2(_05153_),
    .B(_05313_),
    .Y(_18151_));
 OR2x2_ASAP7_75t_R _24487_ (.A(_05268_),
    .B(_05298_),
    .Y(_18162_));
 NAND2x1_ASAP7_75t_R _24488_ (.A(_05272_),
    .B(_05293_),
    .Y(_18167_));
 NAND2x2_ASAP7_75t_R _24489_ (.A(_05254_),
    .B(_05308_),
    .Y(_18168_));
 INVx1_ASAP7_75t_R _24490_ (.A(_18168_),
    .Y(_18225_));
 OAI21x1_ASAP7_75t_R _24491_ (.A1(_01316_),
    .A2(_05176_),
    .B(_05313_),
    .Y(_18181_));
 OR2x2_ASAP7_75t_R _24492_ (.A(_05276_),
    .B(_05298_),
    .Y(_18192_));
 NAND2x1_ASAP7_75t_R _24493_ (.A(_05272_),
    .B(_05314_),
    .Y(_18197_));
 NAND2x2_ASAP7_75t_R _24494_ (.A(_05263_),
    .B(_05308_),
    .Y(_18196_));
 INVx1_ASAP7_75t_R _24495_ (.A(_18196_),
    .Y(_18223_));
 BUFx4f_ASAP7_75t_R _24496_ (.A(_01349_),
    .Y(_05319_));
 OAI21x1_ASAP7_75t_R _24497_ (.A1(_05319_),
    .A2(_05176_),
    .B(_05312_),
    .Y(_18209_));
 OR2x2_ASAP7_75t_R _24498_ (.A(_05284_),
    .B(_05298_),
    .Y(_18219_));
 AND2x2_ASAP7_75t_R _24499_ (.A(_05271_),
    .B(_05309_),
    .Y(_18224_));
 OAI21x1_ASAP7_75t_R _24500_ (.A1(_01382_),
    .A2(_05176_),
    .B(_05312_),
    .Y(_18239_));
 OR2x2_ASAP7_75t_R _24501_ (.A(_05292_),
    .B(_05298_),
    .Y(_18250_));
 BUFx4f_ASAP7_75t_R _24502_ (.A(_01415_),
    .Y(_05320_));
 OAI21x1_ASAP7_75t_R _24503_ (.A1(_05320_),
    .A2(_05176_),
    .B(_05312_),
    .Y(_18266_));
 OR2x2_ASAP7_75t_R _24504_ (.A(_05298_),
    .B(_05303_),
    .Y(_18277_));
 OAI21x1_ASAP7_75t_R _24505_ (.A1(_04868_),
    .A2(_05176_),
    .B(_05312_),
    .Y(_18291_));
 OR2x2_ASAP7_75t_R _24506_ (.A(_05298_),
    .B(_05309_),
    .Y(_18301_));
 OAI21x1_ASAP7_75t_R _24507_ (.A1(_01747_),
    .A2(_05176_),
    .B(_05312_),
    .Y(_18308_));
 INVx3_ASAP7_75t_R _24508_ (.A(_18260_),
    .Y(_18255_));
 INVx1_ASAP7_75t_R _24509_ (.A(_18286_),
    .Y(_18285_));
 AO32x2_ASAP7_75t_R _24510_ (.A1(_13593_),
    .A2(_13394_),
    .A3(_13635_),
    .B1(_13655_),
    .B2(_13391_),
    .Y(_05321_));
 AND5x2_ASAP7_75t_R _24511_ (.A(_14022_),
    .B(_14034_),
    .C(_14068_),
    .D(_04926_),
    .E(_05321_),
    .Y(_05322_));
 INVx1_ASAP7_75t_R _24512_ (.A(_14026_),
    .Y(_05323_));
 AND4x1_ASAP7_75t_R _24513_ (.A(_04930_),
    .B(_13568_),
    .C(_05323_),
    .D(_04938_),
    .Y(_05324_));
 AND3x4_ASAP7_75t_R _24514_ (.A(_01778_),
    .B(_02219_),
    .C(_02221_),
    .Y(_05325_));
 INVx1_ASAP7_75t_R _24515_ (.A(_05325_),
    .Y(_05326_));
 AOI211x1_ASAP7_75t_R _24516_ (.A1(_14065_),
    .A2(_14062_),
    .B(_05065_),
    .C(_14057_),
    .Y(_05327_));
 BUFx4f_ASAP7_75t_R _24517_ (.A(_00791_),
    .Y(_05328_));
 OR2x4_ASAP7_75t_R _24518_ (.A(_01456_),
    .B(_04930_),
    .Y(_05329_));
 NAND3x1_ASAP7_75t_R _24519_ (.A(_05328_),
    .B(_05081_),
    .C(_05329_),
    .Y(_05330_));
 NAND2x1_ASAP7_75t_R _24520_ (.A(_05068_),
    .B(_14812_),
    .Y(_05331_));
 OR3x1_ASAP7_75t_R _24521_ (.A(_00790_),
    .B(_05068_),
    .C(_14812_),
    .Y(_05332_));
 OA211x2_ASAP7_75t_R _24522_ (.A1(_00783_),
    .A2(_05331_),
    .B(_05332_),
    .C(_01455_),
    .Y(_05333_));
 OR2x2_ASAP7_75t_R _24523_ (.A(_13492_),
    .B(_05325_),
    .Y(_05334_));
 OR5x2_ASAP7_75t_R _24524_ (.A(_14065_),
    .B(_05065_),
    .C(_05330_),
    .D(_05333_),
    .E(_05334_),
    .Y(_05335_));
 OA211x2_ASAP7_75t_R _24525_ (.A1(_05326_),
    .A2(_05327_),
    .B(_05335_),
    .C(_05077_),
    .Y(_05336_));
 NOR2x2_ASAP7_75t_R _24526_ (.A(_05061_),
    .B(_04930_),
    .Y(_05337_));
 OR3x1_ASAP7_75t_R _24527_ (.A(_01777_),
    .B(_04931_),
    .C(_05337_),
    .Y(_05338_));
 AO21x1_ASAP7_75t_R _24528_ (.A1(_05075_),
    .A2(_05338_),
    .B(_04933_),
    .Y(_05339_));
 INVx4_ASAP7_75t_R _24529_ (.A(_04931_),
    .Y(_05340_));
 NAND2x1_ASAP7_75t_R _24530_ (.A(_04934_),
    .B(_05340_),
    .Y(_05341_));
 AOI21x1_ASAP7_75t_R _24531_ (.A1(_05339_),
    .A2(_05341_),
    .B(_04936_),
    .Y(_05342_));
 INVx1_ASAP7_75t_R _24532_ (.A(_01931_),
    .Y(_05343_));
 INVx1_ASAP7_75t_R _24533_ (.A(_01932_),
    .Y(_05344_));
 AO22x1_ASAP7_75t_R _24534_ (.A1(net191),
    .A2(_05343_),
    .B1(_05344_),
    .B2(net190),
    .Y(_05345_));
 INVx2_ASAP7_75t_R _24535_ (.A(_01933_),
    .Y(_05346_));
 INVx1_ASAP7_75t_R _24536_ (.A(_01934_),
    .Y(_05347_));
 AO22x1_ASAP7_75t_R _24537_ (.A1(net189),
    .A2(_05346_),
    .B1(_05347_),
    .B2(net188),
    .Y(_05348_));
 INVx1_ASAP7_75t_R _24538_ (.A(_01935_),
    .Y(_05349_));
 INVx1_ASAP7_75t_R _24539_ (.A(_01936_),
    .Y(_05350_));
 AO22x1_ASAP7_75t_R _24540_ (.A1(net187),
    .A2(_05349_),
    .B1(_05350_),
    .B2(net186),
    .Y(_05351_));
 INVx1_ASAP7_75t_R _24541_ (.A(_01937_),
    .Y(_05352_));
 INVx1_ASAP7_75t_R _24542_ (.A(_01946_),
    .Y(_05353_));
 AO22x1_ASAP7_75t_R _24543_ (.A1(net185),
    .A2(_05352_),
    .B1(_05353_),
    .B2(net179),
    .Y(_05354_));
 OR4x2_ASAP7_75t_R _24544_ (.A(_05345_),
    .B(_05348_),
    .C(_05351_),
    .D(_05354_),
    .Y(_05355_));
 INVx1_ASAP7_75t_R _24545_ (.A(_01941_),
    .Y(_05356_));
 AND2x2_ASAP7_75t_R _24546_ (.A(net184),
    .B(_05356_),
    .Y(_05357_));
 INVx1_ASAP7_75t_R _24547_ (.A(_01942_),
    .Y(_05358_));
 INVx1_ASAP7_75t_R _24548_ (.A(_01943_),
    .Y(_05359_));
 AO22x1_ASAP7_75t_R _24549_ (.A1(net183),
    .A2(_05358_),
    .B1(_05359_),
    .B2(net182),
    .Y(_05360_));
 INVx1_ASAP7_75t_R _24550_ (.A(_01944_),
    .Y(_05361_));
 INVx1_ASAP7_75t_R _24551_ (.A(_01945_),
    .Y(_05362_));
 AO22x1_ASAP7_75t_R _24552_ (.A1(net181),
    .A2(_05361_),
    .B1(_05362_),
    .B2(net180),
    .Y(_05363_));
 INVx1_ASAP7_75t_R _24553_ (.A(_01929_),
    .Y(_05364_));
 INVx1_ASAP7_75t_R _24554_ (.A(_01930_),
    .Y(_05365_));
 AO22x1_ASAP7_75t_R _24555_ (.A1(net193),
    .A2(_05364_),
    .B1(_05365_),
    .B2(net192),
    .Y(_05366_));
 OR4x2_ASAP7_75t_R _24556_ (.A(_05357_),
    .B(_05360_),
    .C(_05363_),
    .D(_05366_),
    .Y(_05367_));
 INVx1_ASAP7_75t_R _24557_ (.A(net195),
    .Y(_05368_));
 INVx1_ASAP7_75t_R _24558_ (.A(net178),
    .Y(_05369_));
 OAI22x1_ASAP7_75t_R _24559_ (.A1(_05368_),
    .A2(_01938_),
    .B1(_01940_),
    .B2(_05369_),
    .Y(_05370_));
 INVx1_ASAP7_75t_R _24560_ (.A(_01939_),
    .Y(_05371_));
 AO21x1_ASAP7_75t_R _24561_ (.A1(net196),
    .A2(_05371_),
    .B(net194),
    .Y(_05372_));
 OR2x2_ASAP7_75t_R _24562_ (.A(_05370_),
    .B(_05372_),
    .Y(_05373_));
 AND2x4_ASAP7_75t_R _24563_ (.A(_04932_),
    .B(_05075_),
    .Y(_05374_));
 INVx1_ASAP7_75t_R _24564_ (.A(_01850_),
    .Y(_05375_));
 OA211x2_ASAP7_75t_R _24565_ (.A1(net194),
    .A2(_05375_),
    .B(_02220_),
    .C(_01455_),
    .Y(_05376_));
 AND4x2_ASAP7_75t_R _24566_ (.A(_04936_),
    .B(_05340_),
    .C(_05374_),
    .D(_05376_),
    .Y(_05377_));
 OA31x2_ASAP7_75t_R _24567_ (.A1(_05355_),
    .A2(_05367_),
    .A3(_05373_),
    .B1(_05377_),
    .Y(_05378_));
 INVx2_ASAP7_75t_R _24568_ (.A(_01460_),
    .Y(_05379_));
 AND2x4_ASAP7_75t_R _24569_ (.A(_01780_),
    .B(_04935_),
    .Y(_05380_));
 AND2x2_ASAP7_75t_R _24570_ (.A(_04933_),
    .B(_05380_),
    .Y(_05381_));
 OA211x2_ASAP7_75t_R _24571_ (.A1(net105),
    .A2(_05379_),
    .B(_04931_),
    .C(_05381_),
    .Y(_05382_));
 BUFx4f_ASAP7_75t_R _24572_ (.A(_05382_),
    .Y(_05383_));
 OR4x1_ASAP7_75t_R _24573_ (.A(_05336_),
    .B(_05342_),
    .C(_05378_),
    .D(_05383_),
    .Y(_05384_));
 AO21x2_ASAP7_75t_R _24574_ (.A1(_05322_),
    .A2(_05324_),
    .B(_05384_),
    .Y(_05385_));
 BUFx6f_ASAP7_75t_R _24575_ (.A(_05385_),
    .Y(_05386_));
 BUFx6f_ASAP7_75t_R _24576_ (.A(_05386_),
    .Y(_05387_));
 BUFx6f_ASAP7_75t_R _24577_ (.A(_05387_),
    .Y(_05388_));
 BUFx6f_ASAP7_75t_R _24578_ (.A(_05388_),
    .Y(_05389_));
 BUFx4f_ASAP7_75t_R _24579_ (.A(_05389_),
    .Y(_05390_));
 NAND2x1_ASAP7_75t_R _24580_ (.A(net184),
    .B(_05356_),
    .Y(_05391_));
 NAND2x1_ASAP7_75t_R _24581_ (.A(net182),
    .B(_05359_),
    .Y(_05392_));
 NAND2x1_ASAP7_75t_R _24582_ (.A(net180),
    .B(_05362_),
    .Y(_05393_));
 NAND2x1_ASAP7_75t_R _24583_ (.A(net192),
    .B(_05365_),
    .Y(_05394_));
 NAND2x1_ASAP7_75t_R _24584_ (.A(net190),
    .B(_05344_),
    .Y(_05395_));
 INVx1_ASAP7_75t_R _24585_ (.A(net188),
    .Y(_05396_));
 NAND2x1_ASAP7_75t_R _24586_ (.A(net186),
    .B(_05350_),
    .Y(_05397_));
 AO32x1_ASAP7_75t_R _24587_ (.A1(net185),
    .A2(_05352_),
    .A3(_05397_),
    .B1(net187),
    .B2(_05349_),
    .Y(_05398_));
 OA21x2_ASAP7_75t_R _24588_ (.A1(_05396_),
    .A2(_01934_),
    .B(_05398_),
    .Y(_05399_));
 AO21x1_ASAP7_75t_R _24589_ (.A1(net189),
    .A2(_05346_),
    .B(_05399_),
    .Y(_05400_));
 AO22x1_ASAP7_75t_R _24590_ (.A1(net191),
    .A2(_05343_),
    .B1(_05395_),
    .B2(_05400_),
    .Y(_05401_));
 AO22x1_ASAP7_75t_R _24591_ (.A1(net193),
    .A2(_05364_),
    .B1(_05394_),
    .B2(_05401_),
    .Y(_05402_));
 AO22x1_ASAP7_75t_R _24592_ (.A1(net181),
    .A2(_05361_),
    .B1(_05393_),
    .B2(_05402_),
    .Y(_05403_));
 AO22x1_ASAP7_75t_R _24593_ (.A1(net183),
    .A2(_05358_),
    .B1(_05392_),
    .B2(_05403_),
    .Y(_05404_));
 NOR2x1_ASAP7_75t_R _24594_ (.A(_05355_),
    .B(_05367_),
    .Y(_05405_));
 AO221x1_ASAP7_75t_R _24595_ (.A1(net194),
    .A2(_02220_),
    .B1(_05391_),
    .B2(_05404_),
    .C(_05405_),
    .Y(_05406_));
 AND2x2_ASAP7_75t_R _24596_ (.A(_05378_),
    .B(_05406_),
    .Y(_05407_));
 OR3x4_ASAP7_75t_R _24597_ (.A(_14057_),
    .B(_14065_),
    .C(_05065_),
    .Y(_05408_));
 NAND2x2_ASAP7_75t_R _24598_ (.A(_05077_),
    .B(_05325_),
    .Y(_05409_));
 OR2x4_ASAP7_75t_R _24599_ (.A(_05408_),
    .B(_05409_),
    .Y(_05410_));
 BUFx4f_ASAP7_75t_R _24600_ (.A(_05410_),
    .Y(_05411_));
 BUFx6f_ASAP7_75t_R _24601_ (.A(_05411_),
    .Y(_05412_));
 BUFx6f_ASAP7_75t_R _24602_ (.A(_05412_),
    .Y(_05413_));
 OR2x2_ASAP7_75t_R _24603_ (.A(_05066_),
    .B(_05409_),
    .Y(_05414_));
 BUFx4f_ASAP7_75t_R _24604_ (.A(_05414_),
    .Y(_05415_));
 BUFx4f_ASAP7_75t_R _24605_ (.A(_05415_),
    .Y(_05416_));
 BUFx4f_ASAP7_75t_R _24606_ (.A(_05416_),
    .Y(_05417_));
 BUFx6f_ASAP7_75t_R _24607_ (.A(_05417_),
    .Y(_05418_));
 OAI22x1_ASAP7_75t_R _24608_ (.A1(_01956_),
    .A2(_05413_),
    .B1(_05418_),
    .B2(_02054_),
    .Y(_05419_));
 NOR2x1_ASAP7_75t_R _24609_ (.A(_05407_),
    .B(_05419_),
    .Y(_05420_));
 BUFx4f_ASAP7_75t_R _24610_ (.A(_04931_),
    .Y(_05421_));
 OR2x6_ASAP7_75t_R _24611_ (.A(_05421_),
    .B(_04937_),
    .Y(_05422_));
 BUFx6f_ASAP7_75t_R _24612_ (.A(_05422_),
    .Y(_05423_));
 OR2x2_ASAP7_75t_R _24613_ (.A(_05423_),
    .B(_05126_),
    .Y(_05424_));
 AOI21x1_ASAP7_75t_R _24614_ (.A1(_05322_),
    .A2(_05324_),
    .B(_05384_),
    .Y(_05425_));
 INVx1_ASAP7_75t_R _24615_ (.A(_05374_),
    .Y(_05426_));
 OA31x2_ASAP7_75t_R _24616_ (.A1(_14057_),
    .A2(_14065_),
    .A3(_05065_),
    .B1(_05325_),
    .Y(_05427_));
 OA21x2_ASAP7_75t_R _24617_ (.A1(_04935_),
    .A2(_05427_),
    .B(_04931_),
    .Y(_05428_));
 AO21x1_ASAP7_75t_R _24618_ (.A1(_05066_),
    .A2(_05408_),
    .B(_05409_),
    .Y(_05429_));
 NAND2x2_ASAP7_75t_R _24619_ (.A(_04933_),
    .B(_05380_),
    .Y(_05430_));
 OA211x2_ASAP7_75t_R _24620_ (.A1(_05426_),
    .A2(_05428_),
    .B(_05429_),
    .C(_05430_),
    .Y(_05431_));
 BUFx4f_ASAP7_75t_R _24621_ (.A(_05431_),
    .Y(_05432_));
 OR2x4_ASAP7_75t_R _24622_ (.A(_05425_),
    .B(_05432_),
    .Y(_05433_));
 AO21x2_ASAP7_75t_R _24623_ (.A1(_05420_),
    .A2(_05424_),
    .B(_05433_),
    .Y(_05434_));
 OA21x2_ASAP7_75t_R _24624_ (.A1(_01722_),
    .A2(_05390_),
    .B(_05434_),
    .Y(_05435_));
 INVx1_ASAP7_75t_R _24625_ (.A(_05435_),
    .Y(_18774_));
 OR3x1_ASAP7_75t_R _24626_ (.A(_04933_),
    .B(_04934_),
    .C(_04935_),
    .Y(_05436_));
 OR3x4_ASAP7_75t_R _24627_ (.A(_05355_),
    .B(_05367_),
    .C(_05373_),
    .Y(_05437_));
 NAND2x2_ASAP7_75t_R _24628_ (.A(_05377_),
    .B(_05437_),
    .Y(_05438_));
 INVx1_ASAP7_75t_R _24629_ (.A(_05360_),
    .Y(_05439_));
 INVx1_ASAP7_75t_R _24630_ (.A(net193),
    .Y(_05440_));
 OA21x2_ASAP7_75t_R _24631_ (.A1(_05440_),
    .A2(_01929_),
    .B(_05394_),
    .Y(_05441_));
 AOI22x1_ASAP7_75t_R _24632_ (.A1(net189),
    .A2(_05346_),
    .B1(_05347_),
    .B2(net188),
    .Y(_05442_));
 AO21x1_ASAP7_75t_R _24633_ (.A1(_05442_),
    .A2(_05351_),
    .B(_05345_),
    .Y(_05443_));
 AO21x1_ASAP7_75t_R _24634_ (.A1(_05441_),
    .A2(_05443_),
    .B(_05363_),
    .Y(_05444_));
 NAND2x1_ASAP7_75t_R _24635_ (.A(net194),
    .B(_02220_),
    .Y(_05445_));
 AND2x2_ASAP7_75t_R _24636_ (.A(_05391_),
    .B(_05445_),
    .Y(_05446_));
 OAI21x1_ASAP7_75t_R _24637_ (.A1(_05355_),
    .A2(_05367_),
    .B(_05446_),
    .Y(_05447_));
 AOI21x1_ASAP7_75t_R _24638_ (.A1(_05439_),
    .A2(_05444_),
    .B(_05447_),
    .Y(_05448_));
 AO31x2_ASAP7_75t_R _24639_ (.A1(_13774_),
    .A2(_05080_),
    .A3(_05082_),
    .B(_05079_),
    .Y(_05449_));
 AO21x1_ASAP7_75t_R _24640_ (.A1(_13407_),
    .A2(_05449_),
    .B(_02221_),
    .Y(_05450_));
 OR3x1_ASAP7_75t_R _24641_ (.A(net10),
    .B(_05068_),
    .C(_14812_),
    .Y(_05451_));
 NAND2x1_ASAP7_75t_R _24642_ (.A(net10),
    .B(_05333_),
    .Y(_05452_));
 OR3x4_ASAP7_75t_R _24643_ (.A(_14065_),
    .B(_05065_),
    .C(_05330_),
    .Y(_05453_));
 AO21x1_ASAP7_75t_R _24644_ (.A1(_05451_),
    .A2(_05452_),
    .B(_05453_),
    .Y(_05454_));
 AND2x4_ASAP7_75t_R _24645_ (.A(_05077_),
    .B(_05326_),
    .Y(_05455_));
 NAND2x1_ASAP7_75t_R _24646_ (.A(_05329_),
    .B(_05455_),
    .Y(_05456_));
 AO31x2_ASAP7_75t_R _24647_ (.A1(_05328_),
    .A2(_05450_),
    .A3(_05454_),
    .B(_05456_),
    .Y(_05457_));
 OA211x2_ASAP7_75t_R _24648_ (.A1(_05438_),
    .A2(_05448_),
    .B(_05457_),
    .C(_05430_),
    .Y(_05458_));
 OR4x1_ASAP7_75t_R _24649_ (.A(_04945_),
    .B(_05340_),
    .C(_05325_),
    .D(_05381_),
    .Y(_05459_));
 OA21x2_ASAP7_75t_R _24650_ (.A1(_05421_),
    .A2(_05458_),
    .B(_05459_),
    .Y(_05460_));
 INVx2_ASAP7_75t_R _24651_ (.A(\alu_adder_result_ex[3] ),
    .Y(_05461_));
 OA222x2_ASAP7_75t_R _24652_ (.A1(_05422_),
    .A2(_05461_),
    .B1(_05412_),
    .B2(_01953_),
    .C1(_01461_),
    .C2(_05416_),
    .Y(_05462_));
 OA21x2_ASAP7_75t_R _24653_ (.A1(_05436_),
    .A2(_05460_),
    .B(_05462_),
    .Y(_05463_));
 OA22x2_ASAP7_75t_R _24654_ (.A1(_01719_),
    .A2(_05386_),
    .B1(_05433_),
    .B2(_05463_),
    .Y(_05464_));
 INVx1_ASAP7_75t_R _24655_ (.A(_05464_),
    .Y(_18776_));
 BUFx4f_ASAP7_75t_R _24656_ (.A(_05425_),
    .Y(_05465_));
 BUFx6f_ASAP7_75t_R _24657_ (.A(_05465_),
    .Y(_05466_));
 BUFx6f_ASAP7_75t_R _24658_ (.A(_05466_),
    .Y(_05467_));
 BUFx4f_ASAP7_75t_R _24659_ (.A(_05467_),
    .Y(_05468_));
 BUFx6f_ASAP7_75t_R _24660_ (.A(_00288_),
    .Y(_05469_));
 BUFx4f_ASAP7_75t_R _24661_ (.A(_05469_),
    .Y(_05470_));
 AOI21x1_ASAP7_75t_R _24662_ (.A1(_01743_),
    .A2(_05468_),
    .B(_05470_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 BUFx4f_ASAP7_75t_R _24663_ (.A(_00365_),
    .Y(_05471_));
 INVx4_ASAP7_75t_R _24664_ (.A(_05471_),
    .Y(_05472_));
 BUFx4f_ASAP7_75t_R _24665_ (.A(_00291_),
    .Y(_05473_));
 AND2x2_ASAP7_75t_R _24666_ (.A(_05473_),
    .B(net149),
    .Y(_05474_));
 NOR2x1_ASAP7_75t_R _24667_ (.A(_05473_),
    .B(_01672_),
    .Y(_05475_));
 INVx1_ASAP7_75t_R _24668_ (.A(_01673_),
    .Y(_05476_));
 AOI22x1_ASAP7_75t_R _24669_ (.A1(net150),
    .A2(_05474_),
    .B1(_05475_),
    .B2(_05476_),
    .Y(_05477_));
 INVx1_ASAP7_75t_R _24670_ (.A(_05473_),
    .Y(_05478_));
 INVx2_ASAP7_75t_R _24671_ (.A(net139),
    .Y(_05479_));
 AND2x2_ASAP7_75t_R _24672_ (.A(_05473_),
    .B(_05479_),
    .Y(_05480_));
 AO21x1_ASAP7_75t_R _24673_ (.A1(_05478_),
    .A2(_01712_),
    .B(_05480_),
    .Y(_05481_));
 AND2x2_ASAP7_75t_R _24674_ (.A(_05477_),
    .B(_05481_),
    .Y(_05482_));
 NAND2x2_ASAP7_75t_R _24675_ (.A(_05472_),
    .B(_05482_),
    .Y(_18319_));
 BUFx4f_ASAP7_75t_R _24676_ (.A(_05472_),
    .Y(_05483_));
 BUFx4f_ASAP7_75t_R _24677_ (.A(_05483_),
    .Y(_05484_));
 BUFx4f_ASAP7_75t_R _24678_ (.A(_05473_),
    .Y(_05485_));
 BUFx4f_ASAP7_75t_R _24679_ (.A(_05485_),
    .Y(_05486_));
 BUFx6f_ASAP7_75t_R _24680_ (.A(_05486_),
    .Y(_05487_));
 AND3x1_ASAP7_75t_R _24681_ (.A(_05487_),
    .B(net141),
    .C(net156),
    .Y(_05488_));
 BUFx3_ASAP7_75t_R _24682_ (.A(_05478_),
    .Y(_05489_));
 BUFx3_ASAP7_75t_R _24683_ (.A(_05489_),
    .Y(_05490_));
 OA211x2_ASAP7_75t_R _24684_ (.A1(_01669_),
    .A2(_01680_),
    .B(_01712_),
    .C(_05490_),
    .Y(_05491_));
 NOR2x1_ASAP7_75t_R _24685_ (.A(_05480_),
    .B(_05491_),
    .Y(_05492_));
 OR3x4_ASAP7_75t_R _24686_ (.A(_05484_),
    .B(_05488_),
    .C(_05492_),
    .Y(_05493_));
 AND2x2_ASAP7_75t_R _24687_ (.A(_18319_),
    .B(_05493_),
    .Y(_18606_));
 INVx1_ASAP7_75t_R _24688_ (.A(_18606_),
    .Y(_18318_));
 INVx2_ASAP7_75t_R _24689_ (.A(_18614_),
    .Y(_18607_));
 INVx1_ASAP7_75t_R _24690_ (.A(net198),
    .Y(_05494_));
 INVx1_ASAP7_75t_R _24691_ (.A(net105),
    .Y(_05495_));
 NAND2x1_ASAP7_75t_R _24692_ (.A(_05495_),
    .B(_02209_),
    .Y(_05496_));
 INVx1_ASAP7_75t_R _24693_ (.A(_01815_),
    .Y(_05497_));
 OAI21x1_ASAP7_75t_R _24694_ (.A1(_05437_),
    .A2(_05496_),
    .B(_05497_),
    .Y(net199));
 NAND2x1_ASAP7_75t_R _24695_ (.A(_05494_),
    .B(net199),
    .Y(_00006_));
 INVx1_ASAP7_75t_R _24696_ (.A(_02290_),
    .Y(_18775_));
 INVx1_ASAP7_75t_R _24697_ (.A(_18317_),
    .Y(\cs_registers_i.pc_if_i[2] ));
 BUFx6f_ASAP7_75t_R _24698_ (.A(_05168_),
    .Y(_05498_));
 NAND2x1_ASAP7_75t_R _24699_ (.A(_05498_),
    .B(_05192_),
    .Y(_17347_));
 OA22x2_ASAP7_75t_R _24700_ (.A1(_00792_),
    .A2(_05176_),
    .B1(_05179_),
    .B2(_01019_),
    .Y(_17350_));
 BUFx3_ASAP7_75t_R _24701_ (.A(_05152_),
    .Y(_05499_));
 OA22x2_ASAP7_75t_R _24702_ (.A1(_00798_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_05315_),
    .Y(_17360_));
 NAND2x1_ASAP7_75t_R _24703_ (.A(_05498_),
    .B(_05228_),
    .Y(_17392_));
 OA22x2_ASAP7_75t_R _24704_ (.A1(_00807_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_01184_),
    .Y(_17413_));
 BUFx6f_ASAP7_75t_R _24705_ (.A(_05216_),
    .Y(_05500_));
 NAND2x1_ASAP7_75t_R _24706_ (.A(_05200_),
    .B(_05500_),
    .Y(_17425_));
 BUFx6f_ASAP7_75t_R _24707_ (.A(_05209_),
    .Y(_05501_));
 NAND2x1_ASAP7_75t_R _24708_ (.A(_05501_),
    .B(_05213_),
    .Y(_17448_));
 NAND2x1_ASAP7_75t_R _24709_ (.A(_05498_),
    .B(_05252_),
    .Y(_17457_));
 BUFx6f_ASAP7_75t_R _24710_ (.A(_05233_),
    .Y(_05502_));
 NAND2x1_ASAP7_75t_R _24711_ (.A(_05200_),
    .B(_05502_),
    .Y(_17475_));
 NAND2x1_ASAP7_75t_R _24712_ (.A(_05501_),
    .B(_05220_),
    .Y(_17478_));
 NAND2x1_ASAP7_75t_R _24713_ (.A(_05498_),
    .B(_05260_),
    .Y(_17488_));
 NAND2x1_ASAP7_75t_R _24714_ (.A(_05207_),
    .B(_05502_),
    .Y(_17503_));
 NAND2x1_ASAP7_75t_R _24715_ (.A(_05501_),
    .B(_05228_),
    .Y(_17506_));
 NAND2x1_ASAP7_75t_R _24716_ (.A(_05498_),
    .B(_05269_),
    .Y(_17518_));
 BUFx6f_ASAP7_75t_R _24717_ (.A(_05240_),
    .Y(_05503_));
 NAND2x1_ASAP7_75t_R _24718_ (.A(_05207_),
    .B(_05503_),
    .Y(_17533_));
 NAND2x1_ASAP7_75t_R _24719_ (.A(_05501_),
    .B(_05237_),
    .Y(_17537_));
 NAND2x1_ASAP7_75t_R _24720_ (.A(_05220_),
    .B(_05502_),
    .Y(_17570_));
 NAND2x1_ASAP7_75t_R _24721_ (.A(_05200_),
    .B(_05264_),
    .Y(_17608_));
 NAND2x1_ASAP7_75t_R _24722_ (.A(_05228_),
    .B(_05503_),
    .Y(_17652_));
 NAND2x1_ASAP7_75t_R _24723_ (.A(_05500_),
    .B(_05252_),
    .Y(_17662_));
 BUFx6f_ASAP7_75t_R _24724_ (.A(_05280_),
    .Y(_05504_));
 NAND2x1_ASAP7_75t_R _24725_ (.A(_05200_),
    .B(_05504_),
    .Y(_17690_));
 NAND2x1_ASAP7_75t_R _24726_ (.A(_05237_),
    .B(_05503_),
    .Y(_17701_));
 NAND2x1_ASAP7_75t_R _24727_ (.A(_05501_),
    .B(_05269_),
    .Y(_17710_));
 NAND2x1_ASAP7_75t_R _24728_ (.A(_05503_),
    .B(_05244_),
    .Y(_17754_));
 BUFx6f_ASAP7_75t_R _24729_ (.A(_05288_),
    .Y(_05505_));
 NAND2x1_ASAP7_75t_R _24730_ (.A(_05207_),
    .B(_05505_),
    .Y(_17792_));
 NAND2x1_ASAP7_75t_R _24731_ (.A(_05500_),
    .B(_05277_),
    .Y(_17813_));
 NAND2x1_ASAP7_75t_R _24732_ (.A(_05213_),
    .B(_05505_),
    .Y(_17837_));
 NAND2x1_ASAP7_75t_R _24733_ (.A(_05500_),
    .B(_05285_),
    .Y(_17858_));
 NAND2x1_ASAP7_75t_R _24734_ (.A(_05503_),
    .B(_05269_),
    .Y(_17895_));
 NAND2x1_ASAP7_75t_R _24735_ (.A(_05237_),
    .B(_05504_),
    .Y(_17930_));
 NAND2x1_ASAP7_75t_R _24736_ (.A(_05503_),
    .B(_05277_),
    .Y(_17941_));
 NAND2x1_ASAP7_75t_R _24737_ (.A(_05237_),
    .B(_05505_),
    .Y(_17971_));
 NAND2x1_ASAP7_75t_R _24738_ (.A(_05255_),
    .B(_05277_),
    .Y(_18016_));
 NAND2x1_ASAP7_75t_R _24739_ (.A(_05240_),
    .B(_05293_),
    .Y(_18023_));
 NAND2x1_ASAP7_75t_R _24740_ (.A(_05260_),
    .B(_05504_),
    .Y(_18056_));
 NAND2x1_ASAP7_75t_R _24741_ (.A(_05264_),
    .B(_05277_),
    .Y(_18061_));
 NAND2x1_ASAP7_75t_R _24742_ (.A(_05240_),
    .B(_05314_),
    .Y(_18068_));
 NAND2x1_ASAP7_75t_R _24743_ (.A(_05259_),
    .B(_05505_),
    .Y(_18094_));
 NAND2x1_ASAP7_75t_R _24744_ (.A(_05264_),
    .B(_05285_),
    .Y(_18099_));
 NAND2x2_ASAP7_75t_R _24745_ (.A(_05276_),
    .B(_05504_),
    .Y(_18128_));
 NAND2x1_ASAP7_75t_R _24746_ (.A(_05255_),
    .B(_05314_),
    .Y(_18133_));
 NAND2x1_ASAP7_75t_R _24747_ (.A(_05276_),
    .B(_05505_),
    .Y(_18161_));
 NAND2x1_ASAP7_75t_R _24748_ (.A(_05264_),
    .B(_05314_),
    .Y(_18166_));
 NAND2x1_ASAP7_75t_R _24749_ (.A(_05284_),
    .B(_05505_),
    .Y(_18191_));
 NAND2x1_ASAP7_75t_R _24750_ (.A(_05288_),
    .B(_05314_),
    .Y(_18249_));
 NAND2x2_ASAP7_75t_R _24751_ (.A(_05288_),
    .B(_05309_),
    .Y(_18276_));
 OA22x2_ASAP7_75t_R _24752_ (.A1(_00414_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_00986_),
    .Y(_17348_));
 NAND2x1_ASAP7_75t_R _24753_ (.A(_05498_),
    .B(_05207_),
    .Y(_17354_));
 NAND2x1_ASAP7_75t_R _24754_ (.A(_05498_),
    .B(_05220_),
    .Y(_17377_));
 OA22x2_ASAP7_75t_R _24755_ (.A1(_00804_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_05316_),
    .Y(_17393_));
 NAND2x1_ASAP7_75t_R _24756_ (.A(_05200_),
    .B(_05501_),
    .Y(_17402_));
 NAND2x1_ASAP7_75t_R _24757_ (.A(_05498_),
    .B(_05244_),
    .Y(_17435_));
 NAND2x1_ASAP7_75t_R _24758_ (.A(_05207_),
    .B(_05500_),
    .Y(_17449_));
 OA22x2_ASAP7_75t_R _24759_ (.A1(_00812_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_01250_),
    .Y(_17458_));
 NAND2x1_ASAP7_75t_R _24760_ (.A(_05192_),
    .B(_05503_),
    .Y(_17476_));
 NAND2x1_ASAP7_75t_R _24761_ (.A(_05213_),
    .B(_05500_),
    .Y(_17479_));
 OA22x2_ASAP7_75t_R _24762_ (.A1(_00815_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_05318_),
    .Y(_17489_));
 NAND2x1_ASAP7_75t_R _24763_ (.A(_05200_),
    .B(_05503_),
    .Y(_17504_));
 NAND2x1_ASAP7_75t_R _24764_ (.A(_05500_),
    .B(_05220_),
    .Y(_17507_));
 BUFx4f_ASAP7_75t_R _24765_ (.A(_00818_),
    .Y(_05506_));
 OA22x2_ASAP7_75t_R _24766_ (.A1(_05506_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_01316_),
    .Y(_17519_));
 NAND2x1_ASAP7_75t_R _24767_ (.A(_05500_),
    .B(_05228_),
    .Y(_17538_));
 NAND2x1_ASAP7_75t_R _24768_ (.A(_05498_),
    .B(_05277_),
    .Y(_17554_));
 NAND2x1_ASAP7_75t_R _24769_ (.A(_05213_),
    .B(_05503_),
    .Y(_17571_));
 NAND2x1_ASAP7_75t_R _24770_ (.A(_05501_),
    .B(_05244_),
    .Y(_17578_));
 NAND2x1_ASAP7_75t_R _24771_ (.A(_05498_),
    .B(_05285_),
    .Y(_17593_));
 NAND2x1_ASAP7_75t_R _24772_ (.A(_05228_),
    .B(_05502_),
    .Y(_17613_));
 NAND2x1_ASAP7_75t_R _24773_ (.A(_05501_),
    .B(_05252_),
    .Y(_17620_));
 NAND2x1_ASAP7_75t_R _24774_ (.A(_05168_),
    .B(_05293_),
    .Y(_17634_));
 NAND2x1_ASAP7_75t_R _24775_ (.A(_05168_),
    .B(_05314_),
    .Y(_17676_));
 NAND2x1_ASAP7_75t_R _24776_ (.A(_05192_),
    .B(_05505_),
    .Y(_17691_));
 NAND2x1_ASAP7_75t_R _24777_ (.A(_05500_),
    .B(_05260_),
    .Y(_17711_));
 NAND2x1_ASAP7_75t_R _24778_ (.A(_05207_),
    .B(_05504_),
    .Y(_17744_));
 NAND2x1_ASAP7_75t_R _24779_ (.A(_05501_),
    .B(_05277_),
    .Y(_17766_));
 NAND2x1_ASAP7_75t_R _24780_ (.A(_05502_),
    .B(_05260_),
    .Y(_17804_));
 NAND2x1_ASAP7_75t_R _24781_ (.A(_05502_),
    .B(_05269_),
    .Y(_17849_));
 NAND2x1_ASAP7_75t_R _24782_ (.A(_05228_),
    .B(_05504_),
    .Y(_17885_));
 NAND2x1_ASAP7_75t_R _24783_ (.A(_05209_),
    .B(_05314_),
    .Y(_17906_));
 NAND2x1_ASAP7_75t_R _24784_ (.A(_05228_),
    .B(_05505_),
    .Y(_17931_));
 NAND2x1_ASAP7_75t_R _24785_ (.A(_05216_),
    .B(_05303_),
    .Y(_17952_));
 NAND2x1_ASAP7_75t_R _24786_ (.A(_05502_),
    .B(_05293_),
    .Y(_17983_));
 NAND2x1_ASAP7_75t_R _24787_ (.A(_05252_),
    .B(_05504_),
    .Y(_18012_));
 NAND2x1_ASAP7_75t_R _24788_ (.A(_05264_),
    .B(_05269_),
    .Y(_18017_));
 NAND2x1_ASAP7_75t_R _24789_ (.A(_05252_),
    .B(_05505_),
    .Y(_18057_));
 NAND2x1_ASAP7_75t_R _24790_ (.A(_05268_),
    .B(_05505_),
    .Y(_18129_));
 NAND2x1_ASAP7_75t_R _24791_ (.A(_05264_),
    .B(_05293_),
    .Y(_18134_));
 NAND2x1_ASAP7_75t_R _24792_ (.A(_05280_),
    .B(_05303_),
    .Y(_18220_));
 NAND2x1_ASAP7_75t_R _24793_ (.A(_05168_),
    .B(_05200_),
    .Y(_17352_));
 OA22x2_ASAP7_75t_R _24794_ (.A1(_00795_),
    .A2(_05499_),
    .B1(_05179_),
    .B2(_01052_),
    .Y(_17355_));
 NAND2x1_ASAP7_75t_R _24795_ (.A(_05168_),
    .B(_05213_),
    .Y(_17362_));
 OA22x2_ASAP7_75t_R _24796_ (.A1(_00801_),
    .A2(_05499_),
    .B1(_05178_),
    .B2(_01118_),
    .Y(_17378_));
 NAND2x1_ASAP7_75t_R _24797_ (.A(_05192_),
    .B(_05500_),
    .Y(_17403_));
 NAND2x1_ASAP7_75t_R _24798_ (.A(_05168_),
    .B(_05237_),
    .Y(_17415_));
 NAND2x1_ASAP7_75t_R _24799_ (.A(_05207_),
    .B(_05501_),
    .Y(_17427_));
 OA22x2_ASAP7_75t_R _24800_ (.A1(_00809_),
    .A2(_05499_),
    .B1(_05178_),
    .B2(_05317_),
    .Y(_17436_));
 NAND2x1_ASAP7_75t_R _24801_ (.A(_05213_),
    .B(_05502_),
    .Y(_17535_));
 OA22x2_ASAP7_75t_R _24802_ (.A1(_00821_),
    .A2(_05152_),
    .B1(_05178_),
    .B2(_05319_),
    .Y(_17555_));
 NAND2x1_ASAP7_75t_R _24803_ (.A(_05216_),
    .B(_05237_),
    .Y(_17579_));
 OA22x2_ASAP7_75t_R _24804_ (.A1(_00854_),
    .A2(_05152_),
    .B1(_05178_),
    .B2(_01382_),
    .Y(_17594_));
 NAND2x1_ASAP7_75t_R _24805_ (.A(_05206_),
    .B(_05255_),
    .Y(_17610_));
 NAND2x1_ASAP7_75t_R _24806_ (.A(_05220_),
    .B(_05503_),
    .Y(_17614_));
 NAND2x1_ASAP7_75t_R _24807_ (.A(_05216_),
    .B(_05244_),
    .Y(_17621_));
 OA22x2_ASAP7_75t_R _24808_ (.A1(_00887_),
    .A2(_05152_),
    .B1(_05178_),
    .B2(_05320_),
    .Y(_17635_));
 NAND2x1_ASAP7_75t_R _24809_ (.A(_05502_),
    .B(_05237_),
    .Y(_17654_));
 NAND2x1_ASAP7_75t_R _24810_ (.A(_05209_),
    .B(_05260_),
    .Y(_17664_));
 OA22x2_ASAP7_75t_R _24811_ (.A1(_00920_),
    .A2(_05152_),
    .B1(_05178_),
    .B2(_04868_),
    .Y(_17677_));
 NAND2x1_ASAP7_75t_R _24812_ (.A(_05502_),
    .B(_05244_),
    .Y(_17703_));
 NAND2x1_ASAP7_75t_R _24813_ (.A(_05199_),
    .B(_05288_),
    .Y(_17745_));
 NAND2x1_ASAP7_75t_R _24814_ (.A(_05233_),
    .B(_05252_),
    .Y(_17756_));
 NAND2x1_ASAP7_75t_R _24815_ (.A(_05216_),
    .B(_05269_),
    .Y(_17767_));
 NAND2x1_ASAP7_75t_R _24816_ (.A(_05213_),
    .B(_05504_),
    .Y(_17794_));
 NAND2x1_ASAP7_75t_R _24817_ (.A(_05240_),
    .B(_05252_),
    .Y(_17805_));
 NAND2x1_ASAP7_75t_R _24818_ (.A(_05209_),
    .B(_05285_),
    .Y(_17815_));
 NAND2x1_ASAP7_75t_R _24819_ (.A(_05220_),
    .B(_05504_),
    .Y(_17839_));
 NAND2x1_ASAP7_75t_R _24820_ (.A(_05240_),
    .B(_05260_),
    .Y(_17850_));
 NAND2x1_ASAP7_75t_R _24821_ (.A(_05209_),
    .B(_05293_),
    .Y(_17860_));
 NAND2x1_ASAP7_75t_R _24822_ (.A(_05220_),
    .B(_05288_),
    .Y(_17886_));
 NAND2x1_ASAP7_75t_R _24823_ (.A(_05233_),
    .B(_05276_),
    .Y(_17897_));
 NAND2x1_ASAP7_75t_R _24824_ (.A(_05216_),
    .B(_05293_),
    .Y(_17907_));
 NAND2x1_ASAP7_75t_R _24825_ (.A(_05233_),
    .B(_05285_),
    .Y(_17943_));
 NAND2x1_ASAP7_75t_R _24826_ (.A(_05244_),
    .B(_05504_),
    .Y(_17973_));
 NAND2x1_ASAP7_75t_R _24827_ (.A(_05240_),
    .B(_05285_),
    .Y(_17984_));
 NAND2x1_ASAP7_75t_R _24828_ (.A(_05244_),
    .B(_05288_),
    .Y(_18013_));
 NAND2x1_ASAP7_75t_R _24829_ (.A(_05233_),
    .B(_05303_),
    .Y(_18025_));
 NAND2x1_ASAP7_75t_R _24830_ (.A(_05255_),
    .B(_05284_),
    .Y(_18063_));
 NAND2x1_ASAP7_75t_R _24831_ (.A(_05268_),
    .B(_05280_),
    .Y(_18096_));
 NAND2x1_ASAP7_75t_R _24832_ (.A(_05255_),
    .B(_05292_),
    .Y(_18101_));
 NAND2x1_ASAP7_75t_R _24833_ (.A(_05280_),
    .B(_05284_),
    .Y(_18163_));
 NAND2x1_ASAP7_75t_R _24834_ (.A(_05280_),
    .B(_05292_),
    .Y(_18193_));
 NAND2x1_ASAP7_75t_R _24835_ (.A(_05288_),
    .B(_05292_),
    .Y(_18221_));
 NAND2x2_ASAP7_75t_R _24836_ (.A(_05280_),
    .B(_05309_),
    .Y(_18251_));
 INVx1_ASAP7_75t_R _24837_ (.A(_00233_),
    .Y(_17831_));
 INVx1_ASAP7_75t_R _24838_ (.A(_00239_),
    .Y(_17924_));
 INVx1_ASAP7_75t_R _24839_ (.A(_00242_),
    .Y(_17964_));
 INVx1_ASAP7_75t_R _24840_ (.A(_00266_),
    .Y(_18242_));
 INVx2_ASAP7_75t_R _24841_ (.A(net2011),
    .Y(_18077_));
 INVx1_ASAP7_75t_R _24842_ (.A(_00272_),
    .Y(_18262_));
 INVx1_ASAP7_75t_R _24843_ (.A(_00276_),
    .Y(_18284_));
 INVx1_ASAP7_75t_R _24844_ (.A(_18679_),
    .Y(_18677_));
 INVx1_ASAP7_75t_R _24845_ (.A(_18684_),
    .Y(_18682_));
 INVx1_ASAP7_75t_R _24846_ (.A(_18714_),
    .Y(_18712_));
 INVx1_ASAP7_75t_R _24847_ (.A(_18724_),
    .Y(_18722_));
 INVx1_ASAP7_75t_R _24848_ (.A(_18729_),
    .Y(_18727_));
 INVx1_ASAP7_75t_R _24849_ (.A(_18739_),
    .Y(_18737_));
 INVx1_ASAP7_75t_R _24850_ (.A(_18759_),
    .Y(_18757_));
 INVx4_ASAP7_75t_R _24851_ (.A(_00288_),
    .Y(_05507_));
 BUFx6f_ASAP7_75t_R _24852_ (.A(_00290_),
    .Y(_05508_));
 AO21x1_ASAP7_75t_R _24853_ (.A1(_02226_),
    .A2(_02227_),
    .B(_05508_),
    .Y(_05509_));
 OA21x2_ASAP7_75t_R _24854_ (.A1(_04933_),
    .A2(_05340_),
    .B(_05380_),
    .Y(_05510_));
 OA21x2_ASAP7_75t_R _24855_ (.A1(_05374_),
    .A2(_05510_),
    .B(_00289_),
    .Y(_05511_));
 OAI21x1_ASAP7_75t_R _24856_ (.A1(_05388_),
    .A2(_05509_),
    .B(_05511_),
    .Y(_05512_));
 OR2x4_ASAP7_75t_R _24857_ (.A(_05507_),
    .B(_05512_),
    .Y(_05513_));
 INVx3_ASAP7_75t_R _24858_ (.A(_05513_),
    .Y(_18773_));
 BUFx4f_ASAP7_75t_R _24859_ (.A(_05304_),
    .Y(_05514_));
 BUFx4f_ASAP7_75t_R _24860_ (.A(_05514_),
    .Y(_05515_));
 BUFx4f_ASAP7_75t_R _24861_ (.A(_05515_),
    .Y(_05516_));
 BUFx4f_ASAP7_75t_R _24862_ (.A(_05516_),
    .Y(_05517_));
 BUFx6f_ASAP7_75t_R _24863_ (.A(_05517_),
    .Y(_05518_));
 BUFx16f_ASAP7_75t_R _24864_ (.A(_14922_),
    .Y(_05519_));
 XNOR2x1_ASAP7_75t_R _24865_ (.B(_05519_),
    .Y(_05520_),
    .A(_18614_));
 BUFx3_ASAP7_75t_R _24866_ (.A(_05142_),
    .Y(_05521_));
 BUFx3_ASAP7_75t_R _24867_ (.A(_04870_),
    .Y(_05522_));
 BUFx4f_ASAP7_75t_R _24868_ (.A(_00408_),
    .Y(_05523_));
 BUFx6f_ASAP7_75t_R _24869_ (.A(_00407_),
    .Y(_05524_));
 AND2x4_ASAP7_75t_R _24870_ (.A(_01816_),
    .B(_02217_),
    .Y(_05525_));
 AND3x4_ASAP7_75t_R _24871_ (.A(_05523_),
    .B(_05524_),
    .C(_05525_),
    .Y(_05526_));
 BUFx4f_ASAP7_75t_R _24872_ (.A(_05526_),
    .Y(_05527_));
 NAND2x2_ASAP7_75t_R _24873_ (.A(_13514_),
    .B(_13549_),
    .Y(_05528_));
 AO222x2_ASAP7_75t_R _24874_ (.A1(_05139_),
    .A2(_00414_),
    .B1(_01764_),
    .B2(_05522_),
    .C1(_05527_),
    .C2(_05528_),
    .Y(_05529_));
 BUFx6f_ASAP7_75t_R _24875_ (.A(_05524_),
    .Y(_05530_));
 AND2x2_ASAP7_75t_R _24876_ (.A(_13733_),
    .B(_13768_),
    .Y(_05531_));
 NOR2x1_ASAP7_75t_R _24877_ (.A(_05530_),
    .B(_05531_),
    .Y(_05532_));
 OR3x1_ASAP7_75t_R _24878_ (.A(_05521_),
    .B(_05529_),
    .C(_05532_),
    .Y(_05533_));
 OA21x2_ASAP7_75t_R _24879_ (.A1(_05518_),
    .A2(_05520_),
    .B(_05533_),
    .Y(_18784_));
 BUFx6f_ASAP7_75t_R _24880_ (.A(_05517_),
    .Y(_05534_));
 BUFx3_ASAP7_75t_R _24881_ (.A(_05142_),
    .Y(_05535_));
 BUFx3_ASAP7_75t_R _24882_ (.A(_05525_),
    .Y(_05536_));
 BUFx3_ASAP7_75t_R _24883_ (.A(_05536_),
    .Y(_05537_));
 OR3x1_ASAP7_75t_R _24884_ (.A(_00447_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05538_));
 OAI21x1_ASAP7_75t_R _24885_ (.A1(_18611_),
    .A2(_05534_),
    .B(_05538_),
    .Y(_17345_));
 OR3x1_ASAP7_75t_R _24886_ (.A(_00792_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05539_));
 OAI21x1_ASAP7_75t_R _24887_ (.A1(_18620_),
    .A2(_05534_),
    .B(_05539_),
    .Y(_18786_));
 BUFx3_ASAP7_75t_R _24888_ (.A(_05142_),
    .Y(_05540_));
 BUFx6f_ASAP7_75t_R _24889_ (.A(_05540_),
    .Y(_05541_));
 XNOR2x1_ASAP7_75t_R _24890_ (.B(_05519_),
    .Y(_05542_),
    .A(_18625_));
 BUFx4f_ASAP7_75t_R _24891_ (.A(_05524_),
    .Y(_05543_));
 BUFx4f_ASAP7_75t_R _24892_ (.A(_05523_),
    .Y(_05544_));
 INVx2_ASAP7_75t_R _24893_ (.A(_00795_),
    .Y(_05545_));
 INVx1_ASAP7_75t_R _24894_ (.A(_01750_),
    .Y(_05546_));
 BUFx4f_ASAP7_75t_R _24895_ (.A(_04879_),
    .Y(_05547_));
 OA222x2_ASAP7_75t_R _24896_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05546_),
    .B2(_05536_),
    .C1(_05547_),
    .C2(_14225_),
    .Y(_05548_));
 BUFx3_ASAP7_75t_R _24897_ (.A(_05516_),
    .Y(_05549_));
 OA211x2_ASAP7_75t_R _24898_ (.A1(_05543_),
    .A2(_05204_),
    .B(_05548_),
    .C(_05549_),
    .Y(_05550_));
 AOI21x1_ASAP7_75t_R _24899_ (.A1(_05541_),
    .A2(_05542_),
    .B(_05550_),
    .Y(_18788_));
 OR3x1_ASAP7_75t_R _24900_ (.A(_00798_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05551_));
 OAI21x1_ASAP7_75t_R _24901_ (.A1(_05534_),
    .A2(_18628_),
    .B(_05551_),
    .Y(_18790_));
 XNOR2x1_ASAP7_75t_R _24902_ (.B(_05519_),
    .Y(_05552_),
    .A(_18632_));
 AND2x2_ASAP7_75t_R _24903_ (.A(_15087_),
    .B(_15113_),
    .Y(_05553_));
 NOR2x1_ASAP7_75t_R _24904_ (.A(_05530_),
    .B(_05553_),
    .Y(_05554_));
 BUFx4f_ASAP7_75t_R _24905_ (.A(_05138_),
    .Y(_05555_));
 AO222x2_ASAP7_75t_R _24906_ (.A1(_05555_),
    .A2(_00801_),
    .B1(_01748_),
    .B2(_04870_),
    .C1(_05526_),
    .C2(_14371_),
    .Y(_05556_));
 OR3x1_ASAP7_75t_R _24907_ (.A(_05521_),
    .B(_05554_),
    .C(_05556_),
    .Y(_05557_));
 OA21x2_ASAP7_75t_R _24908_ (.A1(_05518_),
    .A2(_05552_),
    .B(_05557_),
    .Y(_18792_));
 INVx2_ASAP7_75t_R _24909_ (.A(_14426_),
    .Y(_05558_));
 NAND2x2_ASAP7_75t_R _24910_ (.A(_15154_),
    .B(_15179_),
    .Y(_05559_));
 AO222x2_ASAP7_75t_R _24911_ (.A1(_05139_),
    .A2(_00804_),
    .B1(_01746_),
    .B2(_05522_),
    .C1(_05559_),
    .C2(_05109_),
    .Y(_05560_));
 AO21x1_ASAP7_75t_R _24912_ (.A1(_05558_),
    .A2(_05527_),
    .B(_05560_),
    .Y(_05561_));
 BUFx12f_ASAP7_75t_R _24913_ (.A(_14922_),
    .Y(_05562_));
 XNOR2x1_ASAP7_75t_R _24914_ (.B(_05562_),
    .Y(_05563_),
    .A(_18638_));
 AND2x2_ASAP7_75t_R _24915_ (.A(_05563_),
    .B(_05142_),
    .Y(_05564_));
 AO21x1_ASAP7_75t_R _24916_ (.A1(_05517_),
    .A2(_05561_),
    .B(_05564_),
    .Y(_18794_));
 XNOR2x1_ASAP7_75t_R _24917_ (.B(_05519_),
    .Y(_05565_),
    .A(_18645_));
 INVx2_ASAP7_75t_R _24918_ (.A(_00807_),
    .Y(_05566_));
 INVx1_ASAP7_75t_R _24919_ (.A(_01745_),
    .Y(_05567_));
 AND2x2_ASAP7_75t_R _24920_ (.A(_15206_),
    .B(_15234_),
    .Y(_05568_));
 OA222x2_ASAP7_75t_R _24921_ (.A1(_05544_),
    .A2(_05566_),
    .B1(_05567_),
    .B2(_05536_),
    .C1(_05568_),
    .C2(_05524_),
    .Y(_05569_));
 OA211x2_ASAP7_75t_R _24922_ (.A1(_14486_),
    .A2(_05547_),
    .B(_05569_),
    .C(_05549_),
    .Y(_05570_));
 AOI21x1_ASAP7_75t_R _24923_ (.A1(_05541_),
    .A2(_05565_),
    .B(_05570_),
    .Y(_18796_));
 INVx3_ASAP7_75t_R _24924_ (.A(_00809_),
    .Y(_05571_));
 BUFx3_ASAP7_75t_R _24925_ (.A(_05522_),
    .Y(_05572_));
 BUFx4f_ASAP7_75t_R _24926_ (.A(_05142_),
    .Y(_05573_));
 AO21x1_ASAP7_75t_R _24927_ (.A1(_05571_),
    .A2(_05572_),
    .B(_05573_),
    .Y(_05574_));
 OA21x2_ASAP7_75t_R _24928_ (.A1(_05518_),
    .A2(_18647_),
    .B(_05574_),
    .Y(_18798_));
 BUFx3_ASAP7_75t_R _24929_ (.A(_05516_),
    .Y(_05575_));
 XNOR2x1_ASAP7_75t_R _24930_ (.B(_05519_),
    .Y(_05576_),
    .A(_18652_));
 NAND2x1_ASAP7_75t_R _24931_ (.A(_15365_),
    .B(_15390_),
    .Y(_05577_));
 AO22x1_ASAP7_75t_R _24932_ (.A1(_05109_),
    .A2(_05577_),
    .B1(_05522_),
    .B2(_02222_),
    .Y(_05578_));
 INVx2_ASAP7_75t_R _24933_ (.A(_00812_),
    .Y(_05579_));
 OAI22x1_ASAP7_75t_R _24934_ (.A1(_05544_),
    .A2(_05579_),
    .B1(_14603_),
    .B2(_05547_),
    .Y(_05580_));
 OR3x1_ASAP7_75t_R _24935_ (.A(_05521_),
    .B(_05578_),
    .C(_05580_),
    .Y(_05581_));
 OA21x2_ASAP7_75t_R _24936_ (.A1(_05575_),
    .A2(_05576_),
    .B(_05581_),
    .Y(_18800_));
 XNOR2x1_ASAP7_75t_R _24937_ (.B(_05519_),
    .Y(_05582_),
    .A(_18660_));
 INVx2_ASAP7_75t_R _24938_ (.A(_00815_),
    .Y(_05583_));
 INVx1_ASAP7_75t_R _24939_ (.A(_01774_),
    .Y(_05584_));
 BUFx3_ASAP7_75t_R _24940_ (.A(_05525_),
    .Y(_05585_));
 OA222x2_ASAP7_75t_R _24941_ (.A1(_05544_),
    .A2(_05583_),
    .B1(_05584_),
    .B2(_05585_),
    .C1(_05256_),
    .C2(_05524_),
    .Y(_05586_));
 OA211x2_ASAP7_75t_R _24942_ (.A1(_14666_),
    .A2(_05547_),
    .B(_05586_),
    .C(_05549_),
    .Y(_05587_));
 AOI21x1_ASAP7_75t_R _24943_ (.A1(_05541_),
    .A2(_05582_),
    .B(_05587_),
    .Y(_18802_));
 NAND2x1_ASAP7_75t_R _24944_ (.A(_14775_),
    .B(_14803_),
    .Y(_05588_));
 INVx2_ASAP7_75t_R _24945_ (.A(_14723_),
    .Y(_05589_));
 AO222x2_ASAP7_75t_R _24946_ (.A1(_05139_),
    .A2(_05506_),
    .B1(_01773_),
    .B2(_05522_),
    .C1(_05527_),
    .C2(_05589_),
    .Y(_05590_));
 AO21x1_ASAP7_75t_R _24947_ (.A1(_05109_),
    .A2(_05588_),
    .B(_05590_),
    .Y(_05591_));
 XNOR2x1_ASAP7_75t_R _24948_ (.B(_05562_),
    .Y(_05592_),
    .A(_18663_));
 AND2x2_ASAP7_75t_R _24949_ (.A(_05142_),
    .B(_05592_),
    .Y(_05593_));
 AO21x1_ASAP7_75t_R _24950_ (.A1(_05517_),
    .A2(_05591_),
    .B(_05593_),
    .Y(_18804_));
 OR3x1_ASAP7_75t_R _24951_ (.A(_00821_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05594_));
 OAI21x1_ASAP7_75t_R _24952_ (.A1(_18669_),
    .A2(_05534_),
    .B(_05594_),
    .Y(_18806_));
 BUFx12_ASAP7_75t_R _24953_ (.A(_04901_),
    .Y(_05595_));
 XNOR2x1_ASAP7_75t_R _24954_ (.B(_18673_),
    .Y(_05596_),
    .A(_05595_));
 AND2x2_ASAP7_75t_R _24955_ (.A(_15698_),
    .B(_15723_),
    .Y(_05597_));
 INVx2_ASAP7_75t_R _24956_ (.A(_00854_),
    .Y(_05598_));
 INVx1_ASAP7_75t_R _24957_ (.A(_01771_),
    .Y(_05599_));
 OA222x2_ASAP7_75t_R _24958_ (.A1(_05544_),
    .A2(_05598_),
    .B1(_05599_),
    .B2(_05585_),
    .C1(_05547_),
    .C2(_15671_),
    .Y(_05600_));
 OA211x2_ASAP7_75t_R _24959_ (.A1(_05543_),
    .A2(_05597_),
    .B(_05600_),
    .C(_05549_),
    .Y(_05601_));
 AOI21x1_ASAP7_75t_R _24960_ (.A1(_05541_),
    .A2(_05596_),
    .B(_05601_),
    .Y(_18808_));
 XNOR2x1_ASAP7_75t_R _24961_ (.B(_18679_),
    .Y(_05602_),
    .A(_05595_));
 AND2x2_ASAP7_75t_R _24962_ (.A(_15839_),
    .B(_15863_),
    .Y(_05603_));
 INVx3_ASAP7_75t_R _24963_ (.A(_00887_),
    .Y(_05604_));
 INVx1_ASAP7_75t_R _24964_ (.A(_01770_),
    .Y(_05605_));
 OA222x2_ASAP7_75t_R _24965_ (.A1(_05544_),
    .A2(_05604_),
    .B1(_05605_),
    .B2(_05585_),
    .C1(_05547_),
    .C2(_15816_),
    .Y(_05606_));
 OA211x2_ASAP7_75t_R _24966_ (.A1(_05543_),
    .A2(_05603_),
    .B(_05606_),
    .C(_05549_),
    .Y(_05607_));
 AOI21x1_ASAP7_75t_R _24967_ (.A1(_05541_),
    .A2(_05602_),
    .B(_05607_),
    .Y(_18810_));
 XNOR2x1_ASAP7_75t_R _24968_ (.B(_18684_),
    .Y(_05608_),
    .A(_05595_));
 INVx2_ASAP7_75t_R _24969_ (.A(_00920_),
    .Y(_05609_));
 INVx1_ASAP7_75t_R _24970_ (.A(_01769_),
    .Y(_05610_));
 OA222x2_ASAP7_75t_R _24971_ (.A1(_05544_),
    .A2(_05609_),
    .B1(_05610_),
    .B2(_05585_),
    .C1(_05547_),
    .C2(_15950_),
    .Y(_05611_));
 OA211x2_ASAP7_75t_R _24972_ (.A1(_05543_),
    .A2(_05300_),
    .B(_05611_),
    .C(_05549_),
    .Y(_05612_));
 AOI21x1_ASAP7_75t_R _24973_ (.A1(_05541_),
    .A2(_05608_),
    .B(_05612_),
    .Y(_18812_));
 XNOR2x1_ASAP7_75t_R _24974_ (.B(_18688_),
    .Y(_05613_),
    .A(_05595_));
 INVx1_ASAP7_75t_R _24975_ (.A(_05180_),
    .Y(_05614_));
 INVx1_ASAP7_75t_R _24976_ (.A(_01768_),
    .Y(_05615_));
 OA222x2_ASAP7_75t_R _24977_ (.A1(_05544_),
    .A2(_05614_),
    .B1(_05615_),
    .B2(_05585_),
    .C1(_05547_),
    .C2(_16094_),
    .Y(_05616_));
 OA211x2_ASAP7_75t_R _24978_ (.A1(_05543_),
    .A2(_05169_),
    .B(_05616_),
    .C(_05549_),
    .Y(_05617_));
 AOI21x1_ASAP7_75t_R _24979_ (.A1(_05541_),
    .A2(_05613_),
    .B(_05617_),
    .Y(_18814_));
 OR3x1_ASAP7_75t_R _24980_ (.A(_00986_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05618_));
 OAI21x1_ASAP7_75t_R _24981_ (.A1(_05534_),
    .A2(_18694_),
    .B(_05618_),
    .Y(_18816_));
 OR3x1_ASAP7_75t_R _24982_ (.A(_01019_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05619_));
 OAI21x1_ASAP7_75t_R _24983_ (.A1(_05534_),
    .A2(_18699_),
    .B(_05619_),
    .Y(_18818_));
 XNOR2x1_ASAP7_75t_R _24984_ (.B(_18703_),
    .Y(_05620_),
    .A(_05595_));
 AND2x2_ASAP7_75t_R _24985_ (.A(_16489_),
    .B(_16512_),
    .Y(_05621_));
 BUFx4f_ASAP7_75t_R _24986_ (.A(_05523_),
    .Y(_05622_));
 INVx4_ASAP7_75t_R _24987_ (.A(_01052_),
    .Y(_05623_));
 INVx1_ASAP7_75t_R _24988_ (.A(_01765_),
    .Y(_05624_));
 OA222x2_ASAP7_75t_R _24989_ (.A1(_05622_),
    .A2(_05623_),
    .B1(_05624_),
    .B2(_05585_),
    .C1(_04879_),
    .C2(_16466_),
    .Y(_05625_));
 OA211x2_ASAP7_75t_R _24990_ (.A1(_05543_),
    .A2(_05621_),
    .B(_05625_),
    .C(_05549_),
    .Y(_05626_));
 AOI21x1_ASAP7_75t_R _24991_ (.A1(_05541_),
    .A2(_05620_),
    .B(_05626_),
    .Y(_18820_));
 XNOR2x1_ASAP7_75t_R _24992_ (.B(_18708_),
    .Y(_05627_),
    .A(_05519_));
 BUFx3_ASAP7_75t_R _24993_ (.A(_05142_),
    .Y(_05628_));
 BUFx3_ASAP7_75t_R _24994_ (.A(_04870_),
    .Y(_05629_));
 AO222x2_ASAP7_75t_R _24995_ (.A1(_05139_),
    .A2(_05315_),
    .B1(_01763_),
    .B2(_05629_),
    .C1(_05527_),
    .C2(_16592_),
    .Y(_05630_));
 AND2x2_ASAP7_75t_R _24996_ (.A(_16618_),
    .B(_16641_),
    .Y(_05631_));
 NOR2x1_ASAP7_75t_R _24997_ (.A(_05530_),
    .B(_05631_),
    .Y(_05632_));
 OR3x1_ASAP7_75t_R _24998_ (.A(_05628_),
    .B(_05630_),
    .C(_05632_),
    .Y(_05633_));
 OA21x2_ASAP7_75t_R _24999_ (.A1(_05575_),
    .A2(_05627_),
    .B(_05633_),
    .Y(_18822_));
 XNOR2x1_ASAP7_75t_R _25000_ (.B(_18714_),
    .Y(_05634_),
    .A(_05519_));
 AO222x2_ASAP7_75t_R _25001_ (.A1(_05139_),
    .A2(_01118_),
    .B1(_01762_),
    .B2(_05629_),
    .C1(_05527_),
    .C2(_16706_),
    .Y(_05635_));
 NOR2x1_ASAP7_75t_R _25002_ (.A(_05530_),
    .B(_05217_),
    .Y(_05636_));
 OR3x1_ASAP7_75t_R _25003_ (.A(_05628_),
    .B(_05635_),
    .C(_05636_),
    .Y(_05637_));
 OA21x2_ASAP7_75t_R _25004_ (.A1(_05575_),
    .A2(_05634_),
    .B(_05637_),
    .Y(_18824_));
 XNOR2x1_ASAP7_75t_R _25005_ (.B(_18718_),
    .Y(_05638_),
    .A(_05562_));
 AO222x2_ASAP7_75t_R _25006_ (.A1(_05555_),
    .A2(_05316_),
    .B1(_01761_),
    .B2(_05629_),
    .C1(_05527_),
    .C2(_16836_),
    .Y(_05639_));
 NOR2x1_ASAP7_75t_R _25007_ (.A(_05530_),
    .B(_05225_),
    .Y(_05640_));
 OR3x1_ASAP7_75t_R _25008_ (.A(_05628_),
    .B(_05639_),
    .C(_05640_),
    .Y(_05641_));
 OA21x2_ASAP7_75t_R _25009_ (.A1(_05575_),
    .A2(_05638_),
    .B(_05641_),
    .Y(_18826_));
 INVx2_ASAP7_75t_R _25010_ (.A(_01184_),
    .Y(_05642_));
 AO21x1_ASAP7_75t_R _25011_ (.A1(_05642_),
    .A2(_05572_),
    .B(_05573_),
    .Y(_05643_));
 OA21x2_ASAP7_75t_R _25012_ (.A1(_05575_),
    .A2(_18725_),
    .B(_05643_),
    .Y(_18828_));
 OR3x1_ASAP7_75t_R _25013_ (.A(_05317_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05644_));
 OAI21x1_ASAP7_75t_R _25014_ (.A1(_05534_),
    .A2(_18728_),
    .B(_05644_),
    .Y(_18830_));
 INVx2_ASAP7_75t_R _25015_ (.A(_01250_),
    .Y(_05645_));
 AO21x1_ASAP7_75t_R _25016_ (.A1(_05645_),
    .A2(_05572_),
    .B(_05573_),
    .Y(_05646_));
 OA21x2_ASAP7_75t_R _25017_ (.A1(_05575_),
    .A2(_18732_),
    .B(_05646_),
    .Y(_18832_));
 XNOR2x1_ASAP7_75t_R _25018_ (.B(_18739_),
    .Y(_05647_),
    .A(net2007));
 AO222x2_ASAP7_75t_R _25019_ (.A1(_05555_),
    .A2(_05318_),
    .B1(_01757_),
    .B2(_05629_),
    .C1(_05527_),
    .C2(_17316_),
    .Y(_05648_));
 NAND2x2_ASAP7_75t_R _25020_ (.A(_17338_),
    .B(_04279_),
    .Y(_05649_));
 AND2x2_ASAP7_75t_R _25021_ (.A(_05109_),
    .B(_05649_),
    .Y(_05650_));
 OR3x1_ASAP7_75t_R _25022_ (.A(_05628_),
    .B(_05648_),
    .C(_05650_),
    .Y(_05651_));
 OA21x2_ASAP7_75t_R _25023_ (.A1(_05575_),
    .A2(_05647_),
    .B(_05651_),
    .Y(_18834_));
 XNOR2x1_ASAP7_75t_R _25024_ (.B(_18743_),
    .Y(_05652_),
    .A(_05562_));
 AO222x2_ASAP7_75t_R _25025_ (.A1(_05555_),
    .A2(_01316_),
    .B1(_01756_),
    .B2(_05629_),
    .C1(_05527_),
    .C2(_04343_),
    .Y(_05653_));
 NOR2x1_ASAP7_75t_R _25026_ (.A(_05530_),
    .B(_05265_),
    .Y(_05654_));
 OR3x1_ASAP7_75t_R _25027_ (.A(_05628_),
    .B(_05653_),
    .C(_05654_),
    .Y(_05655_));
 OA21x2_ASAP7_75t_R _25028_ (.A1(_05575_),
    .A2(_05652_),
    .B(_05655_),
    .Y(_18836_));
 XNOR2x1_ASAP7_75t_R _25029_ (.B(_18748_),
    .Y(_05656_),
    .A(net2007));
 AO222x2_ASAP7_75t_R _25030_ (.A1(_05555_),
    .A2(_05319_),
    .B1(_01755_),
    .B2(_05629_),
    .C1(_05527_),
    .C2(_04473_),
    .Y(_05657_));
 NOR2x1_ASAP7_75t_R _25031_ (.A(_05530_),
    .B(_05273_),
    .Y(_05658_));
 OR3x1_ASAP7_75t_R _25032_ (.A(_05628_),
    .B(_05657_),
    .C(_05658_),
    .Y(_05659_));
 OA21x2_ASAP7_75t_R _25033_ (.A1(_05575_),
    .A2(_05656_),
    .B(_05659_),
    .Y(_18838_));
 XNOR2x1_ASAP7_75t_R _25034_ (.B(_18753_),
    .Y(_05660_),
    .A(net2007));
 AO222x2_ASAP7_75t_R _25035_ (.A1(_05555_),
    .A2(_01382_),
    .B1(_01754_),
    .B2(_05629_),
    .C1(_05527_),
    .C2(_04583_),
    .Y(_05661_));
 NOR2x1_ASAP7_75t_R _25036_ (.A(_05530_),
    .B(_05281_),
    .Y(_05662_));
 OR3x1_ASAP7_75t_R _25037_ (.A(_05628_),
    .B(_05661_),
    .C(_05662_),
    .Y(_05663_));
 OA21x2_ASAP7_75t_R _25038_ (.A1(_05575_),
    .A2(_05660_),
    .B(_05663_),
    .Y(_18840_));
 BUFx3_ASAP7_75t_R _25039_ (.A(_05516_),
    .Y(_05664_));
 XNOR2x1_ASAP7_75t_R _25040_ (.B(_18759_),
    .Y(_05665_),
    .A(net2007));
 AO222x2_ASAP7_75t_R _25041_ (.A1(_05555_),
    .A2(_05320_),
    .B1(_01752_),
    .B2(_05629_),
    .C1(_05526_),
    .C2(_04697_),
    .Y(_05666_));
 NOR2x1_ASAP7_75t_R _25042_ (.A(_05524_),
    .B(_05289_),
    .Y(_05667_));
 OR3x1_ASAP7_75t_R _25043_ (.A(_05628_),
    .B(_05666_),
    .C(_05667_),
    .Y(_05668_));
 OA21x2_ASAP7_75t_R _25044_ (.A1(_05664_),
    .A2(_05665_),
    .B(_05668_),
    .Y(_18842_));
 AND2x2_ASAP7_75t_R _25045_ (.A(_14071_),
    .B(_18652_),
    .Y(_18849_));
 BUFx6f_ASAP7_75t_R _25046_ (.A(_14736_),
    .Y(_18861_));
 INVx1_ASAP7_75t_R _25047_ (.A(_00169_),
    .Y(_17412_));
 INVx1_ASAP7_75t_R _25048_ (.A(_00173_),
    .Y(_17411_));
 INVx1_ASAP7_75t_R _25049_ (.A(_00217_),
    .Y(_19040_));
 INVx1_ASAP7_75t_R _25050_ (.A(_00218_),
    .Y(_17651_));
 INVx1_ASAP7_75t_R _25051_ (.A(_00221_),
    .Y(_17681_));
 INVx1_ASAP7_75t_R _25052_ (.A(_18038_),
    .Y(_18037_));
 INVx1_ASAP7_75t_R _25053_ (.A(_18079_),
    .Y(_18036_));
 INVx1_ASAP7_75t_R _25054_ (.A(_00257_),
    .Y(_18156_));
 INVx2_ASAP7_75t_R _25055_ (.A(net1968),
    .Y(_18078_));
 INVx3_ASAP7_75t_R _25056_ (.A(_18227_),
    .Y(_18226_));
 INVx1_ASAP7_75t_R _25057_ (.A(net1),
    .Y(_17912_));
 INVx1_ASAP7_75t_R _25058_ (.A(_00278_),
    .Y(_18292_));
 INVx1_ASAP7_75t_R _25059_ (.A(_00279_),
    .Y(_18312_));
 INVx1_ASAP7_75t_R _25060_ (.A(_18668_),
    .Y(_18670_));
 INVx1_ASAP7_75t_R _25061_ (.A(_18673_),
    .Y(_18675_));
 INVx1_ASAP7_75t_R _25062_ (.A(_18688_),
    .Y(_18690_));
 INVx1_ASAP7_75t_R _25063_ (.A(_18693_),
    .Y(_18695_));
 INVx1_ASAP7_75t_R _25064_ (.A(_18698_),
    .Y(_18700_));
 INVx1_ASAP7_75t_R _25065_ (.A(_18703_),
    .Y(_18705_));
 INVx1_ASAP7_75t_R _25066_ (.A(_18708_),
    .Y(_18710_));
 INVx1_ASAP7_75t_R _25067_ (.A(_18718_),
    .Y(_18720_));
 INVx1_ASAP7_75t_R _25068_ (.A(_18733_),
    .Y(_18735_));
 INVx1_ASAP7_75t_R _25069_ (.A(_18743_),
    .Y(_18745_));
 INVx1_ASAP7_75t_R _25070_ (.A(_18748_),
    .Y(_18750_));
 INVx1_ASAP7_75t_R _25071_ (.A(_18753_),
    .Y(_18755_));
 INVx1_ASAP7_75t_R _25072_ (.A(_18779_),
    .Y(_18778_));
 OR3x1_ASAP7_75t_R _25073_ (.A(_00414_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05669_));
 OAI21x1_ASAP7_75t_R _25074_ (.A1(_18615_),
    .A2(_05534_),
    .B(_05669_),
    .Y(_18785_));
 XNOR2x1_ASAP7_75t_R _25075_ (.B(_04901_),
    .Y(_05670_),
    .A(_18608_));
 NAND2x1_ASAP7_75t_R _25076_ (.A(_13901_),
    .B(_13941_),
    .Y(_05671_));
 NAND2x2_ASAP7_75t_R _25077_ (.A(_13821_),
    .B(_13852_),
    .Y(_05672_));
 AO222x2_ASAP7_75t_R _25078_ (.A1(_05138_),
    .A2(_00447_),
    .B1(_01775_),
    .B2(_04870_),
    .C1(_05526_),
    .C2(_05672_),
    .Y(_05673_));
 AO21x1_ASAP7_75t_R _25079_ (.A1(_05109_),
    .A2(_05671_),
    .B(_05673_),
    .Y(_05674_));
 AND2x2_ASAP7_75t_R _25080_ (.A(_05517_),
    .B(_05674_),
    .Y(_05675_));
 AO21x1_ASAP7_75t_R _25081_ (.A1(_05573_),
    .A2(_05670_),
    .B(_05675_),
    .Y(_17346_));
 XNOR2x1_ASAP7_75t_R _25082_ (.B(_05595_),
    .Y(_05676_),
    .A(_18617_));
 INVx2_ASAP7_75t_R _25083_ (.A(_00792_),
    .Y(_05677_));
 INVx1_ASAP7_75t_R _25084_ (.A(_01753_),
    .Y(_05678_));
 OA222x2_ASAP7_75t_R _25085_ (.A1(_05622_),
    .A2(_05677_),
    .B1(_05678_),
    .B2(_05525_),
    .C1(_04879_),
    .C2(_14148_),
    .Y(_05679_));
 OA211x2_ASAP7_75t_R _25086_ (.A1(_05543_),
    .A2(_05196_),
    .B(_05549_),
    .C(_05679_),
    .Y(_05680_));
 AOI21x1_ASAP7_75t_R _25087_ (.A1(_05541_),
    .A2(_05676_),
    .B(_05680_),
    .Y(_18787_));
 OR3x1_ASAP7_75t_R _25088_ (.A(_00795_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05681_));
 OAI21x1_ASAP7_75t_R _25089_ (.A1(_05534_),
    .A2(_18624_),
    .B(_05681_),
    .Y(_18789_));
 XNOR2x1_ASAP7_75t_R _25090_ (.B(_05519_),
    .Y(_05682_),
    .A(_18627_));
 INVx2_ASAP7_75t_R _25091_ (.A(_00798_),
    .Y(_05683_));
 INVx1_ASAP7_75t_R _25092_ (.A(_01749_),
    .Y(_05684_));
 OA222x2_ASAP7_75t_R _25093_ (.A1(_05622_),
    .A2(_05683_),
    .B1(_05684_),
    .B2(_05585_),
    .C1(_05210_),
    .C2(_05524_),
    .Y(_05685_));
 OA211x2_ASAP7_75t_R _25094_ (.A1(_14295_),
    .A2(_05547_),
    .B(_05685_),
    .C(_05516_),
    .Y(_05686_));
 AOI21x1_ASAP7_75t_R _25095_ (.A1(_05541_),
    .A2(_05682_),
    .B(_05686_),
    .Y(_18791_));
 OR3x1_ASAP7_75t_R _25096_ (.A(_00801_),
    .B(_05535_),
    .C(_05537_),
    .Y(_05687_));
 OAI21x1_ASAP7_75t_R _25097_ (.A1(_05518_),
    .A2(_18635_),
    .B(_05687_),
    .Y(_18793_));
 INVx2_ASAP7_75t_R _25098_ (.A(_00804_),
    .Y(_05688_));
 AO21x1_ASAP7_75t_R _25099_ (.A1(_05688_),
    .A2(_05572_),
    .B(_05573_),
    .Y(_05689_));
 OA21x2_ASAP7_75t_R _25100_ (.A1(_05664_),
    .A2(_18637_),
    .B(_05689_),
    .Y(_18795_));
 AO21x1_ASAP7_75t_R _25101_ (.A1(_05566_),
    .A2(_05572_),
    .B(_05573_),
    .Y(_05690_));
 OA21x2_ASAP7_75t_R _25102_ (.A1(_05664_),
    .A2(_18642_),
    .B(_05690_),
    .Y(_18797_));
 XNOR2x1_ASAP7_75t_R _25103_ (.B(_05519_),
    .Y(_05691_),
    .A(_18648_));
 NAND2x2_ASAP7_75t_R _25104_ (.A(_15303_),
    .B(_15332_),
    .Y(_05692_));
 AO22x1_ASAP7_75t_R _25105_ (.A1(_05109_),
    .A2(_05692_),
    .B1(_05522_),
    .B2(_01744_),
    .Y(_05693_));
 OAI22x1_ASAP7_75t_R _25106_ (.A1(_05544_),
    .A2(_05571_),
    .B1(_05230_),
    .B2(_05547_),
    .Y(_05694_));
 OR3x1_ASAP7_75t_R _25107_ (.A(_05628_),
    .B(_05693_),
    .C(_05694_),
    .Y(_05695_));
 OA21x2_ASAP7_75t_R _25108_ (.A1(_05664_),
    .A2(_05691_),
    .B(_05695_),
    .Y(_18799_));
 AO21x1_ASAP7_75t_R _25109_ (.A1(_05579_),
    .A2(_05572_),
    .B(_05540_),
    .Y(_05696_));
 OA21x2_ASAP7_75t_R _25110_ (.A1(_05664_),
    .A2(_18653_),
    .B(_05696_),
    .Y(_18801_));
 AO21x1_ASAP7_75t_R _25111_ (.A1(_05583_),
    .A2(_05572_),
    .B(_05540_),
    .Y(_05697_));
 OA21x2_ASAP7_75t_R _25112_ (.A1(_05664_),
    .A2(_18657_),
    .B(_05697_),
    .Y(_18803_));
 OR3x1_ASAP7_75t_R _25113_ (.A(_05506_),
    .B(_05521_),
    .C(_05536_),
    .Y(_05698_));
 OAI21x1_ASAP7_75t_R _25114_ (.A1(_18664_),
    .A2(_05534_),
    .B(_05698_),
    .Y(_18805_));
 XNOR2x1_ASAP7_75t_R _25115_ (.B(_18668_),
    .Y(_05699_),
    .A(_05595_));
 AND2x2_ASAP7_75t_R _25116_ (.A(_13979_),
    .B(_14013_),
    .Y(_05700_));
 INVx1_ASAP7_75t_R _25117_ (.A(_00821_),
    .Y(_05701_));
 INVx1_ASAP7_75t_R _25118_ (.A(_01772_),
    .Y(_05702_));
 OA222x2_ASAP7_75t_R _25119_ (.A1(_05622_),
    .A2(_05701_),
    .B1(_05702_),
    .B2(_05525_),
    .C1(_04879_),
    .C2(_05261_),
    .Y(_05703_));
 OA211x2_ASAP7_75t_R _25120_ (.A1(_05543_),
    .A2(_05700_),
    .B(_05549_),
    .C(_05703_),
    .Y(_05704_));
 AOI21x1_ASAP7_75t_R _25121_ (.A1(_05573_),
    .A2(_05699_),
    .B(_05704_),
    .Y(_18807_));
 AO21x1_ASAP7_75t_R _25122_ (.A1(_05598_),
    .A2(_05572_),
    .B(_05540_),
    .Y(_05705_));
 OA21x2_ASAP7_75t_R _25123_ (.A1(_05664_),
    .A2(_18672_),
    .B(_05705_),
    .Y(_18809_));
 AO21x1_ASAP7_75t_R _25124_ (.A1(_05604_),
    .A2(_05572_),
    .B(_05540_),
    .Y(_05706_));
 OA21x2_ASAP7_75t_R _25125_ (.A1(_05664_),
    .A2(_18680_),
    .B(_05706_),
    .Y(_18811_));
 OR3x1_ASAP7_75t_R _25126_ (.A(_00920_),
    .B(_05521_),
    .C(_05536_),
    .Y(_05707_));
 OAI21x1_ASAP7_75t_R _25127_ (.A1(_05518_),
    .A2(_18683_),
    .B(_05707_),
    .Y(_18813_));
 AO21x1_ASAP7_75t_R _25128_ (.A1(_05614_),
    .A2(_05572_),
    .B(_05540_),
    .Y(_05708_));
 OA21x2_ASAP7_75t_R _25129_ (.A1(_05664_),
    .A2(_18687_),
    .B(_05708_),
    .Y(_18815_));
 XNOR2x1_ASAP7_75t_R _25130_ (.B(_18693_),
    .Y(_05709_),
    .A(_05595_));
 INVx2_ASAP7_75t_R _25131_ (.A(_00986_),
    .Y(_05710_));
 INVx1_ASAP7_75t_R _25132_ (.A(_01767_),
    .Y(_05711_));
 OA222x2_ASAP7_75t_R _25133_ (.A1(_05622_),
    .A2(_05710_),
    .B1(_05711_),
    .B2(_05585_),
    .C1(_04879_),
    .C2(_16209_),
    .Y(_05712_));
 OA211x2_ASAP7_75t_R _25134_ (.A1(_05543_),
    .A2(_05189_),
    .B(_05712_),
    .C(_05516_),
    .Y(_05713_));
 AOI21x1_ASAP7_75t_R _25135_ (.A1(_05573_),
    .A2(_05709_),
    .B(_05713_),
    .Y(_18817_));
 XNOR2x1_ASAP7_75t_R _25136_ (.B(_18698_),
    .Y(_05714_),
    .A(_05595_));
 AND2x4_ASAP7_75t_R _25137_ (.A(_16377_),
    .B(_16400_),
    .Y(_05715_));
 INVx1_ASAP7_75t_R _25138_ (.A(_01019_),
    .Y(_05716_));
 INVx1_ASAP7_75t_R _25139_ (.A(_01766_),
    .Y(_05717_));
 OA222x2_ASAP7_75t_R _25140_ (.A1(_05622_),
    .A2(_05716_),
    .B1(_05717_),
    .B2(_05585_),
    .C1(_04879_),
    .C2(_16354_),
    .Y(_05718_));
 OA211x2_ASAP7_75t_R _25141_ (.A1(_05530_),
    .A2(_05715_),
    .B(_05718_),
    .C(_05516_),
    .Y(_05719_));
 AOI21x1_ASAP7_75t_R _25142_ (.A1(_05573_),
    .A2(_05714_),
    .B(_05719_),
    .Y(_18819_));
 AO21x1_ASAP7_75t_R _25143_ (.A1(_05623_),
    .A2(_05522_),
    .B(_05540_),
    .Y(_05720_));
 OA21x2_ASAP7_75t_R _25144_ (.A1(_05664_),
    .A2(_18702_),
    .B(_05720_),
    .Y(_18821_));
 OR3x1_ASAP7_75t_R _25145_ (.A(_05315_),
    .B(_05521_),
    .C(_05536_),
    .Y(_05721_));
 OAI21x1_ASAP7_75t_R _25146_ (.A1(_05518_),
    .A2(_18709_),
    .B(_05721_),
    .Y(_18823_));
 INVx2_ASAP7_75t_R _25147_ (.A(_01118_),
    .Y(_05722_));
 AO21x1_ASAP7_75t_R _25148_ (.A1(_05722_),
    .A2(_05522_),
    .B(_05540_),
    .Y(_05723_));
 OA21x2_ASAP7_75t_R _25149_ (.A1(_05517_),
    .A2(_18715_),
    .B(_05723_),
    .Y(_18825_));
 OR3x1_ASAP7_75t_R _25150_ (.A(_05316_),
    .B(_05521_),
    .C(_05536_),
    .Y(_05724_));
 OAI21x1_ASAP7_75t_R _25151_ (.A1(_05518_),
    .A2(_18719_),
    .B(_05724_),
    .Y(_18827_));
 XNOR2x1_ASAP7_75t_R _25152_ (.B(_18724_),
    .Y(_05725_),
    .A(_05595_));
 INVx1_ASAP7_75t_R _25153_ (.A(_01760_),
    .Y(_05726_));
 OA222x2_ASAP7_75t_R _25154_ (.A1(_05622_),
    .A2(_05642_),
    .B1(_05726_),
    .B2(_05585_),
    .C1(_04879_),
    .C2(_16946_),
    .Y(_05727_));
 OA211x2_ASAP7_75t_R _25155_ (.A1(_05530_),
    .A2(_05234_),
    .B(_05727_),
    .C(_05516_),
    .Y(_05728_));
 AOI21x1_ASAP7_75t_R _25156_ (.A1(_05573_),
    .A2(_05725_),
    .B(_05728_),
    .Y(_18829_));
 XNOR2x1_ASAP7_75t_R _25157_ (.B(_18729_),
    .Y(_05729_),
    .A(net2007));
 AO222x2_ASAP7_75t_R _25158_ (.A1(_05555_),
    .A2(_05317_),
    .B1(_01759_),
    .B2(_05629_),
    .C1(_05526_),
    .C2(_17076_),
    .Y(_05730_));
 NOR2x1_ASAP7_75t_R _25159_ (.A(_05524_),
    .B(_05241_),
    .Y(_05731_));
 OR3x1_ASAP7_75t_R _25160_ (.A(_05628_),
    .B(_05730_),
    .C(_05731_),
    .Y(_05732_));
 OA21x2_ASAP7_75t_R _25161_ (.A1(_05517_),
    .A2(_05729_),
    .B(_05732_),
    .Y(_18831_));
 XNOR2x1_ASAP7_75t_R _25162_ (.B(_18733_),
    .Y(_05733_),
    .A(_05562_));
 AO222x2_ASAP7_75t_R _25163_ (.A1(_05555_),
    .A2(_01250_),
    .B1(_01758_),
    .B2(_05629_),
    .C1(_05526_),
    .C2(_17185_),
    .Y(_05734_));
 NOR2x1_ASAP7_75t_R _25164_ (.A(_05524_),
    .B(_05249_),
    .Y(_05735_));
 OR3x1_ASAP7_75t_R _25165_ (.A(_05142_),
    .B(_05734_),
    .C(_05735_),
    .Y(_05736_));
 OA21x2_ASAP7_75t_R _25166_ (.A1(_05517_),
    .A2(_05733_),
    .B(_05736_),
    .Y(_18833_));
 OR3x1_ASAP7_75t_R _25167_ (.A(_05318_),
    .B(_05521_),
    .C(_05536_),
    .Y(_05737_));
 OAI21x1_ASAP7_75t_R _25168_ (.A1(_05518_),
    .A2(_18738_),
    .B(_05737_),
    .Y(_18835_));
 INVx3_ASAP7_75t_R _25169_ (.A(_01316_),
    .Y(_05738_));
 AO21x1_ASAP7_75t_R _25170_ (.A1(_05738_),
    .A2(_05522_),
    .B(_05540_),
    .Y(_05739_));
 OA21x2_ASAP7_75t_R _25171_ (.A1(_05517_),
    .A2(_18742_),
    .B(_05739_),
    .Y(_18837_));
 OR3x1_ASAP7_75t_R _25172_ (.A(_05319_),
    .B(_05521_),
    .C(_05536_),
    .Y(_05740_));
 OAI21x1_ASAP7_75t_R _25173_ (.A1(_05518_),
    .A2(_18749_),
    .B(_05740_),
    .Y(_18839_));
 INVx1_ASAP7_75t_R _25174_ (.A(_01382_),
    .Y(_05741_));
 AO21x1_ASAP7_75t_R _25175_ (.A1(_05741_),
    .A2(_05522_),
    .B(_05540_),
    .Y(_05742_));
 OA21x2_ASAP7_75t_R _25176_ (.A1(_05517_),
    .A2(_18752_),
    .B(_05742_),
    .Y(_18841_));
 OR3x1_ASAP7_75t_R _25177_ (.A(_05320_),
    .B(_05521_),
    .C(_05536_),
    .Y(_05743_));
 OAI21x1_ASAP7_75t_R _25178_ (.A1(_05518_),
    .A2(_18758_),
    .B(_05743_),
    .Y(_18843_));
 INVx1_ASAP7_75t_R _25179_ (.A(_00168_),
    .Y(_17408_));
 INVx1_ASAP7_75t_R _25180_ (.A(_00185_),
    .Y(_17446_));
 INVx1_ASAP7_75t_R _25181_ (.A(_00191_),
    .Y(_17473_));
 INVx1_ASAP7_75t_R _25182_ (.A(_00199_),
    .Y(_18990_));
 INVx1_ASAP7_75t_R _25183_ (.A(_00202_),
    .Y(_17552_));
 INVx1_ASAP7_75t_R _25184_ (.A(_00204_),
    .Y(_17562_));
 INVx1_ASAP7_75t_R _25185_ (.A(_00225_),
    .Y(_17700_));
 INVx1_ASAP7_75t_R _25186_ (.A(_00226_),
    .Y(_17735_));
 AND2x2_ASAP7_75t_R _25187_ (.A(_02214_),
    .B(_05144_),
    .Y(_05744_));
 AOI21x1_ASAP7_75t_R _25188_ (.A1(_02216_),
    .A2(_05145_),
    .B(_05744_),
    .Y(_02352_));
 AND2x2_ASAP7_75t_R _25189_ (.A(_02213_),
    .B(_05144_),
    .Y(_05745_));
 AOI21x1_ASAP7_75t_R _25190_ (.A1(_02214_),
    .A2(_05145_),
    .B(_05745_),
    .Y(_02353_));
 NAND2x1_ASAP7_75t_R _25191_ (.A(_05157_),
    .B(_05158_),
    .Y(_05746_));
 OA21x2_ASAP7_75t_R _25192_ (.A1(_05139_),
    .A2(_05158_),
    .B(_05746_),
    .Y(_02354_));
 NAND2x1_ASAP7_75t_R _25193_ (.A(_05543_),
    .B(_05158_),
    .Y(_05747_));
 OA21x2_ASAP7_75t_R _25194_ (.A1(_05105_),
    .A2(_05158_),
    .B(_05747_),
    .Y(_02355_));
 NAND2x1_ASAP7_75t_R _25195_ (.A(_02218_),
    .B(_05158_),
    .Y(_05748_));
 OA21x2_ASAP7_75t_R _25196_ (.A1(_05133_),
    .A2(_05158_),
    .B(_05748_),
    .Y(_02356_));
 BUFx4f_ASAP7_75t_R _25197_ (.A(_02210_),
    .Y(_05749_));
 INVx2_ASAP7_75t_R _25198_ (.A(_05749_),
    .Y(_05750_));
 BUFx4f_ASAP7_75t_R _25199_ (.A(_00399_),
    .Y(_05751_));
 BUFx4f_ASAP7_75t_R _25200_ (.A(data_gnt_i),
    .Y(_05752_));
 AND2x2_ASAP7_75t_R _25201_ (.A(_01776_),
    .B(_04940_),
    .Y(_05753_));
 AND3x4_ASAP7_75t_R _25202_ (.A(_14026_),
    .B(_04928_),
    .C(_05753_),
    .Y(_05754_));
 AO21x2_ASAP7_75t_R _25203_ (.A1(_13359_),
    .A2(_05754_),
    .B(_13358_),
    .Y(_05755_));
 NAND3x2_ASAP7_75t_R _25204_ (.B(_05752_),
    .C(_05755_),
    .Y(_05756_),
    .A(_05751_));
 AND3x1_ASAP7_75t_R _25205_ (.A(_05751_),
    .B(_05752_),
    .C(_05755_),
    .Y(_05757_));
 BUFx3_ASAP7_75t_R _25206_ (.A(_05757_),
    .Y(_05758_));
 AND3x1_ASAP7_75t_R _25207_ (.A(_13635_),
    .B(_14026_),
    .C(_05758_),
    .Y(_05759_));
 AO21x1_ASAP7_75t_R _25208_ (.A1(_05750_),
    .A2(_05756_),
    .B(_05759_),
    .Y(_02357_));
 INVx1_ASAP7_75t_R _25209_ (.A(_02215_),
    .Y(_05760_));
 AND2x4_ASAP7_75t_R _25210_ (.A(_13585_),
    .B(_14026_),
    .Y(_05761_));
 AND3x1_ASAP7_75t_R _25211_ (.A(_13561_),
    .B(_05758_),
    .C(_05761_),
    .Y(_05762_));
 AO21x1_ASAP7_75t_R _25212_ (.A1(_05760_),
    .A2(_05756_),
    .B(_05762_),
    .Y(_02358_));
 NAND2x2_ASAP7_75t_R _25213_ (.A(_18658_),
    .B(_18663_),
    .Y(_05763_));
 NAND2x2_ASAP7_75t_R _25214_ (.A(_05763_),
    .B(_05085_),
    .Y(_05764_));
 BUFx6f_ASAP7_75t_R _25215_ (.A(_05764_),
    .Y(_05765_));
 BUFx3_ASAP7_75t_R _25216_ (.A(_14307_),
    .Y(_05766_));
 NAND2x2_ASAP7_75t_R _25217_ (.A(_14070_),
    .B(_18632_),
    .Y(_05767_));
 OR4x2_ASAP7_75t_R _25218_ (.A(_14299_),
    .B(_18629_),
    .C(_05766_),
    .D(_05767_),
    .Y(_05768_));
 OR2x4_ASAP7_75t_R _25219_ (.A(_04993_),
    .B(_05768_),
    .Y(_05769_));
 OR3x2_ASAP7_75t_R _25220_ (.A(_05059_),
    .B(_05765_),
    .C(_05769_),
    .Y(_05770_));
 BUFx4f_ASAP7_75t_R _25221_ (.A(_02307_),
    .Y(_05771_));
 BUFx3_ASAP7_75t_R _25222_ (.A(_02309_),
    .Y(_05772_));
 BUFx4f_ASAP7_75t_R _25223_ (.A(_14736_),
    .Y(_05773_));
 AND2x2_ASAP7_75t_R _25224_ (.A(_18609_),
    .B(_05773_),
    .Y(_05774_));
 AO21x1_ASAP7_75t_R _25225_ (.A1(_05772_),
    .A2(_18611_),
    .B(_05774_),
    .Y(_05775_));
 AND4x1_ASAP7_75t_R _25226_ (.A(_05034_),
    .B(_04946_),
    .C(_04948_),
    .D(_02303_),
    .Y(_05776_));
 OAI21x1_ASAP7_75t_R _25227_ (.A1(_14300_),
    .A2(_04999_),
    .B(_05776_),
    .Y(_05777_));
 BUFx6f_ASAP7_75t_R _25228_ (.A(_05777_),
    .Y(_05778_));
 BUFx6f_ASAP7_75t_R _25229_ (.A(_05778_),
    .Y(_05779_));
 BUFx6f_ASAP7_75t_R _25230_ (.A(_05779_),
    .Y(_05780_));
 OR3x2_ASAP7_75t_R _25231_ (.A(_05034_),
    .B(_18852_),
    .C(_05766_),
    .Y(_05781_));
 BUFx6f_ASAP7_75t_R _25232_ (.A(_05781_),
    .Y(_05782_));
 BUFx6f_ASAP7_75t_R _25233_ (.A(_05782_),
    .Y(_05783_));
 BUFx6f_ASAP7_75t_R _25234_ (.A(_05783_),
    .Y(_05784_));
 OAI22x1_ASAP7_75t_R _25235_ (.A1(_00786_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_00787_),
    .Y(_05785_));
 INVx1_ASAP7_75t_R _25236_ (.A(_05030_),
    .Y(_05786_));
 OA21x2_ASAP7_75t_R _25237_ (.A1(_18623_),
    .A2(_05044_),
    .B(_04995_),
    .Y(_05787_));
 OA21x2_ASAP7_75t_R _25238_ (.A1(_04976_),
    .A2(_05787_),
    .B(_04975_),
    .Y(_05788_));
 OA21x2_ASAP7_75t_R _25239_ (.A1(_18623_),
    .A2(_04975_),
    .B(_05022_),
    .Y(_05789_));
 OA21x2_ASAP7_75t_R _25240_ (.A1(_04947_),
    .A2(_05788_),
    .B(_05789_),
    .Y(_05790_));
 OR2x2_ASAP7_75t_R _25241_ (.A(_05037_),
    .B(_05038_),
    .Y(_05791_));
 AND3x1_ASAP7_75t_R _25242_ (.A(_04949_),
    .B(_05022_),
    .C(_05042_),
    .Y(_05792_));
 AND2x2_ASAP7_75t_R _25243_ (.A(_05028_),
    .B(_05039_),
    .Y(_05793_));
 OA31x2_ASAP7_75t_R _25244_ (.A1(_05790_),
    .A2(_05791_),
    .A3(_05792_),
    .B1(_05793_),
    .Y(_05794_));
 AND2x2_ASAP7_75t_R _25245_ (.A(_05786_),
    .B(_05794_),
    .Y(_05795_));
 BUFx3_ASAP7_75t_R _25246_ (.A(_05795_),
    .Y(_05796_));
 OAI22x1_ASAP7_75t_R _25247_ (.A1(_02184_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_02121_),
    .Y(_05797_));
 AND2x2_ASAP7_75t_R _25248_ (.A(_05002_),
    .B(_05794_),
    .Y(_05798_));
 BUFx3_ASAP7_75t_R _25249_ (.A(_05798_),
    .Y(_05799_));
 AND3x4_ASAP7_75t_R _25250_ (.A(_18625_),
    .B(_04975_),
    .C(_04977_),
    .Y(_05800_));
 AND3x1_ASAP7_75t_R _25251_ (.A(_18629_),
    .B(_18658_),
    .C(_18663_),
    .Y(_05801_));
 AND5x2_ASAP7_75t_R _25252_ (.A(_05021_),
    .B(_05022_),
    .C(_05800_),
    .D(_05023_),
    .E(_05801_),
    .Y(_05802_));
 BUFx4f_ASAP7_75t_R _25253_ (.A(_05802_),
    .Y(_05803_));
 BUFx4f_ASAP7_75t_R _25254_ (.A(_05000_),
    .Y(_05804_));
 OR3x1_ASAP7_75t_R _25255_ (.A(_14308_),
    .B(_04987_),
    .C(_05804_),
    .Y(_05805_));
 NOR2x1_ASAP7_75t_R _25256_ (.A(_05034_),
    .B(_05805_),
    .Y(_05806_));
 INVx1_ASAP7_75t_R _25257_ (.A(_01984_),
    .Y(_05807_));
 OR3x1_ASAP7_75t_R _25258_ (.A(_04986_),
    .B(_05009_),
    .C(_05013_),
    .Y(_05808_));
 BUFx4f_ASAP7_75t_R _25259_ (.A(_05808_),
    .Y(_05809_));
 INVx3_ASAP7_75t_R _25260_ (.A(_05809_),
    .Y(_05810_));
 BUFx4f_ASAP7_75t_R _25261_ (.A(_05810_),
    .Y(_05811_));
 AO221x1_ASAP7_75t_R _25262_ (.A1(net107),
    .A2(_05803_),
    .B1(_05806_),
    .B2(_05807_),
    .C(_05811_),
    .Y(_05812_));
 OR4x1_ASAP7_75t_R _25263_ (.A(_14299_),
    .B(_14307_),
    .C(_04987_),
    .D(_05000_),
    .Y(_05813_));
 BUFx6f_ASAP7_75t_R _25264_ (.A(_05813_),
    .Y(_05814_));
 BUFx6f_ASAP7_75t_R _25265_ (.A(_05814_),
    .Y(_05815_));
 OR4x2_ASAP7_75t_R _25266_ (.A(_04948_),
    .B(_14307_),
    .C(_04986_),
    .D(_05000_),
    .Y(_05816_));
 BUFx6f_ASAP7_75t_R _25267_ (.A(_05816_),
    .Y(_05817_));
 OAI22x1_ASAP7_75t_R _25268_ (.A1(_01928_),
    .A2(_05815_),
    .B1(_05817_),
    .B2(_01849_),
    .Y(_05818_));
 OR5x1_ASAP7_75t_R _25269_ (.A(_14299_),
    .B(_18629_),
    .C(_14307_),
    .D(_05767_),
    .E(_04993_),
    .Y(_05819_));
 BUFx3_ASAP7_75t_R _25270_ (.A(_05819_),
    .Y(_05820_));
 BUFx10_ASAP7_75t_R _25271_ (.A(_05820_),
    .Y(_05821_));
 BUFx6f_ASAP7_75t_R _25272_ (.A(_05778_),
    .Y(_05822_));
 AND3x1_ASAP7_75t_R _25273_ (.A(_04948_),
    .B(_18627_),
    .C(_04982_),
    .Y(_05823_));
 OR4x2_ASAP7_75t_R _25274_ (.A(_04983_),
    .B(_05767_),
    .C(_04993_),
    .D(_05823_),
    .Y(_05824_));
 OAI22x1_ASAP7_75t_R _25275_ (.A1(_00788_),
    .A2(_05821_),
    .B1(_05822_),
    .B2(_05824_),
    .Y(_05825_));
 OR5x1_ASAP7_75t_R _25276_ (.A(_14299_),
    .B(_05766_),
    .C(_04952_),
    .D(_04984_),
    .E(_04969_),
    .Y(_05826_));
 BUFx6f_ASAP7_75t_R _25277_ (.A(_05826_),
    .Y(_05827_));
 OR5x2_ASAP7_75t_R _25278_ (.A(_04948_),
    .B(_14307_),
    .C(_04952_),
    .D(_04984_),
    .E(_04969_),
    .Y(_05828_));
 BUFx6f_ASAP7_75t_R _25279_ (.A(_05828_),
    .Y(_05829_));
 BUFx6f_ASAP7_75t_R _25280_ (.A(_05829_),
    .Y(_05830_));
 OAI22x1_ASAP7_75t_R _25281_ (.A1(_02081_),
    .A2(_05827_),
    .B1(_05830_),
    .B2(_02016_),
    .Y(_05831_));
 OR5x2_ASAP7_75t_R _25282_ (.A(_05034_),
    .B(_14307_),
    .C(_04952_),
    .D(_04984_),
    .E(_04969_),
    .Y(_05832_));
 BUFx6f_ASAP7_75t_R _25283_ (.A(_05832_),
    .Y(_05833_));
 BUFx6f_ASAP7_75t_R _25284_ (.A(_05833_),
    .Y(_05834_));
 OR4x2_ASAP7_75t_R _25285_ (.A(_04946_),
    .B(_14307_),
    .C(_04986_),
    .D(_05000_),
    .Y(_05835_));
 BUFx6f_ASAP7_75t_R _25286_ (.A(_05835_),
    .Y(_05836_));
 OAI22x1_ASAP7_75t_R _25287_ (.A1(_02048_),
    .A2(_05834_),
    .B1(_05836_),
    .B2(_01978_),
    .Y(_05837_));
 OR5x2_ASAP7_75t_R _25288_ (.A(_05812_),
    .B(_05818_),
    .C(_05825_),
    .D(_05831_),
    .E(_05837_),
    .Y(_05838_));
 AOI221x1_ASAP7_75t_R _25289_ (.A1(_05785_),
    .A2(_05796_),
    .B1(_05797_),
    .B2(_05799_),
    .C(_05838_),
    .Y(_05839_));
 AOI22x1_ASAP7_75t_R _25290_ (.A1(_05771_),
    .A2(_05775_),
    .B1(_05839_),
    .B2(_18611_),
    .Y(_05840_));
 BUFx6f_ASAP7_75t_R _25291_ (.A(_05840_),
    .Y(_05841_));
 NAND2x1_ASAP7_75t_R _25292_ (.A(_00788_),
    .B(_05770_),
    .Y(_05842_));
 OA21x2_ASAP7_75t_R _25293_ (.A1(_05770_),
    .A2(_05841_),
    .B(_05842_),
    .Y(_02359_));
 INVx1_ASAP7_75t_R _25294_ (.A(_02307_),
    .Y(_05843_));
 BUFx4f_ASAP7_75t_R _25295_ (.A(_05843_),
    .Y(_05844_));
 INVx1_ASAP7_75t_R _25296_ (.A(_02309_),
    .Y(_05845_));
 BUFx3_ASAP7_75t_R _25297_ (.A(_05845_),
    .Y(_05846_));
 NAND2x1_ASAP7_75t_R _25298_ (.A(_18861_),
    .B(_18618_),
    .Y(_05847_));
 OA21x2_ASAP7_75t_R _25299_ (.A1(_05846_),
    .A2(_18618_),
    .B(_05847_),
    .Y(_05848_));
 BUFx6f_ASAP7_75t_R _25300_ (.A(_05778_),
    .Y(_05849_));
 BUFx6f_ASAP7_75t_R _25301_ (.A(_05849_),
    .Y(_05850_));
 BUFx6f_ASAP7_75t_R _25302_ (.A(_05782_),
    .Y(_05851_));
 BUFx6f_ASAP7_75t_R _25303_ (.A(_05851_),
    .Y(_05852_));
 BUFx3_ASAP7_75t_R _25304_ (.A(_02119_),
    .Y(_05853_));
 OAI22x1_ASAP7_75t_R _25305_ (.A1(_02182_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_05853_),
    .Y(_05854_));
 OAI22x1_ASAP7_75t_R _25306_ (.A1(_02187_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_02124_),
    .Y(_05855_));
 OR5x2_ASAP7_75t_R _25307_ (.A(_04946_),
    .B(_14307_),
    .C(_04952_),
    .D(_04984_),
    .E(_04969_),
    .Y(_05856_));
 BUFx6f_ASAP7_75t_R _25308_ (.A(_05856_),
    .Y(_05857_));
 BUFx6f_ASAP7_75t_R _25309_ (.A(_05857_),
    .Y(_05858_));
 OA222x2_ASAP7_75t_R _25310_ (.A1(_01827_),
    .A2(_05817_),
    .B1(_05830_),
    .B2(_01994_),
    .C1(_05858_),
    .C2(_02054_),
    .Y(_05859_));
 INVx1_ASAP7_75t_R _25311_ (.A(_05859_),
    .Y(_05860_));
 OR3x1_ASAP7_75t_R _25312_ (.A(_05034_),
    .B(_01982_),
    .C(_05805_),
    .Y(_05861_));
 OAI21x1_ASAP7_75t_R _25313_ (.A1(_02026_),
    .A2(_05834_),
    .B(_05861_),
    .Y(_05862_));
 OAI22x1_ASAP7_75t_R _25314_ (.A1(_01906_),
    .A2(_05815_),
    .B1(_05827_),
    .B2(_01460_),
    .Y(_05863_));
 NOR2x1_ASAP7_75t_R _25315_ (.A(_01453_),
    .B(_05821_),
    .Y(_05864_));
 AO32x1_ASAP7_75t_R _25316_ (.A1(_05011_),
    .A2(_04999_),
    .A3(_05010_),
    .B1(_05803_),
    .B2(net129),
    .Y(_05865_));
 NOR2x1_ASAP7_75t_R _25317_ (.A(_01956_),
    .B(_05836_),
    .Y(_05866_));
 OR3x1_ASAP7_75t_R _25318_ (.A(_05864_),
    .B(_05865_),
    .C(_05866_),
    .Y(_05867_));
 NOR2x1_ASAP7_75t_R _25319_ (.A(_05824_),
    .B(_05782_),
    .Y(_05868_));
 OR5x1_ASAP7_75t_R _25320_ (.A(_05860_),
    .B(_05862_),
    .C(_05863_),
    .D(_05867_),
    .E(_05868_),
    .Y(_05869_));
 AO221x2_ASAP7_75t_R _25321_ (.A1(_05799_),
    .A2(_05854_),
    .B1(_05855_),
    .B2(_05796_),
    .C(_05869_),
    .Y(_05870_));
 OAI22x1_ASAP7_75t_R _25322_ (.A1(_05844_),
    .A2(_05848_),
    .B1(_05870_),
    .B2(_18618_),
    .Y(_05871_));
 CKINVDCx8_ASAP7_75t_R _25323_ (.A(_05871_),
    .Y(_05872_));
 NAND2x1_ASAP7_75t_R _25324_ (.A(_01453_),
    .B(_05770_),
    .Y(_05873_));
 OA21x2_ASAP7_75t_R _25325_ (.A1(_05770_),
    .A2(_05872_),
    .B(_05873_),
    .Y(_02360_));
 NAND2x2_ASAP7_75t_R _25326_ (.A(_18652_),
    .B(_04968_),
    .Y(_05874_));
 AND2x2_ASAP7_75t_R _25327_ (.A(_05029_),
    .B(_05030_),
    .Y(_05875_));
 AOI211x1_ASAP7_75t_R _25328_ (.A1(_05040_),
    .A2(_05051_),
    .B(_05874_),
    .C(_05875_),
    .Y(_05876_));
 NOR2x2_ASAP7_75t_R _25329_ (.A(_05059_),
    .B(_05765_),
    .Y(_05877_));
 OR3x1_ASAP7_75t_R _25330_ (.A(_18614_),
    .B(_18610_),
    .C(_05054_),
    .Y(_05878_));
 OR3x1_ASAP7_75t_R _25331_ (.A(_14300_),
    .B(_02305_),
    .C(_02304_),
    .Y(_05879_));
 AOI21x1_ASAP7_75t_R _25332_ (.A1(_14071_),
    .A2(_05878_),
    .B(_05879_),
    .Y(_05880_));
 AND3x1_ASAP7_75t_R _25333_ (.A(_05876_),
    .B(_05877_),
    .C(_05880_),
    .Y(_05881_));
 BUFx4f_ASAP7_75t_R _25334_ (.A(_05881_),
    .Y(_05882_));
 BUFx4f_ASAP7_75t_R _25335_ (.A(_05882_),
    .Y(_05883_));
 AO21x1_ASAP7_75t_R _25336_ (.A1(_05040_),
    .A2(_05051_),
    .B(_05874_),
    .Y(_05884_));
 AO21x1_ASAP7_75t_R _25337_ (.A1(_14071_),
    .A2(_05878_),
    .B(_05879_),
    .Y(_05885_));
 OR5x1_ASAP7_75t_R _25338_ (.A(_05875_),
    .B(_05884_),
    .C(_05058_),
    .D(_05764_),
    .E(_05885_),
    .Y(_05886_));
 BUFx4f_ASAP7_75t_R _25339_ (.A(_05886_),
    .Y(_05887_));
 NAND2x2_ASAP7_75t_R _25340_ (.A(_00788_),
    .B(_05887_),
    .Y(_05888_));
 AOI21x1_ASAP7_75t_R _25341_ (.A1(_05040_),
    .A2(_05051_),
    .B(_05874_),
    .Y(_05889_));
 NAND2x1_ASAP7_75t_R _25342_ (.A(_05786_),
    .B(_05889_),
    .Y(_05890_));
 OR4x2_ASAP7_75t_R _25343_ (.A(_05058_),
    .B(_05764_),
    .C(_05890_),
    .D(_05885_),
    .Y(_05891_));
 AND2x6_ASAP7_75t_R _25344_ (.A(_05888_),
    .B(_05891_),
    .Y(_05892_));
 BUFx4f_ASAP7_75t_R _25345_ (.A(_05892_),
    .Y(_05893_));
 AO21x1_ASAP7_75t_R _25346_ (.A1(_05841_),
    .A2(_05883_),
    .B(_05893_),
    .Y(_05894_));
 OR4x1_ASAP7_75t_R _25347_ (.A(_18654_),
    .B(_18658_),
    .C(_18663_),
    .D(_18851_),
    .Y(_05895_));
 BUFx4f_ASAP7_75t_R _25348_ (.A(_05895_),
    .Y(_05896_));
 OR2x2_ASAP7_75t_R _25349_ (.A(_05804_),
    .B(_05896_),
    .Y(_05897_));
 NOR3x1_ASAP7_75t_R _25350_ (.A(_14308_),
    .B(_04983_),
    .C(_05897_),
    .Y(_05898_));
 AND4x1_ASAP7_75t_R _25351_ (.A(_18665_),
    .B(_05028_),
    .C(_05015_),
    .D(_05018_),
    .Y(_05899_));
 NAND3x1_ASAP7_75t_R _25352_ (.A(_18663_),
    .B(_05022_),
    .C(_05023_),
    .Y(_05900_));
 OR3x1_ASAP7_75t_R _25353_ (.A(_18627_),
    .B(_18660_),
    .C(_04992_),
    .Y(_05901_));
 NOR2x1_ASAP7_75t_R _25354_ (.A(_05900_),
    .B(_05901_),
    .Y(_05902_));
 AND3x1_ASAP7_75t_R _25355_ (.A(_18652_),
    .B(_18665_),
    .C(_04968_),
    .Y(_05903_));
 AND5x1_ASAP7_75t_R _25356_ (.A(_04950_),
    .B(_05002_),
    .C(_04989_),
    .D(_05903_),
    .E(_05003_),
    .Y(_05904_));
 AO222x2_ASAP7_75t_R _25357_ (.A1(_05020_),
    .A2(_05899_),
    .B1(_05902_),
    .B2(_05800_),
    .C1(_05904_),
    .C2(_04999_),
    .Y(_05905_));
 OR5x1_ASAP7_75t_R _25358_ (.A(_18654_),
    .B(_18658_),
    .C(_18663_),
    .D(_18851_),
    .E(_04992_),
    .Y(_05906_));
 OR3x1_ASAP7_75t_R _25359_ (.A(_04983_),
    .B(_05767_),
    .C(_05906_),
    .Y(_05907_));
 NOR2x1_ASAP7_75t_R _25360_ (.A(_05823_),
    .B(_05907_),
    .Y(_05908_));
 AOI21x1_ASAP7_75t_R _25361_ (.A1(_04979_),
    .A2(_04985_),
    .B(_05896_),
    .Y(_05909_));
 NOR2x1_ASAP7_75t_R _25362_ (.A(_05009_),
    .B(_05896_),
    .Y(_05910_));
 AND2x2_ASAP7_75t_R _25363_ (.A(_05014_),
    .B(_05910_),
    .Y(_05911_));
 OR5x1_ASAP7_75t_R _25364_ (.A(_05898_),
    .B(_05905_),
    .C(_05908_),
    .D(_05909_),
    .E(_05911_),
    .Y(_05912_));
 AND4x2_ASAP7_75t_R _25365_ (.A(_18660_),
    .B(_05903_),
    .C(_05021_),
    .D(_05056_),
    .Y(_05913_));
 OA31x2_ASAP7_75t_R _25366_ (.A1(_05912_),
    .A2(_05913_),
    .A3(_05876_),
    .B1(_04971_),
    .Y(_05914_));
 AND2x4_ASAP7_75t_R _25367_ (.A(_05763_),
    .B(_05085_),
    .Y(_05915_));
 NAND2x2_ASAP7_75t_R _25368_ (.A(_05914_),
    .B(_05915_),
    .Y(_05916_));
 OR4x2_ASAP7_75t_R _25369_ (.A(_05875_),
    .B(_05884_),
    .C(_05916_),
    .D(_05885_),
    .Y(_05917_));
 BUFx4f_ASAP7_75t_R _25370_ (.A(_05917_),
    .Y(_05918_));
 NAND2x2_ASAP7_75t_R _25371_ (.A(_05888_),
    .B(_05891_),
    .Y(_05919_));
 OA211x2_ASAP7_75t_R _25372_ (.A1(_05841_),
    .A2(_05918_),
    .B(_05919_),
    .C(_00786_),
    .Y(_05920_));
 AO21x1_ASAP7_75t_R _25373_ (.A1(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .A2(_05894_),
    .B(_05920_),
    .Y(_02361_));
 BUFx4f_ASAP7_75t_R _25374_ (.A(_05917_),
    .Y(_05921_));
 BUFx6f_ASAP7_75t_R _25375_ (.A(_05921_),
    .Y(_05922_));
 OR3x1_ASAP7_75t_R _25376_ (.A(_02176_),
    .B(_02187_),
    .C(_02313_),
    .Y(_05923_));
 OR3x2_ASAP7_75t_R _25377_ (.A(_02154_),
    .B(_02165_),
    .C(_05923_),
    .Y(_05924_));
 OR5x1_ASAP7_75t_R _25378_ (.A(_02146_),
    .B(_02147_),
    .C(_02148_),
    .D(_02149_),
    .E(_05924_),
    .Y(_05925_));
 BUFx4f_ASAP7_75t_R _25379_ (.A(_05892_),
    .Y(_05926_));
 AO21x1_ASAP7_75t_R _25380_ (.A1(_05922_),
    .A2(_05925_),
    .B(_05926_),
    .Y(_05927_));
 OR2x4_ASAP7_75t_R _25381_ (.A(_02208_),
    .B(_05925_),
    .Y(_05928_));
 AND2x4_ASAP7_75t_R _25382_ (.A(_05002_),
    .B(_05889_),
    .Y(_05929_));
 BUFx4f_ASAP7_75t_R _25383_ (.A(_05929_),
    .Y(_05930_));
 BUFx3_ASAP7_75t_R _25384_ (.A(_02110_),
    .Y(_05931_));
 OAI22x1_ASAP7_75t_R _25385_ (.A1(_02173_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_05931_),
    .Y(_05932_));
 NAND2x2_ASAP7_75t_R _25386_ (.A(_05930_),
    .B(_05932_),
    .Y(_05933_));
 BUFx6f_ASAP7_75t_R _25387_ (.A(_05782_),
    .Y(_05934_));
 OA22x2_ASAP7_75t_R _25388_ (.A1(_02208_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02145_),
    .Y(_05935_));
 OR5x2_ASAP7_75t_R _25389_ (.A(_04948_),
    .B(_05766_),
    .C(_04952_),
    .D(_04984_),
    .E(_05005_),
    .Y(_05936_));
 BUFx6f_ASAP7_75t_R _25390_ (.A(_05936_),
    .Y(_05937_));
 BUFx4f_ASAP7_75t_R _25391_ (.A(_05025_),
    .Y(_05938_));
 NAND2x1_ASAP7_75t_R _25392_ (.A(net108),
    .B(_05938_),
    .Y(_05939_));
 OA211x2_ASAP7_75t_R _25393_ (.A1(_01467_),
    .A2(_05809_),
    .B(_05939_),
    .C(_05769_),
    .Y(_05940_));
 BUFx6f_ASAP7_75t_R _25394_ (.A(_05814_),
    .Y(_05941_));
 OR5x2_ASAP7_75t_R _25395_ (.A(_04946_),
    .B(_05766_),
    .C(_04952_),
    .D(_04984_),
    .E(_05005_),
    .Y(_05942_));
 BUFx6f_ASAP7_75t_R _25396_ (.A(_05942_),
    .Y(_05943_));
 OR4x2_ASAP7_75t_R _25397_ (.A(_04948_),
    .B(_05766_),
    .C(_04987_),
    .D(_05804_),
    .Y(_05944_));
 BUFx6f_ASAP7_75t_R _25398_ (.A(_05944_),
    .Y(_05945_));
 OA222x2_ASAP7_75t_R _25399_ (.A1(_01927_),
    .A2(_05941_),
    .B1(_05943_),
    .B2(_02074_),
    .C1(_05945_),
    .C2(_01848_),
    .Y(_05946_));
 OA211x2_ASAP7_75t_R _25400_ (.A1(_02015_),
    .A2(_05937_),
    .B(_05940_),
    .C(_05946_),
    .Y(_05947_));
 OR5x2_ASAP7_75t_R _25401_ (.A(_05034_),
    .B(_05766_),
    .C(_04952_),
    .D(_04984_),
    .E(_05005_),
    .Y(_05948_));
 BUFx6f_ASAP7_75t_R _25402_ (.A(_05948_),
    .Y(_05949_));
 OR4x2_ASAP7_75t_R _25403_ (.A(_04946_),
    .B(_14308_),
    .C(_04987_),
    .D(_05804_),
    .Y(_05950_));
 BUFx6f_ASAP7_75t_R _25404_ (.A(_05950_),
    .Y(_05951_));
 OA22x2_ASAP7_75t_R _25405_ (.A1(_02047_),
    .A2(_05949_),
    .B1(_05951_),
    .B2(_01977_),
    .Y(_05952_));
 OA211x2_ASAP7_75t_R _25406_ (.A1(_05890_),
    .A2(_05935_),
    .B(_05947_),
    .C(_05952_),
    .Y(_05953_));
 AND2x2_ASAP7_75t_R _25407_ (.A(_18861_),
    .B(_18657_),
    .Y(_05954_));
 AO21x1_ASAP7_75t_R _25408_ (.A1(_05772_),
    .A2(_18659_),
    .B(_05954_),
    .Y(_05955_));
 AO32x2_ASAP7_75t_R _25409_ (.A1(_18659_),
    .A2(_05933_),
    .A3(_05953_),
    .B1(_05955_),
    .B2(_05771_),
    .Y(_05956_));
 NAND2x1_ASAP7_75t_R _25410_ (.A(_05883_),
    .B(_05956_),
    .Y(_05957_));
 OAI21x1_ASAP7_75t_R _25411_ (.A1(_05883_),
    .A2(_05928_),
    .B(_05957_),
    .Y(_05958_));
 BUFx6f_ASAP7_75t_R _25412_ (.A(_05919_),
    .Y(_05959_));
 AOI22x1_ASAP7_75t_R _25413_ (.A1(_02208_),
    .A2(_05927_),
    .B1(_05958_),
    .B2(_05959_),
    .Y(_02362_));
 BUFx4f_ASAP7_75t_R _25414_ (.A(_02207_),
    .Y(_05960_));
 OR3x1_ASAP7_75t_R _25415_ (.A(_00786_),
    .B(_02187_),
    .C(_02198_),
    .Y(_05961_));
 OR3x1_ASAP7_75t_R _25416_ (.A(_02165_),
    .B(_02176_),
    .C(_05961_),
    .Y(_05962_));
 OR3x2_ASAP7_75t_R _25417_ (.A(_02149_),
    .B(_02154_),
    .C(_05962_),
    .Y(_05963_));
 OR3x2_ASAP7_75t_R _25418_ (.A(_02147_),
    .B(_02148_),
    .C(_05963_),
    .Y(_05964_));
 OR3x4_ASAP7_75t_R _25419_ (.A(_02146_),
    .B(_02208_),
    .C(_05964_),
    .Y(_05965_));
 AO21x1_ASAP7_75t_R _25420_ (.A1(_05922_),
    .A2(_05965_),
    .B(_05926_),
    .Y(_05966_));
 INVx1_ASAP7_75t_R _25421_ (.A(_05960_),
    .Y(_05967_));
 AND4x1_ASAP7_75t_R _25422_ (.A(_05876_),
    .B(_05914_),
    .C(_05915_),
    .D(_05880_),
    .Y(_05968_));
 BUFx4f_ASAP7_75t_R _25423_ (.A(_05968_),
    .Y(_05969_));
 BUFx6f_ASAP7_75t_R _25424_ (.A(_05969_),
    .Y(_05970_));
 NOR2x1_ASAP7_75t_R _25425_ (.A(_05970_),
    .B(_05965_),
    .Y(_05971_));
 AND2x2_ASAP7_75t_R _25426_ (.A(_05773_),
    .B(_18662_),
    .Y(_05972_));
 AO21x1_ASAP7_75t_R _25427_ (.A1(_05772_),
    .A2(_18664_),
    .B(_05972_),
    .Y(_05973_));
 NAND2x2_ASAP7_75t_R _25428_ (.A(_05002_),
    .B(_05889_),
    .Y(_05974_));
 OA22x2_ASAP7_75t_R _25429_ (.A1(_02172_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02109_),
    .Y(_05975_));
 AOI211x1_ASAP7_75t_R _25430_ (.A1(_05040_),
    .A2(_05051_),
    .B(_05874_),
    .C(_05030_),
    .Y(_05976_));
 OAI22x1_ASAP7_75t_R _25431_ (.A1(_05960_),
    .A2(_05779_),
    .B1(_05934_),
    .B2(_02144_),
    .Y(_05977_));
 NAND2x1_ASAP7_75t_R _25432_ (.A(_05976_),
    .B(_05977_),
    .Y(_05978_));
 OR4x1_ASAP7_75t_R _25433_ (.A(_04948_),
    .B(_14307_),
    .C(_05804_),
    .D(_05896_),
    .Y(_05979_));
 BUFx6f_ASAP7_75t_R _25434_ (.A(_05979_),
    .Y(_05980_));
 OA222x2_ASAP7_75t_R _25435_ (.A1(_02046_),
    .A2(_05834_),
    .B1(_05858_),
    .B2(_02073_),
    .C1(_05980_),
    .C2(_01847_),
    .Y(_05981_));
 OR4x1_ASAP7_75t_R _25436_ (.A(_14300_),
    .B(_14308_),
    .C(_05804_),
    .D(_05896_),
    .Y(_05982_));
 BUFx4f_ASAP7_75t_R _25437_ (.A(_05982_),
    .Y(_05983_));
 OA22x2_ASAP7_75t_R _25438_ (.A1(_02014_),
    .A2(_05830_),
    .B1(_05983_),
    .B2(_01926_),
    .Y(_05984_));
 OR4x2_ASAP7_75t_R _25439_ (.A(_04946_),
    .B(_05766_),
    .C(_05804_),
    .D(_05896_),
    .Y(_05985_));
 OA22x2_ASAP7_75t_R _25440_ (.A1(_02080_),
    .A2(_05827_),
    .B1(_05985_),
    .B2(_01976_),
    .Y(_05986_));
 OR3x4_ASAP7_75t_R _25441_ (.A(_05009_),
    .B(_05013_),
    .C(_05896_),
    .Y(_05987_));
 INVx1_ASAP7_75t_R _25442_ (.A(net109),
    .Y(_05988_));
 OR3x4_ASAP7_75t_R _25443_ (.A(_04978_),
    .B(_05900_),
    .C(_05901_),
    .Y(_05989_));
 NAND2x1_ASAP7_75t_R _25444_ (.A(_18625_),
    .B(_04975_),
    .Y(_05990_));
 OR5x2_ASAP7_75t_R _25445_ (.A(_14300_),
    .B(_04966_),
    .C(_05990_),
    .D(_05009_),
    .E(_05896_),
    .Y(_05991_));
 OR3x4_ASAP7_75t_R _25446_ (.A(_04978_),
    .B(_05804_),
    .C(_05896_),
    .Y(_05992_));
 OA222x2_ASAP7_75t_R _25447_ (.A1(_05988_),
    .A2(_05989_),
    .B1(_05991_),
    .B2(_01940_),
    .C1(_05992_),
    .C2(_05369_),
    .Y(_05993_));
 OR4x2_ASAP7_75t_R _25448_ (.A(_14300_),
    .B(_05766_),
    .C(_05009_),
    .D(_05896_),
    .Y(_05994_));
 OR5x2_ASAP7_75t_R _25449_ (.A(_14300_),
    .B(_18629_),
    .C(_05766_),
    .D(_05767_),
    .E(_05906_),
    .Y(_05995_));
 OA21x2_ASAP7_75t_R _25450_ (.A1(_01853_),
    .A2(_05994_),
    .B(_05995_),
    .Y(_05996_));
 OA211x2_ASAP7_75t_R _25451_ (.A1(_00785_),
    .A2(_05987_),
    .B(_05993_),
    .C(_05996_),
    .Y(_05997_));
 AND4x1_ASAP7_75t_R _25452_ (.A(_05981_),
    .B(_05984_),
    .C(_05986_),
    .D(_05997_),
    .Y(_05998_));
 OA211x2_ASAP7_75t_R _25453_ (.A1(_05974_),
    .A2(_05975_),
    .B(_05978_),
    .C(_05998_),
    .Y(_05999_));
 AO22x2_ASAP7_75t_R _25454_ (.A1(_05771_),
    .A2(_05973_),
    .B1(_05999_),
    .B2(_18664_),
    .Y(_06000_));
 AO22x1_ASAP7_75t_R _25455_ (.A1(_05967_),
    .A2(_05971_),
    .B1(_06000_),
    .B2(_05883_),
    .Y(_06001_));
 AOI22x1_ASAP7_75t_R _25456_ (.A1(_05960_),
    .A2(_05966_),
    .B1(_06001_),
    .B2(_05959_),
    .Y(_02363_));
 BUFx6f_ASAP7_75t_R _25457_ (.A(_05892_),
    .Y(_06002_));
 AND2x2_ASAP7_75t_R _25458_ (.A(_18667_),
    .B(_05773_),
    .Y(_06003_));
 AO21x1_ASAP7_75t_R _25459_ (.A1(_05772_),
    .A2(_18669_),
    .B(_06003_),
    .Y(_06004_));
 OAI22x1_ASAP7_75t_R _25460_ (.A1(_02171_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_02108_),
    .Y(_06005_));
 OAI22x1_ASAP7_75t_R _25461_ (.A1(_02206_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_02143_),
    .Y(_06006_));
 BUFx4f_ASAP7_75t_R _25462_ (.A(_05976_),
    .Y(_06007_));
 OA222x2_ASAP7_75t_R _25463_ (.A1(_00783_),
    .A2(_05827_),
    .B1(_05985_),
    .B2(_01975_),
    .C1(_05980_),
    .C2(_01846_),
    .Y(_06008_));
 INVx1_ASAP7_75t_R _25464_ (.A(_06008_),
    .Y(_06009_));
 OAI22x1_ASAP7_75t_R _25465_ (.A1(_02013_),
    .A2(_05830_),
    .B1(_05994_),
    .B2(_01852_),
    .Y(_06010_));
 OAI22x1_ASAP7_75t_R _25466_ (.A1(_01925_),
    .A2(_05983_),
    .B1(_05858_),
    .B2(_02072_),
    .Y(_06011_));
 INVx1_ASAP7_75t_R _25467_ (.A(net110),
    .Y(_06012_));
 OA222x2_ASAP7_75t_R _25468_ (.A1(_06012_),
    .A2(_05989_),
    .B1(_05833_),
    .B2(_02045_),
    .C1(_05987_),
    .C2(_00784_),
    .Y(_06013_));
 INVx1_ASAP7_75t_R _25469_ (.A(_06013_),
    .Y(_06014_));
 OR5x2_ASAP7_75t_R _25470_ (.A(_05913_),
    .B(_06009_),
    .C(_06010_),
    .D(_06011_),
    .E(_06014_),
    .Y(_06015_));
 AOI221x1_ASAP7_75t_R _25471_ (.A1(_05930_),
    .A2(_06005_),
    .B1(_06006_),
    .B2(_06007_),
    .C(_06015_),
    .Y(_06016_));
 AO22x2_ASAP7_75t_R _25472_ (.A1(_05771_),
    .A2(_06004_),
    .B1(_06016_),
    .B2(_18669_),
    .Y(_06017_));
 INVx1_ASAP7_75t_R _25473_ (.A(_02206_),
    .Y(_06018_));
 OR4x1_ASAP7_75t_R _25474_ (.A(_06018_),
    .B(_05960_),
    .C(_05970_),
    .D(_05928_),
    .Y(_06019_));
 OA21x2_ASAP7_75t_R _25475_ (.A1(_05922_),
    .A2(_06017_),
    .B(_06019_),
    .Y(_06020_));
 BUFx6f_ASAP7_75t_R _25476_ (.A(_05887_),
    .Y(_06021_));
 OAI21x1_ASAP7_75t_R _25477_ (.A1(_05960_),
    .A2(_05928_),
    .B(_06021_),
    .Y(_06022_));
 AO21x1_ASAP7_75t_R _25478_ (.A1(_05919_),
    .A2(_06022_),
    .B(_02206_),
    .Y(_06023_));
 OAI21x1_ASAP7_75t_R _25479_ (.A1(_06002_),
    .A2(_06020_),
    .B(_06023_),
    .Y(_02364_));
 INVx1_ASAP7_75t_R _25480_ (.A(_02205_),
    .Y(_06024_));
 BUFx4f_ASAP7_75t_R _25481_ (.A(_05921_),
    .Y(_06025_));
 OR3x1_ASAP7_75t_R _25482_ (.A(_02206_),
    .B(_05960_),
    .C(_05965_),
    .Y(_06026_));
 AO21x1_ASAP7_75t_R _25483_ (.A1(_06025_),
    .A2(_06026_),
    .B(_05893_),
    .Y(_06027_));
 NOR2x1_ASAP7_75t_R _25484_ (.A(_02206_),
    .B(_05960_),
    .Y(_06028_));
 NAND2x1_ASAP7_75t_R _25485_ (.A(_18861_),
    .B(_18672_),
    .Y(_06029_));
 OA21x2_ASAP7_75t_R _25486_ (.A1(_05846_),
    .A2(_18672_),
    .B(_06029_),
    .Y(_06030_));
 OAI22x1_ASAP7_75t_R _25487_ (.A1(_02205_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_02142_),
    .Y(_06031_));
 OAI22x1_ASAP7_75t_R _25488_ (.A1(_02170_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_02107_),
    .Y(_06032_));
 OA222x2_ASAP7_75t_R _25489_ (.A1(_01845_),
    .A2(_05817_),
    .B1(_05827_),
    .B2(_02079_),
    .C1(_05829_),
    .C2(_02012_),
    .Y(_06033_));
 INVx1_ASAP7_75t_R _25490_ (.A(_06033_),
    .Y(_06034_));
 NOR2x1_ASAP7_75t_R _25491_ (.A(_02044_),
    .B(_05834_),
    .Y(_06035_));
 INVx1_ASAP7_75t_R _25492_ (.A(_01468_),
    .Y(_06036_));
 AO22x1_ASAP7_75t_R _25493_ (.A1(net111),
    .A2(_05803_),
    .B1(_05811_),
    .B2(_06036_),
    .Y(_06037_));
 OAI22x1_ASAP7_75t_R _25494_ (.A1(_01924_),
    .A2(_05815_),
    .B1(_05836_),
    .B2(_01974_),
    .Y(_06038_));
 OAI21x1_ASAP7_75t_R _25495_ (.A1(_02071_),
    .A2(_05858_),
    .B(_05821_),
    .Y(_06039_));
 OR5x2_ASAP7_75t_R _25496_ (.A(_06034_),
    .B(_06035_),
    .C(_06037_),
    .D(_06038_),
    .E(_06039_),
    .Y(_06040_));
 AO221x2_ASAP7_75t_R _25497_ (.A1(_05796_),
    .A2(_06031_),
    .B1(_06032_),
    .B2(_05799_),
    .C(_06040_),
    .Y(_06041_));
 OA22x2_ASAP7_75t_R _25498_ (.A1(_05844_),
    .A2(_06030_),
    .B1(_06041_),
    .B2(_18672_),
    .Y(_06042_));
 BUFx4f_ASAP7_75t_R _25499_ (.A(_05969_),
    .Y(_06043_));
 AO32x1_ASAP7_75t_R _25500_ (.A1(_02205_),
    .A2(_05971_),
    .A3(_06028_),
    .B1(_06042_),
    .B2(_06043_),
    .Y(_06044_));
 BUFx3_ASAP7_75t_R _25501_ (.A(_05919_),
    .Y(_06045_));
 AO22x1_ASAP7_75t_R _25502_ (.A1(_06024_),
    .A2(_06027_),
    .B1(_06044_),
    .B2(_06045_),
    .Y(_02365_));
 BUFx3_ASAP7_75t_R _25503_ (.A(_02204_),
    .Y(_06046_));
 BUFx4f_ASAP7_75t_R _25504_ (.A(_05969_),
    .Y(_06047_));
 OR3x4_ASAP7_75t_R _25505_ (.A(_02205_),
    .B(_02206_),
    .C(_05960_),
    .Y(_06048_));
 NOR2x1_ASAP7_75t_R _25506_ (.A(_05928_),
    .B(_06048_),
    .Y(_06049_));
 OA21x2_ASAP7_75t_R _25507_ (.A1(_06047_),
    .A2(_06049_),
    .B(_05919_),
    .Y(_06050_));
 NAND2x1_ASAP7_75t_R _25508_ (.A(_05773_),
    .B(_18680_),
    .Y(_06051_));
 OA21x2_ASAP7_75t_R _25509_ (.A1(_05845_),
    .A2(_18680_),
    .B(_06051_),
    .Y(_06052_));
 OAI22x1_ASAP7_75t_R _25510_ (.A1(_06046_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_02141_),
    .Y(_06053_));
 OAI22x1_ASAP7_75t_R _25511_ (.A1(_02169_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_02106_),
    .Y(_06054_));
 OAI22x1_ASAP7_75t_R _25512_ (.A1(_02043_),
    .A2(_05834_),
    .B1(_05858_),
    .B2(_02070_),
    .Y(_06055_));
 OAI22x1_ASAP7_75t_R _25513_ (.A1(_01844_),
    .A2(_05817_),
    .B1(_05830_),
    .B2(_02011_),
    .Y(_06056_));
 INVx1_ASAP7_75t_R _25514_ (.A(_05835_),
    .Y(_06057_));
 INVx1_ASAP7_75t_R _25515_ (.A(_01973_),
    .Y(_06058_));
 INVx1_ASAP7_75t_R _25516_ (.A(_01469_),
    .Y(_06059_));
 AO222x2_ASAP7_75t_R _25517_ (.A1(net112),
    .A2(_05803_),
    .B1(_06057_),
    .B2(_06058_),
    .C1(_05810_),
    .C2(_06059_),
    .Y(_06060_));
 OAI21x1_ASAP7_75t_R _25518_ (.A1(_01923_),
    .A2(_05941_),
    .B(_05821_),
    .Y(_06061_));
 OR4x2_ASAP7_75t_R _25519_ (.A(_06055_),
    .B(_06056_),
    .C(_06060_),
    .D(_06061_),
    .Y(_06062_));
 AO221x2_ASAP7_75t_R _25520_ (.A1(_05796_),
    .A2(_06053_),
    .B1(_06054_),
    .B2(_05799_),
    .C(_06062_),
    .Y(_06063_));
 OA22x2_ASAP7_75t_R _25521_ (.A1(_05843_),
    .A2(_06052_),
    .B1(_06063_),
    .B2(_18680_),
    .Y(_06064_));
 BUFx10_ASAP7_75t_R _25522_ (.A(_06064_),
    .Y(_06065_));
 AND3x1_ASAP7_75t_R _25523_ (.A(_06046_),
    .B(_05918_),
    .C(_06049_),
    .Y(_06066_));
 AOI21x1_ASAP7_75t_R _25524_ (.A1(_06047_),
    .A2(_06065_),
    .B(_06066_),
    .Y(_06067_));
 OAI22x1_ASAP7_75t_R _25525_ (.A1(_06046_),
    .A2(_06050_),
    .B1(_06067_),
    .B2(_06002_),
    .Y(_02366_));
 INVx1_ASAP7_75t_R _25526_ (.A(_02203_),
    .Y(_06068_));
 OR3x1_ASAP7_75t_R _25527_ (.A(_06046_),
    .B(_05965_),
    .C(_06048_),
    .Y(_06069_));
 AO21x1_ASAP7_75t_R _25528_ (.A1(_06025_),
    .A2(_06069_),
    .B(_05893_),
    .Y(_06070_));
 NOR2x1_ASAP7_75t_R _25529_ (.A(_06046_),
    .B(_06048_),
    .Y(_06071_));
 BUFx3_ASAP7_75t_R _25530_ (.A(_05843_),
    .Y(_06072_));
 BUFx3_ASAP7_75t_R _25531_ (.A(_05845_),
    .Y(_06073_));
 BUFx6f_ASAP7_75t_R _25532_ (.A(_14736_),
    .Y(_06074_));
 NAND2x1_ASAP7_75t_R _25533_ (.A(_06074_),
    .B(_18685_),
    .Y(_06075_));
 OA21x2_ASAP7_75t_R _25534_ (.A1(_06073_),
    .A2(_18685_),
    .B(_06075_),
    .Y(_06076_));
 OAI22x1_ASAP7_75t_R _25535_ (.A1(_02203_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_02140_),
    .Y(_06077_));
 OAI22x1_ASAP7_75t_R _25536_ (.A1(_02168_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_02105_),
    .Y(_06078_));
 OA222x2_ASAP7_75t_R _25537_ (.A1(_01843_),
    .A2(_05817_),
    .B1(_05836_),
    .B2(_01972_),
    .C1(_05827_),
    .C2(_00790_),
    .Y(_06079_));
 INVx1_ASAP7_75t_R _25538_ (.A(_06079_),
    .Y(_06080_));
 NOR2x1_ASAP7_75t_R _25539_ (.A(_02042_),
    .B(_05833_),
    .Y(_06081_));
 INVx1_ASAP7_75t_R _25540_ (.A(_01470_),
    .Y(_06082_));
 AO22x1_ASAP7_75t_R _25541_ (.A1(net113),
    .A2(_05803_),
    .B1(_05811_),
    .B2(_06082_),
    .Y(_06083_));
 OAI22x1_ASAP7_75t_R _25542_ (.A1(_01922_),
    .A2(_05941_),
    .B1(_05857_),
    .B2(_02069_),
    .Y(_06084_));
 OAI21x1_ASAP7_75t_R _25543_ (.A1(_02010_),
    .A2(_05829_),
    .B(_05821_),
    .Y(_06085_));
 OR5x2_ASAP7_75t_R _25544_ (.A(_06080_),
    .B(_06081_),
    .C(_06083_),
    .D(_06084_),
    .E(_06085_),
    .Y(_06086_));
 AO221x2_ASAP7_75t_R _25545_ (.A1(_05796_),
    .A2(_06077_),
    .B1(_06078_),
    .B2(_05799_),
    .C(_06086_),
    .Y(_06087_));
 OA22x2_ASAP7_75t_R _25546_ (.A1(_06072_),
    .A2(_06076_),
    .B1(_06087_),
    .B2(_18685_),
    .Y(_06088_));
 AO32x1_ASAP7_75t_R _25547_ (.A1(_02203_),
    .A2(_05971_),
    .A3(_06071_),
    .B1(_06088_),
    .B2(_06043_),
    .Y(_06089_));
 AO22x1_ASAP7_75t_R _25548_ (.A1(_06068_),
    .A2(_06070_),
    .B1(_06089_),
    .B2(_06045_),
    .Y(_02367_));
 INVx1_ASAP7_75t_R _25549_ (.A(_02202_),
    .Y(_06090_));
 OR4x1_ASAP7_75t_R _25550_ (.A(_02203_),
    .B(_06046_),
    .C(_05928_),
    .D(_06048_),
    .Y(_06091_));
 AO21x1_ASAP7_75t_R _25551_ (.A1(_06025_),
    .A2(_06091_),
    .B(_05893_),
    .Y(_06092_));
 BUFx6f_ASAP7_75t_R _25552_ (.A(_05921_),
    .Y(_06093_));
 NAND2x1_ASAP7_75t_R _25553_ (.A(_05773_),
    .B(_18687_),
    .Y(_06094_));
 OA21x2_ASAP7_75t_R _25554_ (.A1(_06073_),
    .A2(_18687_),
    .B(_06094_),
    .Y(_06095_));
 OAI22x1_ASAP7_75t_R _25555_ (.A1(_02202_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_02139_),
    .Y(_06096_));
 BUFx4f_ASAP7_75t_R _25556_ (.A(_02104_),
    .Y(_06097_));
 OAI22x1_ASAP7_75t_R _25557_ (.A1(_02167_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_06097_),
    .Y(_06098_));
 OA222x2_ASAP7_75t_R _25558_ (.A1(_01842_),
    .A2(_05816_),
    .B1(_05835_),
    .B2(_01971_),
    .C1(_05857_),
    .C2(_02068_),
    .Y(_06099_));
 INVx1_ASAP7_75t_R _25559_ (.A(_06099_),
    .Y(_06100_));
 OAI22x1_ASAP7_75t_R _25560_ (.A1(_02009_),
    .A2(_05829_),
    .B1(_05833_),
    .B2(_02041_),
    .Y(_06101_));
 OAI21x1_ASAP7_75t_R _25561_ (.A1(_01921_),
    .A2(_05941_),
    .B(_05821_),
    .Y(_06102_));
 NOR2x1_ASAP7_75t_R _25562_ (.A(_01471_),
    .B(_05809_),
    .Y(_06103_));
 AOI211x1_ASAP7_75t_R _25563_ (.A1(_14070_),
    .A2(_05009_),
    .B(_04978_),
    .C(_04987_),
    .Y(_06104_));
 BUFx4f_ASAP7_75t_R _25564_ (.A(_06104_),
    .Y(_06105_));
 NOR3x2_ASAP7_75t_R _25565_ (.B(_04978_),
    .C(_05804_),
    .Y(_06106_),
    .A(_04987_));
 AO222x2_ASAP7_75t_R _25566_ (.A1(net114),
    .A2(_05802_),
    .B1(_06105_),
    .B2(_05353_),
    .C1(_06106_),
    .C2(net179),
    .Y(_06107_));
 OR5x2_ASAP7_75t_R _25567_ (.A(_06100_),
    .B(_06101_),
    .C(_06102_),
    .D(_06103_),
    .E(_06107_),
    .Y(_06108_));
 AO221x2_ASAP7_75t_R _25568_ (.A1(_05795_),
    .A2(_06096_),
    .B1(_06098_),
    .B2(_05799_),
    .C(_06108_),
    .Y(_06109_));
 OA22x2_ASAP7_75t_R _25569_ (.A1(_06072_),
    .A2(_06095_),
    .B1(_06109_),
    .B2(_18687_),
    .Y(_06110_));
 BUFx10_ASAP7_75t_R _25570_ (.A(_06110_),
    .Y(_06111_));
 INVx4_ASAP7_75t_R _25571_ (.A(_06111_),
    .Y(_06112_));
 BUFx4f_ASAP7_75t_R _25572_ (.A(_05969_),
    .Y(_06113_));
 OR3x1_ASAP7_75t_R _25573_ (.A(_06090_),
    .B(_06113_),
    .C(_06091_),
    .Y(_06114_));
 OAI21x1_ASAP7_75t_R _25574_ (.A1(_06093_),
    .A2(_06112_),
    .B(_06114_),
    .Y(_06115_));
 AO22x1_ASAP7_75t_R _25575_ (.A1(_06090_),
    .A2(_06092_),
    .B1(_06115_),
    .B2(_06045_),
    .Y(_02368_));
 BUFx4f_ASAP7_75t_R _25576_ (.A(_05918_),
    .Y(_06116_));
 OR5x2_ASAP7_75t_R _25577_ (.A(_02202_),
    .B(_02203_),
    .C(_06046_),
    .D(_05965_),
    .E(_06048_),
    .Y(_06117_));
 AO21x1_ASAP7_75t_R _25578_ (.A1(_06116_),
    .A2(_06117_),
    .B(_05926_),
    .Y(_06118_));
 AND2x2_ASAP7_75t_R _25579_ (.A(_18861_),
    .B(_18692_),
    .Y(_06119_));
 AO21x1_ASAP7_75t_R _25580_ (.A1(_05772_),
    .A2(_18694_),
    .B(_06119_),
    .Y(_06120_));
 BUFx4f_ASAP7_75t_R _25581_ (.A(_02166_),
    .Y(_06121_));
 BUFx3_ASAP7_75t_R _25582_ (.A(_02103_),
    .Y(_06122_));
 OAI22x1_ASAP7_75t_R _25583_ (.A1(_06121_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_06122_),
    .Y(_06123_));
 BUFx4f_ASAP7_75t_R _25584_ (.A(_02138_),
    .Y(_06124_));
 OAI22x1_ASAP7_75t_R _25585_ (.A1(_02201_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_06124_),
    .Y(_06125_));
 OAI22x1_ASAP7_75t_R _25586_ (.A1(_02008_),
    .A2(_05830_),
    .B1(_05980_),
    .B2(_01841_),
    .Y(_06126_));
 OAI22x1_ASAP7_75t_R _25587_ (.A1(_01970_),
    .A2(_05985_),
    .B1(_05858_),
    .B2(_02067_),
    .Y(_06127_));
 INVx1_ASAP7_75t_R _25588_ (.A(net115),
    .Y(_06128_));
 INVx1_ASAP7_75t_R _25589_ (.A(net185),
    .Y(_06129_));
 OA222x2_ASAP7_75t_R _25590_ (.A1(_06128_),
    .A2(_05989_),
    .B1(_05991_),
    .B2(_01937_),
    .C1(_05992_),
    .C2(_06129_),
    .Y(_06130_));
 OAI21x1_ASAP7_75t_R _25591_ (.A1(_01472_),
    .A2(_05987_),
    .B(_06130_),
    .Y(_06131_));
 OAI21x1_ASAP7_75t_R _25592_ (.A1(_01854_),
    .A2(_05994_),
    .B(_05995_),
    .Y(_06132_));
 OAI22x1_ASAP7_75t_R _25593_ (.A1(_02040_),
    .A2(_05834_),
    .B1(_05983_),
    .B2(_01920_),
    .Y(_06133_));
 OR5x2_ASAP7_75t_R _25594_ (.A(_06126_),
    .B(_06127_),
    .C(_06131_),
    .D(_06132_),
    .E(_06133_),
    .Y(_06134_));
 AOI221x1_ASAP7_75t_R _25595_ (.A1(_05930_),
    .A2(_06123_),
    .B1(_06125_),
    .B2(_06007_),
    .C(_06134_),
    .Y(_06135_));
 AOI22x1_ASAP7_75t_R _25596_ (.A1(_05771_),
    .A2(_06120_),
    .B1(_06135_),
    .B2(_18694_),
    .Y(_06136_));
 BUFx10_ASAP7_75t_R _25597_ (.A(_06136_),
    .Y(_06137_));
 OR3x1_ASAP7_75t_R _25598_ (.A(_02201_),
    .B(_05882_),
    .C(_06117_),
    .Y(_06138_));
 OAI21x1_ASAP7_75t_R _25599_ (.A1(_06021_),
    .A2(_06137_),
    .B(_06138_),
    .Y(_06139_));
 AOI22x1_ASAP7_75t_R _25600_ (.A1(_02201_),
    .A2(_06118_),
    .B1(_06139_),
    .B2(_05959_),
    .Y(_02369_));
 OR3x4_ASAP7_75t_R _25601_ (.A(_02201_),
    .B(_02202_),
    .C(_06091_),
    .Y(_06140_));
 AOI21x1_ASAP7_75t_R _25602_ (.A1(_05922_),
    .A2(_06140_),
    .B(_06002_),
    .Y(_06141_));
 INVx1_ASAP7_75t_R _25603_ (.A(_02200_),
    .Y(_06142_));
 OR3x1_ASAP7_75t_R _25604_ (.A(_06142_),
    .B(_06113_),
    .C(_06140_),
    .Y(_06143_));
 BUFx4f_ASAP7_75t_R _25605_ (.A(_05969_),
    .Y(_06144_));
 NAND2x1_ASAP7_75t_R _25606_ (.A(_05773_),
    .B(_18697_),
    .Y(_06145_));
 OA21x2_ASAP7_75t_R _25607_ (.A1(_06073_),
    .A2(_18697_),
    .B(_06145_),
    .Y(_06146_));
 BUFx6f_ASAP7_75t_R _25608_ (.A(_05778_),
    .Y(_06147_));
 BUFx6f_ASAP7_75t_R _25609_ (.A(_05782_),
    .Y(_06148_));
 OAI22x1_ASAP7_75t_R _25610_ (.A1(_02164_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02101_),
    .Y(_06149_));
 OAI22x1_ASAP7_75t_R _25611_ (.A1(_02200_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_02137_),
    .Y(_06150_));
 NOR2x2_ASAP7_75t_R _25612_ (.A(_04993_),
    .B(_05768_),
    .Y(_06151_));
 INVx1_ASAP7_75t_R _25613_ (.A(_01473_),
    .Y(_06152_));
 AO22x1_ASAP7_75t_R _25614_ (.A1(net116),
    .A2(_05938_),
    .B1(_06105_),
    .B2(_05350_),
    .Y(_06153_));
 AO221x1_ASAP7_75t_R _25615_ (.A1(_06152_),
    .A2(_05811_),
    .B1(_06106_),
    .B2(net186),
    .C(_06153_),
    .Y(_06154_));
 OAI22x1_ASAP7_75t_R _25616_ (.A1(_02039_),
    .A2(_05949_),
    .B1(_05937_),
    .B2(_02007_),
    .Y(_06155_));
 OAI22x1_ASAP7_75t_R _25617_ (.A1(_01919_),
    .A2(_05815_),
    .B1(_05943_),
    .B2(_02066_),
    .Y(_06156_));
 OAI22x1_ASAP7_75t_R _25618_ (.A1(_01840_),
    .A2(_05945_),
    .B1(_05951_),
    .B2(_01969_),
    .Y(_06157_));
 OR5x2_ASAP7_75t_R _25619_ (.A(_06151_),
    .B(_06154_),
    .C(_06155_),
    .D(_06156_),
    .E(_06157_),
    .Y(_06158_));
 AO221x2_ASAP7_75t_R _25620_ (.A1(_05929_),
    .A2(_06149_),
    .B1(_06150_),
    .B2(_06007_),
    .C(_06158_),
    .Y(_06159_));
 OA22x2_ASAP7_75t_R _25621_ (.A1(_06072_),
    .A2(_06146_),
    .B1(_06159_),
    .B2(_18697_),
    .Y(_06160_));
 BUFx10_ASAP7_75t_R _25622_ (.A(_06160_),
    .Y(_06161_));
 NAND2x1_ASAP7_75t_R _25623_ (.A(_06144_),
    .B(_06161_),
    .Y(_06162_));
 AO21x1_ASAP7_75t_R _25624_ (.A1(_06143_),
    .A2(_06162_),
    .B(_06002_),
    .Y(_06163_));
 OAI21x1_ASAP7_75t_R _25625_ (.A1(_02200_),
    .A2(_06141_),
    .B(_06163_),
    .Y(_02370_));
 OR3x2_ASAP7_75t_R _25626_ (.A(_02200_),
    .B(_02201_),
    .C(_06117_),
    .Y(_06164_));
 AO21x1_ASAP7_75t_R _25627_ (.A1(_06116_),
    .A2(_06164_),
    .B(_05926_),
    .Y(_06165_));
 AND2x2_ASAP7_75t_R _25628_ (.A(_05773_),
    .B(_18702_),
    .Y(_06166_));
 AO21x1_ASAP7_75t_R _25629_ (.A1(_05772_),
    .A2(_18704_),
    .B(_06166_),
    .Y(_06167_));
 OA22x2_ASAP7_75t_R _25630_ (.A1(_02163_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02100_),
    .Y(_06168_));
 OAI22x1_ASAP7_75t_R _25631_ (.A1(_02199_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02136_),
    .Y(_06169_));
 NAND2x1_ASAP7_75t_R _25632_ (.A(_05976_),
    .B(_06169_),
    .Y(_06170_));
 NAND2x1_ASAP7_75t_R _25633_ (.A(net187),
    .B(_06106_),
    .Y(_06171_));
 AOI22x1_ASAP7_75t_R _25634_ (.A1(net117),
    .A2(_05938_),
    .B1(_06105_),
    .B2(_05349_),
    .Y(_06172_));
 OA211x2_ASAP7_75t_R _25635_ (.A1(_01474_),
    .A2(_05809_),
    .B(_06171_),
    .C(_06172_),
    .Y(_06173_));
 OA22x2_ASAP7_75t_R _25636_ (.A1(_02038_),
    .A2(_05949_),
    .B1(_05937_),
    .B2(_02006_),
    .Y(_06174_));
 OA22x2_ASAP7_75t_R _25637_ (.A1(_01839_),
    .A2(_05945_),
    .B1(_05943_),
    .B2(_02065_),
    .Y(_06175_));
 OA22x2_ASAP7_75t_R _25638_ (.A1(_01918_),
    .A2(_05941_),
    .B1(_05951_),
    .B2(_01968_),
    .Y(_06176_));
 AND5x2_ASAP7_75t_R _25639_ (.A(_05769_),
    .B(_06173_),
    .C(_06174_),
    .D(_06175_),
    .E(_06176_),
    .Y(_06177_));
 OA211x2_ASAP7_75t_R _25640_ (.A1(_05974_),
    .A2(_06168_),
    .B(_06170_),
    .C(_06177_),
    .Y(_06178_));
 AOI22x1_ASAP7_75t_R _25641_ (.A1(_05771_),
    .A2(_06167_),
    .B1(_06178_),
    .B2(_18704_),
    .Y(_06179_));
 BUFx10_ASAP7_75t_R _25642_ (.A(_06179_),
    .Y(_06180_));
 OR3x1_ASAP7_75t_R _25643_ (.A(_02199_),
    .B(_05882_),
    .C(_06164_),
    .Y(_06181_));
 OAI21x1_ASAP7_75t_R _25644_ (.A1(_06021_),
    .A2(_06180_),
    .B(_06181_),
    .Y(_06182_));
 AOI22x1_ASAP7_75t_R _25645_ (.A1(_02199_),
    .A2(_06165_),
    .B1(_06182_),
    .B2(_05959_),
    .Y(_02371_));
 OA22x2_ASAP7_75t_R _25646_ (.A1(_02183_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02120_),
    .Y(_06183_));
 OAI22x1_ASAP7_75t_R _25647_ (.A1(_02198_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02135_),
    .Y(_06184_));
 NAND2x1_ASAP7_75t_R _25648_ (.A(_05976_),
    .B(_06184_),
    .Y(_06185_));
 OR5x2_ASAP7_75t_R _25649_ (.A(_14300_),
    .B(_14308_),
    .C(_04952_),
    .D(_04984_),
    .E(_05005_),
    .Y(_06186_));
 OA22x2_ASAP7_75t_R _25650_ (.A1(_02005_),
    .A2(_05937_),
    .B1(_06186_),
    .B2(_02078_),
    .Y(_06187_));
 OA22x2_ASAP7_75t_R _25651_ (.A1(_01917_),
    .A2(_05815_),
    .B1(_05943_),
    .B2(_00789_),
    .Y(_06188_));
 OR4x2_ASAP7_75t_R _25652_ (.A(_05034_),
    .B(_14308_),
    .C(_04987_),
    .D(_05804_),
    .Y(_06189_));
 OA222x2_ASAP7_75t_R _25653_ (.A1(_01838_),
    .A2(_05945_),
    .B1(_06189_),
    .B2(_01983_),
    .C1(_05951_),
    .C2(_01967_),
    .Y(_06190_));
 NAND2x1_ASAP7_75t_R _25654_ (.A(net118),
    .B(_05938_),
    .Y(_06191_));
 OA21x2_ASAP7_75t_R _25655_ (.A1(_02037_),
    .A2(_05949_),
    .B(_06191_),
    .Y(_06192_));
 AND4x2_ASAP7_75t_R _25656_ (.A(_06187_),
    .B(_06188_),
    .C(_06190_),
    .D(_06192_),
    .Y(_06193_));
 OA211x2_ASAP7_75t_R _25657_ (.A1(_05974_),
    .A2(_06183_),
    .B(_06185_),
    .C(_06193_),
    .Y(_06194_));
 AND2x2_ASAP7_75t_R _25658_ (.A(_18613_),
    .B(_14736_),
    .Y(_06195_));
 AO21x1_ASAP7_75t_R _25659_ (.A1(_05772_),
    .A2(_18615_),
    .B(_06195_),
    .Y(_06196_));
 AND2x2_ASAP7_75t_R _25660_ (.A(_05771_),
    .B(_06196_),
    .Y(_06197_));
 AO21x2_ASAP7_75t_R _25661_ (.A1(_18615_),
    .A2(_06194_),
    .B(_06197_),
    .Y(_06198_));
 OR2x2_ASAP7_75t_R _25662_ (.A(_02314_),
    .B(_05970_),
    .Y(_06199_));
 OA211x2_ASAP7_75t_R _25663_ (.A1(_06093_),
    .A2(_06198_),
    .B(_06199_),
    .C(_05919_),
    .Y(_06200_));
 AOI21x1_ASAP7_75t_R _25664_ (.A1(_02198_),
    .A2(_06002_),
    .B(_06200_),
    .Y(_02372_));
 INVx1_ASAP7_75t_R _25665_ (.A(_02197_),
    .Y(_06201_));
 OR3x1_ASAP7_75t_R _25666_ (.A(_02199_),
    .B(_02200_),
    .C(_06140_),
    .Y(_06202_));
 AO21x1_ASAP7_75t_R _25667_ (.A1(_06025_),
    .A2(_06202_),
    .B(_05892_),
    .Y(_06203_));
 NAND2x1_ASAP7_75t_R _25668_ (.A(_18861_),
    .B(_18707_),
    .Y(_06204_));
 OA21x2_ASAP7_75t_R _25669_ (.A1(_05846_),
    .A2(_18707_),
    .B(_06204_),
    .Y(_06205_));
 OAI22x1_ASAP7_75t_R _25670_ (.A1(_02197_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_02134_),
    .Y(_06206_));
 BUFx3_ASAP7_75t_R _25671_ (.A(_02099_),
    .Y(_06207_));
 OAI22x1_ASAP7_75t_R _25672_ (.A1(_02162_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_06207_),
    .Y(_06208_));
 OAI22x1_ASAP7_75t_R _25673_ (.A1(_01837_),
    .A2(_05980_),
    .B1(_05858_),
    .B2(_02064_),
    .Y(_06209_));
 OAI22x1_ASAP7_75t_R _25674_ (.A1(_02036_),
    .A2(_05833_),
    .B1(_05985_),
    .B2(_01966_),
    .Y(_06210_));
 INVx1_ASAP7_75t_R _25675_ (.A(net119),
    .Y(_06211_));
 OA222x2_ASAP7_75t_R _25676_ (.A1(_06211_),
    .A2(_05989_),
    .B1(_05991_),
    .B2(_01934_),
    .C1(_05987_),
    .C2(_01475_),
    .Y(_06212_));
 OAI21x1_ASAP7_75t_R _25677_ (.A1(_05396_),
    .A2(_05992_),
    .B(_06212_),
    .Y(_06213_));
 OAI22x1_ASAP7_75t_R _25678_ (.A1(_02004_),
    .A2(_05830_),
    .B1(_05983_),
    .B2(_01916_),
    .Y(_06214_));
 OR5x2_ASAP7_75t_R _25679_ (.A(_05913_),
    .B(_06209_),
    .C(_06210_),
    .D(_06213_),
    .E(_06214_),
    .Y(_06215_));
 AO221x2_ASAP7_75t_R _25680_ (.A1(_05976_),
    .A2(_06206_),
    .B1(_06208_),
    .B2(_05929_),
    .C(_06215_),
    .Y(_06216_));
 OA22x2_ASAP7_75t_R _25681_ (.A1(_05844_),
    .A2(_06205_),
    .B1(_06216_),
    .B2(_18707_),
    .Y(_06217_));
 BUFx10_ASAP7_75t_R _25682_ (.A(_06217_),
    .Y(_06218_));
 INVx1_ASAP7_75t_R _25683_ (.A(_06202_),
    .Y(_06219_));
 AND3x1_ASAP7_75t_R _25684_ (.A(_02197_),
    .B(_05921_),
    .C(_06219_),
    .Y(_06220_));
 AO21x1_ASAP7_75t_R _25685_ (.A1(_06047_),
    .A2(_06218_),
    .B(_06220_),
    .Y(_06221_));
 AO22x1_ASAP7_75t_R _25686_ (.A1(_06201_),
    .A2(_06203_),
    .B1(_06221_),
    .B2(_06045_),
    .Y(_02373_));
 BUFx3_ASAP7_75t_R _25687_ (.A(_02196_),
    .Y(_06222_));
 INVx1_ASAP7_75t_R _25688_ (.A(_06222_),
    .Y(_06223_));
 OR3x2_ASAP7_75t_R _25689_ (.A(_02197_),
    .B(_02199_),
    .C(_06164_),
    .Y(_06224_));
 AO21x1_ASAP7_75t_R _25690_ (.A1(_06025_),
    .A2(_06224_),
    .B(_05892_),
    .Y(_06225_));
 NOR2x1_ASAP7_75t_R _25691_ (.A(_05970_),
    .B(_06224_),
    .Y(_06226_));
 NAND2x1_ASAP7_75t_R _25692_ (.A(_06074_),
    .B(_18715_),
    .Y(_06227_));
 OA21x2_ASAP7_75t_R _25693_ (.A1(_05846_),
    .A2(_18715_),
    .B(_06227_),
    .Y(_06228_));
 OAI22x1_ASAP7_75t_R _25694_ (.A1(_06222_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_02133_),
    .Y(_06229_));
 OAI22x1_ASAP7_75t_R _25695_ (.A1(_02161_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_02098_),
    .Y(_06230_));
 OAI22x1_ASAP7_75t_R _25696_ (.A1(_02035_),
    .A2(_05833_),
    .B1(_05857_),
    .B2(_02063_),
    .Y(_06231_));
 OAI22x1_ASAP7_75t_R _25697_ (.A1(_01836_),
    .A2(_05817_),
    .B1(_05836_),
    .B2(_01965_),
    .Y(_06232_));
 OAI22x1_ASAP7_75t_R _25698_ (.A1(_01915_),
    .A2(_05814_),
    .B1(_05829_),
    .B2(_02003_),
    .Y(_06233_));
 OR4x2_ASAP7_75t_R _25699_ (.A(_14300_),
    .B(_14308_),
    .C(_04987_),
    .D(_05009_),
    .Y(_06234_));
 OAI21x1_ASAP7_75t_R _25700_ (.A1(_01855_),
    .A2(_06234_),
    .B(_05820_),
    .Y(_06235_));
 OR4x1_ASAP7_75t_R _25701_ (.A(_06231_),
    .B(_06232_),
    .C(_06233_),
    .D(_06235_),
    .Y(_06236_));
 NOR2x1_ASAP7_75t_R _25702_ (.A(_01476_),
    .B(_05809_),
    .Y(_06237_));
 AO222x2_ASAP7_75t_R _25703_ (.A1(net120),
    .A2(_05803_),
    .B1(_06105_),
    .B2(_05346_),
    .C1(_06106_),
    .C2(net189),
    .Y(_06238_));
 OR3x4_ASAP7_75t_R _25704_ (.A(_06236_),
    .B(_06237_),
    .C(_06238_),
    .Y(_06239_));
 AO221x1_ASAP7_75t_R _25705_ (.A1(_05796_),
    .A2(_06229_),
    .B1(_06230_),
    .B2(_05799_),
    .C(_06239_),
    .Y(_06240_));
 OA22x2_ASAP7_75t_R _25706_ (.A1(_05844_),
    .A2(_06228_),
    .B1(_06240_),
    .B2(_18715_),
    .Y(_06241_));
 AO22x1_ASAP7_75t_R _25707_ (.A1(_06222_),
    .A2(_06226_),
    .B1(_06241_),
    .B2(_06043_),
    .Y(_06242_));
 AO22x1_ASAP7_75t_R _25708_ (.A1(_06223_),
    .A2(_06225_),
    .B1(_06242_),
    .B2(_06045_),
    .Y(_02374_));
 BUFx3_ASAP7_75t_R _25709_ (.A(_02195_),
    .Y(_06243_));
 OR3x1_ASAP7_75t_R _25710_ (.A(_06222_),
    .B(_02197_),
    .C(_06202_),
    .Y(_06244_));
 AO21x1_ASAP7_75t_R _25711_ (.A1(_06116_),
    .A2(_06244_),
    .B(_05926_),
    .Y(_06245_));
 AND2x2_ASAP7_75t_R _25712_ (.A(_06074_),
    .B(_18717_),
    .Y(_06246_));
 AO21x1_ASAP7_75t_R _25713_ (.A1(_05772_),
    .A2(_18719_),
    .B(_06246_),
    .Y(_06247_));
 OA22x2_ASAP7_75t_R _25714_ (.A1(_02160_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_02097_),
    .Y(_06248_));
 OAI22x1_ASAP7_75t_R _25715_ (.A1(_06243_),
    .A2(_05778_),
    .B1(_05851_),
    .B2(_02132_),
    .Y(_06249_));
 NAND2x1_ASAP7_75t_R _25716_ (.A(_05976_),
    .B(_06249_),
    .Y(_06250_));
 OR5x2_ASAP7_75t_R _25717_ (.A(_14300_),
    .B(_04966_),
    .C(_04987_),
    .D(_05990_),
    .E(_05009_),
    .Y(_06251_));
 OAI22x1_ASAP7_75t_R _25718_ (.A1(_01477_),
    .A2(_05809_),
    .B1(_06251_),
    .B2(_01932_),
    .Y(_06252_));
 AOI221x1_ASAP7_75t_R _25719_ (.A1(net121),
    .A2(_05938_),
    .B1(_06106_),
    .B2(net190),
    .C(_06252_),
    .Y(_06253_));
 OA22x2_ASAP7_75t_R _25720_ (.A1(_02034_),
    .A2(_05948_),
    .B1(_05945_),
    .B2(_01835_),
    .Y(_06254_));
 OA22x2_ASAP7_75t_R _25721_ (.A1(_01914_),
    .A2(_05814_),
    .B1(_05942_),
    .B2(_02062_),
    .Y(_06255_));
 OA22x2_ASAP7_75t_R _25722_ (.A1(_02002_),
    .A2(_05936_),
    .B1(_05950_),
    .B2(_01964_),
    .Y(_06256_));
 AND5x2_ASAP7_75t_R _25723_ (.A(_05769_),
    .B(_06253_),
    .C(_06254_),
    .D(_06255_),
    .E(_06256_),
    .Y(_06257_));
 OA211x2_ASAP7_75t_R _25724_ (.A1(_05974_),
    .A2(_06248_),
    .B(_06250_),
    .C(_06257_),
    .Y(_06258_));
 AOI22x1_ASAP7_75t_R _25725_ (.A1(_05771_),
    .A2(_06247_),
    .B1(_06258_),
    .B2(_18719_),
    .Y(_06259_));
 BUFx10_ASAP7_75t_R _25726_ (.A(_06259_),
    .Y(_06260_));
 OR3x1_ASAP7_75t_R _25727_ (.A(_06243_),
    .B(_05882_),
    .C(_06244_),
    .Y(_06261_));
 OAI21x1_ASAP7_75t_R _25728_ (.A1(_06021_),
    .A2(_06260_),
    .B(_06261_),
    .Y(_06262_));
 AOI22x1_ASAP7_75t_R _25729_ (.A1(_06243_),
    .A2(_06245_),
    .B1(_06262_),
    .B2(_05959_),
    .Y(_02375_));
 INVx1_ASAP7_75t_R _25730_ (.A(_02194_),
    .Y(_06263_));
 OR3x1_ASAP7_75t_R _25731_ (.A(_06243_),
    .B(_06222_),
    .C(_06224_),
    .Y(_06264_));
 AO21x1_ASAP7_75t_R _25732_ (.A1(_06025_),
    .A2(_06264_),
    .B(_05892_),
    .Y(_06265_));
 NOR2x1_ASAP7_75t_R _25733_ (.A(_06243_),
    .B(_06222_),
    .Y(_06266_));
 NAND2x1_ASAP7_75t_R _25734_ (.A(_06074_),
    .B(_18725_),
    .Y(_06267_));
 OA21x2_ASAP7_75t_R _25735_ (.A1(_06073_),
    .A2(_18725_),
    .B(_06267_),
    .Y(_06268_));
 OAI22x1_ASAP7_75t_R _25736_ (.A1(_02159_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02096_),
    .Y(_06269_));
 OAI22x1_ASAP7_75t_R _25737_ (.A1(_02194_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02131_),
    .Y(_06270_));
 AO22x1_ASAP7_75t_R _25738_ (.A1(net122),
    .A2(_05938_),
    .B1(_06105_),
    .B2(_05343_),
    .Y(_06271_));
 INVx1_ASAP7_75t_R _25739_ (.A(_01478_),
    .Y(_06272_));
 AO32x1_ASAP7_75t_R _25740_ (.A1(net191),
    .A2(_05800_),
    .A3(_05001_),
    .B1(_05811_),
    .B2(_06272_),
    .Y(_06273_));
 OAI22x1_ASAP7_75t_R _25741_ (.A1(_01913_),
    .A2(_05815_),
    .B1(_05951_),
    .B2(_01963_),
    .Y(_06274_));
 OA22x2_ASAP7_75t_R _25742_ (.A1(_01834_),
    .A2(_05944_),
    .B1(_05937_),
    .B2(_02001_),
    .Y(_06275_));
 OA22x2_ASAP7_75t_R _25743_ (.A1(_02033_),
    .A2(_05949_),
    .B1(_05943_),
    .B2(_02061_),
    .Y(_06276_));
 NAND2x1_ASAP7_75t_R _25744_ (.A(_06275_),
    .B(_06276_),
    .Y(_06277_));
 OR5x2_ASAP7_75t_R _25745_ (.A(_06151_),
    .B(_06271_),
    .C(_06273_),
    .D(_06274_),
    .E(_06277_),
    .Y(_06278_));
 AO221x2_ASAP7_75t_R _25746_ (.A1(_05929_),
    .A2(_06269_),
    .B1(_06270_),
    .B2(_06007_),
    .C(_06278_),
    .Y(_06279_));
 OA22x2_ASAP7_75t_R _25747_ (.A1(_06072_),
    .A2(_06268_),
    .B1(_06279_),
    .B2(_18725_),
    .Y(_06280_));
 AO32x1_ASAP7_75t_R _25748_ (.A1(_02194_),
    .A2(_06226_),
    .A3(_06266_),
    .B1(_06280_),
    .B2(_06043_),
    .Y(_06281_));
 AO22x1_ASAP7_75t_R _25749_ (.A1(_06263_),
    .A2(_06265_),
    .B1(_06281_),
    .B2(_06045_),
    .Y(_02376_));
 INVx1_ASAP7_75t_R _25750_ (.A(_02193_),
    .Y(_06282_));
 OR3x1_ASAP7_75t_R _25751_ (.A(_02194_),
    .B(_06243_),
    .C(_06244_),
    .Y(_06283_));
 AO21x1_ASAP7_75t_R _25752_ (.A1(_06025_),
    .A2(_06283_),
    .B(_05892_),
    .Y(_06284_));
 NAND2x1_ASAP7_75t_R _25753_ (.A(_18861_),
    .B(_18730_),
    .Y(_06285_));
 OA21x2_ASAP7_75t_R _25754_ (.A1(_05846_),
    .A2(_18730_),
    .B(_06285_),
    .Y(_06286_));
 OAI22x1_ASAP7_75t_R _25755_ (.A1(_02193_),
    .A2(_05778_),
    .B1(_05782_),
    .B2(_02130_),
    .Y(_06287_));
 OAI22x1_ASAP7_75t_R _25756_ (.A1(_02158_),
    .A2(_05778_),
    .B1(_05782_),
    .B2(_02095_),
    .Y(_06288_));
 OA222x2_ASAP7_75t_R _25757_ (.A1(_01833_),
    .A2(_05816_),
    .B1(_05835_),
    .B2(_01962_),
    .C1(_05856_),
    .C2(_02060_),
    .Y(_06289_));
 INVx1_ASAP7_75t_R _25758_ (.A(_06289_),
    .Y(_06290_));
 OAI22x1_ASAP7_75t_R _25759_ (.A1(_02000_),
    .A2(_05829_),
    .B1(_05833_),
    .B2(_02032_),
    .Y(_06291_));
 OAI21x1_ASAP7_75t_R _25760_ (.A1(_01912_),
    .A2(_05941_),
    .B(_05821_),
    .Y(_06292_));
 AND2x2_ASAP7_75t_R _25761_ (.A(net192),
    .B(_06106_),
    .Y(_06293_));
 INVx1_ASAP7_75t_R _25762_ (.A(_01479_),
    .Y(_06294_));
 AO222x2_ASAP7_75t_R _25763_ (.A1(net123),
    .A2(_05802_),
    .B1(_06105_),
    .B2(_05365_),
    .C1(_05810_),
    .C2(_06294_),
    .Y(_06295_));
 OR5x2_ASAP7_75t_R _25764_ (.A(_06290_),
    .B(_06291_),
    .C(_06292_),
    .D(_06293_),
    .E(_06295_),
    .Y(_06296_));
 AO221x2_ASAP7_75t_R _25765_ (.A1(_05795_),
    .A2(_06287_),
    .B1(_06288_),
    .B2(_05798_),
    .C(_06296_),
    .Y(_06297_));
 OA22x2_ASAP7_75t_R _25766_ (.A1(_05844_),
    .A2(_06286_),
    .B1(_06297_),
    .B2(_18730_),
    .Y(_06298_));
 BUFx10_ASAP7_75t_R _25767_ (.A(_06298_),
    .Y(_06299_));
 INVx1_ASAP7_75t_R _25768_ (.A(_06283_),
    .Y(_06300_));
 AND3x1_ASAP7_75t_R _25769_ (.A(_02193_),
    .B(_05921_),
    .C(_06300_),
    .Y(_06301_));
 AO21x1_ASAP7_75t_R _25770_ (.A1(_06047_),
    .A2(_06299_),
    .B(_06301_),
    .Y(_06302_));
 AO22x1_ASAP7_75t_R _25771_ (.A1(_06282_),
    .A2(_06284_),
    .B1(_06302_),
    .B2(_06045_),
    .Y(_02377_));
 OR4x1_ASAP7_75t_R _25772_ (.A(_02194_),
    .B(_06243_),
    .C(_06222_),
    .D(_02197_),
    .Y(_06303_));
 OR3x1_ASAP7_75t_R _25773_ (.A(_02193_),
    .B(_02199_),
    .C(_06303_),
    .Y(_06304_));
 OR2x2_ASAP7_75t_R _25774_ (.A(_06164_),
    .B(_06304_),
    .Y(_06305_));
 AO21x1_ASAP7_75t_R _25775_ (.A1(_06116_),
    .A2(_06305_),
    .B(_05926_),
    .Y(_06306_));
 NAND2x1_ASAP7_75t_R _25776_ (.A(_06074_),
    .B(_18732_),
    .Y(_06307_));
 OA21x2_ASAP7_75t_R _25777_ (.A1(_06073_),
    .A2(_18732_),
    .B(_06307_),
    .Y(_06308_));
 OAI22x1_ASAP7_75t_R _25778_ (.A1(_02192_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02129_),
    .Y(_06309_));
 OAI22x1_ASAP7_75t_R _25779_ (.A1(_02157_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_02094_),
    .Y(_06310_));
 INVx1_ASAP7_75t_R _25780_ (.A(_01480_),
    .Y(_06311_));
 AO22x1_ASAP7_75t_R _25781_ (.A1(net124),
    .A2(_05938_),
    .B1(_06105_),
    .B2(_05364_),
    .Y(_06312_));
 AO221x1_ASAP7_75t_R _25782_ (.A1(_06311_),
    .A2(_05811_),
    .B1(_06106_),
    .B2(net193),
    .C(_06312_),
    .Y(_06313_));
 OAI22x1_ASAP7_75t_R _25783_ (.A1(_01911_),
    .A2(_05815_),
    .B1(_05949_),
    .B2(_02031_),
    .Y(_06314_));
 OAI22x1_ASAP7_75t_R _25784_ (.A1(_01832_),
    .A2(_05945_),
    .B1(_05943_),
    .B2(_02059_),
    .Y(_06315_));
 OAI22x1_ASAP7_75t_R _25785_ (.A1(_01999_),
    .A2(_05937_),
    .B1(_05951_),
    .B2(_01961_),
    .Y(_06316_));
 OR5x2_ASAP7_75t_R _25786_ (.A(_06151_),
    .B(_06313_),
    .C(_06314_),
    .D(_06315_),
    .E(_06316_),
    .Y(_06317_));
 AO221x2_ASAP7_75t_R _25787_ (.A1(_06007_),
    .A2(_06309_),
    .B1(_06310_),
    .B2(_05930_),
    .C(_06317_),
    .Y(_06318_));
 OA22x2_ASAP7_75t_R _25788_ (.A1(_06072_),
    .A2(_06308_),
    .B1(_06318_),
    .B2(_18732_),
    .Y(_06319_));
 BUFx10_ASAP7_75t_R _25789_ (.A(_06319_),
    .Y(_06320_));
 AND2x4_ASAP7_75t_R _25790_ (.A(_04971_),
    .B(_05915_),
    .Y(_06321_));
 AND3x1_ASAP7_75t_R _25791_ (.A(_05031_),
    .B(_05889_),
    .C(_06321_),
    .Y(_06322_));
 BUFx6f_ASAP7_75t_R _25792_ (.A(_06322_),
    .Y(_06323_));
 OR3x1_ASAP7_75t_R _25793_ (.A(_02192_),
    .B(_06164_),
    .C(_06304_),
    .Y(_06324_));
 BUFx3_ASAP7_75t_R _25794_ (.A(_06324_),
    .Y(_06325_));
 AO21x1_ASAP7_75t_R _25795_ (.A1(_05880_),
    .A2(_06323_),
    .B(_06325_),
    .Y(_06326_));
 OAI21x1_ASAP7_75t_R _25796_ (.A1(_06021_),
    .A2(_06320_),
    .B(_06326_),
    .Y(_06327_));
 AOI22x1_ASAP7_75t_R _25797_ (.A1(_02192_),
    .A2(_06306_),
    .B1(_06327_),
    .B2(_05959_),
    .Y(_02378_));
 BUFx4f_ASAP7_75t_R _25798_ (.A(_02191_),
    .Y(_06328_));
 OR4x2_ASAP7_75t_R _25799_ (.A(_02192_),
    .B(_02200_),
    .C(_06140_),
    .D(_06304_),
    .Y(_06329_));
 AOI21x1_ASAP7_75t_R _25800_ (.A1(_05922_),
    .A2(_06329_),
    .B(_06002_),
    .Y(_06330_));
 NOR2x1_ASAP7_75t_R _25801_ (.A(_05970_),
    .B(_06329_),
    .Y(_06331_));
 NAND2x1_ASAP7_75t_R _25802_ (.A(_06328_),
    .B(_06331_),
    .Y(_06332_));
 AND2x2_ASAP7_75t_R _25803_ (.A(_05773_),
    .B(_18740_),
    .Y(_06333_));
 AO21x1_ASAP7_75t_R _25804_ (.A1(_05772_),
    .A2(_18738_),
    .B(_06333_),
    .Y(_06334_));
 OAI22x1_ASAP7_75t_R _25805_ (.A1(_02156_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_02093_),
    .Y(_06335_));
 BUFx4f_ASAP7_75t_R _25806_ (.A(_02128_),
    .Y(_06336_));
 OAI22x1_ASAP7_75t_R _25807_ (.A1(_06328_),
    .A2(_05780_),
    .B1(_05784_),
    .B2(_06336_),
    .Y(_06337_));
 AO32x1_ASAP7_75t_R _25808_ (.A1(net180),
    .A2(_05800_),
    .A3(_05001_),
    .B1(_06105_),
    .B2(_05362_),
    .Y(_06338_));
 INVx1_ASAP7_75t_R _25809_ (.A(_01481_),
    .Y(_06339_));
 AO221x1_ASAP7_75t_R _25810_ (.A1(net125),
    .A2(_05938_),
    .B1(_05811_),
    .B2(_06339_),
    .C(_06151_),
    .Y(_06340_));
 OAI22x1_ASAP7_75t_R _25811_ (.A1(_02030_),
    .A2(_05949_),
    .B1(_05937_),
    .B2(_01998_),
    .Y(_06341_));
 OA22x2_ASAP7_75t_R _25812_ (.A1(_01960_),
    .A2(_05951_),
    .B1(_05943_),
    .B2(_02058_),
    .Y(_06342_));
 OA22x2_ASAP7_75t_R _25813_ (.A1(_01910_),
    .A2(_05815_),
    .B1(_05945_),
    .B2(_01831_),
    .Y(_06343_));
 NAND2x1_ASAP7_75t_R _25814_ (.A(_06342_),
    .B(_06343_),
    .Y(_06344_));
 OR4x2_ASAP7_75t_R _25815_ (.A(_06338_),
    .B(_06340_),
    .C(_06341_),
    .D(_06344_),
    .Y(_06345_));
 AOI221x1_ASAP7_75t_R _25816_ (.A1(_05930_),
    .A2(_06335_),
    .B1(_06337_),
    .B2(_06007_),
    .C(_06345_),
    .Y(_06346_));
 AO22x2_ASAP7_75t_R _25817_ (.A1(_05771_),
    .A2(_06334_),
    .B1(_06346_),
    .B2(_18738_),
    .Y(_06347_));
 OR2x2_ASAP7_75t_R _25818_ (.A(_05921_),
    .B(_06347_),
    .Y(_06348_));
 AO21x1_ASAP7_75t_R _25819_ (.A1(_06332_),
    .A2(_06348_),
    .B(_05926_),
    .Y(_06349_));
 OAI21x1_ASAP7_75t_R _25820_ (.A1(_06328_),
    .A2(_06330_),
    .B(_06349_),
    .Y(_02379_));
 BUFx10_ASAP7_75t_R _25821_ (.A(_05887_),
    .Y(_06350_));
 OAI21x1_ASAP7_75t_R _25822_ (.A1(_06328_),
    .A2(_06325_),
    .B(_06350_),
    .Y(_06351_));
 AO21x1_ASAP7_75t_R _25823_ (.A1(_05919_),
    .A2(_06351_),
    .B(_02190_),
    .Y(_06352_));
 INVx1_ASAP7_75t_R _25824_ (.A(_02190_),
    .Y(_06353_));
 OR4x1_ASAP7_75t_R _25825_ (.A(_06353_),
    .B(_06328_),
    .C(_05882_),
    .D(_06325_),
    .Y(_06354_));
 NAND2x1_ASAP7_75t_R _25826_ (.A(_18861_),
    .B(_18742_),
    .Y(_06355_));
 OA21x2_ASAP7_75t_R _25827_ (.A1(_05846_),
    .A2(_18742_),
    .B(_06355_),
    .Y(_06356_));
 OAI22x1_ASAP7_75t_R _25828_ (.A1(_02190_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_02127_),
    .Y(_06357_));
 BUFx4f_ASAP7_75t_R _25829_ (.A(_02155_),
    .Y(_06358_));
 BUFx4f_ASAP7_75t_R _25830_ (.A(_02092_),
    .Y(_06359_));
 OAI22x1_ASAP7_75t_R _25831_ (.A1(_06358_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_06359_),
    .Y(_06360_));
 OA222x2_ASAP7_75t_R _25832_ (.A1(_01830_),
    .A2(_05817_),
    .B1(_05836_),
    .B2(_01959_),
    .C1(_05857_),
    .C2(_02057_),
    .Y(_06361_));
 INVx1_ASAP7_75t_R _25833_ (.A(_06361_),
    .Y(_06362_));
 OAI22x1_ASAP7_75t_R _25834_ (.A1(_01997_),
    .A2(_05830_),
    .B1(_05834_),
    .B2(_02029_),
    .Y(_06363_));
 OAI21x1_ASAP7_75t_R _25835_ (.A1(_01909_),
    .A2(_05941_),
    .B(_05821_),
    .Y(_06364_));
 AND2x2_ASAP7_75t_R _25836_ (.A(net181),
    .B(_06106_),
    .Y(_06365_));
 INVx1_ASAP7_75t_R _25837_ (.A(_00007_),
    .Y(_06366_));
 AO222x2_ASAP7_75t_R _25838_ (.A1(net126),
    .A2(_05803_),
    .B1(_06105_),
    .B2(_05361_),
    .C1(_05810_),
    .C2(_06366_),
    .Y(_06367_));
 OR5x2_ASAP7_75t_R _25839_ (.A(_06362_),
    .B(_06363_),
    .C(_06364_),
    .D(_06365_),
    .E(_06367_),
    .Y(_06368_));
 AO221x2_ASAP7_75t_R _25840_ (.A1(_05796_),
    .A2(_06357_),
    .B1(_06360_),
    .B2(_05799_),
    .C(_06368_),
    .Y(_06369_));
 OAI22x1_ASAP7_75t_R _25841_ (.A1(_05844_),
    .A2(_06356_),
    .B1(_06369_),
    .B2(_18742_),
    .Y(_06370_));
 OR2x2_ASAP7_75t_R _25842_ (.A(_05921_),
    .B(_06370_),
    .Y(_06371_));
 AO21x1_ASAP7_75t_R _25843_ (.A1(_06354_),
    .A2(_06371_),
    .B(_05893_),
    .Y(_06372_));
 NAND2x1_ASAP7_75t_R _25844_ (.A(_06352_),
    .B(_06372_),
    .Y(_02380_));
 INVx1_ASAP7_75t_R _25845_ (.A(_02189_),
    .Y(_06373_));
 OR3x1_ASAP7_75t_R _25846_ (.A(_02190_),
    .B(_06328_),
    .C(_06329_),
    .Y(_06374_));
 AO21x1_ASAP7_75t_R _25847_ (.A1(_05918_),
    .A2(_06374_),
    .B(_05892_),
    .Y(_06375_));
 NOR2x1_ASAP7_75t_R _25848_ (.A(_02190_),
    .B(_06328_),
    .Y(_06376_));
 NAND2x1_ASAP7_75t_R _25849_ (.A(_05773_),
    .B(_18747_),
    .Y(_06377_));
 OA21x2_ASAP7_75t_R _25850_ (.A1(_06073_),
    .A2(_18747_),
    .B(_06377_),
    .Y(_06378_));
 OAI22x1_ASAP7_75t_R _25851_ (.A1(_02189_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02126_),
    .Y(_06379_));
 BUFx3_ASAP7_75t_R _25852_ (.A(_02090_),
    .Y(_06380_));
 OAI22x1_ASAP7_75t_R _25853_ (.A1(_02153_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_06380_),
    .Y(_06381_));
 OA222x2_ASAP7_75t_R _25854_ (.A1(_01996_),
    .A2(_05829_),
    .B1(_05857_),
    .B2(_02056_),
    .C1(_05985_),
    .C2(_01958_),
    .Y(_06382_));
 OR2x2_ASAP7_75t_R _25855_ (.A(_00008_),
    .B(_05987_),
    .Y(_06383_));
 INVx1_ASAP7_75t_R _25856_ (.A(net127),
    .Y(_06384_));
 INVx1_ASAP7_75t_R _25857_ (.A(net182),
    .Y(_06385_));
 OA222x2_ASAP7_75t_R _25858_ (.A1(_06384_),
    .A2(_05989_),
    .B1(_05991_),
    .B2(_01943_),
    .C1(_05992_),
    .C2(_06385_),
    .Y(_06386_));
 OA21x2_ASAP7_75t_R _25859_ (.A1(_01908_),
    .A2(_05983_),
    .B(_05995_),
    .Y(_06387_));
 OA22x2_ASAP7_75t_R _25860_ (.A1(_02028_),
    .A2(_05833_),
    .B1(_05980_),
    .B2(_01829_),
    .Y(_06388_));
 AND5x1_ASAP7_75t_R _25861_ (.A(_06382_),
    .B(_06383_),
    .C(_06386_),
    .D(_06387_),
    .E(_06388_),
    .Y(_06389_));
 INVx1_ASAP7_75t_R _25862_ (.A(_06389_),
    .Y(_06390_));
 AO221x2_ASAP7_75t_R _25863_ (.A1(_05976_),
    .A2(_06379_),
    .B1(_06381_),
    .B2(_05929_),
    .C(_06390_),
    .Y(_06391_));
 OA22x2_ASAP7_75t_R _25864_ (.A1(_06072_),
    .A2(_06378_),
    .B1(_06391_),
    .B2(_18747_),
    .Y(_06392_));
 AO32x1_ASAP7_75t_R _25865_ (.A1(_02189_),
    .A2(_06331_),
    .A3(_06376_),
    .B1(_06392_),
    .B2(_06043_),
    .Y(_06393_));
 AO22x1_ASAP7_75t_R _25866_ (.A1(_06373_),
    .A2(_06375_),
    .B1(_06393_),
    .B2(_05919_),
    .Y(_02381_));
 INVx1_ASAP7_75t_R _25867_ (.A(_02188_),
    .Y(_06394_));
 OR3x2_ASAP7_75t_R _25868_ (.A(_02189_),
    .B(_02190_),
    .C(_06328_),
    .Y(_06395_));
 OR4x1_ASAP7_75t_R _25869_ (.A(_06394_),
    .B(_05882_),
    .C(_06325_),
    .D(_06395_),
    .Y(_06396_));
 NAND2x1_ASAP7_75t_R _25870_ (.A(_14736_),
    .B(_18752_),
    .Y(_06397_));
 OA21x2_ASAP7_75t_R _25871_ (.A1(_05845_),
    .A2(_18752_),
    .B(_06397_),
    .Y(_06398_));
 OAI22x1_ASAP7_75t_R _25872_ (.A1(_02188_),
    .A2(_05777_),
    .B1(_05781_),
    .B2(_02125_),
    .Y(_06399_));
 OAI22x1_ASAP7_75t_R _25873_ (.A1(_02152_),
    .A2(_05778_),
    .B1(_05782_),
    .B2(_02089_),
    .Y(_06400_));
 OA222x2_ASAP7_75t_R _25874_ (.A1(_01828_),
    .A2(_05816_),
    .B1(_05835_),
    .B2(_01957_),
    .C1(_05856_),
    .C2(_02055_),
    .Y(_06401_));
 INVx1_ASAP7_75t_R _25875_ (.A(_06401_),
    .Y(_06402_));
 OAI22x1_ASAP7_75t_R _25876_ (.A1(_01995_),
    .A2(_05828_),
    .B1(_05832_),
    .B2(_02027_),
    .Y(_06403_));
 OAI21x1_ASAP7_75t_R _25877_ (.A1(_01907_),
    .A2(_05814_),
    .B(_05820_),
    .Y(_06404_));
 AND2x2_ASAP7_75t_R _25878_ (.A(net183),
    .B(_06106_),
    .Y(_06405_));
 INVx1_ASAP7_75t_R _25879_ (.A(_00009_),
    .Y(_06406_));
 AO222x2_ASAP7_75t_R _25880_ (.A1(net128),
    .A2(_05802_),
    .B1(_06104_),
    .B2(_05358_),
    .C1(_05810_),
    .C2(_06406_),
    .Y(_06407_));
 OR5x2_ASAP7_75t_R _25881_ (.A(_06402_),
    .B(_06403_),
    .C(_06404_),
    .D(_06405_),
    .E(_06407_),
    .Y(_06408_));
 AO221x2_ASAP7_75t_R _25882_ (.A1(_05795_),
    .A2(_06399_),
    .B1(_06400_),
    .B2(_05798_),
    .C(_06408_),
    .Y(_06409_));
 OA22x2_ASAP7_75t_R _25883_ (.A1(_05843_),
    .A2(_06398_),
    .B1(_06409_),
    .B2(_18752_),
    .Y(_06410_));
 BUFx10_ASAP7_75t_R _25884_ (.A(_06410_),
    .Y(_06411_));
 NAND2x1_ASAP7_75t_R _25885_ (.A(_06144_),
    .B(_06411_),
    .Y(_06412_));
 NAND2x1_ASAP7_75t_R _25886_ (.A(_06396_),
    .B(_06412_),
    .Y(_06413_));
 OA21x2_ASAP7_75t_R _25887_ (.A1(_06325_),
    .A2(_06395_),
    .B(_05887_),
    .Y(_06414_));
 OA21x2_ASAP7_75t_R _25888_ (.A1(_05893_),
    .A2(_06414_),
    .B(_06394_),
    .Y(_06415_));
 AO21x1_ASAP7_75t_R _25889_ (.A1(_05959_),
    .A2(_06413_),
    .B(_06415_),
    .Y(_02382_));
 OR3x1_ASAP7_75t_R _25890_ (.A(_02187_),
    .B(_02313_),
    .C(_06113_),
    .Y(_06416_));
 OAI21x1_ASAP7_75t_R _25891_ (.A1(_05872_),
    .A2(_05922_),
    .B(_06416_),
    .Y(_06417_));
 AO21x1_ASAP7_75t_R _25892_ (.A1(_02313_),
    .A2(_05922_),
    .B(_05926_),
    .Y(_06418_));
 AOI22x1_ASAP7_75t_R _25893_ (.A1(_05959_),
    .A2(_06417_),
    .B1(_06418_),
    .B2(_02187_),
    .Y(_02383_));
 INVx1_ASAP7_75t_R _25894_ (.A(_02186_),
    .Y(_06419_));
 OR2x2_ASAP7_75t_R _25895_ (.A(_02188_),
    .B(_06395_),
    .Y(_06420_));
 OR2x2_ASAP7_75t_R _25896_ (.A(_06329_),
    .B(_06420_),
    .Y(_06421_));
 AO21x1_ASAP7_75t_R _25897_ (.A1(_05918_),
    .A2(_06421_),
    .B(_05892_),
    .Y(_06422_));
 INVx1_ASAP7_75t_R _25898_ (.A(_06420_),
    .Y(_06423_));
 NAND2x1_ASAP7_75t_R _25899_ (.A(_06074_),
    .B(_18760_),
    .Y(_06424_));
 OA21x2_ASAP7_75t_R _25900_ (.A1(_06073_),
    .A2(_18760_),
    .B(_06424_),
    .Y(_06425_));
 OAI22x1_ASAP7_75t_R _25901_ (.A1(_02186_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02123_),
    .Y(_06426_));
 OAI22x1_ASAP7_75t_R _25902_ (.A1(_02151_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02088_),
    .Y(_06427_));
 AND2x2_ASAP7_75t_R _25903_ (.A(_04994_),
    .B(_05056_),
    .Y(_06428_));
 OAI21x1_ASAP7_75t_R _25904_ (.A1(_01941_),
    .A2(_06251_),
    .B(_05827_),
    .Y(_06429_));
 AO21x1_ASAP7_75t_R _25905_ (.A1(net130),
    .A2(_05803_),
    .B(_06429_),
    .Y(_06430_));
 INVx1_ASAP7_75t_R _25906_ (.A(_00010_),
    .Y(_06431_));
 AO32x1_ASAP7_75t_R _25907_ (.A1(net184),
    .A2(_05800_),
    .A3(_05001_),
    .B1(_05811_),
    .B2(_06431_),
    .Y(_06432_));
 OAI22x1_ASAP7_75t_R _25908_ (.A1(_01905_),
    .A2(_05941_),
    .B1(_05834_),
    .B2(_02025_),
    .Y(_06433_));
 OA22x2_ASAP7_75t_R _25909_ (.A1(_01993_),
    .A2(_05829_),
    .B1(_05857_),
    .B2(_02053_),
    .Y(_06434_));
 OA22x2_ASAP7_75t_R _25910_ (.A1(_01826_),
    .A2(_05817_),
    .B1(_05836_),
    .B2(_01955_),
    .Y(_06435_));
 NAND2x1_ASAP7_75t_R _25911_ (.A(_06434_),
    .B(_06435_),
    .Y(_06436_));
 OR5x2_ASAP7_75t_R _25912_ (.A(_06428_),
    .B(_06430_),
    .C(_06432_),
    .D(_06433_),
    .E(_06436_),
    .Y(_06437_));
 AO221x2_ASAP7_75t_R _25913_ (.A1(_05796_),
    .A2(_06426_),
    .B1(_06427_),
    .B2(_05799_),
    .C(_06437_),
    .Y(_06438_));
 OA22x2_ASAP7_75t_R _25914_ (.A1(_06072_),
    .A2(_06425_),
    .B1(_06438_),
    .B2(_18760_),
    .Y(_06439_));
 AO32x1_ASAP7_75t_R _25915_ (.A1(_02186_),
    .A2(_06331_),
    .A3(_06423_),
    .B1(_06439_),
    .B2(_06144_),
    .Y(_06440_));
 AO22x1_ASAP7_75t_R _25916_ (.A1(_06419_),
    .A2(_06422_),
    .B1(_06440_),
    .B2(_05919_),
    .Y(_02384_));
 NOR2x1_ASAP7_75t_R _25917_ (.A(_18865_),
    .B(_18845_),
    .Y(_06441_));
 AO21x1_ASAP7_75t_R _25918_ (.A1(_05772_),
    .A2(_18845_),
    .B(_06441_),
    .Y(_06442_));
 OA22x2_ASAP7_75t_R _25919_ (.A1(_02150_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_02087_),
    .Y(_06443_));
 OAI22x1_ASAP7_75t_R _25920_ (.A1(_02185_),
    .A2(_05849_),
    .B1(_05851_),
    .B2(_02122_),
    .Y(_06444_));
 NAND2x1_ASAP7_75t_R _25921_ (.A(_05976_),
    .B(_06444_),
    .Y(_06445_));
 NAND2x1_ASAP7_75t_R _25922_ (.A(net131),
    .B(_05025_),
    .Y(_06446_));
 OA211x2_ASAP7_75t_R _25923_ (.A1(_00011_),
    .A2(_05809_),
    .B(_06446_),
    .C(_05769_),
    .Y(_06447_));
 OR2x2_ASAP7_75t_R _25924_ (.A(_01954_),
    .B(_05950_),
    .Y(_06448_));
 OA22x2_ASAP7_75t_R _25925_ (.A1(_01825_),
    .A2(_05945_),
    .B1(_05943_),
    .B2(_02052_),
    .Y(_06449_));
 OA22x2_ASAP7_75t_R _25926_ (.A1(_02024_),
    .A2(_05948_),
    .B1(_06189_),
    .B2(_01979_),
    .Y(_06450_));
 OA22x2_ASAP7_75t_R _25927_ (.A1(_01904_),
    .A2(_05941_),
    .B1(_05937_),
    .B2(_01992_),
    .Y(_06451_));
 AND5x2_ASAP7_75t_R _25928_ (.A(_06447_),
    .B(_06448_),
    .C(_06449_),
    .D(_06450_),
    .E(_06451_),
    .Y(_06452_));
 OA211x2_ASAP7_75t_R _25929_ (.A1(_05974_),
    .A2(_06443_),
    .B(_06445_),
    .C(_06452_),
    .Y(_06453_));
 AO22x1_ASAP7_75t_R _25930_ (.A1(_02307_),
    .A2(_06442_),
    .B1(_06453_),
    .B2(_18845_),
    .Y(_06454_));
 BUFx10_ASAP7_75t_R _25931_ (.A(_06454_),
    .Y(_06455_));
 INVx1_ASAP7_75t_R _25932_ (.A(_02185_),
    .Y(_06456_));
 OR3x2_ASAP7_75t_R _25933_ (.A(_02186_),
    .B(_02188_),
    .C(_06395_),
    .Y(_06457_));
 OR4x1_ASAP7_75t_R _25934_ (.A(_06456_),
    .B(_05882_),
    .C(_06325_),
    .D(_06457_),
    .Y(_06458_));
 OA21x2_ASAP7_75t_R _25935_ (.A1(_06021_),
    .A2(_06455_),
    .B(_06458_),
    .Y(_06459_));
 OAI21x1_ASAP7_75t_R _25936_ (.A1(_06325_),
    .A2(_06457_),
    .B(_06021_),
    .Y(_06460_));
 AO21x1_ASAP7_75t_R _25937_ (.A1(_05919_),
    .A2(_06460_),
    .B(_02185_),
    .Y(_06461_));
 OAI21x1_ASAP7_75t_R _25938_ (.A1(_06002_),
    .A2(_06459_),
    .B(_06461_),
    .Y(_02385_));
 INVx1_ASAP7_75t_R _25939_ (.A(_02184_),
    .Y(_06462_));
 OR3x4_ASAP7_75t_R _25940_ (.A(_02185_),
    .B(_06329_),
    .C(_06457_),
    .Y(_06463_));
 AOI22x1_ASAP7_75t_R _25941_ (.A1(_05930_),
    .A2(_05969_),
    .B1(_05891_),
    .B2(_00788_),
    .Y(_06464_));
 BUFx4f_ASAP7_75t_R _25942_ (.A(_06464_),
    .Y(_06465_));
 AO21x1_ASAP7_75t_R _25943_ (.A1(_05918_),
    .A2(_06463_),
    .B(_06465_),
    .Y(_06466_));
 NOR2x1_ASAP7_75t_R _25944_ (.A(_05970_),
    .B(_06463_),
    .Y(_06467_));
 AO22x1_ASAP7_75t_R _25945_ (.A1(_05841_),
    .A2(_06043_),
    .B1(_06467_),
    .B2(_02184_),
    .Y(_06468_));
 AO22x1_ASAP7_75t_R _25946_ (.A1(_05930_),
    .A2(_05969_),
    .B1(_05891_),
    .B2(_00788_),
    .Y(_06469_));
 BUFx4f_ASAP7_75t_R _25947_ (.A(_06469_),
    .Y(_06470_));
 BUFx4f_ASAP7_75t_R _25948_ (.A(_06470_),
    .Y(_06471_));
 AO22x1_ASAP7_75t_R _25949_ (.A1(_06462_),
    .A2(_06466_),
    .B1(_06468_),
    .B2(_06471_),
    .Y(_02386_));
 BUFx6f_ASAP7_75t_R _25950_ (.A(_06470_),
    .Y(_06472_));
 OR3x4_ASAP7_75t_R _25951_ (.A(_02185_),
    .B(_06325_),
    .C(_06457_),
    .Y(_06473_));
 AOI21x1_ASAP7_75t_R _25952_ (.A1(_05880_),
    .A2(_06323_),
    .B(_06473_),
    .Y(_06474_));
 AOI21x1_ASAP7_75t_R _25953_ (.A1(_18615_),
    .A2(_06194_),
    .B(_06197_),
    .Y(_06475_));
 AO32x1_ASAP7_75t_R _25954_ (.A1(_02183_),
    .A2(_06462_),
    .A3(_06474_),
    .B1(_06475_),
    .B2(_05882_),
    .Y(_06476_));
 OAI21x1_ASAP7_75t_R _25955_ (.A1(_02184_),
    .A2(_06473_),
    .B(_06021_),
    .Y(_06477_));
 AOI21x1_ASAP7_75t_R _25956_ (.A1(_06471_),
    .A2(_06477_),
    .B(_02183_),
    .Y(_06478_));
 AO21x1_ASAP7_75t_R _25957_ (.A1(_06472_),
    .A2(_06476_),
    .B(_06478_),
    .Y(_02387_));
 OR3x1_ASAP7_75t_R _25958_ (.A(_02183_),
    .B(_02184_),
    .C(_06463_),
    .Y(_06479_));
 BUFx4f_ASAP7_75t_R _25959_ (.A(_06464_),
    .Y(_06480_));
 AO21x1_ASAP7_75t_R _25960_ (.A1(_06116_),
    .A2(_06479_),
    .B(_06480_),
    .Y(_06481_));
 OR3x2_ASAP7_75t_R _25961_ (.A(_02182_),
    .B(_02183_),
    .C(_02184_),
    .Y(_06482_));
 INVx1_ASAP7_75t_R _25962_ (.A(_06482_),
    .Y(_06483_));
 AO22x1_ASAP7_75t_R _25963_ (.A1(_05871_),
    .A2(_05883_),
    .B1(_06467_),
    .B2(_06483_),
    .Y(_06484_));
 AOI22x1_ASAP7_75t_R _25964_ (.A1(_02182_),
    .A2(_06481_),
    .B1(_06484_),
    .B2(_06472_),
    .Y(_02388_));
 NAND2x1_ASAP7_75t_R _25965_ (.A(_06074_),
    .B(_18622_),
    .Y(_06485_));
 OA21x2_ASAP7_75t_R _25966_ (.A1(_06073_),
    .A2(_18622_),
    .B(_06485_),
    .Y(_06486_));
 OAI22x1_ASAP7_75t_R _25967_ (.A1(_02176_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02113_),
    .Y(_06487_));
 BUFx3_ASAP7_75t_R _25968_ (.A(_02118_),
    .Y(_06488_));
 OAI22x1_ASAP7_75t_R _25969_ (.A1(_02181_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_06488_),
    .Y(_06489_));
 OA22x2_ASAP7_75t_R _25970_ (.A1(_02023_),
    .A2(_05833_),
    .B1(_05857_),
    .B2(_01461_),
    .Y(_06490_));
 OR4x1_ASAP7_75t_R _25971_ (.A(_05034_),
    .B(_01981_),
    .C(_14308_),
    .D(_05897_),
    .Y(_06491_));
 OA211x2_ASAP7_75t_R _25972_ (.A1(_01991_),
    .A2(_05830_),
    .B(_06490_),
    .C(_06491_),
    .Y(_06492_));
 INVx1_ASAP7_75t_R _25973_ (.A(net132),
    .Y(_06493_));
 OA222x2_ASAP7_75t_R _25974_ (.A1(_06493_),
    .A2(_05989_),
    .B1(_05991_),
    .B2(_01938_),
    .C1(_05992_),
    .C2(_05368_),
    .Y(_06494_));
 OA22x2_ASAP7_75t_R _25975_ (.A1(_01953_),
    .A2(_05985_),
    .B1(_05980_),
    .B2(_01824_),
    .Y(_06495_));
 OA211x2_ASAP7_75t_R _25976_ (.A1(_01850_),
    .A2(_05994_),
    .B(_06495_),
    .C(_05995_),
    .Y(_06496_));
 OA211x2_ASAP7_75t_R _25977_ (.A1(_01903_),
    .A2(_05983_),
    .B(_06494_),
    .C(_06496_),
    .Y(_06497_));
 NAND2x1_ASAP7_75t_R _25978_ (.A(_06492_),
    .B(_06497_),
    .Y(_06498_));
 AO221x2_ASAP7_75t_R _25979_ (.A1(_06007_),
    .A2(_06487_),
    .B1(_06489_),
    .B2(_05929_),
    .C(_06498_),
    .Y(_06499_));
 OA22x2_ASAP7_75t_R _25980_ (.A1(_06072_),
    .A2(_06486_),
    .B1(_06499_),
    .B2(_18622_),
    .Y(_06500_));
 AO32x1_ASAP7_75t_R _25981_ (.A1(_02181_),
    .A2(_06474_),
    .A3(_06483_),
    .B1(_06500_),
    .B2(_06047_),
    .Y(_06501_));
 OAI21x1_ASAP7_75t_R _25982_ (.A1(_06473_),
    .A2(_06482_),
    .B(_06350_),
    .Y(_06502_));
 AOI21x1_ASAP7_75t_R _25983_ (.A1(_06471_),
    .A2(_06502_),
    .B(_02181_),
    .Y(_06503_));
 AO21x1_ASAP7_75t_R _25984_ (.A1(_06472_),
    .A2(_06501_),
    .B(_06503_),
    .Y(_02389_));
 OR3x1_ASAP7_75t_R _25985_ (.A(_02181_),
    .B(_06463_),
    .C(_06482_),
    .Y(_06504_));
 AO21x1_ASAP7_75t_R _25986_ (.A1(_06116_),
    .A2(_06504_),
    .B(_06480_),
    .Y(_06505_));
 NAND2x1_ASAP7_75t_R _25987_ (.A(_18861_),
    .B(_18630_),
    .Y(_06506_));
 OA21x2_ASAP7_75t_R _25988_ (.A1(_05846_),
    .A2(_18630_),
    .B(_06506_),
    .Y(_06507_));
 OAI22x1_ASAP7_75t_R _25989_ (.A1(_02180_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02117_),
    .Y(_06508_));
 OAI22x1_ASAP7_75t_R _25990_ (.A1(_02165_),
    .A2(_05822_),
    .B1(_05934_),
    .B2(_02102_),
    .Y(_06509_));
 NOR2x1_ASAP7_75t_R _25991_ (.A(_02022_),
    .B(_05949_),
    .Y(_06510_));
 AO21x1_ASAP7_75t_R _25992_ (.A1(net133),
    .A2(_05938_),
    .B(_06151_),
    .Y(_06511_));
 OAI22x1_ASAP7_75t_R _25993_ (.A1(_01823_),
    .A2(_05945_),
    .B1(_05943_),
    .B2(_01462_),
    .Y(_06512_));
 OA222x2_ASAP7_75t_R _25994_ (.A1(_01902_),
    .A2(_05814_),
    .B1(_05936_),
    .B2(_01990_),
    .C1(_05950_),
    .C2(_01952_),
    .Y(_06513_));
 OAI21x1_ASAP7_75t_R _25995_ (.A1(_01980_),
    .A2(_06189_),
    .B(_06513_),
    .Y(_06514_));
 OR4x2_ASAP7_75t_R _25996_ (.A(_06510_),
    .B(_06511_),
    .C(_06512_),
    .D(_06514_),
    .Y(_06515_));
 AO221x2_ASAP7_75t_R _25997_ (.A1(_05929_),
    .A2(_06508_),
    .B1(_06509_),
    .B2(_05976_),
    .C(_06515_),
    .Y(_06516_));
 OAI22x1_ASAP7_75t_R _25998_ (.A1(_05844_),
    .A2(_06507_),
    .B1(_06516_),
    .B2(_18630_),
    .Y(_06517_));
 OR3x2_ASAP7_75t_R _25999_ (.A(_02180_),
    .B(_02181_),
    .C(_06482_),
    .Y(_06518_));
 INVx1_ASAP7_75t_R _26000_ (.A(_06518_),
    .Y(_06519_));
 AO22x1_ASAP7_75t_R _26001_ (.A1(_05883_),
    .A2(_06517_),
    .B1(_06519_),
    .B2(_06467_),
    .Y(_06520_));
 AOI22x1_ASAP7_75t_R _26002_ (.A1(_02180_),
    .A2(_06505_),
    .B1(_06520_),
    .B2(_06472_),
    .Y(_02390_));
 NAND2x1_ASAP7_75t_R _26003_ (.A(_18861_),
    .B(_18633_),
    .Y(_06521_));
 OA21x2_ASAP7_75t_R _26004_ (.A1(_05846_),
    .A2(_18633_),
    .B(_06521_),
    .Y(_06522_));
 BUFx3_ASAP7_75t_R _26005_ (.A(_02116_),
    .Y(_06523_));
 OAI22x1_ASAP7_75t_R _26006_ (.A1(_02179_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_06523_),
    .Y(_06524_));
 OAI22x1_ASAP7_75t_R _26007_ (.A1(_02154_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_02091_),
    .Y(_06525_));
 OA222x2_ASAP7_75t_R _26008_ (.A1(_02021_),
    .A2(_05949_),
    .B1(_05937_),
    .B2(_01989_),
    .C1(_01463_),
    .C2(_05943_),
    .Y(_06526_));
 NAND2x1_ASAP7_75t_R _26009_ (.A(net134),
    .B(_05938_),
    .Y(_06527_));
 OA211x2_ASAP7_75t_R _26010_ (.A1(_01901_),
    .A2(_05941_),
    .B(_06527_),
    .C(_05769_),
    .Y(_06528_));
 OR2x2_ASAP7_75t_R _26011_ (.A(_01822_),
    .B(_05945_),
    .Y(_06529_));
 OA211x2_ASAP7_75t_R _26012_ (.A1(_01951_),
    .A2(_05951_),
    .B(_06528_),
    .C(_06529_),
    .Y(_06530_));
 NAND2x2_ASAP7_75t_R _26013_ (.A(_06526_),
    .B(_06530_),
    .Y(_06531_));
 AO221x2_ASAP7_75t_R _26014_ (.A1(_05930_),
    .A2(_06524_),
    .B1(_06525_),
    .B2(_06007_),
    .C(_06531_),
    .Y(_06532_));
 OA22x2_ASAP7_75t_R _26015_ (.A1(_05844_),
    .A2(_06522_),
    .B1(_06532_),
    .B2(_18633_),
    .Y(_06533_));
 BUFx10_ASAP7_75t_R _26016_ (.A(_06533_),
    .Y(_06534_));
 BUFx3_ASAP7_75t_R _26017_ (.A(_05970_),
    .Y(_06535_));
 AO32x1_ASAP7_75t_R _26018_ (.A1(_02179_),
    .A2(_06474_),
    .A3(_06519_),
    .B1(_06534_),
    .B2(_06535_),
    .Y(_06536_));
 NOR2x1_ASAP7_75t_R _26019_ (.A(_06473_),
    .B(_06518_),
    .Y(_06537_));
 OA21x2_ASAP7_75t_R _26020_ (.A1(_06113_),
    .A2(_06537_),
    .B(_06470_),
    .Y(_06538_));
 NOR2x1_ASAP7_75t_R _26021_ (.A(_02179_),
    .B(_06538_),
    .Y(_06539_));
 AO21x1_ASAP7_75t_R _26022_ (.A1(_06472_),
    .A2(_06536_),
    .B(_06539_),
    .Y(_02391_));
 INVx1_ASAP7_75t_R _26023_ (.A(_02178_),
    .Y(_06540_));
 OR3x1_ASAP7_75t_R _26024_ (.A(_02179_),
    .B(_06463_),
    .C(_06518_),
    .Y(_06541_));
 BUFx4f_ASAP7_75t_R _26025_ (.A(_06541_),
    .Y(_06542_));
 AO21x1_ASAP7_75t_R _26026_ (.A1(_05918_),
    .A2(_06542_),
    .B(_06465_),
    .Y(_06543_));
 NOR2x1_ASAP7_75t_R _26027_ (.A(_05970_),
    .B(_06542_),
    .Y(_06544_));
 NAND2x1_ASAP7_75t_R _26028_ (.A(_06074_),
    .B(_18637_),
    .Y(_06545_));
 OA21x2_ASAP7_75t_R _26029_ (.A1(_05846_),
    .A2(_18637_),
    .B(_06545_),
    .Y(_06546_));
 BUFx4f_ASAP7_75t_R _26030_ (.A(_02086_),
    .Y(_06547_));
 OAI22x1_ASAP7_75t_R _26031_ (.A1(_02149_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_06547_),
    .Y(_06548_));
 OAI22x1_ASAP7_75t_R _26032_ (.A1(_02178_),
    .A2(_05850_),
    .B1(_05852_),
    .B2(_02115_),
    .Y(_06549_));
 OA222x2_ASAP7_75t_R _26033_ (.A1(_01950_),
    .A2(_05985_),
    .B1(_05980_),
    .B2(_01821_),
    .C1(_01464_),
    .C2(_05858_),
    .Y(_06550_));
 INVx1_ASAP7_75t_R _26034_ (.A(net135),
    .Y(_06551_));
 OR2x2_ASAP7_75t_R _26035_ (.A(_01988_),
    .B(_05829_),
    .Y(_06552_));
 OA22x2_ASAP7_75t_R _26036_ (.A1(_02077_),
    .A2(_05827_),
    .B1(_05832_),
    .B2(_02020_),
    .Y(_06553_));
 OA211x2_ASAP7_75t_R _26037_ (.A1(_01900_),
    .A2(_05983_),
    .B(_05995_),
    .C(_06553_),
    .Y(_06554_));
 OA211x2_ASAP7_75t_R _26038_ (.A1(_06551_),
    .A2(_05989_),
    .B(_06552_),
    .C(_06554_),
    .Y(_06555_));
 NAND2x1_ASAP7_75t_R _26039_ (.A(_06550_),
    .B(_06555_),
    .Y(_06556_));
 AO221x2_ASAP7_75t_R _26040_ (.A1(_06007_),
    .A2(_06548_),
    .B1(_06549_),
    .B2(_05930_),
    .C(_06556_),
    .Y(_06557_));
 OA22x2_ASAP7_75t_R _26041_ (.A1(_05844_),
    .A2(_06546_),
    .B1(_06557_),
    .B2(_18637_),
    .Y(_06558_));
 BUFx6f_ASAP7_75t_R _26042_ (.A(_06558_),
    .Y(_06559_));
 AO22x1_ASAP7_75t_R _26043_ (.A1(_02178_),
    .A2(_06544_),
    .B1(_06559_),
    .B2(_06043_),
    .Y(_06560_));
 AO22x1_ASAP7_75t_R _26044_ (.A1(_06540_),
    .A2(_06543_),
    .B1(_06560_),
    .B2(_06471_),
    .Y(_02392_));
 BUFx4f_ASAP7_75t_R _26045_ (.A(_06470_),
    .Y(_06561_));
 AND5x2_ASAP7_75t_R _26046_ (.A(_14071_),
    .B(_05031_),
    .C(_05023_),
    .D(_05052_),
    .E(_06321_),
    .Y(_06562_));
 OR3x1_ASAP7_75t_R _26047_ (.A(_02179_),
    .B(_06473_),
    .C(_06518_),
    .Y(_06563_));
 BUFx6f_ASAP7_75t_R _26048_ (.A(_06563_),
    .Y(_06564_));
 AOI21x1_ASAP7_75t_R _26049_ (.A1(_05880_),
    .A2(_06562_),
    .B(_06564_),
    .Y(_06565_));
 NAND2x1_ASAP7_75t_R _26050_ (.A(_06074_),
    .B(_18642_),
    .Y(_06566_));
 OA21x2_ASAP7_75t_R _26051_ (.A1(_05846_),
    .A2(_18642_),
    .B(_06566_),
    .Y(_06567_));
 BUFx3_ASAP7_75t_R _26052_ (.A(_02114_),
    .Y(_06568_));
 OAI22x1_ASAP7_75t_R _26053_ (.A1(_02177_),
    .A2(_05849_),
    .B1(_05783_),
    .B2(_06568_),
    .Y(_06569_));
 OAI22x1_ASAP7_75t_R _26054_ (.A1(_02148_),
    .A2(_05779_),
    .B1(_05783_),
    .B2(_02085_),
    .Y(_06570_));
 OAI22x1_ASAP7_75t_R _26055_ (.A1(_02076_),
    .A2(_05827_),
    .B1(_05834_),
    .B2(_02019_),
    .Y(_06571_));
 NOR2x1_ASAP7_75t_R _26056_ (.A(_01899_),
    .B(_05814_),
    .Y(_06572_));
 AO221x1_ASAP7_75t_R _26057_ (.A1(net136),
    .A2(_05803_),
    .B1(_06105_),
    .B2(_05371_),
    .C(_06572_),
    .Y(_06573_));
 OAI21x1_ASAP7_75t_R _26058_ (.A1(_01851_),
    .A2(_06234_),
    .B(_05821_),
    .Y(_06574_));
 OAI22x1_ASAP7_75t_R _26059_ (.A1(_01949_),
    .A2(_05836_),
    .B1(_05857_),
    .B2(_02051_),
    .Y(_06575_));
 INVx1_ASAP7_75t_R _26060_ (.A(net196),
    .Y(_06576_));
 OR3x1_ASAP7_75t_R _26061_ (.A(_04948_),
    .B(_01820_),
    .C(_14308_),
    .Y(_06577_));
 OA21x2_ASAP7_75t_R _26062_ (.A1(_06576_),
    .A2(_04978_),
    .B(_06577_),
    .Y(_06578_));
 INVx1_ASAP7_75t_R _26063_ (.A(_05001_),
    .Y(_06579_));
 OAI22x1_ASAP7_75t_R _26064_ (.A1(_01987_),
    .A2(_05829_),
    .B1(_06578_),
    .B2(_06579_),
    .Y(_06580_));
 OR5x2_ASAP7_75t_R _26065_ (.A(_06571_),
    .B(_06573_),
    .C(_06574_),
    .D(_06575_),
    .E(_06580_),
    .Y(_06581_));
 AO221x2_ASAP7_75t_R _26066_ (.A1(_05798_),
    .A2(_06569_),
    .B1(_06570_),
    .B2(_05796_),
    .C(_06581_),
    .Y(_06582_));
 OA22x2_ASAP7_75t_R _26067_ (.A1(_05844_),
    .A2(_06567_),
    .B1(_06582_),
    .B2(_18642_),
    .Y(_06583_));
 BUFx6f_ASAP7_75t_R _26068_ (.A(_06583_),
    .Y(_06584_));
 AO32x1_ASAP7_75t_R _26069_ (.A1(_02177_),
    .A2(_06540_),
    .A3(_06565_),
    .B1(_06584_),
    .B2(_06535_),
    .Y(_06585_));
 OAI21x1_ASAP7_75t_R _26070_ (.A1(_02178_),
    .A2(_06564_),
    .B(_06350_),
    .Y(_06586_));
 AOI21x1_ASAP7_75t_R _26071_ (.A1(_06471_),
    .A2(_06586_),
    .B(_02177_),
    .Y(_06587_));
 AO21x1_ASAP7_75t_R _26072_ (.A1(_06561_),
    .A2(_06585_),
    .B(_06587_),
    .Y(_02393_));
 BUFx6f_ASAP7_75t_R _26073_ (.A(_06500_),
    .Y(_06588_));
 INVx1_ASAP7_75t_R _26074_ (.A(_05961_),
    .Y(_06589_));
 AND3x1_ASAP7_75t_R _26075_ (.A(_02176_),
    .B(_05921_),
    .C(_06589_),
    .Y(_06590_));
 AO21x1_ASAP7_75t_R _26076_ (.A1(_06047_),
    .A2(_06588_),
    .B(_06590_),
    .Y(_06591_));
 AO21x1_ASAP7_75t_R _26077_ (.A1(_06093_),
    .A2(_05961_),
    .B(_05893_),
    .Y(_06592_));
 INVx1_ASAP7_75t_R _26078_ (.A(_02176_),
    .Y(_06593_));
 AO22x1_ASAP7_75t_R _26079_ (.A1(_05959_),
    .A2(_06591_),
    .B1(_06592_),
    .B2(_06593_),
    .Y(_02394_));
 OR3x1_ASAP7_75t_R _26080_ (.A(_02177_),
    .B(_02178_),
    .C(_06542_),
    .Y(_06594_));
 AO21x1_ASAP7_75t_R _26081_ (.A1(_06116_),
    .A2(_06594_),
    .B(_06480_),
    .Y(_06595_));
 NAND2x1_ASAP7_75t_R _26082_ (.A(_05773_),
    .B(_18647_),
    .Y(_06596_));
 OA21x2_ASAP7_75t_R _26083_ (.A1(_06073_),
    .A2(_18647_),
    .B(_06596_),
    .Y(_06597_));
 OAI22x1_ASAP7_75t_R _26084_ (.A1(_02147_),
    .A2(_05778_),
    .B1(_05782_),
    .B2(_02084_),
    .Y(_06598_));
 OAI22x1_ASAP7_75t_R _26085_ (.A1(_02175_),
    .A2(_05778_),
    .B1(_05782_),
    .B2(_02112_),
    .Y(_06599_));
 INVx1_ASAP7_75t_R _26086_ (.A(_01465_),
    .Y(_06600_));
 NOR2x1_ASAP7_75t_R _26087_ (.A(_01986_),
    .B(_05828_),
    .Y(_06601_));
 AO221x1_ASAP7_75t_R _26088_ (.A1(net137),
    .A2(_05802_),
    .B1(_05810_),
    .B2(_06600_),
    .C(_06601_),
    .Y(_06602_));
 OAI22x1_ASAP7_75t_R _26089_ (.A1(_01898_),
    .A2(_05814_),
    .B1(_05827_),
    .B2(_02075_),
    .Y(_06603_));
 OAI22x1_ASAP7_75t_R _26090_ (.A1(_02018_),
    .A2(_05833_),
    .B1(_05857_),
    .B2(_02050_),
    .Y(_06604_));
 OAI22x1_ASAP7_75t_R _26091_ (.A1(_01819_),
    .A2(_05817_),
    .B1(_05836_),
    .B2(_01948_),
    .Y(_06605_));
 OR5x2_ASAP7_75t_R _26092_ (.A(_06428_),
    .B(_06602_),
    .C(_06603_),
    .D(_06604_),
    .E(_06605_),
    .Y(_06606_));
 AO221x2_ASAP7_75t_R _26093_ (.A1(_05795_),
    .A2(_06598_),
    .B1(_06599_),
    .B2(_05798_),
    .C(_06606_),
    .Y(_06607_));
 OA22x2_ASAP7_75t_R _26094_ (.A1(_06072_),
    .A2(_06597_),
    .B1(_06607_),
    .B2(_18647_),
    .Y(_06608_));
 BUFx6f_ASAP7_75t_R _26095_ (.A(_06608_),
    .Y(_06609_));
 INVx3_ASAP7_75t_R _26096_ (.A(_06609_),
    .Y(_06610_));
 OR3x2_ASAP7_75t_R _26097_ (.A(_02175_),
    .B(_02177_),
    .C(_02178_),
    .Y(_06611_));
 INVx1_ASAP7_75t_R _26098_ (.A(_06611_),
    .Y(_06612_));
 AO22x1_ASAP7_75t_R _26099_ (.A1(_05883_),
    .A2(_06610_),
    .B1(_06612_),
    .B2(_06544_),
    .Y(_06613_));
 AOI22x1_ASAP7_75t_R _26100_ (.A1(_02175_),
    .A2(_06595_),
    .B1(_06613_),
    .B2(_06472_),
    .Y(_02395_));
 NAND2x1_ASAP7_75t_R _26101_ (.A(_06074_),
    .B(_18653_),
    .Y(_06614_));
 OA21x2_ASAP7_75t_R _26102_ (.A1(_06073_),
    .A2(_18653_),
    .B(_06614_),
    .Y(_06615_));
 OAI22x1_ASAP7_75t_R _26103_ (.A1(_02146_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02083_),
    .Y(_06616_));
 OAI22x1_ASAP7_75t_R _26104_ (.A1(_02174_),
    .A2(_06147_),
    .B1(_06148_),
    .B2(_02111_),
    .Y(_06617_));
 OAI22x1_ASAP7_75t_R _26105_ (.A1(_01818_),
    .A2(_05817_),
    .B1(_05830_),
    .B2(_01985_),
    .Y(_06618_));
 OAI22x1_ASAP7_75t_R _26106_ (.A1(_02017_),
    .A2(_05834_),
    .B1(_05836_),
    .B2(_01947_),
    .Y(_06619_));
 NOR2x1_ASAP7_75t_R _26107_ (.A(_02049_),
    .B(_05858_),
    .Y(_06620_));
 INVx1_ASAP7_75t_R _26108_ (.A(_01466_),
    .Y(_06621_));
 AO22x1_ASAP7_75t_R _26109_ (.A1(net138),
    .A2(_05803_),
    .B1(_05811_),
    .B2(_06621_),
    .Y(_06622_));
 OAI21x1_ASAP7_75t_R _26110_ (.A1(_01897_),
    .A2(_05815_),
    .B(_05821_),
    .Y(_06623_));
 OR5x2_ASAP7_75t_R _26111_ (.A(_06618_),
    .B(_06619_),
    .C(_06620_),
    .D(_06622_),
    .E(_06623_),
    .Y(_06624_));
 AO221x2_ASAP7_75t_R _26112_ (.A1(_05796_),
    .A2(_06616_),
    .B1(_06617_),
    .B2(_05799_),
    .C(_06624_),
    .Y(_06625_));
 OA22x2_ASAP7_75t_R _26113_ (.A1(_06072_),
    .A2(_06615_),
    .B1(_06625_),
    .B2(_18653_),
    .Y(_06626_));
 BUFx6f_ASAP7_75t_R _26114_ (.A(_06626_),
    .Y(_06627_));
 AO32x1_ASAP7_75t_R _26115_ (.A1(_02174_),
    .A2(_06565_),
    .A3(_06612_),
    .B1(_06627_),
    .B2(_06535_),
    .Y(_06628_));
 BUFx6f_ASAP7_75t_R _26116_ (.A(_06470_),
    .Y(_06629_));
 OAI21x1_ASAP7_75t_R _26117_ (.A1(_06564_),
    .A2(_06611_),
    .B(_06350_),
    .Y(_06630_));
 AOI21x1_ASAP7_75t_R _26118_ (.A1(_06629_),
    .A2(_06630_),
    .B(_02174_),
    .Y(_06631_));
 AO21x1_ASAP7_75t_R _26119_ (.A1(_06561_),
    .A2(_06628_),
    .B(_06631_),
    .Y(_02396_));
 OR3x1_ASAP7_75t_R _26120_ (.A(_02174_),
    .B(_06542_),
    .C(_06611_),
    .Y(_06632_));
 AO21x1_ASAP7_75t_R _26121_ (.A1(_06116_),
    .A2(_06632_),
    .B(_06480_),
    .Y(_06633_));
 AND3x1_ASAP7_75t_R _26122_ (.A(_18659_),
    .B(_05933_),
    .C(_05953_),
    .Y(_06634_));
 AOI21x1_ASAP7_75t_R _26123_ (.A1(_05771_),
    .A2(_05955_),
    .B(_06634_),
    .Y(_06635_));
 OR3x2_ASAP7_75t_R _26124_ (.A(_02173_),
    .B(_02174_),
    .C(_06611_),
    .Y(_06636_));
 OR3x1_ASAP7_75t_R _26125_ (.A(_06144_),
    .B(_06542_),
    .C(_06636_),
    .Y(_06637_));
 OAI21x1_ASAP7_75t_R _26126_ (.A1(_06021_),
    .A2(_06635_),
    .B(_06637_),
    .Y(_06638_));
 AOI22x1_ASAP7_75t_R _26127_ (.A1(_02173_),
    .A2(_06633_),
    .B1(_06638_),
    .B2(_06472_),
    .Y(_02397_));
 INVx6_ASAP7_75t_R _26128_ (.A(_06000_),
    .Y(_06639_));
 NOR2x1_ASAP7_75t_R _26129_ (.A(_06564_),
    .B(_06636_),
    .Y(_06640_));
 AND3x1_ASAP7_75t_R _26130_ (.A(_02172_),
    .B(_05921_),
    .C(_06640_),
    .Y(_06641_));
 AO21x1_ASAP7_75t_R _26131_ (.A1(_06047_),
    .A2(_06639_),
    .B(_06641_),
    .Y(_06642_));
 OA21x2_ASAP7_75t_R _26132_ (.A1(_06113_),
    .A2(_06640_),
    .B(_06470_),
    .Y(_06643_));
 NOR2x1_ASAP7_75t_R _26133_ (.A(_02172_),
    .B(_06643_),
    .Y(_06644_));
 AO21x1_ASAP7_75t_R _26134_ (.A1(_06561_),
    .A2(_06642_),
    .B(_06644_),
    .Y(_02398_));
 OR3x1_ASAP7_75t_R _26135_ (.A(_02172_),
    .B(_06542_),
    .C(_06636_),
    .Y(_06645_));
 AO21x1_ASAP7_75t_R _26136_ (.A1(_06116_),
    .A2(_06645_),
    .B(_06480_),
    .Y(_06646_));
 OR3x2_ASAP7_75t_R _26137_ (.A(_02171_),
    .B(_02172_),
    .C(_06636_),
    .Y(_06647_));
 INVx1_ASAP7_75t_R _26138_ (.A(_06647_),
    .Y(_06648_));
 AO22x1_ASAP7_75t_R _26139_ (.A1(_05883_),
    .A2(_06017_),
    .B1(_06544_),
    .B2(_06648_),
    .Y(_06649_));
 AOI22x1_ASAP7_75t_R _26140_ (.A1(_02171_),
    .A2(_06646_),
    .B1(_06649_),
    .B2(_06472_),
    .Y(_02399_));
 BUFx6f_ASAP7_75t_R _26141_ (.A(_06042_),
    .Y(_06650_));
 AO32x1_ASAP7_75t_R _26142_ (.A1(_02170_),
    .A2(_06565_),
    .A3(_06648_),
    .B1(_06535_),
    .B2(_06650_),
    .Y(_06651_));
 OAI21x1_ASAP7_75t_R _26143_ (.A1(_06564_),
    .A2(_06647_),
    .B(_06350_),
    .Y(_06652_));
 AOI21x1_ASAP7_75t_R _26144_ (.A1(_06629_),
    .A2(_06652_),
    .B(_02170_),
    .Y(_06653_));
 AO21x1_ASAP7_75t_R _26145_ (.A1(_06561_),
    .A2(_06651_),
    .B(_06653_),
    .Y(_02400_));
 OR3x1_ASAP7_75t_R _26146_ (.A(_02170_),
    .B(_06542_),
    .C(_06647_),
    .Y(_06654_));
 AO21x1_ASAP7_75t_R _26147_ (.A1(_06116_),
    .A2(_06654_),
    .B(_06465_),
    .Y(_06655_));
 INVx2_ASAP7_75t_R _26148_ (.A(_06065_),
    .Y(_06656_));
 OR3x2_ASAP7_75t_R _26149_ (.A(_02169_),
    .B(_02170_),
    .C(_06647_),
    .Y(_06657_));
 INVx1_ASAP7_75t_R _26150_ (.A(_06657_),
    .Y(_06658_));
 AO22x1_ASAP7_75t_R _26151_ (.A1(_05883_),
    .A2(_06656_),
    .B1(_06544_),
    .B2(_06658_),
    .Y(_06659_));
 AOI22x1_ASAP7_75t_R _26152_ (.A1(_02169_),
    .A2(_06655_),
    .B1(_06659_),
    .B2(_06472_),
    .Y(_02401_));
 BUFx10_ASAP7_75t_R _26153_ (.A(_06088_),
    .Y(_06660_));
 AO32x1_ASAP7_75t_R _26154_ (.A1(_02168_),
    .A2(_06565_),
    .A3(_06658_),
    .B1(_06535_),
    .B2(_06660_),
    .Y(_06661_));
 OAI21x1_ASAP7_75t_R _26155_ (.A1(_06564_),
    .A2(_06657_),
    .B(_06350_),
    .Y(_06662_));
 AOI21x1_ASAP7_75t_R _26156_ (.A1(_06629_),
    .A2(_06662_),
    .B(_02168_),
    .Y(_06663_));
 AO21x1_ASAP7_75t_R _26157_ (.A1(_06561_),
    .A2(_06661_),
    .B(_06663_),
    .Y(_02402_));
 OR3x1_ASAP7_75t_R _26158_ (.A(_02168_),
    .B(_06542_),
    .C(_06657_),
    .Y(_06664_));
 AO21x1_ASAP7_75t_R _26159_ (.A1(_06093_),
    .A2(_06664_),
    .B(_06465_),
    .Y(_06665_));
 OR3x4_ASAP7_75t_R _26160_ (.A(_02167_),
    .B(_02168_),
    .C(_06657_),
    .Y(_06666_));
 OR2x2_ASAP7_75t_R _26161_ (.A(_06541_),
    .B(_06666_),
    .Y(_06667_));
 BUFx4f_ASAP7_75t_R _26162_ (.A(_06667_),
    .Y(_06668_));
 NOR2x2_ASAP7_75t_R _26163_ (.A(_05970_),
    .B(_06668_),
    .Y(_06669_));
 AO21x1_ASAP7_75t_R _26164_ (.A1(_05883_),
    .A2(_06112_),
    .B(_06669_),
    .Y(_06670_));
 AOI22x1_ASAP7_75t_R _26165_ (.A1(_02167_),
    .A2(_06665_),
    .B1(_06670_),
    .B2(_06472_),
    .Y(_02403_));
 NOR2x2_ASAP7_75t_R _26166_ (.A(_06564_),
    .B(_06666_),
    .Y(_06671_));
 OA21x2_ASAP7_75t_R _26167_ (.A1(_06047_),
    .A2(_06671_),
    .B(_06470_),
    .Y(_06672_));
 AND2x2_ASAP7_75t_R _26168_ (.A(_05887_),
    .B(_06671_),
    .Y(_06673_));
 AOI22x1_ASAP7_75t_R _26169_ (.A1(_06047_),
    .A2(_06137_),
    .B1(_06673_),
    .B2(_06121_),
    .Y(_06674_));
 OAI22x1_ASAP7_75t_R _26170_ (.A1(_06121_),
    .A2(_06672_),
    .B1(_06674_),
    .B2(_06480_),
    .Y(_02404_));
 INVx1_ASAP7_75t_R _26171_ (.A(_02165_),
    .Y(_06675_));
 OR3x1_ASAP7_75t_R _26172_ (.A(_06675_),
    .B(_06113_),
    .C(_05923_),
    .Y(_06676_));
 OAI21x1_ASAP7_75t_R _26173_ (.A1(_06093_),
    .A2(_06517_),
    .B(_06676_),
    .Y(_06677_));
 AO21x1_ASAP7_75t_R _26174_ (.A1(_06025_),
    .A2(_05923_),
    .B(_05893_),
    .Y(_06678_));
 AO22x1_ASAP7_75t_R _26175_ (.A1(_06045_),
    .A2(_06677_),
    .B1(_06678_),
    .B2(_06675_),
    .Y(_02405_));
 OAI21x1_ASAP7_75t_R _26176_ (.A1(_06121_),
    .A2(_06668_),
    .B(_05887_),
    .Y(_06679_));
 AO21x1_ASAP7_75t_R _26177_ (.A1(_06470_),
    .A2(_06679_),
    .B(_02164_),
    .Y(_06680_));
 INVx1_ASAP7_75t_R _26178_ (.A(_02164_),
    .Y(_06681_));
 OR2x2_ASAP7_75t_R _26179_ (.A(_05969_),
    .B(_06668_),
    .Y(_06682_));
 OR3x1_ASAP7_75t_R _26180_ (.A(_06681_),
    .B(_06121_),
    .C(_06682_),
    .Y(_06683_));
 AO21x1_ASAP7_75t_R _26181_ (.A1(_06162_),
    .A2(_06683_),
    .B(_06465_),
    .Y(_06684_));
 NAND2x1_ASAP7_75t_R _26182_ (.A(_06680_),
    .B(_06684_),
    .Y(_02406_));
 NOR2x1_ASAP7_75t_R _26183_ (.A(_02164_),
    .B(_06121_),
    .Y(_06685_));
 AO32x1_ASAP7_75t_R _26184_ (.A1(_02163_),
    .A2(_06673_),
    .A3(_06685_),
    .B1(_06535_),
    .B2(_06180_),
    .Y(_06686_));
 AO21x1_ASAP7_75t_R _26185_ (.A1(_06671_),
    .A2(_06685_),
    .B(_06144_),
    .Y(_06687_));
 AOI21x1_ASAP7_75t_R _26186_ (.A1(_06629_),
    .A2(_06687_),
    .B(_02163_),
    .Y(_06688_));
 AO21x1_ASAP7_75t_R _26187_ (.A1(_06561_),
    .A2(_06686_),
    .B(_06688_),
    .Y(_02407_));
 OR3x4_ASAP7_75t_R _26188_ (.A(_02163_),
    .B(_02164_),
    .C(_06121_),
    .Y(_06689_));
 INVx1_ASAP7_75t_R _26189_ (.A(_06689_),
    .Y(_06690_));
 AO32x1_ASAP7_75t_R _26190_ (.A1(_02162_),
    .A2(_06669_),
    .A3(_06690_),
    .B1(_06535_),
    .B2(_06218_),
    .Y(_06691_));
 OAI21x1_ASAP7_75t_R _26191_ (.A1(_06668_),
    .A2(_06689_),
    .B(_06350_),
    .Y(_06692_));
 AOI21x1_ASAP7_75t_R _26192_ (.A1(_06629_),
    .A2(_06692_),
    .B(_02162_),
    .Y(_06693_));
 AO21x1_ASAP7_75t_R _26193_ (.A1(_06561_),
    .A2(_06691_),
    .B(_06693_),
    .Y(_02408_));
 NOR2x1_ASAP7_75t_R _26194_ (.A(_02162_),
    .B(_06689_),
    .Y(_06694_));
 BUFx10_ASAP7_75t_R _26195_ (.A(_06241_),
    .Y(_06695_));
 AO32x1_ASAP7_75t_R _26196_ (.A1(_02161_),
    .A2(_06673_),
    .A3(_06694_),
    .B1(_06535_),
    .B2(_06695_),
    .Y(_06696_));
 AO21x1_ASAP7_75t_R _26197_ (.A1(_06671_),
    .A2(_06694_),
    .B(_06144_),
    .Y(_06697_));
 AOI21x1_ASAP7_75t_R _26198_ (.A1(_06629_),
    .A2(_06697_),
    .B(_02161_),
    .Y(_06698_));
 AO21x1_ASAP7_75t_R _26199_ (.A1(_06561_),
    .A2(_06696_),
    .B(_06698_),
    .Y(_02409_));
 OR3x4_ASAP7_75t_R _26200_ (.A(_02161_),
    .B(_02162_),
    .C(_06689_),
    .Y(_06699_));
 INVx1_ASAP7_75t_R _26201_ (.A(_06699_),
    .Y(_06700_));
 AO32x1_ASAP7_75t_R _26202_ (.A1(_02160_),
    .A2(_06669_),
    .A3(_06700_),
    .B1(_06535_),
    .B2(_06260_),
    .Y(_06701_));
 OAI21x1_ASAP7_75t_R _26203_ (.A1(_06668_),
    .A2(_06699_),
    .B(_06350_),
    .Y(_06702_));
 AOI21x1_ASAP7_75t_R _26204_ (.A1(_06629_),
    .A2(_06702_),
    .B(_02160_),
    .Y(_06703_));
 AO21x1_ASAP7_75t_R _26205_ (.A1(_06561_),
    .A2(_06701_),
    .B(_06703_),
    .Y(_02410_));
 NOR2x1_ASAP7_75t_R _26206_ (.A(_02160_),
    .B(_06699_),
    .Y(_06704_));
 BUFx12_ASAP7_75t_R _26207_ (.A(_06280_),
    .Y(_06705_));
 AO32x1_ASAP7_75t_R _26208_ (.A1(_02159_),
    .A2(_06673_),
    .A3(_06704_),
    .B1(_06535_),
    .B2(_06705_),
    .Y(_06706_));
 AO21x1_ASAP7_75t_R _26209_ (.A1(_06671_),
    .A2(_06704_),
    .B(_06144_),
    .Y(_06707_));
 AOI21x1_ASAP7_75t_R _26210_ (.A1(_06629_),
    .A2(_06707_),
    .B(_02159_),
    .Y(_06708_));
 AO21x1_ASAP7_75t_R _26211_ (.A1(_06561_),
    .A2(_06706_),
    .B(_06708_),
    .Y(_02411_));
 OR3x4_ASAP7_75t_R _26212_ (.A(_02159_),
    .B(_02160_),
    .C(_06699_),
    .Y(_06709_));
 INVx1_ASAP7_75t_R _26213_ (.A(_06709_),
    .Y(_06710_));
 AO32x1_ASAP7_75t_R _26214_ (.A1(_02158_),
    .A2(_06669_),
    .A3(_06710_),
    .B1(_06043_),
    .B2(_06298_),
    .Y(_06711_));
 OAI21x1_ASAP7_75t_R _26215_ (.A1(_06668_),
    .A2(_06709_),
    .B(_06350_),
    .Y(_06712_));
 AOI21x1_ASAP7_75t_R _26216_ (.A1(_06629_),
    .A2(_06712_),
    .B(_02158_),
    .Y(_06713_));
 AO21x1_ASAP7_75t_R _26217_ (.A1(_06471_),
    .A2(_06711_),
    .B(_06713_),
    .Y(_02412_));
 NOR2x1_ASAP7_75t_R _26218_ (.A(_02158_),
    .B(_06709_),
    .Y(_06714_));
 AO32x1_ASAP7_75t_R _26219_ (.A1(_02157_),
    .A2(_06673_),
    .A3(_06714_),
    .B1(_06043_),
    .B2(_06320_),
    .Y(_06715_));
 AO21x1_ASAP7_75t_R _26220_ (.A1(_06671_),
    .A2(_06714_),
    .B(_06144_),
    .Y(_06716_));
 AOI21x1_ASAP7_75t_R _26221_ (.A1(_06629_),
    .A2(_06716_),
    .B(_02157_),
    .Y(_06717_));
 AO21x1_ASAP7_75t_R _26222_ (.A1(_06471_),
    .A2(_06715_),
    .B(_06717_),
    .Y(_02413_));
 INVx1_ASAP7_75t_R _26223_ (.A(_02156_),
    .Y(_06718_));
 OR3x1_ASAP7_75t_R _26224_ (.A(_02157_),
    .B(_02158_),
    .C(_06709_),
    .Y(_06719_));
 OR3x1_ASAP7_75t_R _26225_ (.A(_06542_),
    .B(_06666_),
    .C(_06719_),
    .Y(_06720_));
 AO21x1_ASAP7_75t_R _26226_ (.A1(_06093_),
    .A2(_06720_),
    .B(_06465_),
    .Y(_06721_));
 OR3x1_ASAP7_75t_R _26227_ (.A(_06718_),
    .B(_06682_),
    .C(_06719_),
    .Y(_06722_));
 AOI21x1_ASAP7_75t_R _26228_ (.A1(_06348_),
    .A2(_06722_),
    .B(_06480_),
    .Y(_06723_));
 AO21x1_ASAP7_75t_R _26229_ (.A1(_06718_),
    .A2(_06721_),
    .B(_06723_),
    .Y(_02414_));
 OR2x2_ASAP7_75t_R _26230_ (.A(_02156_),
    .B(_06719_),
    .Y(_06724_));
 OR3x4_ASAP7_75t_R _26231_ (.A(_06564_),
    .B(_06666_),
    .C(_06724_),
    .Y(_06725_));
 AOI21x1_ASAP7_75t_R _26232_ (.A1(_05922_),
    .A2(_06725_),
    .B(_06480_),
    .Y(_06726_));
 INVx1_ASAP7_75t_R _26233_ (.A(_06358_),
    .Y(_06727_));
 OR3x1_ASAP7_75t_R _26234_ (.A(_06727_),
    .B(_06113_),
    .C(_06725_),
    .Y(_06728_));
 AO21x1_ASAP7_75t_R _26235_ (.A1(_06371_),
    .A2(_06728_),
    .B(_06480_),
    .Y(_06729_));
 OAI21x1_ASAP7_75t_R _26236_ (.A1(_06358_),
    .A2(_06726_),
    .B(_06729_),
    .Y(_02415_));
 AND5x1_ASAP7_75t_R _26237_ (.A(_02154_),
    .B(_06675_),
    .C(_06593_),
    .D(_05921_),
    .E(_06589_),
    .Y(_06730_));
 AO21x1_ASAP7_75t_R _26238_ (.A1(_06047_),
    .A2(_06534_),
    .B(_06730_),
    .Y(_06731_));
 AO21x1_ASAP7_75t_R _26239_ (.A1(_06025_),
    .A2(_05962_),
    .B(_05893_),
    .Y(_06732_));
 INVx1_ASAP7_75t_R _26240_ (.A(_02154_),
    .Y(_06733_));
 AO22x1_ASAP7_75t_R _26241_ (.A1(_06045_),
    .A2(_06731_),
    .B1(_06732_),
    .B2(_06733_),
    .Y(_02416_));
 INVx1_ASAP7_75t_R _26242_ (.A(_02153_),
    .Y(_06734_));
 OR3x1_ASAP7_75t_R _26243_ (.A(_06358_),
    .B(_06668_),
    .C(_06724_),
    .Y(_06735_));
 AO21x1_ASAP7_75t_R _26244_ (.A1(_05918_),
    .A2(_06735_),
    .B(_06465_),
    .Y(_06736_));
 NOR2x1_ASAP7_75t_R _26245_ (.A(_06358_),
    .B(_06724_),
    .Y(_06737_));
 BUFx10_ASAP7_75t_R _26246_ (.A(_06392_),
    .Y(_06738_));
 AO32x1_ASAP7_75t_R _26247_ (.A1(_02153_),
    .A2(_06669_),
    .A3(_06737_),
    .B1(_06144_),
    .B2(_06738_),
    .Y(_06739_));
 AO22x1_ASAP7_75t_R _26248_ (.A1(_06734_),
    .A2(_06736_),
    .B1(_06739_),
    .B2(_06471_),
    .Y(_02417_));
 INVx1_ASAP7_75t_R _26249_ (.A(_02152_),
    .Y(_06740_));
 OR3x1_ASAP7_75t_R _26250_ (.A(_02153_),
    .B(_06358_),
    .C(_06725_),
    .Y(_06741_));
 AO21x1_ASAP7_75t_R _26251_ (.A1(_06093_),
    .A2(_06741_),
    .B(_06465_),
    .Y(_06742_));
 OR5x1_ASAP7_75t_R _26252_ (.A(_06740_),
    .B(_02153_),
    .C(_06358_),
    .D(_05970_),
    .E(_06725_),
    .Y(_06743_));
 AOI21x1_ASAP7_75t_R _26253_ (.A1(_06412_),
    .A2(_06743_),
    .B(_06480_),
    .Y(_06744_));
 AO21x1_ASAP7_75t_R _26254_ (.A1(_06740_),
    .A2(_06742_),
    .B(_06744_),
    .Y(_02418_));
 INVx1_ASAP7_75t_R _26255_ (.A(_02151_),
    .Y(_06745_));
 OR4x1_ASAP7_75t_R _26256_ (.A(_02152_),
    .B(_02153_),
    .C(_06358_),
    .D(_06724_),
    .Y(_06746_));
 OR3x1_ASAP7_75t_R _26257_ (.A(_06542_),
    .B(_06666_),
    .C(_06746_),
    .Y(_06747_));
 AO21x1_ASAP7_75t_R _26258_ (.A1(_05918_),
    .A2(_06747_),
    .B(_06465_),
    .Y(_06748_));
 INVx1_ASAP7_75t_R _26259_ (.A(_06746_),
    .Y(_06749_));
 BUFx10_ASAP7_75t_R _26260_ (.A(_06439_),
    .Y(_06750_));
 AO32x1_ASAP7_75t_R _26261_ (.A1(_02151_),
    .A2(_06669_),
    .A3(_06749_),
    .B1(_06144_),
    .B2(_06750_),
    .Y(_06751_));
 AO22x1_ASAP7_75t_R _26262_ (.A1(_06745_),
    .A2(_06748_),
    .B1(_06751_),
    .B2(_06471_),
    .Y(_02419_));
 INVx1_ASAP7_75t_R _26263_ (.A(_02150_),
    .Y(_06752_));
 OR5x1_ASAP7_75t_R _26264_ (.A(_02151_),
    .B(_02152_),
    .C(_02153_),
    .D(_06358_),
    .E(_06725_),
    .Y(_06753_));
 AO21x1_ASAP7_75t_R _26265_ (.A1(_05918_),
    .A2(_06753_),
    .B(_06465_),
    .Y(_06754_));
 OR3x1_ASAP7_75t_R _26266_ (.A(_06752_),
    .B(_06113_),
    .C(_06753_),
    .Y(_06755_));
 OAI21x1_ASAP7_75t_R _26267_ (.A1(_06093_),
    .A2(_06455_),
    .B(_06755_),
    .Y(_06756_));
 AO22x1_ASAP7_75t_R _26268_ (.A1(_06752_),
    .A2(_06754_),
    .B1(_06756_),
    .B2(_06471_),
    .Y(_02420_));
 AO21x1_ASAP7_75t_R _26269_ (.A1(_06093_),
    .A2(_05924_),
    .B(_05926_),
    .Y(_06757_));
 OR3x1_ASAP7_75t_R _26270_ (.A(_02149_),
    .B(_05882_),
    .C(_05924_),
    .Y(_06758_));
 OAI21x1_ASAP7_75t_R _26271_ (.A1(_06021_),
    .A2(_06559_),
    .B(_06758_),
    .Y(_06759_));
 AOI22x1_ASAP7_75t_R _26272_ (.A1(_02149_),
    .A2(_06757_),
    .B1(_06759_),
    .B2(_05959_),
    .Y(_02421_));
 NOR2x1_ASAP7_75t_R _26273_ (.A(_06113_),
    .B(_05963_),
    .Y(_06760_));
 AO22x1_ASAP7_75t_R _26274_ (.A1(_06043_),
    .A2(_06583_),
    .B1(_06760_),
    .B2(_02148_),
    .Y(_06761_));
 AO21x1_ASAP7_75t_R _26275_ (.A1(_06025_),
    .A2(_05963_),
    .B(_05893_),
    .Y(_06762_));
 INVx1_ASAP7_75t_R _26276_ (.A(_02148_),
    .Y(_06763_));
 AO22x1_ASAP7_75t_R _26277_ (.A1(_06045_),
    .A2(_06761_),
    .B1(_06762_),
    .B2(_06763_),
    .Y(_02422_));
 INVx1_ASAP7_75t_R _26278_ (.A(_02147_),
    .Y(_06764_));
 OR3x1_ASAP7_75t_R _26279_ (.A(_02148_),
    .B(_02149_),
    .C(_05924_),
    .Y(_06765_));
 OR3x1_ASAP7_75t_R _26280_ (.A(_06764_),
    .B(_06113_),
    .C(_06765_),
    .Y(_06766_));
 OA21x2_ASAP7_75t_R _26281_ (.A1(_06093_),
    .A2(_06610_),
    .B(_06766_),
    .Y(_06767_));
 AOI21x1_ASAP7_75t_R _26282_ (.A1(_05922_),
    .A2(_06765_),
    .B(_06002_),
    .Y(_06768_));
 OAI22x1_ASAP7_75t_R _26283_ (.A1(_06002_),
    .A2(_06767_),
    .B1(_06768_),
    .B2(_02147_),
    .Y(_02423_));
 INVx1_ASAP7_75t_R _26284_ (.A(_02146_),
    .Y(_06769_));
 AOI21x1_ASAP7_75t_R _26285_ (.A1(_05922_),
    .A2(_05964_),
    .B(_05926_),
    .Y(_06770_));
 OR3x1_ASAP7_75t_R _26286_ (.A(_02146_),
    .B(_05882_),
    .C(_05964_),
    .Y(_06771_));
 OA21x2_ASAP7_75t_R _26287_ (.A1(_06350_),
    .A2(_06627_),
    .B(_06771_),
    .Y(_06772_));
 OA22x2_ASAP7_75t_R _26288_ (.A1(_06769_),
    .A2(_06770_),
    .B1(_06772_),
    .B2(_06002_),
    .Y(_02424_));
 XNOR2x1_ASAP7_75t_R _26289_ (.B(_04975_),
    .Y(_06773_),
    .A(_04976_));
 AND4x1_ASAP7_75t_R _26290_ (.A(_02305_),
    .B(_02304_),
    .C(_18608_),
    .D(_14070_),
    .Y(_06774_));
 AOI211x1_ASAP7_75t_R _26291_ (.A1(_13367_),
    .A2(_13553_),
    .B(_18610_),
    .C(_18617_),
    .Y(_06775_));
 XNOR2x1_ASAP7_75t_R _26292_ (.B(_06775_),
    .Y(_06776_),
    .A(_18623_));
 AND3x2_ASAP7_75t_R _26293_ (.A(_06773_),
    .B(_06774_),
    .C(_06776_),
    .Y(_06777_));
 BUFx6f_ASAP7_75t_R _26294_ (.A(_06777_),
    .Y(_06778_));
 AND3x4_ASAP7_75t_R _26295_ (.A(_05974_),
    .B(_06323_),
    .C(_06778_),
    .Y(_06779_));
 AND3x1_ASAP7_75t_R _26296_ (.A(_14026_),
    .B(_04925_),
    .C(_04926_),
    .Y(_06780_));
 NAND2x1_ASAP7_75t_R _26297_ (.A(_13368_),
    .B(_04923_),
    .Y(_06781_));
 INVx1_ASAP7_75t_R _26298_ (.A(_04923_),
    .Y(_06782_));
 AO32x1_ASAP7_75t_R _26299_ (.A1(_02218_),
    .A2(_16286_),
    .A3(_05149_),
    .B1(_06780_),
    .B2(_06782_),
    .Y(_06783_));
 OR3x1_ASAP7_75t_R _26300_ (.A(_13570_),
    .B(_05304_),
    .C(_05321_),
    .Y(_06784_));
 AND3x1_ASAP7_75t_R _26301_ (.A(_04927_),
    .B(_06783_),
    .C(_06784_),
    .Y(_06785_));
 AO21x1_ASAP7_75t_R _26302_ (.A1(_01776_),
    .A2(_05322_),
    .B(_06785_),
    .Y(_06786_));
 AO32x2_ASAP7_75t_R _26303_ (.A1(_13407_),
    .A2(_06780_),
    .A3(_06781_),
    .B1(_06786_),
    .B2(_04940_),
    .Y(_06787_));
 INVx1_ASAP7_75t_R _26304_ (.A(_01451_),
    .Y(_06788_));
 AND3x2_ASAP7_75t_R _26305_ (.A(_13568_),
    .B(_13570_),
    .C(_14894_),
    .Y(_06789_));
 AOI211x1_ASAP7_75t_R _26306_ (.A1(_13585_),
    .A2(_14019_),
    .B(_13624_),
    .C(_13621_),
    .Y(_06790_));
 AOI211x1_ASAP7_75t_R _26307_ (.A1(_13571_),
    .A2(_13594_),
    .B(_14906_),
    .C(_06790_),
    .Y(_06791_));
 AND4x1_ASAP7_75t_R _26308_ (.A(_14887_),
    .B(_14891_),
    .C(_14897_),
    .D(_06791_),
    .Y(_06792_));
 BUFx3_ASAP7_75t_R _26309_ (.A(_06792_),
    .Y(_06793_));
 BUFx3_ASAP7_75t_R _26310_ (.A(_01450_),
    .Y(_06794_));
 AND2x2_ASAP7_75t_R _26311_ (.A(net1990),
    .B(_06794_),
    .Y(_06795_));
 OAI22x1_ASAP7_75t_R _26312_ (.A1(net1996),
    .A2(_14904_),
    .B1(_06793_),
    .B2(_06795_),
    .Y(_06796_));
 NAND2x2_ASAP7_75t_R _26313_ (.A(_06789_),
    .B(_06796_),
    .Y(_06797_));
 NAND2x2_ASAP7_75t_R _26314_ (.A(_13571_),
    .B(_14894_),
    .Y(_06798_));
 AOI211x1_ASAP7_75t_R _26315_ (.A1(_14904_),
    .A2(_06793_),
    .B(_06798_),
    .C(net1990),
    .Y(_06799_));
 INVx1_ASAP7_75t_R _26316_ (.A(net1995),
    .Y(_06800_));
 AO32x1_ASAP7_75t_R _26317_ (.A1(_06800_),
    .A2(_06789_),
    .A3(_06793_),
    .B1(_14919_),
    .B2(_15251_),
    .Y(_06801_));
 NOR2x2_ASAP7_75t_R _26318_ (.A(_06799_),
    .B(_06801_),
    .Y(_06802_));
 XOR2x1_ASAP7_75t_R _26319_ (.A(_18845_),
    .Y(_06803_),
    .B(_06802_));
 AND5x1_ASAP7_75t_R _26320_ (.A(_01451_),
    .B(_04899_),
    .C(_04905_),
    .D(_04906_),
    .E(_06797_),
    .Y(_06804_));
 AO33x2_ASAP7_75t_R _26321_ (.A1(_06788_),
    .A2(_06797_),
    .A3(_06803_),
    .B1(_06804_),
    .B2(_04890_),
    .B3(_04887_),
    .Y(_06805_));
 AND3x1_ASAP7_75t_R _26322_ (.A(_01451_),
    .B(_04897_),
    .C(_06797_),
    .Y(_06806_));
 OA31x2_ASAP7_75t_R _26323_ (.A1(_04900_),
    .A2(_04902_),
    .A3(_04907_),
    .B1(_06806_),
    .Y(_06807_));
 OR2x4_ASAP7_75t_R _26324_ (.A(_06805_),
    .B(_06807_),
    .Y(_06808_));
 AND2x2_ASAP7_75t_R _26325_ (.A(_04899_),
    .B(_05110_),
    .Y(_06809_));
 INVx2_ASAP7_75t_R _26326_ (.A(_02295_),
    .Y(_06810_));
 NAND2x1_ASAP7_75t_R _26327_ (.A(_06810_),
    .B(_06789_),
    .Y(_06811_));
 OA21x2_ASAP7_75t_R _26328_ (.A1(_15262_),
    .A2(_06795_),
    .B(_06811_),
    .Y(_06812_));
 NAND2x1_ASAP7_75t_R _26329_ (.A(net1990),
    .B(_06794_),
    .Y(_06813_));
 AND2x2_ASAP7_75t_R _26330_ (.A(_06800_),
    .B(_14904_),
    .Y(_06814_));
 AOI22x1_ASAP7_75t_R _26331_ (.A1(_14912_),
    .A2(_06813_),
    .B1(_06814_),
    .B2(_06793_),
    .Y(_06815_));
 OA22x2_ASAP7_75t_R _26332_ (.A1(_06793_),
    .A2(_06812_),
    .B1(_06815_),
    .B2(_06798_),
    .Y(_06816_));
 AND3x1_ASAP7_75t_R _26333_ (.A(_01451_),
    .B(_04899_),
    .C(_06816_),
    .Y(_06817_));
 NAND2x1_ASAP7_75t_R _26334_ (.A(_04887_),
    .B(_04890_),
    .Y(_06818_));
 XNOR2x1_ASAP7_75t_R _26335_ (.B(_06802_),
    .Y(_06819_),
    .A(_18845_));
 AND5x1_ASAP7_75t_R _26336_ (.A(_01451_),
    .B(_04897_),
    .C(_04905_),
    .D(_04906_),
    .E(_06816_),
    .Y(_06820_));
 AO33x2_ASAP7_75t_R _26337_ (.A1(_06788_),
    .A2(_06816_),
    .A3(_06819_),
    .B1(_06820_),
    .B2(_04890_),
    .B3(_04887_),
    .Y(_06821_));
 AO221x2_ASAP7_75t_R _26338_ (.A1(_01451_),
    .A2(_06809_),
    .B1(_06817_),
    .B2(_06818_),
    .C(_06821_),
    .Y(_06822_));
 OR3x4_ASAP7_75t_R _26339_ (.A(_02295_),
    .B(_14904_),
    .C(_06798_),
    .Y(_06823_));
 NAND3x2_ASAP7_75t_R _26340_ (.B(_06797_),
    .C(_06823_),
    .Y(_06824_),
    .A(_06816_));
 OAI21x1_ASAP7_75t_R _26341_ (.A1(_06808_),
    .A2(_06822_),
    .B(_06824_),
    .Y(_06825_));
 AND3x1_ASAP7_75t_R _26342_ (.A(_13570_),
    .B(_04928_),
    .C(_05753_),
    .Y(_06826_));
 AND4x2_ASAP7_75t_R _26343_ (.A(_05135_),
    .B(_05136_),
    .C(_06825_),
    .D(_06826_),
    .Y(_06827_));
 OAI21x1_ASAP7_75t_R _26344_ (.A1(_06808_),
    .A2(_06822_),
    .B(_06823_),
    .Y(_06828_));
 OA211x2_ASAP7_75t_R _26345_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_05131_),
    .B(_06828_),
    .C(_06826_),
    .Y(_06829_));
 NOR3x2_ASAP7_75t_R _26346_ (.B(_06827_),
    .C(_06829_),
    .Y(_06830_),
    .A(_06787_));
 BUFx12_ASAP7_75t_R _26347_ (.A(_06830_),
    .Y(_06831_));
 AND3x1_ASAP7_75t_R _26348_ (.A(_02310_),
    .B(_18658_),
    .C(_18663_),
    .Y(_06832_));
 OAI21x1_ASAP7_75t_R _26349_ (.A1(_05058_),
    .A2(_06832_),
    .B(_14071_),
    .Y(_06833_));
 NAND2x1_ASAP7_75t_R _26350_ (.A(_04921_),
    .B(_04923_),
    .Y(_06834_));
 AND3x1_ASAP7_75t_R _26351_ (.A(_01453_),
    .B(_06834_),
    .C(_05084_),
    .Y(_06835_));
 AND3x4_ASAP7_75t_R _26352_ (.A(_05097_),
    .B(_06833_),
    .C(_06835_),
    .Y(_06836_));
 NAND2x2_ASAP7_75t_R _26353_ (.A(_06323_),
    .B(_06778_),
    .Y(_06837_));
 AND3x4_ASAP7_75t_R _26354_ (.A(_06831_),
    .B(_06836_),
    .C(_06837_),
    .Y(_06838_));
 AO31x2_ASAP7_75t_R _26355_ (.A1(_06831_),
    .A2(_06836_),
    .A3(_06837_),
    .B(_06779_),
    .Y(_06839_));
 BUFx6f_ASAP7_75t_R _26356_ (.A(_06839_),
    .Y(_06840_));
 NOR2x1_ASAP7_75t_R _26357_ (.A(_00787_),
    .B(_06840_),
    .Y(_06841_));
 AO221x1_ASAP7_75t_R _26358_ (.A1(_05841_),
    .A2(_06779_),
    .B1(_06838_),
    .B2(_00787_),
    .C(_06841_),
    .Y(_02425_));
 AND4x1_ASAP7_75t_R _26359_ (.A(_04971_),
    .B(_05031_),
    .C(_05794_),
    .D(_05915_),
    .Y(_06842_));
 NAND2x2_ASAP7_75t_R _26360_ (.A(_06842_),
    .B(_06778_),
    .Y(_06843_));
 BUFx6f_ASAP7_75t_R _26361_ (.A(_06843_),
    .Y(_06844_));
 BUFx6f_ASAP7_75t_R _26362_ (.A(_06844_),
    .Y(_06845_));
 OR4x2_ASAP7_75t_R _26363_ (.A(_02083_),
    .B(_02084_),
    .C(_02085_),
    .D(_06547_),
    .Y(_06846_));
 OR2x2_ASAP7_75t_R _26364_ (.A(_02145_),
    .B(_06846_),
    .Y(_06847_));
 AND3x4_ASAP7_75t_R _26365_ (.A(_05876_),
    .B(_06321_),
    .C(_06777_),
    .Y(_06848_));
 BUFx4f_ASAP7_75t_R _26366_ (.A(_06848_),
    .Y(_06849_));
 OR3x1_ASAP7_75t_R _26367_ (.A(_02113_),
    .B(_02124_),
    .C(_02311_),
    .Y(_06850_));
 OR3x4_ASAP7_75t_R _26368_ (.A(_02091_),
    .B(_02102_),
    .C(_06850_),
    .Y(_06851_));
 OR2x4_ASAP7_75t_R _26369_ (.A(_06849_),
    .B(_06851_),
    .Y(_06852_));
 OA22x2_ASAP7_75t_R _26370_ (.A1(_06635_),
    .A2(_06845_),
    .B1(_06847_),
    .B2(_06852_),
    .Y(_06853_));
 NAND2x1_ASAP7_75t_R _26371_ (.A(_06830_),
    .B(_06836_),
    .Y(_06854_));
 BUFx4f_ASAP7_75t_R _26372_ (.A(_06854_),
    .Y(_06855_));
 NAND2x2_ASAP7_75t_R _26373_ (.A(_05974_),
    .B(_06848_),
    .Y(_06856_));
 OA21x2_ASAP7_75t_R _26374_ (.A1(_06855_),
    .A2(_06849_),
    .B(_06856_),
    .Y(_06857_));
 INVx1_ASAP7_75t_R _26375_ (.A(_06846_),
    .Y(_06858_));
 BUFx10_ASAP7_75t_R _26376_ (.A(_06831_),
    .Y(_06859_));
 OR2x2_ASAP7_75t_R _26377_ (.A(_02102_),
    .B(_06850_),
    .Y(_06860_));
 NOR2x1_ASAP7_75t_R _26378_ (.A(_02091_),
    .B(_06860_),
    .Y(_06861_));
 AND4x2_ASAP7_75t_R _26379_ (.A(_06844_),
    .B(_06859_),
    .C(_06836_),
    .D(_06861_),
    .Y(_06862_));
 BUFx6f_ASAP7_75t_R _26380_ (.A(_06856_),
    .Y(_06863_));
 NAND2x1_ASAP7_75t_R _26381_ (.A(_02145_),
    .B(_06863_),
    .Y(_06864_));
 AO21x1_ASAP7_75t_R _26382_ (.A1(_06858_),
    .A2(_06862_),
    .B(_06864_),
    .Y(_06865_));
 OA21x2_ASAP7_75t_R _26383_ (.A1(_06853_),
    .A2(_06857_),
    .B(_06865_),
    .Y(_02426_));
 BUFx4f_ASAP7_75t_R _26384_ (.A(_06857_),
    .Y(_06866_));
 BUFx6f_ASAP7_75t_R _26385_ (.A(_06844_),
    .Y(_06867_));
 OR3x1_ASAP7_75t_R _26386_ (.A(_00787_),
    .B(_02124_),
    .C(_02135_),
    .Y(_06868_));
 OR2x2_ASAP7_75t_R _26387_ (.A(_02113_),
    .B(_06868_),
    .Y(_06869_));
 OR3x4_ASAP7_75t_R _26388_ (.A(_02091_),
    .B(_02102_),
    .C(_06869_),
    .Y(_06870_));
 OR4x1_ASAP7_75t_R _26389_ (.A(_02144_),
    .B(_06849_),
    .C(_06847_),
    .D(_06870_),
    .Y(_06871_));
 OA21x2_ASAP7_75t_R _26390_ (.A1(_06639_),
    .A2(_06867_),
    .B(_06871_),
    .Y(_06872_));
 NOR2x1_ASAP7_75t_R _26391_ (.A(_02145_),
    .B(_06846_),
    .Y(_06873_));
 INVx1_ASAP7_75t_R _26392_ (.A(_06870_),
    .Y(_06874_));
 AND4x2_ASAP7_75t_R _26393_ (.A(_06844_),
    .B(_06831_),
    .C(_06836_),
    .D(_06874_),
    .Y(_06875_));
 NAND2x1_ASAP7_75t_R _26394_ (.A(_02144_),
    .B(_06863_),
    .Y(_06876_));
 AO21x1_ASAP7_75t_R _26395_ (.A1(_06873_),
    .A2(_06875_),
    .B(_06876_),
    .Y(_06877_));
 OA21x2_ASAP7_75t_R _26396_ (.A1(_06866_),
    .A2(_06872_),
    .B(_06877_),
    .Y(_02427_));
 BUFx4f_ASAP7_75t_R _26397_ (.A(_06856_),
    .Y(_06878_));
 AND2x2_ASAP7_75t_R _26398_ (.A(_02143_),
    .B(_06878_),
    .Y(_06879_));
 AND2x2_ASAP7_75t_R _26399_ (.A(_06323_),
    .B(_06778_),
    .Y(_06880_));
 BUFx4f_ASAP7_75t_R _26400_ (.A(_06880_),
    .Y(_06881_));
 OR5x1_ASAP7_75t_R _26401_ (.A(_02144_),
    .B(_06855_),
    .C(_06881_),
    .D(_06851_),
    .E(_06847_),
    .Y(_06882_));
 INVx5_ASAP7_75t_R _26402_ (.A(_06017_),
    .Y(_06883_));
 OR4x2_ASAP7_75t_R _26403_ (.A(_02143_),
    .B(_02144_),
    .C(_02145_),
    .D(_06846_),
    .Y(_06884_));
 OAI22x1_ASAP7_75t_R _26404_ (.A1(_06883_),
    .A2(_06867_),
    .B1(_06852_),
    .B2(_06884_),
    .Y(_06885_));
 AOI22x1_ASAP7_75t_R _26405_ (.A1(_06879_),
    .A2(_06882_),
    .B1(_06885_),
    .B2(_06840_),
    .Y(_02428_));
 BUFx4f_ASAP7_75t_R _26406_ (.A(_06843_),
    .Y(_06886_));
 OR2x4_ASAP7_75t_R _26407_ (.A(_06848_),
    .B(_06870_),
    .Y(_06887_));
 OR3x1_ASAP7_75t_R _26408_ (.A(_02142_),
    .B(_06884_),
    .C(_06887_),
    .Y(_06888_));
 OA21x2_ASAP7_75t_R _26409_ (.A1(_06650_),
    .A2(_06886_),
    .B(_06888_),
    .Y(_06889_));
 INVx1_ASAP7_75t_R _26410_ (.A(_06884_),
    .Y(_06890_));
 NAND2x1_ASAP7_75t_R _26411_ (.A(_02142_),
    .B(_06863_),
    .Y(_06891_));
 AO21x1_ASAP7_75t_R _26412_ (.A1(_06875_),
    .A2(_06890_),
    .B(_06891_),
    .Y(_06892_));
 OA21x2_ASAP7_75t_R _26413_ (.A1(_06866_),
    .A2(_06889_),
    .B(_06892_),
    .Y(_02429_));
 BUFx6f_ASAP7_75t_R _26414_ (.A(_06848_),
    .Y(_06893_));
 OR3x1_ASAP7_75t_R _26415_ (.A(_02141_),
    .B(_02142_),
    .C(_06884_),
    .Y(_06894_));
 OR3x1_ASAP7_75t_R _26416_ (.A(_06893_),
    .B(_06851_),
    .C(_06894_),
    .Y(_06895_));
 OA21x2_ASAP7_75t_R _26417_ (.A1(_06065_),
    .A2(_06886_),
    .B(_06895_),
    .Y(_06896_));
 NOR2x1_ASAP7_75t_R _26418_ (.A(_02142_),
    .B(_06884_),
    .Y(_06897_));
 NAND2x1_ASAP7_75t_R _26419_ (.A(_02141_),
    .B(_06863_),
    .Y(_06898_));
 AO21x1_ASAP7_75t_R _26420_ (.A1(_06862_),
    .A2(_06897_),
    .B(_06898_),
    .Y(_06899_));
 OA21x2_ASAP7_75t_R _26421_ (.A1(_06866_),
    .A2(_06896_),
    .B(_06899_),
    .Y(_02430_));
 AND2x2_ASAP7_75t_R _26422_ (.A(_02140_),
    .B(_06878_),
    .Y(_06900_));
 BUFx4f_ASAP7_75t_R _26423_ (.A(_06854_),
    .Y(_06901_));
 BUFx3_ASAP7_75t_R _26424_ (.A(_06880_),
    .Y(_06902_));
 OR4x1_ASAP7_75t_R _26425_ (.A(_06901_),
    .B(_06902_),
    .C(_06870_),
    .D(_06894_),
    .Y(_06903_));
 OR2x4_ASAP7_75t_R _26426_ (.A(_02140_),
    .B(_06894_),
    .Y(_06904_));
 OAI22x1_ASAP7_75t_R _26427_ (.A1(_06660_),
    .A2(_06844_),
    .B1(_06887_),
    .B2(_06904_),
    .Y(_06905_));
 AND2x2_ASAP7_75t_R _26428_ (.A(_06839_),
    .B(_06905_),
    .Y(_06906_));
 AOI21x1_ASAP7_75t_R _26429_ (.A1(_06900_),
    .A2(_06903_),
    .B(_06906_),
    .Y(_02431_));
 BUFx4f_ASAP7_75t_R _26430_ (.A(_06880_),
    .Y(_06907_));
 OR3x4_ASAP7_75t_R _26431_ (.A(_02139_),
    .B(_06851_),
    .C(_06904_),
    .Y(_06908_));
 OA22x2_ASAP7_75t_R _26432_ (.A1(_06111_),
    .A2(_06845_),
    .B1(_06907_),
    .B2(_06908_),
    .Y(_06909_));
 INVx1_ASAP7_75t_R _26433_ (.A(_06904_),
    .Y(_06910_));
 NAND2x1_ASAP7_75t_R _26434_ (.A(_02139_),
    .B(_06863_),
    .Y(_06911_));
 AO21x1_ASAP7_75t_R _26435_ (.A1(_06862_),
    .A2(_06910_),
    .B(_06911_),
    .Y(_06912_));
 OA21x2_ASAP7_75t_R _26436_ (.A1(_06866_),
    .A2(_06909_),
    .B(_06912_),
    .Y(_02432_));
 BUFx4f_ASAP7_75t_R _26437_ (.A(_06849_),
    .Y(_06913_));
 OAI21x1_ASAP7_75t_R _26438_ (.A1(_06901_),
    .A2(_06913_),
    .B(_06878_),
    .Y(_06914_));
 NAND3x2_ASAP7_75t_R _26439_ (.B(_06321_),
    .C(_06778_),
    .Y(_06915_),
    .A(_05876_));
 OR3x2_ASAP7_75t_R _26440_ (.A(_02139_),
    .B(_06870_),
    .C(_06904_),
    .Y(_06916_));
 OR2x2_ASAP7_75t_R _26441_ (.A(_06848_),
    .B(_06916_),
    .Y(_06917_));
 OAI22x1_ASAP7_75t_R _26442_ (.A1(_06137_),
    .A2(_06915_),
    .B1(_06917_),
    .B2(_06124_),
    .Y(_06918_));
 BUFx4f_ASAP7_75t_R _26443_ (.A(_06880_),
    .Y(_06919_));
 NAND2x1_ASAP7_75t_R _26444_ (.A(_05974_),
    .B(_06919_),
    .Y(_06920_));
 OA211x2_ASAP7_75t_R _26445_ (.A1(_06901_),
    .A2(_06917_),
    .B(_06920_),
    .C(_06124_),
    .Y(_06921_));
 AOI21x1_ASAP7_75t_R _26446_ (.A1(_06914_),
    .A2(_06918_),
    .B(_06921_),
    .Y(_02433_));
 AND2x2_ASAP7_75t_R _26447_ (.A(_02137_),
    .B(_06878_),
    .Y(_06922_));
 OR4x1_ASAP7_75t_R _26448_ (.A(_06124_),
    .B(_06901_),
    .C(_06881_),
    .D(_06908_),
    .Y(_06923_));
 OR4x1_ASAP7_75t_R _26449_ (.A(_02137_),
    .B(_06124_),
    .C(_06893_),
    .D(_06908_),
    .Y(_06924_));
 OAI21x1_ASAP7_75t_R _26450_ (.A1(_06161_),
    .A2(_06867_),
    .B(_06924_),
    .Y(_06925_));
 AOI22x1_ASAP7_75t_R _26451_ (.A1(_06922_),
    .A2(_06923_),
    .B1(_06925_),
    .B2(_06840_),
    .Y(_02434_));
 AND2x2_ASAP7_75t_R _26452_ (.A(_02136_),
    .B(_06878_),
    .Y(_06926_));
 OR5x1_ASAP7_75t_R _26453_ (.A(_02137_),
    .B(_06124_),
    .C(_06855_),
    .D(_06919_),
    .E(_06916_),
    .Y(_06927_));
 OR4x1_ASAP7_75t_R _26454_ (.A(_02136_),
    .B(_02137_),
    .C(_06124_),
    .D(_06917_),
    .Y(_06928_));
 OAI21x1_ASAP7_75t_R _26455_ (.A1(_06180_),
    .A2(_06867_),
    .B(_06928_),
    .Y(_06929_));
 AOI22x1_ASAP7_75t_R _26456_ (.A1(_06926_),
    .A2(_06927_),
    .B1(_06929_),
    .B2(_06840_),
    .Y(_02435_));
 BUFx6f_ASAP7_75t_R _26457_ (.A(_06837_),
    .Y(_06930_));
 OR2x2_ASAP7_75t_R _26458_ (.A(_02312_),
    .B(_06849_),
    .Y(_06931_));
 OA211x2_ASAP7_75t_R _26459_ (.A1(_06198_),
    .A2(_06930_),
    .B(_06839_),
    .C(_06931_),
    .Y(_06932_));
 AOI21x1_ASAP7_75t_R _26460_ (.A1(_02135_),
    .A2(_06866_),
    .B(_06932_),
    .Y(_02436_));
 OR4x1_ASAP7_75t_R _26461_ (.A(_02134_),
    .B(_02136_),
    .C(_02137_),
    .D(_06124_),
    .Y(_06933_));
 OR3x1_ASAP7_75t_R _26462_ (.A(_06893_),
    .B(_06908_),
    .C(_06933_),
    .Y(_06934_));
 OA21x2_ASAP7_75t_R _26463_ (.A1(_06218_),
    .A2(_06886_),
    .B(_06934_),
    .Y(_06935_));
 OR5x1_ASAP7_75t_R _26464_ (.A(_02136_),
    .B(_02137_),
    .C(_06124_),
    .D(_06893_),
    .E(_06908_),
    .Y(_06936_));
 AND2x2_ASAP7_75t_R _26465_ (.A(_02134_),
    .B(_06856_),
    .Y(_06937_));
 OAI21x1_ASAP7_75t_R _26466_ (.A1(_06901_),
    .A2(_06936_),
    .B(_06937_),
    .Y(_06938_));
 OA21x2_ASAP7_75t_R _26467_ (.A1(_06866_),
    .A2(_06935_),
    .B(_06938_),
    .Y(_02437_));
 AND2x2_ASAP7_75t_R _26468_ (.A(_02133_),
    .B(_06878_),
    .Y(_06939_));
 BUFx3_ASAP7_75t_R _26469_ (.A(_06880_),
    .Y(_06940_));
 OR4x1_ASAP7_75t_R _26470_ (.A(_06901_),
    .B(_06940_),
    .C(_06916_),
    .D(_06933_),
    .Y(_06941_));
 OR2x2_ASAP7_75t_R _26471_ (.A(_02133_),
    .B(_06933_),
    .Y(_06942_));
 OR2x2_ASAP7_75t_R _26472_ (.A(_06916_),
    .B(_06942_),
    .Y(_06943_));
 OAI22x1_ASAP7_75t_R _26473_ (.A1(_06695_),
    .A2(_06867_),
    .B1(_06907_),
    .B2(_06943_),
    .Y(_06944_));
 AOI22x1_ASAP7_75t_R _26474_ (.A1(_06939_),
    .A2(_06941_),
    .B1(_06944_),
    .B2(_06840_),
    .Y(_02438_));
 OR2x2_ASAP7_75t_R _26475_ (.A(_06908_),
    .B(_06942_),
    .Y(_06945_));
 OR3x1_ASAP7_75t_R _26476_ (.A(_02132_),
    .B(_06893_),
    .C(_06945_),
    .Y(_06946_));
 OA21x2_ASAP7_75t_R _26477_ (.A1(_06260_),
    .A2(_06886_),
    .B(_06946_),
    .Y(_06947_));
 INVx1_ASAP7_75t_R _26478_ (.A(_06945_),
    .Y(_06948_));
 NAND2x1_ASAP7_75t_R _26479_ (.A(_02132_),
    .B(_06863_),
    .Y(_06949_));
 AO21x1_ASAP7_75t_R _26480_ (.A1(_06838_),
    .A2(_06948_),
    .B(_06949_),
    .Y(_06950_));
 OA21x2_ASAP7_75t_R _26481_ (.A1(_06866_),
    .A2(_06947_),
    .B(_06950_),
    .Y(_02439_));
 AND2x2_ASAP7_75t_R _26482_ (.A(_02131_),
    .B(_06878_),
    .Y(_06951_));
 OR4x1_ASAP7_75t_R _26483_ (.A(_02132_),
    .B(_06855_),
    .C(_06881_),
    .D(_06943_),
    .Y(_06952_));
 OR2x2_ASAP7_75t_R _26484_ (.A(_02131_),
    .B(_02132_),
    .Y(_06953_));
 OR3x1_ASAP7_75t_R _26485_ (.A(_06881_),
    .B(_06943_),
    .C(_06953_),
    .Y(_06954_));
 OAI21x1_ASAP7_75t_R _26486_ (.A1(_06705_),
    .A2(_06867_),
    .B(_06954_),
    .Y(_06955_));
 AOI22x1_ASAP7_75t_R _26487_ (.A1(_06951_),
    .A2(_06952_),
    .B1(_06955_),
    .B2(_06840_),
    .Y(_02440_));
 AND2x2_ASAP7_75t_R _26488_ (.A(_02130_),
    .B(_06878_),
    .Y(_06956_));
 OR4x1_ASAP7_75t_R _26489_ (.A(_06901_),
    .B(_06940_),
    .C(_06945_),
    .D(_06953_),
    .Y(_06957_));
 OR4x1_ASAP7_75t_R _26490_ (.A(_02130_),
    .B(_06913_),
    .C(_06945_),
    .D(_06953_),
    .Y(_06958_));
 OAI21x1_ASAP7_75t_R _26491_ (.A1(_06299_),
    .A2(_06867_),
    .B(_06958_),
    .Y(_06959_));
 AOI22x1_ASAP7_75t_R _26492_ (.A1(_06956_),
    .A2(_06957_),
    .B1(_06959_),
    .B2(_06840_),
    .Y(_02441_));
 OR5x2_ASAP7_75t_R _26493_ (.A(_02130_),
    .B(_02139_),
    .C(_06904_),
    .D(_06942_),
    .E(_06953_),
    .Y(_06960_));
 OR3x1_ASAP7_75t_R _26494_ (.A(_02129_),
    .B(_06870_),
    .C(_06960_),
    .Y(_06961_));
 BUFx3_ASAP7_75t_R _26495_ (.A(_06961_),
    .Y(_06962_));
 OR2x2_ASAP7_75t_R _26496_ (.A(_06848_),
    .B(_06962_),
    .Y(_06963_));
 OA21x2_ASAP7_75t_R _26497_ (.A1(_06320_),
    .A2(_06886_),
    .B(_06963_),
    .Y(_06964_));
 INVx1_ASAP7_75t_R _26498_ (.A(_06960_),
    .Y(_06965_));
 NAND2x1_ASAP7_75t_R _26499_ (.A(_02129_),
    .B(_06863_),
    .Y(_06966_));
 AO21x1_ASAP7_75t_R _26500_ (.A1(_06875_),
    .A2(_06965_),
    .B(_06966_),
    .Y(_06967_));
 OA21x2_ASAP7_75t_R _26501_ (.A1(_06866_),
    .A2(_06964_),
    .B(_06967_),
    .Y(_02442_));
 INVx3_ASAP7_75t_R _26502_ (.A(_06347_),
    .Y(_06968_));
 OR3x4_ASAP7_75t_R _26503_ (.A(_02129_),
    .B(_06851_),
    .C(_06960_),
    .Y(_06969_));
 OR2x2_ASAP7_75t_R _26504_ (.A(_06849_),
    .B(_06969_),
    .Y(_06970_));
 OAI22x1_ASAP7_75t_R _26505_ (.A1(_06968_),
    .A2(_06915_),
    .B1(_06970_),
    .B2(_06336_),
    .Y(_06971_));
 OA211x2_ASAP7_75t_R _26506_ (.A1(_06901_),
    .A2(_06970_),
    .B(_06920_),
    .C(_06336_),
    .Y(_06972_));
 AOI21x1_ASAP7_75t_R _26507_ (.A1(_06914_),
    .A2(_06971_),
    .B(_06972_),
    .Y(_02443_));
 NOR2x1_ASAP7_75t_R _26508_ (.A(_02127_),
    .B(_06779_),
    .Y(_06973_));
 OR4x1_ASAP7_75t_R _26509_ (.A(_06336_),
    .B(_06855_),
    .C(_06919_),
    .D(_06962_),
    .Y(_06974_));
 NOR2x1_ASAP7_75t_R _26510_ (.A(_06370_),
    .B(_06930_),
    .Y(_06975_));
 INVx1_ASAP7_75t_R _26511_ (.A(_06336_),
    .Y(_06976_));
 INVx1_ASAP7_75t_R _26512_ (.A(_06962_),
    .Y(_06977_));
 NAND2x1_ASAP7_75t_R _26513_ (.A(_06562_),
    .B(_06778_),
    .Y(_06978_));
 AND4x1_ASAP7_75t_R _26514_ (.A(_02127_),
    .B(_06976_),
    .C(_06977_),
    .D(_06978_),
    .Y(_06979_));
 OA21x2_ASAP7_75t_R _26515_ (.A1(_06975_),
    .A2(_06979_),
    .B(_06839_),
    .Y(_06980_));
 AO21x1_ASAP7_75t_R _26516_ (.A1(_06973_),
    .A2(_06974_),
    .B(_06980_),
    .Y(_02444_));
 AND2x2_ASAP7_75t_R _26517_ (.A(_02126_),
    .B(_06878_),
    .Y(_06981_));
 OR5x1_ASAP7_75t_R _26518_ (.A(_02127_),
    .B(_06336_),
    .C(_06855_),
    .D(_06919_),
    .E(_06969_),
    .Y(_06982_));
 OR3x2_ASAP7_75t_R _26519_ (.A(_02126_),
    .B(_02127_),
    .C(_06336_),
    .Y(_06983_));
 OR3x1_ASAP7_75t_R _26520_ (.A(_06913_),
    .B(_06969_),
    .C(_06983_),
    .Y(_06984_));
 OAI21x1_ASAP7_75t_R _26521_ (.A1(_06738_),
    .A2(_06867_),
    .B(_06984_),
    .Y(_06985_));
 AOI22x1_ASAP7_75t_R _26522_ (.A1(_06981_),
    .A2(_06982_),
    .B1(_06985_),
    .B2(_06840_),
    .Y(_02445_));
 NOR2x1_ASAP7_75t_R _26523_ (.A(_02125_),
    .B(_06779_),
    .Y(_06986_));
 OR4x1_ASAP7_75t_R _26524_ (.A(_06855_),
    .B(_06881_),
    .C(_06962_),
    .D(_06983_),
    .Y(_06987_));
 NOR2x1_ASAP7_75t_R _26525_ (.A(_06849_),
    .B(_06962_),
    .Y(_06988_));
 INVx1_ASAP7_75t_R _26526_ (.A(_06983_),
    .Y(_06989_));
 AO32x1_ASAP7_75t_R _26527_ (.A1(_02125_),
    .A2(_06988_),
    .A3(_06989_),
    .B1(_06410_),
    .B2(_06919_),
    .Y(_06990_));
 AND2x2_ASAP7_75t_R _26528_ (.A(_06839_),
    .B(_06990_),
    .Y(_06991_));
 AO21x1_ASAP7_75t_R _26529_ (.A1(_06986_),
    .A2(_06987_),
    .B(_06991_),
    .Y(_02446_));
 OR3x1_ASAP7_75t_R _26530_ (.A(_02124_),
    .B(_02311_),
    .C(_06893_),
    .Y(_06992_));
 OA21x2_ASAP7_75t_R _26531_ (.A1(_05872_),
    .A2(_06886_),
    .B(_06992_),
    .Y(_06993_));
 INVx1_ASAP7_75t_R _26532_ (.A(_02311_),
    .Y(_06994_));
 NAND2x1_ASAP7_75t_R _26533_ (.A(_02124_),
    .B(_06863_),
    .Y(_06995_));
 AO21x1_ASAP7_75t_R _26534_ (.A1(_06994_),
    .A2(_06838_),
    .B(_06995_),
    .Y(_06996_));
 OA21x2_ASAP7_75t_R _26535_ (.A1(_06866_),
    .A2(_06993_),
    .B(_06996_),
    .Y(_02447_));
 OR3x4_ASAP7_75t_R _26536_ (.A(_02123_),
    .B(_02125_),
    .C(_06983_),
    .Y(_06997_));
 OA22x2_ASAP7_75t_R _26537_ (.A1(_06750_),
    .A2(_06845_),
    .B1(_06970_),
    .B2(_06997_),
    .Y(_06998_));
 OR3x1_ASAP7_75t_R _26538_ (.A(_02125_),
    .B(_06969_),
    .C(_06983_),
    .Y(_06999_));
 INVx1_ASAP7_75t_R _26539_ (.A(_06999_),
    .Y(_07000_));
 NAND2x1_ASAP7_75t_R _26540_ (.A(_02123_),
    .B(_06856_),
    .Y(_07001_));
 AO21x1_ASAP7_75t_R _26541_ (.A1(_06838_),
    .A2(_07000_),
    .B(_07001_),
    .Y(_07002_));
 OA21x2_ASAP7_75t_R _26542_ (.A1(_06866_),
    .A2(_06998_),
    .B(_07002_),
    .Y(_02448_));
 NOR2x1_ASAP7_75t_R _26543_ (.A(_02122_),
    .B(_06779_),
    .Y(_07003_));
 OR4x1_ASAP7_75t_R _26544_ (.A(_06855_),
    .B(_06881_),
    .C(_06962_),
    .D(_06997_),
    .Y(_07004_));
 INVx1_ASAP7_75t_R _26545_ (.A(_02122_),
    .Y(_07005_));
 OR3x1_ASAP7_75t_R _26546_ (.A(_07005_),
    .B(_06963_),
    .C(_06997_),
    .Y(_07006_));
 OAI21x1_ASAP7_75t_R _26547_ (.A1(_06455_),
    .A2(_06930_),
    .B(_07006_),
    .Y(_07007_));
 AND2x2_ASAP7_75t_R _26548_ (.A(_06839_),
    .B(_07007_),
    .Y(_07008_));
 AO21x1_ASAP7_75t_R _26549_ (.A1(_07003_),
    .A2(_07004_),
    .B(_07008_),
    .Y(_02449_));
 INVx1_ASAP7_75t_R _26550_ (.A(_02121_),
    .Y(_07009_));
 OR3x1_ASAP7_75t_R _26551_ (.A(_02122_),
    .B(_06969_),
    .C(_06997_),
    .Y(_07010_));
 INVx1_ASAP7_75t_R _26552_ (.A(_07010_),
    .Y(_07011_));
 AND3x1_ASAP7_75t_R _26553_ (.A(_05914_),
    .B(_05915_),
    .C(_06777_),
    .Y(_07012_));
 NAND2x1_ASAP7_75t_R _26554_ (.A(_06007_),
    .B(_07012_),
    .Y(_07013_));
 AO32x1_ASAP7_75t_R _26555_ (.A1(_06830_),
    .A2(_06836_),
    .A3(_07013_),
    .B1(_07012_),
    .B2(_05930_),
    .Y(_07014_));
 BUFx6f_ASAP7_75t_R _26556_ (.A(_07014_),
    .Y(_07015_));
 OAI21x1_ASAP7_75t_R _26557_ (.A1(_06913_),
    .A2(_07011_),
    .B(_07015_),
    .Y(_07016_));
 AND3x1_ASAP7_75t_R _26558_ (.A(_02121_),
    .B(_06930_),
    .C(_07011_),
    .Y(_07017_));
 AO21x1_ASAP7_75t_R _26559_ (.A1(_05841_),
    .A2(_06907_),
    .B(_07017_),
    .Y(_07018_));
 BUFx3_ASAP7_75t_R _26560_ (.A(_07015_),
    .Y(_07019_));
 AO22x1_ASAP7_75t_R _26561_ (.A1(_07009_),
    .A2(_07016_),
    .B1(_07018_),
    .B2(_07019_),
    .Y(_02450_));
 BUFx4f_ASAP7_75t_R _26562_ (.A(_07015_),
    .Y(_07020_));
 INVx1_ASAP7_75t_R _26563_ (.A(_02120_),
    .Y(_07021_));
 OR3x2_ASAP7_75t_R _26564_ (.A(_02121_),
    .B(_02122_),
    .C(_06997_),
    .Y(_07022_));
 OR3x1_ASAP7_75t_R _26565_ (.A(_07021_),
    .B(_06963_),
    .C(_07022_),
    .Y(_07023_));
 OAI21x1_ASAP7_75t_R _26566_ (.A1(_06198_),
    .A2(_06930_),
    .B(_07023_),
    .Y(_07024_));
 BUFx6f_ASAP7_75t_R _26567_ (.A(_07015_),
    .Y(_07025_));
 OAI21x1_ASAP7_75t_R _26568_ (.A1(_06962_),
    .A2(_07022_),
    .B(_06886_),
    .Y(_07026_));
 AOI21x1_ASAP7_75t_R _26569_ (.A1(_07025_),
    .A2(_07026_),
    .B(_02120_),
    .Y(_07027_));
 AO21x1_ASAP7_75t_R _26570_ (.A1(_07020_),
    .A2(_07024_),
    .B(_07027_),
    .Y(_02451_));
 OR3x4_ASAP7_75t_R _26571_ (.A(_02120_),
    .B(_06969_),
    .C(_07022_),
    .Y(_07028_));
 NOR2x1_ASAP7_75t_R _26572_ (.A(_06893_),
    .B(_07028_),
    .Y(_07029_));
 AO32x1_ASAP7_75t_R _26573_ (.A1(_05872_),
    .A2(_06323_),
    .A3(_06778_),
    .B1(_07029_),
    .B2(_05853_),
    .Y(_07030_));
 BUFx6f_ASAP7_75t_R _26574_ (.A(_06843_),
    .Y(_07031_));
 NAND2x1_ASAP7_75t_R _26575_ (.A(_07031_),
    .B(_07028_),
    .Y(_07032_));
 AOI21x1_ASAP7_75t_R _26576_ (.A1(_07025_),
    .A2(_07032_),
    .B(_05853_),
    .Y(_07033_));
 AO21x1_ASAP7_75t_R _26577_ (.A1(_07020_),
    .A2(_07030_),
    .B(_07033_),
    .Y(_02452_));
 INVx1_ASAP7_75t_R _26578_ (.A(_05853_),
    .Y(_07034_));
 OR3x1_ASAP7_75t_R _26579_ (.A(_02120_),
    .B(_06962_),
    .C(_07022_),
    .Y(_07035_));
 INVx2_ASAP7_75t_R _26580_ (.A(_07035_),
    .Y(_07036_));
 AND2x2_ASAP7_75t_R _26581_ (.A(_06978_),
    .B(_07036_),
    .Y(_07037_));
 AO32x1_ASAP7_75t_R _26582_ (.A1(_06488_),
    .A2(_07034_),
    .A3(_07037_),
    .B1(_06881_),
    .B2(_06588_),
    .Y(_07038_));
 AO21x1_ASAP7_75t_R _26583_ (.A1(_07034_),
    .A2(_07036_),
    .B(_06913_),
    .Y(_07039_));
 AOI21x1_ASAP7_75t_R _26584_ (.A1(_07025_),
    .A2(_07039_),
    .B(_06488_),
    .Y(_07040_));
 AO21x1_ASAP7_75t_R _26585_ (.A1(_07020_),
    .A2(_07038_),
    .B(_07040_),
    .Y(_02453_));
 NOR2x1_ASAP7_75t_R _26586_ (.A(_06488_),
    .B(_05853_),
    .Y(_07041_));
 CKINVDCx5p33_ASAP7_75t_R _26587_ (.A(_06517_),
    .Y(_07042_));
 AO32x1_ASAP7_75t_R _26588_ (.A1(_02117_),
    .A2(_07029_),
    .A3(_07041_),
    .B1(_07042_),
    .B2(_06902_),
    .Y(_07043_));
 OR3x1_ASAP7_75t_R _26589_ (.A(_06488_),
    .B(_05853_),
    .C(_07028_),
    .Y(_07044_));
 NAND2x1_ASAP7_75t_R _26590_ (.A(_07031_),
    .B(_07044_),
    .Y(_07045_));
 AOI21x1_ASAP7_75t_R _26591_ (.A1(_07025_),
    .A2(_07045_),
    .B(_02117_),
    .Y(_07046_));
 AO21x1_ASAP7_75t_R _26592_ (.A1(_07020_),
    .A2(_07043_),
    .B(_07046_),
    .Y(_02454_));
 OR3x2_ASAP7_75t_R _26593_ (.A(_02117_),
    .B(_06488_),
    .C(_05853_),
    .Y(_07047_));
 INVx1_ASAP7_75t_R _26594_ (.A(_07047_),
    .Y(_07048_));
 AO32x1_ASAP7_75t_R _26595_ (.A1(_06523_),
    .A2(_07037_),
    .A3(_07048_),
    .B1(_06534_),
    .B2(_06902_),
    .Y(_07049_));
 AO21x1_ASAP7_75t_R _26596_ (.A1(_07036_),
    .A2(_07048_),
    .B(_06913_),
    .Y(_07050_));
 AOI21x1_ASAP7_75t_R _26597_ (.A1(_07025_),
    .A2(_07050_),
    .B(_06523_),
    .Y(_07051_));
 AO21x1_ASAP7_75t_R _26598_ (.A1(_07020_),
    .A2(_07049_),
    .B(_07051_),
    .Y(_02455_));
 NOR2x1_ASAP7_75t_R _26599_ (.A(_06523_),
    .B(_07047_),
    .Y(_07052_));
 AO32x1_ASAP7_75t_R _26600_ (.A1(_02115_),
    .A2(_07029_),
    .A3(_07052_),
    .B1(_06559_),
    .B2(_06902_),
    .Y(_07053_));
 OR3x1_ASAP7_75t_R _26601_ (.A(_06523_),
    .B(_07028_),
    .C(_07047_),
    .Y(_07054_));
 NAND2x1_ASAP7_75t_R _26602_ (.A(_07031_),
    .B(_07054_),
    .Y(_07055_));
 AOI21x1_ASAP7_75t_R _26603_ (.A1(_07025_),
    .A2(_07055_),
    .B(_02115_),
    .Y(_07056_));
 AO21x1_ASAP7_75t_R _26604_ (.A1(_07020_),
    .A2(_07053_),
    .B(_07056_),
    .Y(_02456_));
 OR3x2_ASAP7_75t_R _26605_ (.A(_02115_),
    .B(_06523_),
    .C(_07047_),
    .Y(_07057_));
 INVx1_ASAP7_75t_R _26606_ (.A(_07057_),
    .Y(_07058_));
 AO32x1_ASAP7_75t_R _26607_ (.A1(_06568_),
    .A2(_07037_),
    .A3(_07058_),
    .B1(_06583_),
    .B2(_06902_),
    .Y(_07059_));
 AO21x1_ASAP7_75t_R _26608_ (.A1(_07036_),
    .A2(_07058_),
    .B(_06913_),
    .Y(_07060_));
 AOI21x1_ASAP7_75t_R _26609_ (.A1(_07025_),
    .A2(_07060_),
    .B(_06568_),
    .Y(_07061_));
 AO21x1_ASAP7_75t_R _26610_ (.A1(_07020_),
    .A2(_07059_),
    .B(_07061_),
    .Y(_02457_));
 OR2x2_ASAP7_75t_R _26611_ (.A(_06849_),
    .B(_06869_),
    .Y(_07062_));
 OA21x2_ASAP7_75t_R _26612_ (.A1(_06588_),
    .A2(_06886_),
    .B(_07062_),
    .Y(_07063_));
 INVx1_ASAP7_75t_R _26613_ (.A(_06868_),
    .Y(_07064_));
 NAND2x1_ASAP7_75t_R _26614_ (.A(_02113_),
    .B(_06856_),
    .Y(_07065_));
 AO21x1_ASAP7_75t_R _26615_ (.A1(_06838_),
    .A2(_07064_),
    .B(_07065_),
    .Y(_07066_));
 OA21x2_ASAP7_75t_R _26616_ (.A1(_06857_),
    .A2(_07063_),
    .B(_07066_),
    .Y(_02458_));
 NOR2x1_ASAP7_75t_R _26617_ (.A(_06568_),
    .B(_07057_),
    .Y(_07067_));
 AO32x1_ASAP7_75t_R _26618_ (.A1(_02112_),
    .A2(_07029_),
    .A3(_07067_),
    .B1(_06609_),
    .B2(_06902_),
    .Y(_07068_));
 OR3x1_ASAP7_75t_R _26619_ (.A(_06568_),
    .B(_07028_),
    .C(_07057_),
    .Y(_07069_));
 NAND2x1_ASAP7_75t_R _26620_ (.A(_07031_),
    .B(_07069_),
    .Y(_07070_));
 AOI21x1_ASAP7_75t_R _26621_ (.A1(_07025_),
    .A2(_07070_),
    .B(_02112_),
    .Y(_07071_));
 AO21x1_ASAP7_75t_R _26622_ (.A1(_07020_),
    .A2(_07068_),
    .B(_07071_),
    .Y(_02459_));
 OR3x1_ASAP7_75t_R _26623_ (.A(_02112_),
    .B(_06568_),
    .C(_07057_),
    .Y(_07072_));
 INVx1_ASAP7_75t_R _26624_ (.A(_07072_),
    .Y(_07073_));
 AO32x1_ASAP7_75t_R _26625_ (.A1(_02111_),
    .A2(_07037_),
    .A3(_07073_),
    .B1(_06627_),
    .B2(_06902_),
    .Y(_07074_));
 BUFx6f_ASAP7_75t_R _26626_ (.A(_07015_),
    .Y(_07075_));
 AO21x1_ASAP7_75t_R _26627_ (.A1(_07036_),
    .A2(_07073_),
    .B(_06913_),
    .Y(_07076_));
 AOI21x1_ASAP7_75t_R _26628_ (.A1(_07075_),
    .A2(_07076_),
    .B(_02111_),
    .Y(_07077_));
 AO21x1_ASAP7_75t_R _26629_ (.A1(_07020_),
    .A2(_07074_),
    .B(_07077_),
    .Y(_02460_));
 INVx1_ASAP7_75t_R _26630_ (.A(_05931_),
    .Y(_07078_));
 OR3x2_ASAP7_75t_R _26631_ (.A(_02111_),
    .B(_07028_),
    .C(_07072_),
    .Y(_07079_));
 INVx1_ASAP7_75t_R _26632_ (.A(_07079_),
    .Y(_07080_));
 OAI21x1_ASAP7_75t_R _26633_ (.A1(_06907_),
    .A2(_07080_),
    .B(_07015_),
    .Y(_07081_));
 NOR2x1_ASAP7_75t_R _26634_ (.A(_06849_),
    .B(_07079_),
    .Y(_07082_));
 AO32x1_ASAP7_75t_R _26635_ (.A1(_06635_),
    .A2(_06323_),
    .A3(_06778_),
    .B1(_07082_),
    .B2(_05931_),
    .Y(_07083_));
 AO22x1_ASAP7_75t_R _26636_ (.A1(_07078_),
    .A2(_07081_),
    .B1(_07083_),
    .B2(_07025_),
    .Y(_02461_));
 OR3x4_ASAP7_75t_R _26637_ (.A(_02111_),
    .B(_07035_),
    .C(_07072_),
    .Y(_07084_));
 NOR2x1_ASAP7_75t_R _26638_ (.A(_06893_),
    .B(_07084_),
    .Y(_07085_));
 AO32x1_ASAP7_75t_R _26639_ (.A1(_02109_),
    .A2(_07078_),
    .A3(_07085_),
    .B1(_06881_),
    .B2(_06639_),
    .Y(_07086_));
 OAI21x1_ASAP7_75t_R _26640_ (.A1(_05931_),
    .A2(_07084_),
    .B(_06845_),
    .Y(_07087_));
 AOI21x1_ASAP7_75t_R _26641_ (.A1(_07075_),
    .A2(_07087_),
    .B(_02109_),
    .Y(_07088_));
 AO21x1_ASAP7_75t_R _26642_ (.A1(_07020_),
    .A2(_07086_),
    .B(_07088_),
    .Y(_02462_));
 BUFx4f_ASAP7_75t_R _26643_ (.A(_07015_),
    .Y(_07089_));
 NOR2x1_ASAP7_75t_R _26644_ (.A(_02109_),
    .B(_05931_),
    .Y(_07090_));
 AO32x1_ASAP7_75t_R _26645_ (.A1(_02108_),
    .A2(_07082_),
    .A3(_07090_),
    .B1(_06883_),
    .B2(_06902_),
    .Y(_07091_));
 AO21x1_ASAP7_75t_R _26646_ (.A1(_07080_),
    .A2(_07090_),
    .B(_06913_),
    .Y(_07092_));
 AOI21x1_ASAP7_75t_R _26647_ (.A1(_07075_),
    .A2(_07092_),
    .B(_02108_),
    .Y(_07093_));
 AO21x1_ASAP7_75t_R _26648_ (.A1(_07089_),
    .A2(_07091_),
    .B(_07093_),
    .Y(_02463_));
 OR3x4_ASAP7_75t_R _26649_ (.A(_02108_),
    .B(_02109_),
    .C(_05931_),
    .Y(_07094_));
 INVx1_ASAP7_75t_R _26650_ (.A(_07094_),
    .Y(_07095_));
 AO32x1_ASAP7_75t_R _26651_ (.A1(_02107_),
    .A2(_07085_),
    .A3(_07095_),
    .B1(_06650_),
    .B2(_06902_),
    .Y(_07096_));
 OAI21x1_ASAP7_75t_R _26652_ (.A1(_07084_),
    .A2(_07094_),
    .B(_06845_),
    .Y(_07097_));
 AOI21x1_ASAP7_75t_R _26653_ (.A1(_07075_),
    .A2(_07097_),
    .B(_02107_),
    .Y(_07098_));
 AO21x1_ASAP7_75t_R _26654_ (.A1(_07089_),
    .A2(_07096_),
    .B(_07098_),
    .Y(_02464_));
 NOR2x1_ASAP7_75t_R _26655_ (.A(_02107_),
    .B(_07094_),
    .Y(_07099_));
 AO32x1_ASAP7_75t_R _26656_ (.A1(_02106_),
    .A2(_07082_),
    .A3(_07099_),
    .B1(_06065_),
    .B2(_06940_),
    .Y(_07100_));
 AO21x1_ASAP7_75t_R _26657_ (.A1(_07080_),
    .A2(_07099_),
    .B(_06913_),
    .Y(_07101_));
 AOI21x1_ASAP7_75t_R _26658_ (.A1(_07075_),
    .A2(_07101_),
    .B(_02106_),
    .Y(_07102_));
 AO21x1_ASAP7_75t_R _26659_ (.A1(_07089_),
    .A2(_07100_),
    .B(_07102_),
    .Y(_02465_));
 OR3x2_ASAP7_75t_R _26660_ (.A(_02106_),
    .B(_02107_),
    .C(_07094_),
    .Y(_07103_));
 INVx1_ASAP7_75t_R _26661_ (.A(_07103_),
    .Y(_07104_));
 AO32x1_ASAP7_75t_R _26662_ (.A1(_02105_),
    .A2(_07085_),
    .A3(_07104_),
    .B1(_06660_),
    .B2(_06940_),
    .Y(_07105_));
 OAI21x1_ASAP7_75t_R _26663_ (.A1(_07084_),
    .A2(_07103_),
    .B(_06845_),
    .Y(_07106_));
 AOI21x1_ASAP7_75t_R _26664_ (.A1(_07075_),
    .A2(_07106_),
    .B(_02105_),
    .Y(_07107_));
 AO21x1_ASAP7_75t_R _26665_ (.A1(_07089_),
    .A2(_07105_),
    .B(_07107_),
    .Y(_02466_));
 OR3x1_ASAP7_75t_R _26666_ (.A(_02105_),
    .B(_07079_),
    .C(_07103_),
    .Y(_07108_));
 BUFx3_ASAP7_75t_R _26667_ (.A(_07108_),
    .Y(_07109_));
 NOR2x1_ASAP7_75t_R _26668_ (.A(_06893_),
    .B(_07109_),
    .Y(_07110_));
 AO32x1_ASAP7_75t_R _26669_ (.A1(_06111_),
    .A2(_06323_),
    .A3(_06778_),
    .B1(_07110_),
    .B2(_06097_),
    .Y(_07111_));
 NAND2x1_ASAP7_75t_R _26670_ (.A(_07031_),
    .B(_07109_),
    .Y(_07112_));
 AOI21x1_ASAP7_75t_R _26671_ (.A1(_07075_),
    .A2(_07112_),
    .B(_06097_),
    .Y(_07113_));
 AO21x1_ASAP7_75t_R _26672_ (.A1(_07089_),
    .A2(_07111_),
    .B(_07113_),
    .Y(_02467_));
 INVx1_ASAP7_75t_R _26673_ (.A(_06097_),
    .Y(_07114_));
 OR3x4_ASAP7_75t_R _26674_ (.A(_02105_),
    .B(_07084_),
    .C(_07103_),
    .Y(_07115_));
 NOR2x1_ASAP7_75t_R _26675_ (.A(_06893_),
    .B(_07115_),
    .Y(_07116_));
 AO32x1_ASAP7_75t_R _26676_ (.A1(_06122_),
    .A2(_07114_),
    .A3(_07116_),
    .B1(_06881_),
    .B2(_06136_),
    .Y(_07117_));
 OAI21x1_ASAP7_75t_R _26677_ (.A1(_06097_),
    .A2(_07115_),
    .B(_06845_),
    .Y(_07118_));
 AOI21x1_ASAP7_75t_R _26678_ (.A1(_07075_),
    .A2(_07118_),
    .B(_06122_),
    .Y(_07119_));
 AO21x1_ASAP7_75t_R _26679_ (.A1(_07089_),
    .A2(_07117_),
    .B(_07119_),
    .Y(_02468_));
 OR2x2_ASAP7_75t_R _26680_ (.A(_06849_),
    .B(_06860_),
    .Y(_07120_));
 OA21x2_ASAP7_75t_R _26681_ (.A1(_07042_),
    .A2(_06886_),
    .B(_07120_),
    .Y(_07121_));
 INVx1_ASAP7_75t_R _26682_ (.A(_06850_),
    .Y(_07122_));
 NAND2x1_ASAP7_75t_R _26683_ (.A(_02102_),
    .B(_06856_),
    .Y(_07123_));
 AO21x1_ASAP7_75t_R _26684_ (.A1(_06838_),
    .A2(_07122_),
    .B(_07123_),
    .Y(_07124_));
 OA21x2_ASAP7_75t_R _26685_ (.A1(_06857_),
    .A2(_07121_),
    .B(_07124_),
    .Y(_02469_));
 NOR2x1_ASAP7_75t_R _26686_ (.A(_06122_),
    .B(_06097_),
    .Y(_07125_));
 AO32x1_ASAP7_75t_R _26687_ (.A1(_02101_),
    .A2(_07110_),
    .A3(_07125_),
    .B1(_06161_),
    .B2(_06940_),
    .Y(_07126_));
 OR3x1_ASAP7_75t_R _26688_ (.A(_06122_),
    .B(_06097_),
    .C(_07109_),
    .Y(_07127_));
 NAND2x1_ASAP7_75t_R _26689_ (.A(_07031_),
    .B(_07127_),
    .Y(_07128_));
 AOI21x1_ASAP7_75t_R _26690_ (.A1(_07075_),
    .A2(_07128_),
    .B(_02101_),
    .Y(_07129_));
 AO21x1_ASAP7_75t_R _26691_ (.A1(_07089_),
    .A2(_07126_),
    .B(_07129_),
    .Y(_02470_));
 OR3x1_ASAP7_75t_R _26692_ (.A(_02101_),
    .B(_06122_),
    .C(_06097_),
    .Y(_07130_));
 INVx1_ASAP7_75t_R _26693_ (.A(_07130_),
    .Y(_07131_));
 AO32x1_ASAP7_75t_R _26694_ (.A1(_02100_),
    .A2(_07116_),
    .A3(_07131_),
    .B1(_06179_),
    .B2(_06940_),
    .Y(_07132_));
 OAI21x1_ASAP7_75t_R _26695_ (.A1(_07115_),
    .A2(_07130_),
    .B(_06845_),
    .Y(_07133_));
 AOI21x1_ASAP7_75t_R _26696_ (.A1(_07075_),
    .A2(_07133_),
    .B(_02100_),
    .Y(_07134_));
 AO21x1_ASAP7_75t_R _26697_ (.A1(_07089_),
    .A2(_07132_),
    .B(_07134_),
    .Y(_02471_));
 OR2x4_ASAP7_75t_R _26698_ (.A(_02100_),
    .B(_07130_),
    .Y(_07135_));
 INVx1_ASAP7_75t_R _26699_ (.A(_07135_),
    .Y(_07136_));
 AO32x1_ASAP7_75t_R _26700_ (.A1(_06207_),
    .A2(_07110_),
    .A3(_07136_),
    .B1(_06217_),
    .B2(_06940_),
    .Y(_07137_));
 BUFx6f_ASAP7_75t_R _26701_ (.A(_07015_),
    .Y(_07138_));
 OAI21x1_ASAP7_75t_R _26702_ (.A1(_07109_),
    .A2(_07135_),
    .B(_06845_),
    .Y(_07139_));
 AOI21x1_ASAP7_75t_R _26703_ (.A1(_07138_),
    .A2(_07139_),
    .B(_06207_),
    .Y(_07140_));
 AO21x1_ASAP7_75t_R _26704_ (.A1(_07089_),
    .A2(_07137_),
    .B(_07140_),
    .Y(_02472_));
 NOR2x1_ASAP7_75t_R _26705_ (.A(_06207_),
    .B(_07135_),
    .Y(_07141_));
 AO32x1_ASAP7_75t_R _26706_ (.A1(_02098_),
    .A2(_07116_),
    .A3(_07141_),
    .B1(_06695_),
    .B2(_06940_),
    .Y(_07142_));
 OR3x1_ASAP7_75t_R _26707_ (.A(_06207_),
    .B(_07115_),
    .C(_07135_),
    .Y(_07143_));
 NAND2x1_ASAP7_75t_R _26708_ (.A(_07031_),
    .B(_07143_),
    .Y(_07144_));
 AOI21x1_ASAP7_75t_R _26709_ (.A1(_07138_),
    .A2(_07144_),
    .B(_02098_),
    .Y(_07145_));
 AO21x1_ASAP7_75t_R _26710_ (.A1(_07089_),
    .A2(_07142_),
    .B(_07145_),
    .Y(_02473_));
 OR3x2_ASAP7_75t_R _26711_ (.A(_02098_),
    .B(_06207_),
    .C(_07135_),
    .Y(_07146_));
 INVx1_ASAP7_75t_R _26712_ (.A(_07146_),
    .Y(_07147_));
 AO32x1_ASAP7_75t_R _26713_ (.A1(_02097_),
    .A2(_07110_),
    .A3(_07147_),
    .B1(_06260_),
    .B2(_06940_),
    .Y(_07148_));
 OAI21x1_ASAP7_75t_R _26714_ (.A1(_07109_),
    .A2(_07146_),
    .B(_06845_),
    .Y(_07149_));
 AOI21x1_ASAP7_75t_R _26715_ (.A1(_07138_),
    .A2(_07149_),
    .B(_02097_),
    .Y(_07150_));
 AO21x1_ASAP7_75t_R _26716_ (.A1(_07019_),
    .A2(_07148_),
    .B(_07150_),
    .Y(_02474_));
 INVx1_ASAP7_75t_R _26717_ (.A(_02096_),
    .Y(_07151_));
 OR3x1_ASAP7_75t_R _26718_ (.A(_02097_),
    .B(_07115_),
    .C(_07146_),
    .Y(_07152_));
 INVx1_ASAP7_75t_R _26719_ (.A(_07152_),
    .Y(_07153_));
 OAI21x1_ASAP7_75t_R _26720_ (.A1(_06907_),
    .A2(_07153_),
    .B(_07015_),
    .Y(_07154_));
 AND3x1_ASAP7_75t_R _26721_ (.A(_02096_),
    .B(_06837_),
    .C(_07153_),
    .Y(_07155_));
 AO21x1_ASAP7_75t_R _26722_ (.A1(_06705_),
    .A2(_06907_),
    .B(_07155_),
    .Y(_07156_));
 AO22x1_ASAP7_75t_R _26723_ (.A1(_07151_),
    .A2(_07154_),
    .B1(_07156_),
    .B2(_07025_),
    .Y(_02475_));
 OR4x1_ASAP7_75t_R _26724_ (.A(_02096_),
    .B(_02097_),
    .C(_07109_),
    .D(_07146_),
    .Y(_07157_));
 INVx1_ASAP7_75t_R _26725_ (.A(_07157_),
    .Y(_07158_));
 AND3x1_ASAP7_75t_R _26726_ (.A(_02095_),
    .B(_06930_),
    .C(_07158_),
    .Y(_07159_));
 AO21x1_ASAP7_75t_R _26727_ (.A1(_06299_),
    .A2(_06907_),
    .B(_07159_),
    .Y(_07160_));
 AO21x1_ASAP7_75t_R _26728_ (.A1(_06323_),
    .A2(_06778_),
    .B(_07158_),
    .Y(_07161_));
 AOI21x1_ASAP7_75t_R _26729_ (.A1(_07138_),
    .A2(_07161_),
    .B(_02095_),
    .Y(_07162_));
 AO21x1_ASAP7_75t_R _26730_ (.A1(_07019_),
    .A2(_07160_),
    .B(_07162_),
    .Y(_02476_));
 OR3x2_ASAP7_75t_R _26731_ (.A(_02095_),
    .B(_02096_),
    .C(_07152_),
    .Y(_07163_));
 INVx1_ASAP7_75t_R _26732_ (.A(_07163_),
    .Y(_07164_));
 AND3x1_ASAP7_75t_R _26733_ (.A(_02094_),
    .B(_06930_),
    .C(_07164_),
    .Y(_07165_));
 AO21x1_ASAP7_75t_R _26734_ (.A1(_06320_),
    .A2(_06907_),
    .B(_07165_),
    .Y(_07166_));
 NAND2x1_ASAP7_75t_R _26735_ (.A(_07031_),
    .B(_07163_),
    .Y(_07167_));
 AOI21x1_ASAP7_75t_R _26736_ (.A1(_07138_),
    .A2(_07167_),
    .B(_02094_),
    .Y(_07168_));
 AO21x1_ASAP7_75t_R _26737_ (.A1(_07019_),
    .A2(_07166_),
    .B(_07168_),
    .Y(_02477_));
 INVx1_ASAP7_75t_R _26738_ (.A(_02093_),
    .Y(_07169_));
 OR3x2_ASAP7_75t_R _26739_ (.A(_02094_),
    .B(_02095_),
    .C(_07157_),
    .Y(_07170_));
 OR3x1_ASAP7_75t_R _26740_ (.A(_07169_),
    .B(_06919_),
    .C(_07170_),
    .Y(_07171_));
 OAI21x1_ASAP7_75t_R _26741_ (.A1(_06347_),
    .A2(_06930_),
    .B(_07171_),
    .Y(_07172_));
 NAND2x1_ASAP7_75t_R _26742_ (.A(_07031_),
    .B(_07170_),
    .Y(_07173_));
 AOI21x1_ASAP7_75t_R _26743_ (.A1(_07138_),
    .A2(_07173_),
    .B(_02093_),
    .Y(_07174_));
 AO21x1_ASAP7_75t_R _26744_ (.A1(_07019_),
    .A2(_07172_),
    .B(_07174_),
    .Y(_02478_));
 OR3x4_ASAP7_75t_R _26745_ (.A(_02093_),
    .B(_02094_),
    .C(_07163_),
    .Y(_07175_));
 NOR2x1_ASAP7_75t_R _26746_ (.A(_06919_),
    .B(_07175_),
    .Y(_07176_));
 AO21x1_ASAP7_75t_R _26747_ (.A1(_06359_),
    .A2(_07176_),
    .B(_06975_),
    .Y(_07177_));
 NAND2x1_ASAP7_75t_R _26748_ (.A(_07031_),
    .B(_07175_),
    .Y(_07178_));
 AOI21x1_ASAP7_75t_R _26749_ (.A1(_07138_),
    .A2(_07178_),
    .B(_06359_),
    .Y(_07179_));
 AO21x1_ASAP7_75t_R _26750_ (.A1(_07019_),
    .A2(_07177_),
    .B(_07179_),
    .Y(_02479_));
 AND2x2_ASAP7_75t_R _26751_ (.A(_02091_),
    .B(_06863_),
    .Y(_07180_));
 OR4x1_ASAP7_75t_R _26752_ (.A(_02102_),
    .B(_06855_),
    .C(_06881_),
    .D(_06869_),
    .Y(_07181_));
 OAI21x1_ASAP7_75t_R _26753_ (.A1(_06534_),
    .A2(_06867_),
    .B(_06887_),
    .Y(_07182_));
 AOI22x1_ASAP7_75t_R _26754_ (.A1(_07180_),
    .A2(_07181_),
    .B1(_07182_),
    .B2(_06840_),
    .Y(_02480_));
 INVx1_ASAP7_75t_R _26755_ (.A(_06380_),
    .Y(_07183_));
 OR3x2_ASAP7_75t_R _26756_ (.A(_06359_),
    .B(_02093_),
    .C(_07170_),
    .Y(_07184_));
 NOR3x1_ASAP7_75t_R _26757_ (.A(_07183_),
    .B(_06919_),
    .C(_07184_),
    .Y(_07185_));
 AO21x1_ASAP7_75t_R _26758_ (.A1(_06738_),
    .A2(_06907_),
    .B(_07185_),
    .Y(_07186_));
 NAND2x1_ASAP7_75t_R _26759_ (.A(_06844_),
    .B(_07184_),
    .Y(_07187_));
 AOI21x1_ASAP7_75t_R _26760_ (.A1(_07138_),
    .A2(_07187_),
    .B(_06380_),
    .Y(_07188_));
 AO21x1_ASAP7_75t_R _26761_ (.A1(_07019_),
    .A2(_07186_),
    .B(_07188_),
    .Y(_02481_));
 NOR2x1_ASAP7_75t_R _26762_ (.A(_06380_),
    .B(_06359_),
    .Y(_07189_));
 AO32x1_ASAP7_75t_R _26763_ (.A1(_02089_),
    .A2(_07176_),
    .A3(_07189_),
    .B1(_06411_),
    .B2(_06940_),
    .Y(_07190_));
 OR3x1_ASAP7_75t_R _26764_ (.A(_06380_),
    .B(_06359_),
    .C(_07175_),
    .Y(_07191_));
 NAND2x1_ASAP7_75t_R _26765_ (.A(_06844_),
    .B(_07191_),
    .Y(_07192_));
 AOI21x1_ASAP7_75t_R _26766_ (.A1(_07138_),
    .A2(_07192_),
    .B(_02089_),
    .Y(_07193_));
 AO21x1_ASAP7_75t_R _26767_ (.A1(_07019_),
    .A2(_07190_),
    .B(_07193_),
    .Y(_02482_));
 OR5x2_ASAP7_75t_R _26768_ (.A(_02089_),
    .B(_06380_),
    .C(_06359_),
    .D(_02093_),
    .E(_07170_),
    .Y(_07194_));
 INVx1_ASAP7_75t_R _26769_ (.A(_07194_),
    .Y(_07195_));
 AND3x1_ASAP7_75t_R _26770_ (.A(_02088_),
    .B(_06930_),
    .C(_07195_),
    .Y(_07196_));
 AO21x1_ASAP7_75t_R _26771_ (.A1(_06750_),
    .A2(_06907_),
    .B(_07196_),
    .Y(_07197_));
 NAND2x1_ASAP7_75t_R _26772_ (.A(_06844_),
    .B(_07194_),
    .Y(_07198_));
 AOI21x1_ASAP7_75t_R _26773_ (.A1(_07138_),
    .A2(_07198_),
    .B(_02088_),
    .Y(_07199_));
 AO21x1_ASAP7_75t_R _26774_ (.A1(_07019_),
    .A2(_07197_),
    .B(_07199_),
    .Y(_02483_));
 INVx1_ASAP7_75t_R _26775_ (.A(_02087_),
    .Y(_07200_));
 OR5x1_ASAP7_75t_R _26776_ (.A(_02088_),
    .B(_02089_),
    .C(_06380_),
    .D(_06359_),
    .E(_07175_),
    .Y(_07201_));
 OR3x1_ASAP7_75t_R _26777_ (.A(_07200_),
    .B(_06919_),
    .C(_07201_),
    .Y(_07202_));
 OAI21x1_ASAP7_75t_R _26778_ (.A1(_06455_),
    .A2(_06930_),
    .B(_07202_),
    .Y(_07203_));
 NAND2x1_ASAP7_75t_R _26779_ (.A(_06844_),
    .B(_07201_),
    .Y(_07204_));
 AOI21x1_ASAP7_75t_R _26780_ (.A1(_07015_),
    .A2(_07204_),
    .B(_02087_),
    .Y(_07205_));
 AO21x1_ASAP7_75t_R _26781_ (.A1(_07019_),
    .A2(_07203_),
    .B(_07205_),
    .Y(_02484_));
 OAI22x1_ASAP7_75t_R _26782_ (.A1(_06559_),
    .A2(_06915_),
    .B1(_06852_),
    .B2(_06547_),
    .Y(_07206_));
 OA211x2_ASAP7_75t_R _26783_ (.A1(_06901_),
    .A2(_06852_),
    .B(_06920_),
    .C(_06547_),
    .Y(_07207_));
 AOI21x1_ASAP7_75t_R _26784_ (.A1(_06914_),
    .A2(_07206_),
    .B(_07207_),
    .Y(_02485_));
 OR3x1_ASAP7_75t_R _26785_ (.A(_02085_),
    .B(_06547_),
    .C(_06887_),
    .Y(_07208_));
 OA21x2_ASAP7_75t_R _26786_ (.A1(_06584_),
    .A2(_06886_),
    .B(_07208_),
    .Y(_07209_));
 INVx1_ASAP7_75t_R _26787_ (.A(_06547_),
    .Y(_07210_));
 NAND2x1_ASAP7_75t_R _26788_ (.A(_02085_),
    .B(_06856_),
    .Y(_07211_));
 AO21x1_ASAP7_75t_R _26789_ (.A1(_07210_),
    .A2(_06875_),
    .B(_07211_),
    .Y(_07212_));
 OA21x2_ASAP7_75t_R _26790_ (.A1(_06857_),
    .A2(_07209_),
    .B(_07212_),
    .Y(_02486_));
 AND2x2_ASAP7_75t_R _26791_ (.A(_02084_),
    .B(_06863_),
    .Y(_07213_));
 OR5x1_ASAP7_75t_R _26792_ (.A(_02085_),
    .B(_06547_),
    .C(_06855_),
    .D(_06919_),
    .E(_06851_),
    .Y(_07214_));
 OR3x1_ASAP7_75t_R _26793_ (.A(_02084_),
    .B(_02085_),
    .C(_06547_),
    .Y(_07215_));
 OAI22x1_ASAP7_75t_R _26794_ (.A1(_06609_),
    .A2(_06867_),
    .B1(_07215_),
    .B2(_06852_),
    .Y(_07216_));
 AOI22x1_ASAP7_75t_R _26795_ (.A1(_07213_),
    .A2(_07214_),
    .B1(_07216_),
    .B2(_06840_),
    .Y(_02487_));
 AND2x2_ASAP7_75t_R _26796_ (.A(_02083_),
    .B(_06878_),
    .Y(_07217_));
 OR4x1_ASAP7_75t_R _26797_ (.A(_06901_),
    .B(_06902_),
    .C(_07215_),
    .D(_06870_),
    .Y(_07218_));
 OAI22x1_ASAP7_75t_R _26798_ (.A1(_06627_),
    .A2(_06844_),
    .B1(_06846_),
    .B2(_06887_),
    .Y(_07219_));
 AND2x2_ASAP7_75t_R _26799_ (.A(_06839_),
    .B(_07219_),
    .Y(_07220_));
 AOI21x1_ASAP7_75t_R _26800_ (.A1(_07217_),
    .A2(_07218_),
    .B(_07220_),
    .Y(_02488_));
 OA21x2_ASAP7_75t_R _26801_ (.A1(_00783_),
    .A2(_05331_),
    .B(_05332_),
    .Y(_07221_));
 NOR3x2_ASAP7_75t_R _26802_ (.B(_07221_),
    .C(_05430_),
    .Y(_07222_),
    .A(_05421_));
 AO21x1_ASAP7_75t_R _26803_ (.A1(_07221_),
    .A2(_05455_),
    .B(_07222_),
    .Y(_07223_));
 OR2x4_ASAP7_75t_R _26804_ (.A(_15811_),
    .B(_05453_),
    .Y(_07224_));
 OR2x2_ASAP7_75t_R _26805_ (.A(_05378_),
    .B(_05383_),
    .Y(_07225_));
 BUFx4f_ASAP7_75t_R _26806_ (.A(_07225_),
    .Y(_07226_));
 AO221x2_ASAP7_75t_R _26807_ (.A1(_04945_),
    .A2(_07223_),
    .B1(_07224_),
    .B2(_05455_),
    .C(_07226_),
    .Y(_07227_));
 NOR2x1_ASAP7_75t_R _26808_ (.A(_02081_),
    .B(_05418_),
    .Y(_07228_));
 INVx1_ASAP7_75t_R _26809_ (.A(_01853_),
    .Y(_07229_));
 BUFx6f_ASAP7_75t_R _26810_ (.A(_05413_),
    .Y(_07230_));
 NAND2x1_ASAP7_75t_R _26811_ (.A(_14812_),
    .B(_07230_),
    .Y(_07231_));
 OA211x2_ASAP7_75t_R _26812_ (.A1(_07229_),
    .A2(_07230_),
    .B(_05418_),
    .C(_07231_),
    .Y(_07232_));
 OR3x1_ASAP7_75t_R _26813_ (.A(_07227_),
    .B(_07228_),
    .C(_07232_),
    .Y(_02489_));
 NOR2x1_ASAP7_75t_R _26814_ (.A(_02078_),
    .B(_05418_),
    .Y(_07233_));
 INVx1_ASAP7_75t_R _26815_ (.A(_01852_),
    .Y(_07234_));
 NAND2x1_ASAP7_75t_R _26816_ (.A(_05068_),
    .B(_07230_),
    .Y(_07235_));
 OA211x2_ASAP7_75t_R _26817_ (.A1(_07234_),
    .A2(_07230_),
    .B(_05418_),
    .C(_07235_),
    .Y(_07236_));
 OR3x1_ASAP7_75t_R _26818_ (.A(_07227_),
    .B(_07233_),
    .C(_07236_),
    .Y(_02490_));
 OR3x1_ASAP7_75t_R _26819_ (.A(_05059_),
    .B(_05765_),
    .C(_06186_),
    .Y(_07237_));
 BUFx4f_ASAP7_75t_R _26820_ (.A(_07237_),
    .Y(_07238_));
 NAND2x1_ASAP7_75t_R _26821_ (.A(_02080_),
    .B(_07238_),
    .Y(_07239_));
 OA21x2_ASAP7_75t_R _26822_ (.A1(_06639_),
    .A2(_07238_),
    .B(_07239_),
    .Y(_02492_));
 NAND2x1_ASAP7_75t_R _26823_ (.A(_00783_),
    .B(_07238_),
    .Y(_07240_));
 OA21x2_ASAP7_75t_R _26824_ (.A1(_06883_),
    .A2(_07238_),
    .B(_07240_),
    .Y(_02493_));
 NAND2x1_ASAP7_75t_R _26825_ (.A(_02079_),
    .B(_07238_),
    .Y(_07241_));
 OA21x2_ASAP7_75t_R _26826_ (.A1(_06650_),
    .A2(_07238_),
    .B(_07241_),
    .Y(_02494_));
 NAND2x1_ASAP7_75t_R _26827_ (.A(_00790_),
    .B(_07238_),
    .Y(_07242_));
 OA21x2_ASAP7_75t_R _26828_ (.A1(_06660_),
    .A2(_07238_),
    .B(_07242_),
    .Y(_02495_));
 NAND2x1_ASAP7_75t_R _26829_ (.A(_01460_),
    .B(_07238_),
    .Y(_07243_));
 OA21x2_ASAP7_75t_R _26830_ (.A1(_05872_),
    .A2(_07238_),
    .B(_07243_),
    .Y(_02497_));
 AOI21x1_ASAP7_75t_R _26831_ (.A1(_04945_),
    .A2(_07222_),
    .B(_05383_),
    .Y(_07244_));
 BUFx6f_ASAP7_75t_R _26832_ (.A(_07244_),
    .Y(_07245_));
 AOI22x1_ASAP7_75t_R _26833_ (.A1(_05379_),
    .A2(_05383_),
    .B1(_07245_),
    .B2(_02077_),
    .Y(_02498_));
 INVx1_ASAP7_75t_R _26834_ (.A(_02076_),
    .Y(_07246_));
 AO32x1_ASAP7_75t_R _26835_ (.A1(net105),
    .A2(_01460_),
    .A3(_05383_),
    .B1(_07245_),
    .B2(_07246_),
    .Y(_02499_));
 INVx1_ASAP7_75t_R _26836_ (.A(_02075_),
    .Y(_07247_));
 AO32x1_ASAP7_75t_R _26837_ (.A1(_05379_),
    .A2(_05421_),
    .A3(_05381_),
    .B1(_07245_),
    .B2(_07247_),
    .Y(_02500_));
 NOR2x2_ASAP7_75t_R _26838_ (.A(_05916_),
    .B(_05858_),
    .Y(_07248_));
 BUFx3_ASAP7_75t_R _26839_ (.A(_07248_),
    .Y(_07249_));
 AO21x1_ASAP7_75t_R _26840_ (.A1(_04945_),
    .A2(_07222_),
    .B(_05383_),
    .Y(_07250_));
 BUFx6f_ASAP7_75t_R _26841_ (.A(_07250_),
    .Y(_07251_));
 NOR2x2_ASAP7_75t_R _26842_ (.A(_07251_),
    .B(_07248_),
    .Y(_07252_));
 BUFx4f_ASAP7_75t_R _26843_ (.A(_07252_),
    .Y(_07253_));
 INVx1_ASAP7_75t_R _26844_ (.A(_02074_),
    .Y(_07254_));
 BUFx3_ASAP7_75t_R _26845_ (.A(_01681_),
    .Y(_07255_));
 BUFx3_ASAP7_75t_R _26846_ (.A(_07226_),
    .Y(_07256_));
 NOR2x2_ASAP7_75t_R _26847_ (.A(_05378_),
    .B(_05383_),
    .Y(_07257_));
 BUFx3_ASAP7_75t_R _26848_ (.A(_07257_),
    .Y(_07258_));
 AND2x2_ASAP7_75t_R _26849_ (.A(_00039_),
    .B(_07258_),
    .Y(_07259_));
 AO21x2_ASAP7_75t_R _26850_ (.A1(_07255_),
    .A2(_07256_),
    .B(_07259_),
    .Y(_07260_));
 NOR2x1_ASAP7_75t_R _26851_ (.A(_07245_),
    .B(_07260_),
    .Y(_07261_));
 AO221x1_ASAP7_75t_R _26852_ (.A1(_06635_),
    .A2(_07249_),
    .B1(_07253_),
    .B2(_07254_),
    .C(_07261_),
    .Y(_02501_));
 INVx1_ASAP7_75t_R _26853_ (.A(_02073_),
    .Y(_07262_));
 BUFx4f_ASAP7_75t_R _26854_ (.A(_07226_),
    .Y(_07263_));
 AND2x2_ASAP7_75t_R _26855_ (.A(_00042_),
    .B(_07257_),
    .Y(_07264_));
 AO21x2_ASAP7_75t_R _26856_ (.A1(_01709_),
    .A2(_07263_),
    .B(_07264_),
    .Y(_07265_));
 NOR2x1_ASAP7_75t_R _26857_ (.A(_07245_),
    .B(_07265_),
    .Y(_07266_));
 AO221x1_ASAP7_75t_R _26858_ (.A1(_06639_),
    .A2(_07249_),
    .B1(_07253_),
    .B2(_07262_),
    .C(_07266_),
    .Y(_02502_));
 INVx1_ASAP7_75t_R _26859_ (.A(_02072_),
    .Y(_07267_));
 AND2x2_ASAP7_75t_R _26860_ (.A(_00044_),
    .B(_07257_),
    .Y(_07268_));
 AO21x2_ASAP7_75t_R _26861_ (.A1(_01708_),
    .A2(_07263_),
    .B(_07268_),
    .Y(_07269_));
 NOR2x1_ASAP7_75t_R _26862_ (.A(_07245_),
    .B(_07269_),
    .Y(_07270_));
 AO221x1_ASAP7_75t_R _26863_ (.A1(_06883_),
    .A2(_07249_),
    .B1(_07253_),
    .B2(_07267_),
    .C(_07270_),
    .Y(_02503_));
 INVx1_ASAP7_75t_R _26864_ (.A(_02071_),
    .Y(_07271_));
 AND2x2_ASAP7_75t_R _26865_ (.A(_00046_),
    .B(_07258_),
    .Y(_07272_));
 AO21x2_ASAP7_75t_R _26866_ (.A1(_01707_),
    .A2(_07256_),
    .B(_07272_),
    .Y(_07273_));
 NOR2x1_ASAP7_75t_R _26867_ (.A(_07245_),
    .B(_07273_),
    .Y(_07274_));
 AO221x1_ASAP7_75t_R _26868_ (.A1(_06650_),
    .A2(_07249_),
    .B1(_07253_),
    .B2(_07271_),
    .C(_07274_),
    .Y(_02504_));
 INVx1_ASAP7_75t_R _26869_ (.A(_02070_),
    .Y(_07275_));
 BUFx3_ASAP7_75t_R _26870_ (.A(_01706_),
    .Y(_07276_));
 AND2x2_ASAP7_75t_R _26871_ (.A(_00048_),
    .B(_07257_),
    .Y(_07277_));
 AO21x1_ASAP7_75t_R _26872_ (.A1(_07276_),
    .A2(_07263_),
    .B(_07277_),
    .Y(_07278_));
 NOR2x1_ASAP7_75t_R _26873_ (.A(_07245_),
    .B(_07278_),
    .Y(_07279_));
 AO221x1_ASAP7_75t_R _26874_ (.A1(_06065_),
    .A2(_07249_),
    .B1(_07253_),
    .B2(_07275_),
    .C(_07279_),
    .Y(_02505_));
 BUFx4f_ASAP7_75t_R _26875_ (.A(_07252_),
    .Y(_07280_));
 INVx1_ASAP7_75t_R _26876_ (.A(_02069_),
    .Y(_07281_));
 AND2x2_ASAP7_75t_R _26877_ (.A(_00050_),
    .B(_07258_),
    .Y(_07282_));
 AO21x2_ASAP7_75t_R _26878_ (.A1(_01705_),
    .A2(_07256_),
    .B(_07282_),
    .Y(_07283_));
 NOR2x1_ASAP7_75t_R _26879_ (.A(_07245_),
    .B(_07283_),
    .Y(_07284_));
 AO221x1_ASAP7_75t_R _26880_ (.A1(_06660_),
    .A2(_07249_),
    .B1(_07280_),
    .B2(_07281_),
    .C(_07284_),
    .Y(_02506_));
 INVx1_ASAP7_75t_R _26881_ (.A(_02068_),
    .Y(_07285_));
 BUFx3_ASAP7_75t_R _26882_ (.A(_01704_),
    .Y(_07286_));
 AND2x2_ASAP7_75t_R _26883_ (.A(_00051_),
    .B(_07257_),
    .Y(_07287_));
 AO21x2_ASAP7_75t_R _26884_ (.A1(_07286_),
    .A2(_07226_),
    .B(_07287_),
    .Y(_07288_));
 NOR2x1_ASAP7_75t_R _26885_ (.A(_07245_),
    .B(_07288_),
    .Y(_07289_));
 AO221x1_ASAP7_75t_R _26886_ (.A1(_06111_),
    .A2(_07249_),
    .B1(_07280_),
    .B2(_07285_),
    .C(_07289_),
    .Y(_02507_));
 INVx1_ASAP7_75t_R _26887_ (.A(_02067_),
    .Y(_07290_));
 BUFx6f_ASAP7_75t_R _26888_ (.A(_07244_),
    .Y(_07291_));
 BUFx6f_ASAP7_75t_R _26889_ (.A(_07291_),
    .Y(_07292_));
 BUFx3_ASAP7_75t_R _26890_ (.A(_01703_),
    .Y(_07293_));
 AND2x2_ASAP7_75t_R _26891_ (.A(_00052_),
    .B(_07258_),
    .Y(_07294_));
 AO21x2_ASAP7_75t_R _26892_ (.A1(_07293_),
    .A2(_07256_),
    .B(_07294_),
    .Y(_07295_));
 NOR2x1_ASAP7_75t_R _26893_ (.A(_07292_),
    .B(_07295_),
    .Y(_07296_));
 AO221x1_ASAP7_75t_R _26894_ (.A1(_06137_),
    .A2(_07249_),
    .B1(_07280_),
    .B2(_07290_),
    .C(_07296_),
    .Y(_02508_));
 INVx1_ASAP7_75t_R _26895_ (.A(_02066_),
    .Y(_07297_));
 AND2x2_ASAP7_75t_R _26896_ (.A(_00053_),
    .B(_07258_),
    .Y(_07298_));
 AO21x2_ASAP7_75t_R _26897_ (.A1(_01702_),
    .A2(_07256_),
    .B(_07298_),
    .Y(_07299_));
 NOR2x1_ASAP7_75t_R _26898_ (.A(_07292_),
    .B(_07299_),
    .Y(_07300_));
 AO221x1_ASAP7_75t_R _26899_ (.A1(_06161_),
    .A2(_07249_),
    .B1(_07280_),
    .B2(_07297_),
    .C(_07300_),
    .Y(_02509_));
 INVx1_ASAP7_75t_R _26900_ (.A(_02065_),
    .Y(_07301_));
 BUFx4f_ASAP7_75t_R _26901_ (.A(_01701_),
    .Y(_07302_));
 AND2x2_ASAP7_75t_R _26902_ (.A(_00054_),
    .B(_07258_),
    .Y(_07303_));
 AO21x2_ASAP7_75t_R _26903_ (.A1(_07302_),
    .A2(_07256_),
    .B(_07303_),
    .Y(_07304_));
 NOR2x1_ASAP7_75t_R _26904_ (.A(_07292_),
    .B(_07304_),
    .Y(_07305_));
 AO221x1_ASAP7_75t_R _26905_ (.A1(_06180_),
    .A2(_07249_),
    .B1(_07280_),
    .B2(_07301_),
    .C(_07305_),
    .Y(_02510_));
 BUFx4f_ASAP7_75t_R _26906_ (.A(_07248_),
    .Y(_07306_));
 INVx1_ASAP7_75t_R _26907_ (.A(_00789_),
    .Y(_07307_));
 BUFx4f_ASAP7_75t_R _26908_ (.A(_05471_),
    .Y(_07308_));
 BUFx4f_ASAP7_75t_R _26909_ (.A(_07308_),
    .Y(_07309_));
 BUFx4f_ASAP7_75t_R _26910_ (.A(_07309_),
    .Y(_07310_));
 BUFx3_ASAP7_75t_R _26911_ (.A(_07310_),
    .Y(_07311_));
 BUFx3_ASAP7_75t_R _26912_ (.A(_07311_),
    .Y(_07312_));
 BUFx4f_ASAP7_75t_R _26913_ (.A(_07312_),
    .Y(_07313_));
 BUFx3_ASAP7_75t_R _26914_ (.A(_07257_),
    .Y(_07314_));
 AND2x2_ASAP7_75t_R _26915_ (.A(_01544_),
    .B(_07314_),
    .Y(_07315_));
 AO21x1_ASAP7_75t_R _26916_ (.A1(_07313_),
    .A2(_07263_),
    .B(_07315_),
    .Y(_07316_));
 NOR2x1_ASAP7_75t_R _26917_ (.A(_07292_),
    .B(_07316_),
    .Y(_07317_));
 AO221x1_ASAP7_75t_R _26918_ (.A1(_06475_),
    .A2(_07306_),
    .B1(_07280_),
    .B2(_07307_),
    .C(_07317_),
    .Y(_02511_));
 INVx1_ASAP7_75t_R _26919_ (.A(_02064_),
    .Y(_07318_));
 AND2x2_ASAP7_75t_R _26920_ (.A(_00055_),
    .B(_07258_),
    .Y(_07319_));
 AO21x2_ASAP7_75t_R _26921_ (.A1(_01700_),
    .A2(_07256_),
    .B(_07319_),
    .Y(_07320_));
 NOR2x1_ASAP7_75t_R _26922_ (.A(_07292_),
    .B(_07320_),
    .Y(_07321_));
 AO221x1_ASAP7_75t_R _26923_ (.A1(_06218_),
    .A2(_07306_),
    .B1(_07280_),
    .B2(_07318_),
    .C(_07321_),
    .Y(_02512_));
 INVx1_ASAP7_75t_R _26924_ (.A(_02063_),
    .Y(_07322_));
 BUFx4f_ASAP7_75t_R _26925_ (.A(_07248_),
    .Y(_07323_));
 BUFx4f_ASAP7_75t_R _26926_ (.A(_07226_),
    .Y(_07324_));
 NAND2x1_ASAP7_75t_R _26927_ (.A(_01699_),
    .B(_07324_),
    .Y(_07325_));
 OA21x2_ASAP7_75t_R _26928_ (.A1(_16752_),
    .A2(_07256_),
    .B(_07325_),
    .Y(_07326_));
 AO22x1_ASAP7_75t_R _26929_ (.A1(_06695_),
    .A2(_07323_),
    .B1(_07326_),
    .B2(_07251_),
    .Y(_07327_));
 AO21x1_ASAP7_75t_R _26930_ (.A1(_07322_),
    .A2(_07253_),
    .B(_07327_),
    .Y(_02513_));
 INVx1_ASAP7_75t_R _26931_ (.A(_02062_),
    .Y(_07328_));
 AND2x2_ASAP7_75t_R _26932_ (.A(_00057_),
    .B(_07257_),
    .Y(_07329_));
 AO21x2_ASAP7_75t_R _26933_ (.A1(_01698_),
    .A2(_07226_),
    .B(_07329_),
    .Y(_07330_));
 NOR2x1_ASAP7_75t_R _26934_ (.A(_07292_),
    .B(_07330_),
    .Y(_07331_));
 AO221x1_ASAP7_75t_R _26935_ (.A1(_06260_),
    .A2(_07306_),
    .B1(_07280_),
    .B2(_07328_),
    .C(_07331_),
    .Y(_02514_));
 INVx1_ASAP7_75t_R _26936_ (.A(_02061_),
    .Y(_07332_));
 BUFx4f_ASAP7_75t_R _26937_ (.A(_01697_),
    .Y(_07333_));
 AND2x2_ASAP7_75t_R _26938_ (.A(_00058_),
    .B(_07258_),
    .Y(_07334_));
 AO21x2_ASAP7_75t_R _26939_ (.A1(_07333_),
    .A2(_07256_),
    .B(_07334_),
    .Y(_07335_));
 NOR2x1_ASAP7_75t_R _26940_ (.A(_07292_),
    .B(_07335_),
    .Y(_07336_));
 AO221x1_ASAP7_75t_R _26941_ (.A1(_06705_),
    .A2(_07306_),
    .B1(_07280_),
    .B2(_07332_),
    .C(_07336_),
    .Y(_02515_));
 INVx1_ASAP7_75t_R _26942_ (.A(_02060_),
    .Y(_07337_));
 AND2x2_ASAP7_75t_R _26943_ (.A(_00059_),
    .B(_07258_),
    .Y(_07338_));
 AO21x2_ASAP7_75t_R _26944_ (.A1(_01696_),
    .A2(_07324_),
    .B(_07338_),
    .Y(_07339_));
 NOR2x1_ASAP7_75t_R _26945_ (.A(_07292_),
    .B(_07339_),
    .Y(_07340_));
 AO221x1_ASAP7_75t_R _26946_ (.A1(_06299_),
    .A2(_07306_),
    .B1(_07280_),
    .B2(_07337_),
    .C(_07340_),
    .Y(_02516_));
 BUFx4f_ASAP7_75t_R _26947_ (.A(_07252_),
    .Y(_07341_));
 INVx1_ASAP7_75t_R _26948_ (.A(_02059_),
    .Y(_07342_));
 AND2x2_ASAP7_75t_R _26949_ (.A(_00060_),
    .B(_07257_),
    .Y(_07343_));
 AO21x1_ASAP7_75t_R _26950_ (.A1(_01695_),
    .A2(_07226_),
    .B(_07343_),
    .Y(_07344_));
 NOR2x1_ASAP7_75t_R _26951_ (.A(_07292_),
    .B(_07344_),
    .Y(_07345_));
 AO221x1_ASAP7_75t_R _26952_ (.A1(_06320_),
    .A2(_07306_),
    .B1(_07341_),
    .B2(_07342_),
    .C(_07345_),
    .Y(_02517_));
 AND2x2_ASAP7_75t_R _26953_ (.A(_00061_),
    .B(_07314_),
    .Y(_07346_));
 AO21x1_ASAP7_75t_R _26954_ (.A1(_01694_),
    .A2(_07263_),
    .B(_07346_),
    .Y(_07347_));
 AO22x1_ASAP7_75t_R _26955_ (.A1(_06347_),
    .A2(_07323_),
    .B1(_07347_),
    .B2(_07251_),
    .Y(_07348_));
 AOI21x1_ASAP7_75t_R _26956_ (.A1(_02058_),
    .A2(_07253_),
    .B(_07348_),
    .Y(_02518_));
 AND2x2_ASAP7_75t_R _26957_ (.A(_00062_),
    .B(_07257_),
    .Y(_07349_));
 AO21x1_ASAP7_75t_R _26958_ (.A1(_01693_),
    .A2(_07263_),
    .B(_07349_),
    .Y(_07350_));
 AO22x1_ASAP7_75t_R _26959_ (.A1(_06370_),
    .A2(_07323_),
    .B1(_07350_),
    .B2(_07251_),
    .Y(_07351_));
 AOI21x1_ASAP7_75t_R _26960_ (.A1(_02057_),
    .A2(_07253_),
    .B(_07351_),
    .Y(_02519_));
 INVx1_ASAP7_75t_R _26961_ (.A(_02056_),
    .Y(_07352_));
 AND2x2_ASAP7_75t_R _26962_ (.A(_00063_),
    .B(_07258_),
    .Y(_07353_));
 AO21x2_ASAP7_75t_R _26963_ (.A1(_01692_),
    .A2(_07324_),
    .B(_07353_),
    .Y(_07354_));
 NOR2x1_ASAP7_75t_R _26964_ (.A(_07292_),
    .B(_07354_),
    .Y(_07355_));
 AO221x1_ASAP7_75t_R _26965_ (.A1(_06738_),
    .A2(_07306_),
    .B1(_07341_),
    .B2(_07352_),
    .C(_07355_),
    .Y(_02520_));
 INVx1_ASAP7_75t_R _26966_ (.A(_02055_),
    .Y(_07356_));
 AND2x2_ASAP7_75t_R _26967_ (.A(_00064_),
    .B(_07314_),
    .Y(_07357_));
 AO21x2_ASAP7_75t_R _26968_ (.A1(_01691_),
    .A2(_07324_),
    .B(_07357_),
    .Y(_07358_));
 NOR2x1_ASAP7_75t_R _26969_ (.A(_07291_),
    .B(_07358_),
    .Y(_07359_));
 AO221x1_ASAP7_75t_R _26970_ (.A1(_06411_),
    .A2(_07306_),
    .B1(_07341_),
    .B2(_07356_),
    .C(_07359_),
    .Y(_02521_));
 INVx1_ASAP7_75t_R _26971_ (.A(_02054_),
    .Y(_07360_));
 AND2x2_ASAP7_75t_R _26972_ (.A(_00012_),
    .B(_07314_),
    .Y(_07361_));
 AO21x1_ASAP7_75t_R _26973_ (.A1(_18317_),
    .A2(_07263_),
    .B(_07361_),
    .Y(_07362_));
 NOR2x1_ASAP7_75t_R _26974_ (.A(_07291_),
    .B(_07362_),
    .Y(_07363_));
 AO221x1_ASAP7_75t_R _26975_ (.A1(_05872_),
    .A2(_07306_),
    .B1(_07341_),
    .B2(_07360_),
    .C(_07363_),
    .Y(_02522_));
 INVx1_ASAP7_75t_R _26976_ (.A(_02053_),
    .Y(_07364_));
 AND2x2_ASAP7_75t_R _26977_ (.A(_00065_),
    .B(_07314_),
    .Y(_07365_));
 AO21x2_ASAP7_75t_R _26978_ (.A1(_01690_),
    .A2(_07324_),
    .B(_07365_),
    .Y(_07366_));
 NOR2x1_ASAP7_75t_R _26979_ (.A(_07291_),
    .B(_07366_),
    .Y(_07367_));
 AO221x1_ASAP7_75t_R _26980_ (.A1(_06750_),
    .A2(_07306_),
    .B1(_07341_),
    .B2(_07364_),
    .C(_07367_),
    .Y(_02523_));
 INVx1_ASAP7_75t_R _26981_ (.A(_02052_),
    .Y(_07368_));
 INVx3_ASAP7_75t_R _26982_ (.A(_06455_),
    .Y(_07369_));
 NAND2x1_ASAP7_75t_R _26983_ (.A(_01688_),
    .B(_07263_),
    .Y(_07370_));
 OA21x2_ASAP7_75t_R _26984_ (.A1(_04864_),
    .A2(_07324_),
    .B(_07370_),
    .Y(_07371_));
 AO22x1_ASAP7_75t_R _26985_ (.A1(_07369_),
    .A2(_07323_),
    .B1(_07371_),
    .B2(_07251_),
    .Y(_07372_));
 AO21x1_ASAP7_75t_R _26986_ (.A1(_07368_),
    .A2(_07253_),
    .B(_07372_),
    .Y(_02524_));
 INVx1_ASAP7_75t_R _26987_ (.A(_01461_),
    .Y(_07373_));
 AND2x2_ASAP7_75t_R _26988_ (.A(_00020_),
    .B(_07314_),
    .Y(_07374_));
 AO21x2_ASAP7_75t_R _26989_ (.A1(_01689_),
    .A2(_07263_),
    .B(_07374_),
    .Y(_07375_));
 NOR2x1_ASAP7_75t_R _26990_ (.A(_07291_),
    .B(_07375_),
    .Y(_07376_));
 AO221x1_ASAP7_75t_R _26991_ (.A1(_06588_),
    .A2(_07323_),
    .B1(_07341_),
    .B2(_07373_),
    .C(_07376_),
    .Y(_02525_));
 INVx1_ASAP7_75t_R _26992_ (.A(_01462_),
    .Y(_07377_));
 BUFx4f_ASAP7_75t_R _26993_ (.A(_01687_),
    .Y(_07378_));
 AND2x2_ASAP7_75t_R _26994_ (.A(_00023_),
    .B(_07314_),
    .Y(_07379_));
 AO21x1_ASAP7_75t_R _26995_ (.A1(_07378_),
    .A2(_07263_),
    .B(_07379_),
    .Y(_07380_));
 NOR2x1_ASAP7_75t_R _26996_ (.A(_07291_),
    .B(_07380_),
    .Y(_07381_));
 AO221x1_ASAP7_75t_R _26997_ (.A1(_07042_),
    .A2(_07323_),
    .B1(_07341_),
    .B2(_07377_),
    .C(_07381_),
    .Y(_02526_));
 INVx1_ASAP7_75t_R _26998_ (.A(_01463_),
    .Y(_07382_));
 BUFx3_ASAP7_75t_R _26999_ (.A(_01686_),
    .Y(_07383_));
 NAND2x1_ASAP7_75t_R _27000_ (.A(_07383_),
    .B(_07324_),
    .Y(_07384_));
 OA21x2_ASAP7_75t_R _27001_ (.A1(_15116_),
    .A2(_07256_),
    .B(_07384_),
    .Y(_07385_));
 AO22x1_ASAP7_75t_R _27002_ (.A1(_06534_),
    .A2(_07248_),
    .B1(_07385_),
    .B2(_07251_),
    .Y(_07386_));
 AO21x1_ASAP7_75t_R _27003_ (.A1(_07382_),
    .A2(_07253_),
    .B(_07386_),
    .Y(_02527_));
 INVx1_ASAP7_75t_R _27004_ (.A(_01464_),
    .Y(_07387_));
 AND2x2_ASAP7_75t_R _27005_ (.A(_00028_),
    .B(_07314_),
    .Y(_07388_));
 AO21x2_ASAP7_75t_R _27006_ (.A1(_01685_),
    .A2(_07324_),
    .B(_07388_),
    .Y(_07389_));
 NOR2x1_ASAP7_75t_R _27007_ (.A(_07291_),
    .B(_07389_),
    .Y(_07390_));
 AO221x1_ASAP7_75t_R _27008_ (.A1(_06559_),
    .A2(_07323_),
    .B1(_07341_),
    .B2(_07387_),
    .C(_07390_),
    .Y(_02528_));
 INVx1_ASAP7_75t_R _27009_ (.A(_02051_),
    .Y(_07391_));
 BUFx4f_ASAP7_75t_R _27010_ (.A(_01684_),
    .Y(_07392_));
 AND2x2_ASAP7_75t_R _27011_ (.A(_00030_),
    .B(_07314_),
    .Y(_07393_));
 AO21x1_ASAP7_75t_R _27012_ (.A1(_07392_),
    .A2(_07324_),
    .B(_07393_),
    .Y(_07394_));
 NOR2x1_ASAP7_75t_R _27013_ (.A(_07291_),
    .B(_07394_),
    .Y(_07395_));
 AO221x1_ASAP7_75t_R _27014_ (.A1(_06584_),
    .A2(_07323_),
    .B1(_07341_),
    .B2(_07391_),
    .C(_07395_),
    .Y(_02529_));
 INVx1_ASAP7_75t_R _27015_ (.A(_02050_),
    .Y(_07396_));
 BUFx4f_ASAP7_75t_R _27016_ (.A(_01683_),
    .Y(_07397_));
 AND2x2_ASAP7_75t_R _27017_ (.A(_00033_),
    .B(_07257_),
    .Y(_07398_));
 AO21x1_ASAP7_75t_R _27018_ (.A1(_07397_),
    .A2(_07226_),
    .B(_07398_),
    .Y(_07399_));
 NOR2x1_ASAP7_75t_R _27019_ (.A(_07291_),
    .B(_07399_),
    .Y(_07400_));
 AO221x1_ASAP7_75t_R _27020_ (.A1(_06609_),
    .A2(_07323_),
    .B1(_07341_),
    .B2(_07396_),
    .C(_07400_),
    .Y(_02530_));
 INVx1_ASAP7_75t_R _27021_ (.A(_02049_),
    .Y(_07401_));
 AND2x2_ASAP7_75t_R _27022_ (.A(_00036_),
    .B(_07314_),
    .Y(_07402_));
 AO21x1_ASAP7_75t_R _27023_ (.A1(_01682_),
    .A2(_07324_),
    .B(_07402_),
    .Y(_07403_));
 NOR2x1_ASAP7_75t_R _27024_ (.A(_07291_),
    .B(_07403_),
    .Y(_07404_));
 AO221x1_ASAP7_75t_R _27025_ (.A1(_06627_),
    .A2(_07323_),
    .B1(_07252_),
    .B2(_07401_),
    .C(_07404_),
    .Y(_02531_));
 OR3x1_ASAP7_75t_R _27026_ (.A(_05059_),
    .B(_05765_),
    .C(_05949_),
    .Y(_07405_));
 BUFx6f_ASAP7_75t_R _27027_ (.A(_07405_),
    .Y(_07406_));
 BUFx4f_ASAP7_75t_R _27028_ (.A(_07406_),
    .Y(_07407_));
 BUFx6f_ASAP7_75t_R _27029_ (.A(_07406_),
    .Y(_07408_));
 NAND2x1_ASAP7_75t_R _27030_ (.A(_02048_),
    .B(_07408_),
    .Y(_07409_));
 OA21x2_ASAP7_75t_R _27031_ (.A1(_05841_),
    .A2(_07407_),
    .B(_07409_),
    .Y(_02532_));
 NAND2x1_ASAP7_75t_R _27032_ (.A(_02047_),
    .B(_07408_),
    .Y(_07410_));
 OA21x2_ASAP7_75t_R _27033_ (.A1(_06635_),
    .A2(_07407_),
    .B(_07410_),
    .Y(_02533_));
 NAND2x1_ASAP7_75t_R _27034_ (.A(_02046_),
    .B(_07408_),
    .Y(_07411_));
 OA21x2_ASAP7_75t_R _27035_ (.A1(_06639_),
    .A2(_07407_),
    .B(_07411_),
    .Y(_02534_));
 NAND2x1_ASAP7_75t_R _27036_ (.A(_02045_),
    .B(_07408_),
    .Y(_07412_));
 OA21x2_ASAP7_75t_R _27037_ (.A1(_06883_),
    .A2(_07407_),
    .B(_07412_),
    .Y(_02535_));
 NAND2x1_ASAP7_75t_R _27038_ (.A(_02044_),
    .B(_07408_),
    .Y(_07413_));
 OA21x2_ASAP7_75t_R _27039_ (.A1(_06650_),
    .A2(_07407_),
    .B(_07413_),
    .Y(_02536_));
 NAND2x1_ASAP7_75t_R _27040_ (.A(_02043_),
    .B(_07408_),
    .Y(_07414_));
 OA21x2_ASAP7_75t_R _27041_ (.A1(_06065_),
    .A2(_07407_),
    .B(_07414_),
    .Y(_02537_));
 NAND2x1_ASAP7_75t_R _27042_ (.A(_02042_),
    .B(_07408_),
    .Y(_07415_));
 OA21x2_ASAP7_75t_R _27043_ (.A1(_06660_),
    .A2(_07407_),
    .B(_07415_),
    .Y(_02538_));
 NAND2x1_ASAP7_75t_R _27044_ (.A(_02041_),
    .B(_07408_),
    .Y(_07416_));
 OA21x2_ASAP7_75t_R _27045_ (.A1(_06111_),
    .A2(_07407_),
    .B(_07416_),
    .Y(_02539_));
 BUFx6f_ASAP7_75t_R _27046_ (.A(_07406_),
    .Y(_07417_));
 NAND2x1_ASAP7_75t_R _27047_ (.A(_02040_),
    .B(_07417_),
    .Y(_07418_));
 OA21x2_ASAP7_75t_R _27048_ (.A1(_06137_),
    .A2(_07407_),
    .B(_07418_),
    .Y(_02540_));
 NAND2x1_ASAP7_75t_R _27049_ (.A(_02039_),
    .B(_07417_),
    .Y(_07419_));
 OA21x2_ASAP7_75t_R _27050_ (.A1(_06161_),
    .A2(_07407_),
    .B(_07419_),
    .Y(_02541_));
 BUFx4f_ASAP7_75t_R _27051_ (.A(_07406_),
    .Y(_07420_));
 NAND2x1_ASAP7_75t_R _27052_ (.A(_02038_),
    .B(_07417_),
    .Y(_07421_));
 OA21x2_ASAP7_75t_R _27053_ (.A1(_06180_),
    .A2(_07420_),
    .B(_07421_),
    .Y(_02542_));
 NAND2x1_ASAP7_75t_R _27054_ (.A(_02037_),
    .B(_07417_),
    .Y(_07422_));
 OA21x2_ASAP7_75t_R _27055_ (.A1(_06475_),
    .A2(_07420_),
    .B(_07422_),
    .Y(_02543_));
 NAND2x1_ASAP7_75t_R _27056_ (.A(_02036_),
    .B(_07417_),
    .Y(_07423_));
 OA21x2_ASAP7_75t_R _27057_ (.A1(_06218_),
    .A2(_07420_),
    .B(_07423_),
    .Y(_02544_));
 NAND2x1_ASAP7_75t_R _27058_ (.A(_02035_),
    .B(_07417_),
    .Y(_07424_));
 OA21x2_ASAP7_75t_R _27059_ (.A1(_06695_),
    .A2(_07420_),
    .B(_07424_),
    .Y(_02545_));
 NAND2x1_ASAP7_75t_R _27060_ (.A(_02034_),
    .B(_07417_),
    .Y(_07425_));
 OA21x2_ASAP7_75t_R _27061_ (.A1(_06260_),
    .A2(_07420_),
    .B(_07425_),
    .Y(_02546_));
 NAND2x1_ASAP7_75t_R _27062_ (.A(_02033_),
    .B(_07417_),
    .Y(_07426_));
 OA21x2_ASAP7_75t_R _27063_ (.A1(_06705_),
    .A2(_07420_),
    .B(_07426_),
    .Y(_02547_));
 NAND2x1_ASAP7_75t_R _27064_ (.A(_02032_),
    .B(_07417_),
    .Y(_07427_));
 OA21x2_ASAP7_75t_R _27065_ (.A1(_06299_),
    .A2(_07420_),
    .B(_07427_),
    .Y(_02548_));
 NAND2x1_ASAP7_75t_R _27066_ (.A(_02031_),
    .B(_07417_),
    .Y(_07428_));
 OA21x2_ASAP7_75t_R _27067_ (.A1(_06320_),
    .A2(_07420_),
    .B(_07428_),
    .Y(_02549_));
 BUFx6f_ASAP7_75t_R _27068_ (.A(_07406_),
    .Y(_07429_));
 NAND2x1_ASAP7_75t_R _27069_ (.A(_02030_),
    .B(_07429_),
    .Y(_07430_));
 OA21x2_ASAP7_75t_R _27070_ (.A1(_06968_),
    .A2(_07420_),
    .B(_07430_),
    .Y(_02550_));
 INVx2_ASAP7_75t_R _27071_ (.A(_06370_),
    .Y(_07431_));
 NAND2x1_ASAP7_75t_R _27072_ (.A(_02029_),
    .B(_07429_),
    .Y(_07432_));
 OA21x2_ASAP7_75t_R _27073_ (.A1(_07431_),
    .A2(_07420_),
    .B(_07432_),
    .Y(_02551_));
 BUFx4f_ASAP7_75t_R _27074_ (.A(_07406_),
    .Y(_07433_));
 NAND2x1_ASAP7_75t_R _27075_ (.A(_02028_),
    .B(_07429_),
    .Y(_07434_));
 OA21x2_ASAP7_75t_R _27076_ (.A1(_06738_),
    .A2(_07433_),
    .B(_07434_),
    .Y(_02552_));
 NAND2x1_ASAP7_75t_R _27077_ (.A(_02027_),
    .B(_07429_),
    .Y(_07435_));
 OA21x2_ASAP7_75t_R _27078_ (.A1(_06411_),
    .A2(_07433_),
    .B(_07435_),
    .Y(_02553_));
 NAND2x1_ASAP7_75t_R _27079_ (.A(_02026_),
    .B(_07429_),
    .Y(_07436_));
 OA21x2_ASAP7_75t_R _27080_ (.A1(_05872_),
    .A2(_07433_),
    .B(_07436_),
    .Y(_02554_));
 NAND2x1_ASAP7_75t_R _27081_ (.A(_02025_),
    .B(_07429_),
    .Y(_07437_));
 OA21x2_ASAP7_75t_R _27082_ (.A1(_06750_),
    .A2(_07433_),
    .B(_07437_),
    .Y(_02555_));
 NAND2x1_ASAP7_75t_R _27083_ (.A(_02024_),
    .B(_07429_),
    .Y(_07438_));
 OA21x2_ASAP7_75t_R _27084_ (.A1(_07369_),
    .A2(_07433_),
    .B(_07438_),
    .Y(_02556_));
 NAND2x1_ASAP7_75t_R _27085_ (.A(_02023_),
    .B(_07429_),
    .Y(_07439_));
 OA21x2_ASAP7_75t_R _27086_ (.A1(_06588_),
    .A2(_07433_),
    .B(_07439_),
    .Y(_02557_));
 NAND2x1_ASAP7_75t_R _27087_ (.A(_02022_),
    .B(_07429_),
    .Y(_07440_));
 OA21x2_ASAP7_75t_R _27088_ (.A1(_07042_),
    .A2(_07433_),
    .B(_07440_),
    .Y(_02558_));
 NAND2x1_ASAP7_75t_R _27089_ (.A(_02021_),
    .B(_07429_),
    .Y(_07441_));
 OA21x2_ASAP7_75t_R _27090_ (.A1(_06534_),
    .A2(_07433_),
    .B(_07441_),
    .Y(_02559_));
 NAND2x1_ASAP7_75t_R _27091_ (.A(_02020_),
    .B(_07406_),
    .Y(_07442_));
 OA21x2_ASAP7_75t_R _27092_ (.A1(_06559_),
    .A2(_07433_),
    .B(_07442_),
    .Y(_02560_));
 NAND2x1_ASAP7_75t_R _27093_ (.A(_02019_),
    .B(_07406_),
    .Y(_07443_));
 OA21x2_ASAP7_75t_R _27094_ (.A1(_06584_),
    .A2(_07433_),
    .B(_07443_),
    .Y(_02561_));
 NAND2x1_ASAP7_75t_R _27095_ (.A(_02018_),
    .B(_07406_),
    .Y(_07444_));
 OA21x2_ASAP7_75t_R _27096_ (.A1(_06609_),
    .A2(_07408_),
    .B(_07444_),
    .Y(_02562_));
 NAND2x1_ASAP7_75t_R _27097_ (.A(_02017_),
    .B(_07406_),
    .Y(_07445_));
 OA21x2_ASAP7_75t_R _27098_ (.A1(_06627_),
    .A2(_07408_),
    .B(_07445_),
    .Y(_02563_));
 OR3x1_ASAP7_75t_R _27099_ (.A(_05059_),
    .B(_05765_),
    .C(_05937_),
    .Y(_07446_));
 BUFx6f_ASAP7_75t_R _27100_ (.A(_07446_),
    .Y(_07447_));
 BUFx4f_ASAP7_75t_R _27101_ (.A(_07447_),
    .Y(_07448_));
 BUFx6f_ASAP7_75t_R _27102_ (.A(_07447_),
    .Y(_07449_));
 NAND2x1_ASAP7_75t_R _27103_ (.A(_02016_),
    .B(_07449_),
    .Y(_07450_));
 OA21x2_ASAP7_75t_R _27104_ (.A1(_05841_),
    .A2(_07448_),
    .B(_07450_),
    .Y(_02564_));
 NAND2x1_ASAP7_75t_R _27105_ (.A(_02015_),
    .B(_07449_),
    .Y(_07451_));
 OA21x2_ASAP7_75t_R _27106_ (.A1(_06635_),
    .A2(_07448_),
    .B(_07451_),
    .Y(_02565_));
 NAND2x1_ASAP7_75t_R _27107_ (.A(_02014_),
    .B(_07449_),
    .Y(_07452_));
 OA21x2_ASAP7_75t_R _27108_ (.A1(_06639_),
    .A2(_07448_),
    .B(_07452_),
    .Y(_02566_));
 NAND2x1_ASAP7_75t_R _27109_ (.A(_02013_),
    .B(_07449_),
    .Y(_07453_));
 OA21x2_ASAP7_75t_R _27110_ (.A1(_06883_),
    .A2(_07448_),
    .B(_07453_),
    .Y(_02567_));
 NAND2x1_ASAP7_75t_R _27111_ (.A(_02012_),
    .B(_07449_),
    .Y(_07454_));
 OA21x2_ASAP7_75t_R _27112_ (.A1(_06650_),
    .A2(_07448_),
    .B(_07454_),
    .Y(_02568_));
 NAND2x1_ASAP7_75t_R _27113_ (.A(_02011_),
    .B(_07449_),
    .Y(_07455_));
 OA21x2_ASAP7_75t_R _27114_ (.A1(_06065_),
    .A2(_07448_),
    .B(_07455_),
    .Y(_02569_));
 NAND2x1_ASAP7_75t_R _27115_ (.A(_02010_),
    .B(_07449_),
    .Y(_07456_));
 OA21x2_ASAP7_75t_R _27116_ (.A1(_06660_),
    .A2(_07448_),
    .B(_07456_),
    .Y(_02570_));
 NAND2x1_ASAP7_75t_R _27117_ (.A(_02009_),
    .B(_07449_),
    .Y(_07457_));
 OA21x2_ASAP7_75t_R _27118_ (.A1(_06111_),
    .A2(_07448_),
    .B(_07457_),
    .Y(_02571_));
 BUFx6f_ASAP7_75t_R _27119_ (.A(_07447_),
    .Y(_07458_));
 NAND2x1_ASAP7_75t_R _27120_ (.A(_02008_),
    .B(_07458_),
    .Y(_07459_));
 OA21x2_ASAP7_75t_R _27121_ (.A1(_06137_),
    .A2(_07448_),
    .B(_07459_),
    .Y(_02572_));
 NAND2x1_ASAP7_75t_R _27122_ (.A(_02007_),
    .B(_07458_),
    .Y(_07460_));
 OA21x2_ASAP7_75t_R _27123_ (.A1(_06161_),
    .A2(_07448_),
    .B(_07460_),
    .Y(_02573_));
 BUFx4f_ASAP7_75t_R _27124_ (.A(_07447_),
    .Y(_07461_));
 NAND2x1_ASAP7_75t_R _27125_ (.A(_02006_),
    .B(_07458_),
    .Y(_07462_));
 OA21x2_ASAP7_75t_R _27126_ (.A1(_06180_),
    .A2(_07461_),
    .B(_07462_),
    .Y(_02574_));
 NAND2x1_ASAP7_75t_R _27127_ (.A(_02005_),
    .B(_07458_),
    .Y(_07463_));
 OA21x2_ASAP7_75t_R _27128_ (.A1(_06475_),
    .A2(_07461_),
    .B(_07463_),
    .Y(_02575_));
 NAND2x1_ASAP7_75t_R _27129_ (.A(_02004_),
    .B(_07458_),
    .Y(_07464_));
 OA21x2_ASAP7_75t_R _27130_ (.A1(_06218_),
    .A2(_07461_),
    .B(_07464_),
    .Y(_02576_));
 NAND2x1_ASAP7_75t_R _27131_ (.A(_02003_),
    .B(_07458_),
    .Y(_07465_));
 OA21x2_ASAP7_75t_R _27132_ (.A1(_06695_),
    .A2(_07461_),
    .B(_07465_),
    .Y(_02577_));
 NAND2x1_ASAP7_75t_R _27133_ (.A(_02002_),
    .B(_07458_),
    .Y(_07466_));
 OA21x2_ASAP7_75t_R _27134_ (.A1(_06260_),
    .A2(_07461_),
    .B(_07466_),
    .Y(_02578_));
 NAND2x1_ASAP7_75t_R _27135_ (.A(_02001_),
    .B(_07458_),
    .Y(_07467_));
 OA21x2_ASAP7_75t_R _27136_ (.A1(_06705_),
    .A2(_07461_),
    .B(_07467_),
    .Y(_02579_));
 NAND2x1_ASAP7_75t_R _27137_ (.A(_02000_),
    .B(_07458_),
    .Y(_07468_));
 OA21x2_ASAP7_75t_R _27138_ (.A1(_06299_),
    .A2(_07461_),
    .B(_07468_),
    .Y(_02580_));
 NAND2x1_ASAP7_75t_R _27139_ (.A(_01999_),
    .B(_07458_),
    .Y(_07469_));
 OA21x2_ASAP7_75t_R _27140_ (.A1(_06320_),
    .A2(_07461_),
    .B(_07469_),
    .Y(_02581_));
 BUFx6f_ASAP7_75t_R _27141_ (.A(_07447_),
    .Y(_07470_));
 NAND2x1_ASAP7_75t_R _27142_ (.A(_01998_),
    .B(_07470_),
    .Y(_07471_));
 OA21x2_ASAP7_75t_R _27143_ (.A1(_06968_),
    .A2(_07461_),
    .B(_07471_),
    .Y(_02582_));
 NAND2x1_ASAP7_75t_R _27144_ (.A(_01997_),
    .B(_07470_),
    .Y(_07472_));
 OA21x2_ASAP7_75t_R _27145_ (.A1(_07431_),
    .A2(_07461_),
    .B(_07472_),
    .Y(_02583_));
 BUFx4f_ASAP7_75t_R _27146_ (.A(_07447_),
    .Y(_07473_));
 NAND2x1_ASAP7_75t_R _27147_ (.A(_01996_),
    .B(_07470_),
    .Y(_07474_));
 OA21x2_ASAP7_75t_R _27148_ (.A1(_06738_),
    .A2(_07473_),
    .B(_07474_),
    .Y(_02584_));
 NAND2x1_ASAP7_75t_R _27149_ (.A(_01995_),
    .B(_07470_),
    .Y(_07475_));
 OA21x2_ASAP7_75t_R _27150_ (.A1(_06411_),
    .A2(_07473_),
    .B(_07475_),
    .Y(_02585_));
 NAND2x1_ASAP7_75t_R _27151_ (.A(_01994_),
    .B(_07470_),
    .Y(_07476_));
 OA21x2_ASAP7_75t_R _27152_ (.A1(_05872_),
    .A2(_07473_),
    .B(_07476_),
    .Y(_02586_));
 NAND2x1_ASAP7_75t_R _27153_ (.A(_01993_),
    .B(_07470_),
    .Y(_07477_));
 OA21x2_ASAP7_75t_R _27154_ (.A1(_06750_),
    .A2(_07473_),
    .B(_07477_),
    .Y(_02587_));
 NAND2x1_ASAP7_75t_R _27155_ (.A(_01992_),
    .B(_07470_),
    .Y(_07478_));
 OA21x2_ASAP7_75t_R _27156_ (.A1(_07369_),
    .A2(_07473_),
    .B(_07478_),
    .Y(_02588_));
 NAND2x1_ASAP7_75t_R _27157_ (.A(_01991_),
    .B(_07470_),
    .Y(_07479_));
 OA21x2_ASAP7_75t_R _27158_ (.A1(_06588_),
    .A2(_07473_),
    .B(_07479_),
    .Y(_02589_));
 NAND2x1_ASAP7_75t_R _27159_ (.A(_01990_),
    .B(_07470_),
    .Y(_07480_));
 OA21x2_ASAP7_75t_R _27160_ (.A1(_07042_),
    .A2(_07473_),
    .B(_07480_),
    .Y(_02590_));
 NAND2x1_ASAP7_75t_R _27161_ (.A(_01989_),
    .B(_07470_),
    .Y(_07481_));
 OA21x2_ASAP7_75t_R _27162_ (.A1(_06534_),
    .A2(_07473_),
    .B(_07481_),
    .Y(_02591_));
 NAND2x1_ASAP7_75t_R _27163_ (.A(_01988_),
    .B(_07447_),
    .Y(_07482_));
 OA21x2_ASAP7_75t_R _27164_ (.A1(_06559_),
    .A2(_07473_),
    .B(_07482_),
    .Y(_02592_));
 NAND2x1_ASAP7_75t_R _27165_ (.A(_01987_),
    .B(_07447_),
    .Y(_07483_));
 OA21x2_ASAP7_75t_R _27166_ (.A1(_06584_),
    .A2(_07473_),
    .B(_07483_),
    .Y(_02593_));
 NAND2x1_ASAP7_75t_R _27167_ (.A(_01986_),
    .B(_07447_),
    .Y(_07484_));
 OA21x2_ASAP7_75t_R _27168_ (.A1(_06609_),
    .A2(_07449_),
    .B(_07484_),
    .Y(_02594_));
 NAND2x1_ASAP7_75t_R _27169_ (.A(_01985_),
    .B(_07447_),
    .Y(_07485_));
 OA21x2_ASAP7_75t_R _27170_ (.A1(_06627_),
    .A2(_07449_),
    .B(_07485_),
    .Y(_02595_));
 OR2x4_ASAP7_75t_R _27171_ (.A(_05058_),
    .B(_05765_),
    .Y(_07486_));
 NAND3x2_ASAP7_75t_R _27172_ (.B(_07227_),
    .C(_07244_),
    .Y(_07487_),
    .A(_04945_));
 OR3x4_ASAP7_75t_R _27173_ (.A(_02220_),
    .B(_05408_),
    .C(_05409_),
    .Y(_07488_));
 AND2x6_ASAP7_75t_R _27174_ (.A(_07487_),
    .B(_07488_),
    .Y(_07489_));
 OA21x2_ASAP7_75t_R _27175_ (.A1(_07486_),
    .A2(_06189_),
    .B(_07489_),
    .Y(_07490_));
 BUFx4f_ASAP7_75t_R _27176_ (.A(_07489_),
    .Y(_07491_));
 INVx1_ASAP7_75t_R _27177_ (.A(_05328_),
    .Y(_07492_));
 AO221x2_ASAP7_75t_R _27178_ (.A1(_01778_),
    .A2(_02221_),
    .B1(_05449_),
    .B2(_13407_),
    .C(_07492_),
    .Y(_07493_));
 AND3x1_ASAP7_75t_R _27179_ (.A(_05329_),
    .B(_05454_),
    .C(_07493_),
    .Y(_07494_));
 INVx1_ASAP7_75t_R _27180_ (.A(_07494_),
    .Y(_07495_));
 AO21x1_ASAP7_75t_R _27181_ (.A1(_05455_),
    .A2(_07495_),
    .B(_05407_),
    .Y(_07496_));
 AND3x1_ASAP7_75t_R _27182_ (.A(_04945_),
    .B(_07227_),
    .C(_07244_),
    .Y(_07497_));
 BUFx6f_ASAP7_75t_R _27183_ (.A(_07497_),
    .Y(_07498_));
 BUFx6f_ASAP7_75t_R _27184_ (.A(_07498_),
    .Y(_07499_));
 BUFx6f_ASAP7_75t_R _27185_ (.A(_07488_),
    .Y(_07500_));
 NOR2x1_ASAP7_75t_R _27186_ (.A(_01896_),
    .B(_07500_),
    .Y(_07501_));
 AO221x1_ASAP7_75t_R _27187_ (.A1(_05840_),
    .A2(_07491_),
    .B1(_07496_),
    .B2(_07499_),
    .C(_07501_),
    .Y(_07502_));
 NAND2x1_ASAP7_75t_R _27188_ (.A(_01984_),
    .B(_07490_),
    .Y(_07503_));
 OA21x2_ASAP7_75t_R _27189_ (.A1(_07490_),
    .A2(_07502_),
    .B(_07503_),
    .Y(_02596_));
 OAI21x1_ASAP7_75t_R _27190_ (.A1(_07486_),
    .A2(_06189_),
    .B(_07489_),
    .Y(_07504_));
 AND2x2_ASAP7_75t_R _27191_ (.A(_06198_),
    .B(_07491_),
    .Y(_07505_));
 OR2x2_ASAP7_75t_R _27192_ (.A(_05438_),
    .B(_05448_),
    .Y(_07506_));
 NOR2x2_ASAP7_75t_R _27193_ (.A(_02220_),
    .B(_05413_),
    .Y(_07507_));
 AO32x1_ASAP7_75t_R _27194_ (.A1(_05457_),
    .A2(_07506_),
    .A3(_07498_),
    .B1(_07507_),
    .B2(_01895_),
    .Y(_07508_));
 OR3x1_ASAP7_75t_R _27195_ (.A(_07490_),
    .B(_07505_),
    .C(_07508_),
    .Y(_07509_));
 OAI21x1_ASAP7_75t_R _27196_ (.A1(_01983_),
    .A2(_07504_),
    .B(_07509_),
    .Y(_02597_));
 AND2x2_ASAP7_75t_R _27197_ (.A(_05871_),
    .B(_07491_),
    .Y(_07510_));
 OR3x1_ASAP7_75t_R _27198_ (.A(_05355_),
    .B(_05367_),
    .C(_05370_),
    .Y(_07511_));
 NOR2x1_ASAP7_75t_R _27199_ (.A(_05345_),
    .B(_05348_),
    .Y(_07512_));
 OR2x2_ASAP7_75t_R _27200_ (.A(_05363_),
    .B(_05366_),
    .Y(_07513_));
 OA211x2_ASAP7_75t_R _27201_ (.A1(_07512_),
    .A2(_07513_),
    .B(_05446_),
    .C(_05439_),
    .Y(_07514_));
 AO21x1_ASAP7_75t_R _27202_ (.A1(_07511_),
    .A2(_07514_),
    .B(_05438_),
    .Y(_07515_));
 OR2x2_ASAP7_75t_R _27203_ (.A(_05456_),
    .B(_07493_),
    .Y(_07516_));
 AO32x1_ASAP7_75t_R _27204_ (.A1(_07498_),
    .A2(_07515_),
    .A3(_07516_),
    .B1(_07507_),
    .B2(_01894_),
    .Y(_07517_));
 OR3x1_ASAP7_75t_R _27205_ (.A(_07490_),
    .B(_07510_),
    .C(_07517_),
    .Y(_07518_));
 OAI21x1_ASAP7_75t_R _27206_ (.A1(_01982_),
    .A2(_07504_),
    .B(_07518_),
    .Y(_02598_));
 INVx1_ASAP7_75t_R _27207_ (.A(_01981_),
    .Y(_07519_));
 NAND2x2_ASAP7_75t_R _27208_ (.A(_07487_),
    .B(_07488_),
    .Y(_07520_));
 INVx1_ASAP7_75t_R _27209_ (.A(_01893_),
    .Y(_07521_));
 NOR2x1_ASAP7_75t_R _27210_ (.A(_05360_),
    .B(_07513_),
    .Y(_07522_));
 OR3x1_ASAP7_75t_R _27211_ (.A(_05369_),
    .B(_01940_),
    .C(_05355_),
    .Y(_07523_));
 AND3x1_ASAP7_75t_R _27212_ (.A(_07522_),
    .B(_05446_),
    .C(_07523_),
    .Y(_07524_));
 NOR2x1_ASAP7_75t_R _27213_ (.A(_05438_),
    .B(_07524_),
    .Y(_07525_));
 INVx1_ASAP7_75t_R _27214_ (.A(_05453_),
    .Y(_07526_));
 AND3x1_ASAP7_75t_R _27215_ (.A(_15510_),
    .B(_07526_),
    .C(_05455_),
    .Y(_07527_));
 OA33x2_ASAP7_75t_R _27216_ (.A1(_02220_),
    .A2(_07521_),
    .A3(_07230_),
    .B1(_07487_),
    .B2(_07525_),
    .B3(_07527_),
    .Y(_07528_));
 OA211x2_ASAP7_75t_R _27217_ (.A1(_06588_),
    .A2(_07520_),
    .B(_07504_),
    .C(_07528_),
    .Y(_07529_));
 AO21x1_ASAP7_75t_R _27218_ (.A1(_07519_),
    .A2(_07490_),
    .B(_07529_),
    .Y(_02599_));
 AND2x2_ASAP7_75t_R _27219_ (.A(_06517_),
    .B(_07489_),
    .Y(_07530_));
 AO21x1_ASAP7_75t_R _27220_ (.A1(_05405_),
    .A2(_05445_),
    .B(_05438_),
    .Y(_07531_));
 AO22x1_ASAP7_75t_R _27221_ (.A1(_01892_),
    .A2(_07507_),
    .B1(_07531_),
    .B2(_07499_),
    .Y(_07532_));
 OR3x1_ASAP7_75t_R _27222_ (.A(_07490_),
    .B(_07530_),
    .C(_07532_),
    .Y(_07533_));
 OAI21x1_ASAP7_75t_R _27223_ (.A1(_01980_),
    .A2(_07504_),
    .B(_07533_),
    .Y(_02600_));
 BUFx4f_ASAP7_75t_R _27224_ (.A(_07520_),
    .Y(_07534_));
 BUFx4f_ASAP7_75t_R _27225_ (.A(_07488_),
    .Y(_07535_));
 OA21x2_ASAP7_75t_R _27226_ (.A1(_01891_),
    .A2(_07535_),
    .B(_05438_),
    .Y(_07536_));
 OA211x2_ASAP7_75t_R _27227_ (.A1(_06455_),
    .A2(_07534_),
    .B(_07504_),
    .C(_07536_),
    .Y(_07537_));
 AOI21x1_ASAP7_75t_R _27228_ (.A1(_01979_),
    .A2(_07490_),
    .B(_07537_),
    .Y(_02601_));
 BUFx6f_ASAP7_75t_R _27229_ (.A(_07488_),
    .Y(_07538_));
 OAI21x1_ASAP7_75t_R _27230_ (.A1(_07486_),
    .A2(_05951_),
    .B(_07489_),
    .Y(_07539_));
 BUFx4f_ASAP7_75t_R _27231_ (.A(_07539_),
    .Y(_07540_));
 OAI22x1_ASAP7_75t_R _27232_ (.A1(_01887_),
    .A2(_07538_),
    .B1(_07540_),
    .B2(_01978_),
    .Y(_02602_));
 OA21x2_ASAP7_75t_R _27233_ (.A1(_07486_),
    .A2(_05951_),
    .B(_07489_),
    .Y(_07541_));
 BUFx6f_ASAP7_75t_R _27234_ (.A(_07541_),
    .Y(_07542_));
 BUFx4f_ASAP7_75t_R _27235_ (.A(_07542_),
    .Y(_07543_));
 BUFx3_ASAP7_75t_R _27236_ (.A(_07489_),
    .Y(_07544_));
 BUFx6f_ASAP7_75t_R _27237_ (.A(_07487_),
    .Y(_07545_));
 BUFx6f_ASAP7_75t_R _27238_ (.A(_07545_),
    .Y(_07546_));
 OAI22x1_ASAP7_75t_R _27239_ (.A1(_07260_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01886_),
    .Y(_07547_));
 AO21x1_ASAP7_75t_R _27240_ (.A1(_06635_),
    .A2(_07544_),
    .B(_07547_),
    .Y(_07548_));
 BUFx4f_ASAP7_75t_R _27241_ (.A(_07541_),
    .Y(_07549_));
 NAND2x1_ASAP7_75t_R _27242_ (.A(_01977_),
    .B(_07549_),
    .Y(_07550_));
 OA21x2_ASAP7_75t_R _27243_ (.A1(_07543_),
    .A2(_07548_),
    .B(_07550_),
    .Y(_02603_));
 BUFx6f_ASAP7_75t_R _27244_ (.A(_07542_),
    .Y(_07551_));
 BUFx10_ASAP7_75t_R _27245_ (.A(_07487_),
    .Y(_07552_));
 OA22x2_ASAP7_75t_R _27246_ (.A1(_07265_),
    .A2(_07552_),
    .B1(_07535_),
    .B2(_01885_),
    .Y(_07553_));
 OA211x2_ASAP7_75t_R _27247_ (.A1(_06000_),
    .A2(_07534_),
    .B(_07540_),
    .C(_07553_),
    .Y(_07554_));
 AOI21x1_ASAP7_75t_R _27248_ (.A1(_01976_),
    .A2(_07551_),
    .B(_07554_),
    .Y(_02604_));
 OA22x2_ASAP7_75t_R _27249_ (.A1(_07269_),
    .A2(_07552_),
    .B1(_07535_),
    .B2(_01884_),
    .Y(_07555_));
 OA211x2_ASAP7_75t_R _27250_ (.A1(_06017_),
    .A2(_07534_),
    .B(_07540_),
    .C(_07555_),
    .Y(_07556_));
 AOI21x1_ASAP7_75t_R _27251_ (.A1(_01975_),
    .A2(_07551_),
    .B(_07556_),
    .Y(_02605_));
 OAI22x1_ASAP7_75t_R _27252_ (.A1(_07273_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01883_),
    .Y(_07557_));
 AO21x1_ASAP7_75t_R _27253_ (.A1(_06650_),
    .A2(_07544_),
    .B(_07557_),
    .Y(_07558_));
 NAND2x1_ASAP7_75t_R _27254_ (.A(_01974_),
    .B(_07549_),
    .Y(_07559_));
 OA21x2_ASAP7_75t_R _27255_ (.A1(_07543_),
    .A2(_07558_),
    .B(_07559_),
    .Y(_02606_));
 OA22x2_ASAP7_75t_R _27256_ (.A1(_07278_),
    .A2(_07545_),
    .B1(_07535_),
    .B2(_01882_),
    .Y(_07560_));
 OA211x2_ASAP7_75t_R _27257_ (.A1(_06656_),
    .A2(_07534_),
    .B(_07540_),
    .C(_07560_),
    .Y(_07561_));
 AOI21x1_ASAP7_75t_R _27258_ (.A1(_01973_),
    .A2(_07551_),
    .B(_07561_),
    .Y(_02607_));
 OAI22x1_ASAP7_75t_R _27259_ (.A1(_07283_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01881_),
    .Y(_07562_));
 AO21x1_ASAP7_75t_R _27260_ (.A1(_06660_),
    .A2(_07544_),
    .B(_07562_),
    .Y(_07563_));
 BUFx6f_ASAP7_75t_R _27261_ (.A(_07541_),
    .Y(_07564_));
 NAND2x1_ASAP7_75t_R _27262_ (.A(_01972_),
    .B(_07564_),
    .Y(_07565_));
 OA21x2_ASAP7_75t_R _27263_ (.A1(_07543_),
    .A2(_07563_),
    .B(_07565_),
    .Y(_02608_));
 OA22x2_ASAP7_75t_R _27264_ (.A1(_07288_),
    .A2(_07545_),
    .B1(_07535_),
    .B2(_01880_),
    .Y(_07566_));
 OA211x2_ASAP7_75t_R _27265_ (.A1(_06112_),
    .A2(_07534_),
    .B(_07540_),
    .C(_07566_),
    .Y(_07567_));
 AOI21x1_ASAP7_75t_R _27266_ (.A1(_01971_),
    .A2(_07551_),
    .B(_07567_),
    .Y(_02609_));
 OAI22x1_ASAP7_75t_R _27267_ (.A1(_07295_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01879_),
    .Y(_07568_));
 AO21x1_ASAP7_75t_R _27268_ (.A1(_06137_),
    .A2(_07544_),
    .B(_07568_),
    .Y(_07569_));
 NAND2x1_ASAP7_75t_R _27269_ (.A(_01970_),
    .B(_07564_),
    .Y(_07570_));
 OA21x2_ASAP7_75t_R _27270_ (.A1(_07543_),
    .A2(_07569_),
    .B(_07570_),
    .Y(_02610_));
 OAI22x1_ASAP7_75t_R _27271_ (.A1(_07299_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01878_),
    .Y(_07571_));
 AO21x1_ASAP7_75t_R _27272_ (.A1(_06161_),
    .A2(_07544_),
    .B(_07571_),
    .Y(_07572_));
 NAND2x1_ASAP7_75t_R _27273_ (.A(_01969_),
    .B(_07564_),
    .Y(_07573_));
 OA21x2_ASAP7_75t_R _27274_ (.A1(_07543_),
    .A2(_07572_),
    .B(_07573_),
    .Y(_02611_));
 OAI22x1_ASAP7_75t_R _27275_ (.A1(_07304_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01877_),
    .Y(_07574_));
 AO21x1_ASAP7_75t_R _27276_ (.A1(_06180_),
    .A2(_07544_),
    .B(_07574_),
    .Y(_07575_));
 NAND2x1_ASAP7_75t_R _27277_ (.A(_01968_),
    .B(_07564_),
    .Y(_07576_));
 OA21x2_ASAP7_75t_R _27278_ (.A1(_07543_),
    .A2(_07575_),
    .B(_07576_),
    .Y(_02612_));
 AO22x1_ASAP7_75t_R _27279_ (.A1(_07316_),
    .A2(_07498_),
    .B1(_07507_),
    .B2(_01876_),
    .Y(_07577_));
 OR3x1_ASAP7_75t_R _27280_ (.A(_07505_),
    .B(_07542_),
    .C(_07577_),
    .Y(_07578_));
 OAI21x1_ASAP7_75t_R _27281_ (.A1(_01967_),
    .A2(_07540_),
    .B(_07578_),
    .Y(_02613_));
 OAI22x1_ASAP7_75t_R _27282_ (.A1(_07320_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01875_),
    .Y(_07579_));
 AO21x1_ASAP7_75t_R _27283_ (.A1(_06218_),
    .A2(_07544_),
    .B(_07579_),
    .Y(_07580_));
 NAND2x1_ASAP7_75t_R _27284_ (.A(_01966_),
    .B(_07564_),
    .Y(_07581_));
 OA21x2_ASAP7_75t_R _27285_ (.A1(_07543_),
    .A2(_07580_),
    .B(_07581_),
    .Y(_02614_));
 NOR2x1_ASAP7_75t_R _27286_ (.A(_01874_),
    .B(_07500_),
    .Y(_07582_));
 AO221x1_ASAP7_75t_R _27287_ (.A1(_07326_),
    .A2(_07499_),
    .B1(_07491_),
    .B2(_06241_),
    .C(_07582_),
    .Y(_07583_));
 NAND2x1_ASAP7_75t_R _27288_ (.A(_01965_),
    .B(_07564_),
    .Y(_07584_));
 OA21x2_ASAP7_75t_R _27289_ (.A1(_07543_),
    .A2(_07583_),
    .B(_07584_),
    .Y(_02615_));
 INVx1_ASAP7_75t_R _27290_ (.A(_06259_),
    .Y(_07585_));
 OA22x2_ASAP7_75t_R _27291_ (.A1(_07330_),
    .A2(_07545_),
    .B1(_07535_),
    .B2(_01873_),
    .Y(_07586_));
 OA211x2_ASAP7_75t_R _27292_ (.A1(_07585_),
    .A2(_07534_),
    .B(_07540_),
    .C(_07586_),
    .Y(_07587_));
 AOI21x1_ASAP7_75t_R _27293_ (.A1(_01964_),
    .A2(_07551_),
    .B(_07587_),
    .Y(_02616_));
 OAI22x1_ASAP7_75t_R _27294_ (.A1(_07335_),
    .A2(_07546_),
    .B1(_07538_),
    .B2(_01872_),
    .Y(_07588_));
 AO21x1_ASAP7_75t_R _27295_ (.A1(_06705_),
    .A2(_07544_),
    .B(_07588_),
    .Y(_07589_));
 NAND2x1_ASAP7_75t_R _27296_ (.A(_01963_),
    .B(_07564_),
    .Y(_07590_));
 OA21x2_ASAP7_75t_R _27297_ (.A1(_07543_),
    .A2(_07589_),
    .B(_07590_),
    .Y(_02617_));
 OAI22x1_ASAP7_75t_R _27298_ (.A1(_07339_),
    .A2(_07552_),
    .B1(_07500_),
    .B2(_01871_),
    .Y(_07591_));
 AO21x1_ASAP7_75t_R _27299_ (.A1(_06299_),
    .A2(_07544_),
    .B(_07591_),
    .Y(_07592_));
 NAND2x1_ASAP7_75t_R _27300_ (.A(_01962_),
    .B(_07564_),
    .Y(_07593_));
 OA21x2_ASAP7_75t_R _27301_ (.A1(_07543_),
    .A2(_07592_),
    .B(_07593_),
    .Y(_02618_));
 INVx1_ASAP7_75t_R _27302_ (.A(_06319_),
    .Y(_07594_));
 OA22x2_ASAP7_75t_R _27303_ (.A1(_07344_),
    .A2(_07545_),
    .B1(_07535_),
    .B2(_01870_),
    .Y(_07595_));
 OA211x2_ASAP7_75t_R _27304_ (.A1(_07594_),
    .A2(_07534_),
    .B(_07540_),
    .C(_07595_),
    .Y(_07596_));
 AOI21x1_ASAP7_75t_R _27305_ (.A1(_01961_),
    .A2(_07551_),
    .B(_07596_),
    .Y(_02619_));
 OA22x2_ASAP7_75t_R _27306_ (.A1(_07347_),
    .A2(_07545_),
    .B1(_07535_),
    .B2(_01869_),
    .Y(_07597_));
 OA211x2_ASAP7_75t_R _27307_ (.A1(_06347_),
    .A2(_07534_),
    .B(_07539_),
    .C(_07597_),
    .Y(_07598_));
 AOI21x1_ASAP7_75t_R _27308_ (.A1(_01960_),
    .A2(_07551_),
    .B(_07598_),
    .Y(_02620_));
 OA22x2_ASAP7_75t_R _27309_ (.A1(_07350_),
    .A2(_07545_),
    .B1(_07535_),
    .B2(_01868_),
    .Y(_07599_));
 OA211x2_ASAP7_75t_R _27310_ (.A1(_06370_),
    .A2(_07534_),
    .B(_07539_),
    .C(_07599_),
    .Y(_07600_));
 AOI21x1_ASAP7_75t_R _27311_ (.A1(_01959_),
    .A2(_07551_),
    .B(_07600_),
    .Y(_02621_));
 OAI22x1_ASAP7_75t_R _27312_ (.A1(_07354_),
    .A2(_07552_),
    .B1(_07500_),
    .B2(_01867_),
    .Y(_07601_));
 AO21x1_ASAP7_75t_R _27313_ (.A1(_06738_),
    .A2(_07544_),
    .B(_07601_),
    .Y(_07602_));
 NAND2x1_ASAP7_75t_R _27314_ (.A(_01958_),
    .B(_07564_),
    .Y(_07603_));
 OA21x2_ASAP7_75t_R _27315_ (.A1(_07549_),
    .A2(_07602_),
    .B(_07603_),
    .Y(_02622_));
 OAI22x1_ASAP7_75t_R _27316_ (.A1(_07358_),
    .A2(_07552_),
    .B1(_07500_),
    .B2(_01866_),
    .Y(_07604_));
 AO21x1_ASAP7_75t_R _27317_ (.A1(_06411_),
    .A2(_07491_),
    .B(_07604_),
    .Y(_07605_));
 NAND2x1_ASAP7_75t_R _27318_ (.A(_01957_),
    .B(_07564_),
    .Y(_07606_));
 OA21x2_ASAP7_75t_R _27319_ (.A1(_07549_),
    .A2(_07605_),
    .B(_07606_),
    .Y(_02623_));
 AO22x1_ASAP7_75t_R _27320_ (.A1(_07362_),
    .A2(_07498_),
    .B1(_07507_),
    .B2(_01865_),
    .Y(_07607_));
 OR3x1_ASAP7_75t_R _27321_ (.A(_07510_),
    .B(_07542_),
    .C(_07607_),
    .Y(_07608_));
 OAI21x1_ASAP7_75t_R _27322_ (.A1(_01956_),
    .A2(_07540_),
    .B(_07608_),
    .Y(_02624_));
 OAI22x1_ASAP7_75t_R _27323_ (.A1(_07366_),
    .A2(_07552_),
    .B1(_07500_),
    .B2(_01864_),
    .Y(_07609_));
 AO21x1_ASAP7_75t_R _27324_ (.A1(_06750_),
    .A2(_07491_),
    .B(_07609_),
    .Y(_07610_));
 NAND2x1_ASAP7_75t_R _27325_ (.A(_01955_),
    .B(_07542_),
    .Y(_07611_));
 OA21x2_ASAP7_75t_R _27326_ (.A1(_07549_),
    .A2(_07610_),
    .B(_07611_),
    .Y(_02625_));
 INVx1_ASAP7_75t_R _27327_ (.A(_01863_),
    .Y(_07612_));
 AOI22x1_ASAP7_75t_R _27328_ (.A1(_07371_),
    .A2(_07499_),
    .B1(_07507_),
    .B2(_07612_),
    .Y(_07613_));
 OA211x2_ASAP7_75t_R _27329_ (.A1(_06455_),
    .A2(_07534_),
    .B(_07539_),
    .C(_07613_),
    .Y(_07614_));
 AOI21x1_ASAP7_75t_R _27330_ (.A1(_01954_),
    .A2(_07551_),
    .B(_07614_),
    .Y(_02626_));
 INVx1_ASAP7_75t_R _27331_ (.A(_01953_),
    .Y(_07615_));
 AOI22x1_ASAP7_75t_R _27332_ (.A1(_07375_),
    .A2(_07498_),
    .B1(_07507_),
    .B2(_01862_),
    .Y(_07616_));
 OA211x2_ASAP7_75t_R _27333_ (.A1(_06500_),
    .A2(_07520_),
    .B(_07539_),
    .C(_07616_),
    .Y(_07617_));
 AO21x1_ASAP7_75t_R _27334_ (.A1(_07615_),
    .A2(_07549_),
    .B(_07617_),
    .Y(_02627_));
 AO22x1_ASAP7_75t_R _27335_ (.A1(_07380_),
    .A2(_07498_),
    .B1(_07507_),
    .B2(_01861_),
    .Y(_07618_));
 OR3x1_ASAP7_75t_R _27336_ (.A(_07530_),
    .B(_07542_),
    .C(_07618_),
    .Y(_07619_));
 OAI21x1_ASAP7_75t_R _27337_ (.A1(_01952_),
    .A2(_07540_),
    .B(_07619_),
    .Y(_02628_));
 NOR2x1_ASAP7_75t_R _27338_ (.A(_01860_),
    .B(_07500_),
    .Y(_07620_));
 AO221x1_ASAP7_75t_R _27339_ (.A1(_07385_),
    .A2(_07499_),
    .B1(_07491_),
    .B2(_06534_),
    .C(_07620_),
    .Y(_07621_));
 NAND2x1_ASAP7_75t_R _27340_ (.A(_01951_),
    .B(_07542_),
    .Y(_07622_));
 OA21x2_ASAP7_75t_R _27341_ (.A1(_07549_),
    .A2(_07621_),
    .B(_07622_),
    .Y(_02629_));
 OAI22x1_ASAP7_75t_R _27342_ (.A1(_07389_),
    .A2(_07552_),
    .B1(_07500_),
    .B2(_01859_),
    .Y(_07623_));
 AO21x1_ASAP7_75t_R _27343_ (.A1(_06559_),
    .A2(_07491_),
    .B(_07623_),
    .Y(_07624_));
 NAND2x1_ASAP7_75t_R _27344_ (.A(_01950_),
    .B(_07542_),
    .Y(_07625_));
 OA21x2_ASAP7_75t_R _27345_ (.A1(_07549_),
    .A2(_07624_),
    .B(_07625_),
    .Y(_02630_));
 OAI22x1_ASAP7_75t_R _27346_ (.A1(_07394_),
    .A2(_07552_),
    .B1(_07500_),
    .B2(_01858_),
    .Y(_07626_));
 AO21x1_ASAP7_75t_R _27347_ (.A1(_06584_),
    .A2(_07491_),
    .B(_07626_),
    .Y(_07627_));
 NAND2x1_ASAP7_75t_R _27348_ (.A(_01949_),
    .B(_07542_),
    .Y(_07628_));
 OA21x2_ASAP7_75t_R _27349_ (.A1(_07549_),
    .A2(_07627_),
    .B(_07628_),
    .Y(_02631_));
 OA22x2_ASAP7_75t_R _27350_ (.A1(_07399_),
    .A2(_07545_),
    .B1(_07535_),
    .B2(_01857_),
    .Y(_07629_));
 OA211x2_ASAP7_75t_R _27351_ (.A1(_06610_),
    .A2(_07520_),
    .B(_07539_),
    .C(_07629_),
    .Y(_07630_));
 AOI21x1_ASAP7_75t_R _27352_ (.A1(_01948_),
    .A2(_07551_),
    .B(_07630_),
    .Y(_02632_));
 OAI22x1_ASAP7_75t_R _27353_ (.A1(_07403_),
    .A2(_07552_),
    .B1(_07500_),
    .B2(_01856_),
    .Y(_07631_));
 AO21x1_ASAP7_75t_R _27354_ (.A1(_06627_),
    .A2(_07491_),
    .B(_07631_),
    .Y(_07632_));
 NAND2x1_ASAP7_75t_R _27355_ (.A(_01947_),
    .B(_07542_),
    .Y(_07633_));
 OA21x2_ASAP7_75t_R _27356_ (.A1(_07549_),
    .A2(_07632_),
    .B(_07633_),
    .Y(_02633_));
 OR3x1_ASAP7_75t_R _27357_ (.A(_05059_),
    .B(_05765_),
    .C(_06251_),
    .Y(_07634_));
 BUFx6f_ASAP7_75t_R _27358_ (.A(_07634_),
    .Y(_07635_));
 BUFx4f_ASAP7_75t_R _27359_ (.A(_07635_),
    .Y(_07636_));
 BUFx4f_ASAP7_75t_R _27360_ (.A(_07635_),
    .Y(_07637_));
 NAND2x1_ASAP7_75t_R _27361_ (.A(_01946_),
    .B(_07637_),
    .Y(_07638_));
 OA21x2_ASAP7_75t_R _27362_ (.A1(_06111_),
    .A2(_07636_),
    .B(_07638_),
    .Y(_02634_));
 NAND2x1_ASAP7_75t_R _27363_ (.A(_01945_),
    .B(_07637_),
    .Y(_07639_));
 OA21x2_ASAP7_75t_R _27364_ (.A1(_06968_),
    .A2(_07636_),
    .B(_07639_),
    .Y(_02635_));
 BUFx6f_ASAP7_75t_R _27365_ (.A(_07635_),
    .Y(_07640_));
 NAND2x1_ASAP7_75t_R _27366_ (.A(_01944_),
    .B(_07640_),
    .Y(_07641_));
 OA21x2_ASAP7_75t_R _27367_ (.A1(_07431_),
    .A2(_07636_),
    .B(_07641_),
    .Y(_02636_));
 NAND2x1_ASAP7_75t_R _27368_ (.A(_01943_),
    .B(_07640_),
    .Y(_07642_));
 OA21x2_ASAP7_75t_R _27369_ (.A1(_06738_),
    .A2(_07636_),
    .B(_07642_),
    .Y(_02637_));
 NAND2x1_ASAP7_75t_R _27370_ (.A(_01942_),
    .B(_07640_),
    .Y(_07643_));
 OA21x2_ASAP7_75t_R _27371_ (.A1(_06411_),
    .A2(_07636_),
    .B(_07643_),
    .Y(_02638_));
 NAND2x1_ASAP7_75t_R _27372_ (.A(_01941_),
    .B(_07640_),
    .Y(_07644_));
 OA21x2_ASAP7_75t_R _27373_ (.A1(_06750_),
    .A2(_07636_),
    .B(_07644_),
    .Y(_02639_));
 NAND2x1_ASAP7_75t_R _27374_ (.A(_01940_),
    .B(_07640_),
    .Y(_07645_));
 OA21x2_ASAP7_75t_R _27375_ (.A1(_06639_),
    .A2(_07636_),
    .B(_07645_),
    .Y(_02640_));
 NAND2x1_ASAP7_75t_R _27376_ (.A(_01939_),
    .B(_07640_),
    .Y(_07646_));
 OA21x2_ASAP7_75t_R _27377_ (.A1(_06584_),
    .A2(_07636_),
    .B(_07646_),
    .Y(_02641_));
 NAND2x1_ASAP7_75t_R _27378_ (.A(_01938_),
    .B(_07640_),
    .Y(_07647_));
 OA21x2_ASAP7_75t_R _27379_ (.A1(_06588_),
    .A2(_07636_),
    .B(_07647_),
    .Y(_02642_));
 NAND2x1_ASAP7_75t_R _27380_ (.A(_01937_),
    .B(_07640_),
    .Y(_07648_));
 OA21x2_ASAP7_75t_R _27381_ (.A1(_06137_),
    .A2(_07636_),
    .B(_07648_),
    .Y(_02643_));
 NAND2x1_ASAP7_75t_R _27382_ (.A(_01936_),
    .B(_07640_),
    .Y(_07649_));
 OA21x2_ASAP7_75t_R _27383_ (.A1(_06161_),
    .A2(_07637_),
    .B(_07649_),
    .Y(_02644_));
 NAND2x1_ASAP7_75t_R _27384_ (.A(_01935_),
    .B(_07640_),
    .Y(_07650_));
 OA21x2_ASAP7_75t_R _27385_ (.A1(_06180_),
    .A2(_07637_),
    .B(_07650_),
    .Y(_02645_));
 NAND2x1_ASAP7_75t_R _27386_ (.A(_01934_),
    .B(_07635_),
    .Y(_07651_));
 OA21x2_ASAP7_75t_R _27387_ (.A1(_06218_),
    .A2(_07637_),
    .B(_07651_),
    .Y(_02646_));
 NAND2x1_ASAP7_75t_R _27388_ (.A(_01933_),
    .B(_07635_),
    .Y(_07652_));
 OA21x2_ASAP7_75t_R _27389_ (.A1(_06695_),
    .A2(_07637_),
    .B(_07652_),
    .Y(_02647_));
 NAND2x1_ASAP7_75t_R _27390_ (.A(_01932_),
    .B(_07635_),
    .Y(_07653_));
 OA21x2_ASAP7_75t_R _27391_ (.A1(_06260_),
    .A2(_07637_),
    .B(_07653_),
    .Y(_02648_));
 NAND2x1_ASAP7_75t_R _27392_ (.A(_01931_),
    .B(_07635_),
    .Y(_07654_));
 OA21x2_ASAP7_75t_R _27393_ (.A1(_06705_),
    .A2(_07637_),
    .B(_07654_),
    .Y(_02649_));
 NAND2x1_ASAP7_75t_R _27394_ (.A(_01930_),
    .B(_07635_),
    .Y(_07655_));
 OA21x2_ASAP7_75t_R _27395_ (.A1(_06299_),
    .A2(_07637_),
    .B(_07655_),
    .Y(_02650_));
 NAND2x1_ASAP7_75t_R _27396_ (.A(_01929_),
    .B(_07635_),
    .Y(_07656_));
 OA21x2_ASAP7_75t_R _27397_ (.A1(_06320_),
    .A2(_07637_),
    .B(_07656_),
    .Y(_02651_));
 OR3x1_ASAP7_75t_R _27398_ (.A(_05059_),
    .B(_05765_),
    .C(_05815_),
    .Y(_07657_));
 BUFx6f_ASAP7_75t_R _27399_ (.A(_07657_),
    .Y(_07658_));
 BUFx4f_ASAP7_75t_R _27400_ (.A(_07658_),
    .Y(_07659_));
 BUFx6f_ASAP7_75t_R _27401_ (.A(_07658_),
    .Y(_07660_));
 NAND2x1_ASAP7_75t_R _27402_ (.A(_01928_),
    .B(_07660_),
    .Y(_07661_));
 OA21x2_ASAP7_75t_R _27403_ (.A1(_05841_),
    .A2(_07659_),
    .B(_07661_),
    .Y(_02652_));
 NAND2x1_ASAP7_75t_R _27404_ (.A(_01927_),
    .B(_07660_),
    .Y(_07662_));
 OA21x2_ASAP7_75t_R _27405_ (.A1(_06635_),
    .A2(_07659_),
    .B(_07662_),
    .Y(_02653_));
 NAND2x1_ASAP7_75t_R _27406_ (.A(_01926_),
    .B(_07660_),
    .Y(_07663_));
 OA21x2_ASAP7_75t_R _27407_ (.A1(_06639_),
    .A2(_07659_),
    .B(_07663_),
    .Y(_02654_));
 NAND2x1_ASAP7_75t_R _27408_ (.A(_01925_),
    .B(_07660_),
    .Y(_07664_));
 OA21x2_ASAP7_75t_R _27409_ (.A1(_06883_),
    .A2(_07659_),
    .B(_07664_),
    .Y(_02655_));
 NAND2x1_ASAP7_75t_R _27410_ (.A(_01924_),
    .B(_07660_),
    .Y(_07665_));
 OA21x2_ASAP7_75t_R _27411_ (.A1(_06650_),
    .A2(_07659_),
    .B(_07665_),
    .Y(_02656_));
 NAND2x1_ASAP7_75t_R _27412_ (.A(_01923_),
    .B(_07660_),
    .Y(_07666_));
 OA21x2_ASAP7_75t_R _27413_ (.A1(_06065_),
    .A2(_07659_),
    .B(_07666_),
    .Y(_02657_));
 NAND2x1_ASAP7_75t_R _27414_ (.A(_01922_),
    .B(_07660_),
    .Y(_07667_));
 OA21x2_ASAP7_75t_R _27415_ (.A1(_06660_),
    .A2(_07659_),
    .B(_07667_),
    .Y(_02658_));
 NAND2x1_ASAP7_75t_R _27416_ (.A(_01921_),
    .B(_07660_),
    .Y(_07668_));
 OA21x2_ASAP7_75t_R _27417_ (.A1(_06111_),
    .A2(_07659_),
    .B(_07668_),
    .Y(_02659_));
 BUFx6f_ASAP7_75t_R _27418_ (.A(_07658_),
    .Y(_07669_));
 NAND2x1_ASAP7_75t_R _27419_ (.A(_01920_),
    .B(_07669_),
    .Y(_07670_));
 OA21x2_ASAP7_75t_R _27420_ (.A1(_06137_),
    .A2(_07659_),
    .B(_07670_),
    .Y(_02660_));
 NAND2x1_ASAP7_75t_R _27421_ (.A(_01919_),
    .B(_07669_),
    .Y(_07671_));
 OA21x2_ASAP7_75t_R _27422_ (.A1(_06161_),
    .A2(_07659_),
    .B(_07671_),
    .Y(_02661_));
 BUFx4f_ASAP7_75t_R _27423_ (.A(_07658_),
    .Y(_07672_));
 NAND2x1_ASAP7_75t_R _27424_ (.A(_01918_),
    .B(_07669_),
    .Y(_07673_));
 OA21x2_ASAP7_75t_R _27425_ (.A1(_06180_),
    .A2(_07672_),
    .B(_07673_),
    .Y(_02662_));
 NAND2x1_ASAP7_75t_R _27426_ (.A(_01917_),
    .B(_07669_),
    .Y(_07674_));
 OA21x2_ASAP7_75t_R _27427_ (.A1(_06475_),
    .A2(_07672_),
    .B(_07674_),
    .Y(_02663_));
 NAND2x1_ASAP7_75t_R _27428_ (.A(_01916_),
    .B(_07669_),
    .Y(_07675_));
 OA21x2_ASAP7_75t_R _27429_ (.A1(_06218_),
    .A2(_07672_),
    .B(_07675_),
    .Y(_02664_));
 NAND2x1_ASAP7_75t_R _27430_ (.A(_01915_),
    .B(_07669_),
    .Y(_07676_));
 OA21x2_ASAP7_75t_R _27431_ (.A1(_06695_),
    .A2(_07672_),
    .B(_07676_),
    .Y(_02665_));
 NAND2x1_ASAP7_75t_R _27432_ (.A(_01914_),
    .B(_07669_),
    .Y(_07677_));
 OA21x2_ASAP7_75t_R _27433_ (.A1(_06260_),
    .A2(_07672_),
    .B(_07677_),
    .Y(_02666_));
 NAND2x1_ASAP7_75t_R _27434_ (.A(_01913_),
    .B(_07669_),
    .Y(_07678_));
 OA21x2_ASAP7_75t_R _27435_ (.A1(_06705_),
    .A2(_07672_),
    .B(_07678_),
    .Y(_02667_));
 NAND2x1_ASAP7_75t_R _27436_ (.A(_01912_),
    .B(_07669_),
    .Y(_07679_));
 OA21x2_ASAP7_75t_R _27437_ (.A1(_06299_),
    .A2(_07672_),
    .B(_07679_),
    .Y(_02668_));
 NAND2x1_ASAP7_75t_R _27438_ (.A(_01911_),
    .B(_07669_),
    .Y(_07680_));
 OA21x2_ASAP7_75t_R _27439_ (.A1(_06320_),
    .A2(_07672_),
    .B(_07680_),
    .Y(_02669_));
 BUFx6f_ASAP7_75t_R _27440_ (.A(_07658_),
    .Y(_07681_));
 NAND2x1_ASAP7_75t_R _27441_ (.A(_01910_),
    .B(_07681_),
    .Y(_07682_));
 OA21x2_ASAP7_75t_R _27442_ (.A1(_06968_),
    .A2(_07672_),
    .B(_07682_),
    .Y(_02670_));
 NAND2x1_ASAP7_75t_R _27443_ (.A(_01909_),
    .B(_07681_),
    .Y(_07683_));
 OA21x2_ASAP7_75t_R _27444_ (.A1(_07431_),
    .A2(_07672_),
    .B(_07683_),
    .Y(_02671_));
 BUFx4f_ASAP7_75t_R _27445_ (.A(_07658_),
    .Y(_07684_));
 NAND2x1_ASAP7_75t_R _27446_ (.A(_01908_),
    .B(_07681_),
    .Y(_07685_));
 OA21x2_ASAP7_75t_R _27447_ (.A1(_06738_),
    .A2(_07684_),
    .B(_07685_),
    .Y(_02672_));
 NAND2x1_ASAP7_75t_R _27448_ (.A(_01907_),
    .B(_07681_),
    .Y(_07686_));
 OA21x2_ASAP7_75t_R _27449_ (.A1(_06411_),
    .A2(_07684_),
    .B(_07686_),
    .Y(_02673_));
 NAND2x1_ASAP7_75t_R _27450_ (.A(_01906_),
    .B(_07681_),
    .Y(_07687_));
 OA21x2_ASAP7_75t_R _27451_ (.A1(_05872_),
    .A2(_07684_),
    .B(_07687_),
    .Y(_02674_));
 NAND2x1_ASAP7_75t_R _27452_ (.A(_01905_),
    .B(_07681_),
    .Y(_07688_));
 OA21x2_ASAP7_75t_R _27453_ (.A1(_06750_),
    .A2(_07684_),
    .B(_07688_),
    .Y(_02675_));
 NAND2x1_ASAP7_75t_R _27454_ (.A(_01904_),
    .B(_07681_),
    .Y(_07689_));
 OA21x2_ASAP7_75t_R _27455_ (.A1(_07369_),
    .A2(_07684_),
    .B(_07689_),
    .Y(_02676_));
 NAND2x1_ASAP7_75t_R _27456_ (.A(_01903_),
    .B(_07681_),
    .Y(_07690_));
 OA21x2_ASAP7_75t_R _27457_ (.A1(_06588_),
    .A2(_07684_),
    .B(_07690_),
    .Y(_02677_));
 NAND2x1_ASAP7_75t_R _27458_ (.A(_01902_),
    .B(_07681_),
    .Y(_07691_));
 OA21x2_ASAP7_75t_R _27459_ (.A1(_07042_),
    .A2(_07684_),
    .B(_07691_),
    .Y(_02678_));
 NAND2x1_ASAP7_75t_R _27460_ (.A(_01901_),
    .B(_07681_),
    .Y(_07692_));
 OA21x2_ASAP7_75t_R _27461_ (.A1(_06534_),
    .A2(_07684_),
    .B(_07692_),
    .Y(_02679_));
 NAND2x1_ASAP7_75t_R _27462_ (.A(_01900_),
    .B(_07658_),
    .Y(_07693_));
 OA21x2_ASAP7_75t_R _27463_ (.A1(_06559_),
    .A2(_07684_),
    .B(_07693_),
    .Y(_02680_));
 NAND2x1_ASAP7_75t_R _27464_ (.A(_01899_),
    .B(_07658_),
    .Y(_07694_));
 OA21x2_ASAP7_75t_R _27465_ (.A1(_06584_),
    .A2(_07684_),
    .B(_07694_),
    .Y(_02681_));
 NAND2x1_ASAP7_75t_R _27466_ (.A(_01898_),
    .B(_07658_),
    .Y(_07695_));
 OA21x2_ASAP7_75t_R _27467_ (.A1(_06609_),
    .A2(_07660_),
    .B(_07695_),
    .Y(_02682_));
 NAND2x1_ASAP7_75t_R _27468_ (.A(_01897_),
    .B(_07658_),
    .Y(_07696_));
 OA21x2_ASAP7_75t_R _27469_ (.A1(_06627_),
    .A2(_07660_),
    .B(_07696_),
    .Y(_02683_));
 BUFx6f_ASAP7_75t_R _27470_ (.A(_07546_),
    .Y(_07697_));
 BUFx4f_ASAP7_75t_R _27471_ (.A(_07552_),
    .Y(_07698_));
 NAND2x1_ASAP7_75t_R _27472_ (.A(_01896_),
    .B(_07698_),
    .Y(_07699_));
 OA21x2_ASAP7_75t_R _27473_ (.A1(_05807_),
    .A2(_07697_),
    .B(_07699_),
    .Y(_02684_));
 BUFx6f_ASAP7_75t_R _27474_ (.A(_07545_),
    .Y(_07700_));
 BUFx10_ASAP7_75t_R _27475_ (.A(_07700_),
    .Y(_07701_));
 BUFx4f_ASAP7_75t_R _27476_ (.A(_07498_),
    .Y(_07702_));
 AND2x2_ASAP7_75t_R _27477_ (.A(_01983_),
    .B(_07702_),
    .Y(_07703_));
 AOI21x1_ASAP7_75t_R _27478_ (.A1(_01895_),
    .A2(_07701_),
    .B(_07703_),
    .Y(_02685_));
 AND2x2_ASAP7_75t_R _27479_ (.A(_01982_),
    .B(_07702_),
    .Y(_07704_));
 AOI21x1_ASAP7_75t_R _27480_ (.A1(_01894_),
    .A2(_07701_),
    .B(_07704_),
    .Y(_02686_));
 NAND2x1_ASAP7_75t_R _27481_ (.A(_01981_),
    .B(_07702_),
    .Y(_07705_));
 OA21x2_ASAP7_75t_R _27482_ (.A1(_07521_),
    .A2(_07702_),
    .B(_07705_),
    .Y(_02687_));
 BUFx4f_ASAP7_75t_R _27483_ (.A(_07499_),
    .Y(_07706_));
 AND2x2_ASAP7_75t_R _27484_ (.A(_01980_),
    .B(_07706_),
    .Y(_07707_));
 AOI21x1_ASAP7_75t_R _27485_ (.A1(_01892_),
    .A2(_07701_),
    .B(_07707_),
    .Y(_02688_));
 AND2x2_ASAP7_75t_R _27486_ (.A(_01979_),
    .B(_07706_),
    .Y(_07708_));
 AOI21x1_ASAP7_75t_R _27487_ (.A1(_01891_),
    .A2(_07701_),
    .B(_07708_),
    .Y(_02689_));
 INVx1_ASAP7_75t_R _27488_ (.A(_01890_),
    .Y(_07709_));
 NAND2x1_ASAP7_75t_R _27489_ (.A(_01853_),
    .B(_07702_),
    .Y(_07710_));
 OA21x2_ASAP7_75t_R _27490_ (.A1(_07709_),
    .A2(_07702_),
    .B(_07710_),
    .Y(_02690_));
 NAND2x1_ASAP7_75t_R _27491_ (.A(_01889_),
    .B(_07698_),
    .Y(_07711_));
 OA21x2_ASAP7_75t_R _27492_ (.A1(_07234_),
    .A2(_07697_),
    .B(_07711_),
    .Y(_02691_));
 AND2x2_ASAP7_75t_R _27493_ (.A(_01851_),
    .B(_07706_),
    .Y(_07712_));
 AOI21x1_ASAP7_75t_R _27494_ (.A1(_01888_),
    .A2(_07701_),
    .B(_07712_),
    .Y(_02692_));
 AND2x2_ASAP7_75t_R _27495_ (.A(_01978_),
    .B(_07706_),
    .Y(_07713_));
 AOI21x1_ASAP7_75t_R _27496_ (.A1(_01887_),
    .A2(_07701_),
    .B(_07713_),
    .Y(_02693_));
 AND2x2_ASAP7_75t_R _27497_ (.A(_01977_),
    .B(_07706_),
    .Y(_07714_));
 AOI21x1_ASAP7_75t_R _27498_ (.A1(_01886_),
    .A2(_07701_),
    .B(_07714_),
    .Y(_02694_));
 AND2x2_ASAP7_75t_R _27499_ (.A(_01976_),
    .B(_07706_),
    .Y(_07715_));
 AOI21x1_ASAP7_75t_R _27500_ (.A1(_01885_),
    .A2(_07701_),
    .B(_07715_),
    .Y(_02695_));
 AND2x2_ASAP7_75t_R _27501_ (.A(_01975_),
    .B(_07706_),
    .Y(_07716_));
 AOI21x1_ASAP7_75t_R _27502_ (.A1(_01884_),
    .A2(_07701_),
    .B(_07716_),
    .Y(_02696_));
 AND2x2_ASAP7_75t_R _27503_ (.A(_01974_),
    .B(_07706_),
    .Y(_07717_));
 AOI21x1_ASAP7_75t_R _27504_ (.A1(_01883_),
    .A2(_07701_),
    .B(_07717_),
    .Y(_02697_));
 NAND2x1_ASAP7_75t_R _27505_ (.A(_01882_),
    .B(_07698_),
    .Y(_07718_));
 OA21x2_ASAP7_75t_R _27506_ (.A1(_06058_),
    .A2(_07697_),
    .B(_07718_),
    .Y(_02698_));
 BUFx6f_ASAP7_75t_R _27507_ (.A(_07700_),
    .Y(_07719_));
 AND2x2_ASAP7_75t_R _27508_ (.A(_01972_),
    .B(_07706_),
    .Y(_07720_));
 AOI21x1_ASAP7_75t_R _27509_ (.A1(_01881_),
    .A2(_07719_),
    .B(_07720_),
    .Y(_02699_));
 AND2x2_ASAP7_75t_R _27510_ (.A(_01971_),
    .B(_07706_),
    .Y(_07721_));
 AOI21x1_ASAP7_75t_R _27511_ (.A1(_01880_),
    .A2(_07719_),
    .B(_07721_),
    .Y(_02700_));
 BUFx3_ASAP7_75t_R _27512_ (.A(_07499_),
    .Y(_07722_));
 AND2x2_ASAP7_75t_R _27513_ (.A(_01970_),
    .B(_07722_),
    .Y(_07723_));
 AOI21x1_ASAP7_75t_R _27514_ (.A1(_01879_),
    .A2(_07719_),
    .B(_07723_),
    .Y(_02701_));
 AND2x2_ASAP7_75t_R _27515_ (.A(_01969_),
    .B(_07722_),
    .Y(_07724_));
 AOI21x1_ASAP7_75t_R _27516_ (.A1(_01878_),
    .A2(_07719_),
    .B(_07724_),
    .Y(_02702_));
 AND2x2_ASAP7_75t_R _27517_ (.A(_01968_),
    .B(_07722_),
    .Y(_07725_));
 AOI21x1_ASAP7_75t_R _27518_ (.A1(_01877_),
    .A2(_07719_),
    .B(_07725_),
    .Y(_02703_));
 AND2x2_ASAP7_75t_R _27519_ (.A(_01967_),
    .B(_07722_),
    .Y(_07726_));
 AOI21x1_ASAP7_75t_R _27520_ (.A1(_01876_),
    .A2(_07719_),
    .B(_07726_),
    .Y(_02704_));
 AND2x2_ASAP7_75t_R _27521_ (.A(_01966_),
    .B(_07722_),
    .Y(_07727_));
 AOI21x1_ASAP7_75t_R _27522_ (.A1(_01875_),
    .A2(_07719_),
    .B(_07727_),
    .Y(_02705_));
 AND2x2_ASAP7_75t_R _27523_ (.A(_01965_),
    .B(_07722_),
    .Y(_07728_));
 AOI21x1_ASAP7_75t_R _27524_ (.A1(_01874_),
    .A2(_07719_),
    .B(_07728_),
    .Y(_02706_));
 AND2x2_ASAP7_75t_R _27525_ (.A(_01964_),
    .B(_07722_),
    .Y(_07729_));
 AOI21x1_ASAP7_75t_R _27526_ (.A1(_01873_),
    .A2(_07719_),
    .B(_07729_),
    .Y(_02707_));
 AND2x2_ASAP7_75t_R _27527_ (.A(_01963_),
    .B(_07722_),
    .Y(_07730_));
 AOI21x1_ASAP7_75t_R _27528_ (.A1(_01872_),
    .A2(_07719_),
    .B(_07730_),
    .Y(_02708_));
 BUFx6f_ASAP7_75t_R _27529_ (.A(_07700_),
    .Y(_07731_));
 AND2x2_ASAP7_75t_R _27530_ (.A(_01962_),
    .B(_07722_),
    .Y(_07732_));
 AOI21x1_ASAP7_75t_R _27531_ (.A1(_01871_),
    .A2(_07731_),
    .B(_07732_),
    .Y(_02709_));
 AND2x2_ASAP7_75t_R _27532_ (.A(_01961_),
    .B(_07722_),
    .Y(_07733_));
 AOI21x1_ASAP7_75t_R _27533_ (.A1(_01870_),
    .A2(_07731_),
    .B(_07733_),
    .Y(_02710_));
 BUFx4f_ASAP7_75t_R _27534_ (.A(_07498_),
    .Y(_07734_));
 AND2x2_ASAP7_75t_R _27535_ (.A(_01960_),
    .B(_07734_),
    .Y(_07735_));
 AOI21x1_ASAP7_75t_R _27536_ (.A1(_01869_),
    .A2(_07731_),
    .B(_07735_),
    .Y(_02711_));
 AND2x2_ASAP7_75t_R _27537_ (.A(_01959_),
    .B(_07734_),
    .Y(_07736_));
 AOI21x1_ASAP7_75t_R _27538_ (.A1(_01868_),
    .A2(_07731_),
    .B(_07736_),
    .Y(_02712_));
 AND2x2_ASAP7_75t_R _27539_ (.A(_01958_),
    .B(_07734_),
    .Y(_07737_));
 AOI21x1_ASAP7_75t_R _27540_ (.A1(_01867_),
    .A2(_07731_),
    .B(_07737_),
    .Y(_02713_));
 AND2x2_ASAP7_75t_R _27541_ (.A(_01957_),
    .B(_07734_),
    .Y(_07738_));
 AOI21x1_ASAP7_75t_R _27542_ (.A1(_01866_),
    .A2(_07731_),
    .B(_07738_),
    .Y(_02714_));
 AND2x2_ASAP7_75t_R _27543_ (.A(_01956_),
    .B(_07734_),
    .Y(_07739_));
 AOI21x1_ASAP7_75t_R _27544_ (.A1(_01865_),
    .A2(_07731_),
    .B(_07739_),
    .Y(_02715_));
 AND2x2_ASAP7_75t_R _27545_ (.A(_01955_),
    .B(_07734_),
    .Y(_07740_));
 AOI21x1_ASAP7_75t_R _27546_ (.A1(_01864_),
    .A2(_07731_),
    .B(_07740_),
    .Y(_02716_));
 NAND2x1_ASAP7_75t_R _27547_ (.A(_01954_),
    .B(_07702_),
    .Y(_07741_));
 OA21x2_ASAP7_75t_R _27548_ (.A1(_07612_),
    .A2(_07702_),
    .B(_07741_),
    .Y(_02717_));
 NAND2x1_ASAP7_75t_R _27549_ (.A(_01862_),
    .B(_07698_),
    .Y(_07742_));
 OA21x2_ASAP7_75t_R _27550_ (.A1(_07615_),
    .A2(_07697_),
    .B(_07742_),
    .Y(_02718_));
 AND2x2_ASAP7_75t_R _27551_ (.A(_01952_),
    .B(_07734_),
    .Y(_07743_));
 AOI21x1_ASAP7_75t_R _27552_ (.A1(_01861_),
    .A2(_07731_),
    .B(_07743_),
    .Y(_02719_));
 AND2x2_ASAP7_75t_R _27553_ (.A(_01951_),
    .B(_07734_),
    .Y(_07744_));
 AOI21x1_ASAP7_75t_R _27554_ (.A1(_01860_),
    .A2(_07731_),
    .B(_07744_),
    .Y(_02720_));
 AND2x2_ASAP7_75t_R _27555_ (.A(_01950_),
    .B(_07734_),
    .Y(_07745_));
 AOI21x1_ASAP7_75t_R _27556_ (.A1(_01859_),
    .A2(_07697_),
    .B(_07745_),
    .Y(_02721_));
 AND2x2_ASAP7_75t_R _27557_ (.A(_01949_),
    .B(_07734_),
    .Y(_07746_));
 AOI21x1_ASAP7_75t_R _27558_ (.A1(_01858_),
    .A2(_07697_),
    .B(_07746_),
    .Y(_02722_));
 AND2x2_ASAP7_75t_R _27559_ (.A(_01948_),
    .B(_07499_),
    .Y(_07747_));
 AOI21x1_ASAP7_75t_R _27560_ (.A1(_01857_),
    .A2(_07697_),
    .B(_07747_),
    .Y(_02723_));
 AND2x2_ASAP7_75t_R _27561_ (.A(_01947_),
    .B(_07499_),
    .Y(_07748_));
 AOI21x1_ASAP7_75t_R _27562_ (.A1(_01856_),
    .A2(_07697_),
    .B(_07748_),
    .Y(_02724_));
 NOR2x2_ASAP7_75t_R _27563_ (.A(_05916_),
    .B(_05994_),
    .Y(_07749_));
 NOR2x1_ASAP7_75t_R _27564_ (.A(_01855_),
    .B(_07749_),
    .Y(_07750_));
 AO21x1_ASAP7_75t_R _27565_ (.A1(_06695_),
    .A2(_07749_),
    .B(_07750_),
    .Y(_02725_));
 NOR2x1_ASAP7_75t_R _27566_ (.A(_01854_),
    .B(_07749_),
    .Y(_07751_));
 AO21x1_ASAP7_75t_R _27567_ (.A1(_06137_),
    .A2(_07749_),
    .B(_07751_),
    .Y(_02726_));
 NAND2x2_ASAP7_75t_R _27568_ (.A(_07230_),
    .B(_07545_),
    .Y(_07752_));
 AND3x1_ASAP7_75t_R _27569_ (.A(_06000_),
    .B(_06017_),
    .C(_07749_),
    .Y(_07753_));
 NOR2x1_ASAP7_75t_R _27570_ (.A(_07752_),
    .B(_07753_),
    .Y(_07754_));
 OR3x4_ASAP7_75t_R _27571_ (.A(_05059_),
    .B(_05765_),
    .C(_06234_),
    .Y(_07755_));
 NAND2x1_ASAP7_75t_R _27572_ (.A(_01853_),
    .B(_07755_),
    .Y(_07756_));
 AO222x2_ASAP7_75t_R _27573_ (.A1(\cs_registers_i.priv_lvl_q[0] ),
    .A2(_07702_),
    .B1(_07754_),
    .B2(_07756_),
    .C1(_07507_),
    .C2(_07709_),
    .Y(_02727_));
 NAND2x1_ASAP7_75t_R _27574_ (.A(_01852_),
    .B(_07755_),
    .Y(_07757_));
 OAI22x1_ASAP7_75t_R _27575_ (.A1(_05068_),
    .A2(_07700_),
    .B1(_07538_),
    .B2(_01889_),
    .Y(_07758_));
 AO21x1_ASAP7_75t_R _27576_ (.A1(_07754_),
    .A2(_07757_),
    .B(_07758_),
    .Y(_02728_));
 NOR2x1_ASAP7_75t_R _27577_ (.A(_06584_),
    .B(_07755_),
    .Y(_07759_));
 AO21x1_ASAP7_75t_R _27578_ (.A1(_01851_),
    .A2(_07755_),
    .B(_07759_),
    .Y(_07760_));
 INVx1_ASAP7_75t_R _27579_ (.A(_02220_),
    .Y(_07761_));
 AND3x1_ASAP7_75t_R _27580_ (.A(_07761_),
    .B(_01888_),
    .C(_05418_),
    .Y(_07762_));
 OA22x2_ASAP7_75t_R _27581_ (.A1(_01850_),
    .A2(_07700_),
    .B1(_07762_),
    .B2(_07230_),
    .Y(_07763_));
 OAI21x1_ASAP7_75t_R _27582_ (.A1(_07752_),
    .A2(_07760_),
    .B(_07763_),
    .Y(_02729_));
 AND5x2_ASAP7_75t_R _27583_ (.A(_18853_),
    .B(_18665_),
    .C(_05023_),
    .D(_05060_),
    .E(_05085_),
    .Y(_07764_));
 OAI21x1_ASAP7_75t_R _27584_ (.A1(_18658_),
    .A2(_05009_),
    .B(_14071_),
    .Y(_07765_));
 NAND2x1_ASAP7_75t_R _27585_ (.A(_07764_),
    .B(_07765_),
    .Y(_07766_));
 AO21x1_ASAP7_75t_R _27586_ (.A1(_07764_),
    .A2(_07765_),
    .B(_05375_),
    .Y(_07767_));
 OAI21x1_ASAP7_75t_R _27587_ (.A1(_06588_),
    .A2(_07766_),
    .B(_07767_),
    .Y(_07768_));
 OAI22x1_ASAP7_75t_R _27588_ (.A1(_01851_),
    .A2(_07230_),
    .B1(_07752_),
    .B2(_07768_),
    .Y(_02730_));
 NOR2x2_ASAP7_75t_R _27589_ (.A(_05980_),
    .B(_05916_),
    .Y(_07769_));
 BUFx4f_ASAP7_75t_R _27590_ (.A(_07769_),
    .Y(_07770_));
 BUFx6f_ASAP7_75t_R _27591_ (.A(_07769_),
    .Y(_07771_));
 NOR2x1_ASAP7_75t_R _27592_ (.A(_01849_),
    .B(_07771_),
    .Y(_07772_));
 AO21x1_ASAP7_75t_R _27593_ (.A1(_05841_),
    .A2(_07770_),
    .B(_07772_),
    .Y(_07773_));
 BUFx3_ASAP7_75t_R _27594_ (.A(_05329_),
    .Y(_07774_));
 BUFx4f_ASAP7_75t_R _27595_ (.A(_07493_),
    .Y(_07775_));
 INVx3_ASAP7_75t_R _27596_ (.A(_13417_),
    .Y(_07776_));
 BUFx3_ASAP7_75t_R _27597_ (.A(_07776_),
    .Y(_07777_));
 BUFx3_ASAP7_75t_R _27598_ (.A(_13417_),
    .Y(_07778_));
 AND2x2_ASAP7_75t_R _27599_ (.A(_07778_),
    .B(_13380_),
    .Y(_07779_));
 AO21x1_ASAP7_75t_R _27600_ (.A1(_07777_),
    .A2(_01545_),
    .B(_07779_),
    .Y(_07780_));
 BUFx4f_ASAP7_75t_R _27601_ (.A(_05328_),
    .Y(_07781_));
 OAI22x1_ASAP7_75t_R _27602_ (.A1(_01543_),
    .A2(_07775_),
    .B1(_07780_),
    .B2(_07781_),
    .Y(_07782_));
 AND4x1_ASAP7_75t_R _27603_ (.A(_07774_),
    .B(_05455_),
    .C(_07499_),
    .D(_07782_),
    .Y(_07783_));
 AO21x1_ASAP7_75t_R _27604_ (.A1(_07697_),
    .A2(_07773_),
    .B(_07783_),
    .Y(_02731_));
 NOR2x1_ASAP7_75t_R _27605_ (.A(_01848_),
    .B(_07770_),
    .Y(_07784_));
 AOI21x1_ASAP7_75t_R _27606_ (.A1(_06635_),
    .A2(_07770_),
    .B(_07784_),
    .Y(_07785_));
 NAND2x1_ASAP7_75t_R _27607_ (.A(_05077_),
    .B(_05326_),
    .Y(_07786_));
 BUFx4f_ASAP7_75t_R _27608_ (.A(_01554_),
    .Y(_07787_));
 OR4x2_ASAP7_75t_R _27609_ (.A(_00012_),
    .B(_07787_),
    .C(_00020_),
    .D(_01544_),
    .Y(_07788_));
 OR3x1_ASAP7_75t_R _27610_ (.A(_00023_),
    .B(_00026_),
    .C(_07788_),
    .Y(_07789_));
 OR2x2_ASAP7_75t_R _27611_ (.A(_00028_),
    .B(_07789_),
    .Y(_07790_));
 OR4x2_ASAP7_75t_R _27612_ (.A(_00030_),
    .B(_00033_),
    .C(_00036_),
    .D(_07790_),
    .Y(_07791_));
 XNOR2x1_ASAP7_75t_R _27613_ (.B(_07791_),
    .Y(_07792_),
    .A(_00039_));
 BUFx3_ASAP7_75t_R _27614_ (.A(_05061_),
    .Y(_07793_));
 BUFx3_ASAP7_75t_R _27615_ (.A(_04930_),
    .Y(_07794_));
 BUFx3_ASAP7_75t_R _27616_ (.A(_07493_),
    .Y(_07795_));
 AND2x2_ASAP7_75t_R _27617_ (.A(_07778_),
    .B(_14050_),
    .Y(_07796_));
 AO21x1_ASAP7_75t_R _27618_ (.A1(_07777_),
    .A2(_00038_),
    .B(_07796_),
    .Y(_07797_));
 OA222x2_ASAP7_75t_R _27619_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01542_),
    .C1(_07797_),
    .C2(_07781_),
    .Y(_07798_));
 AO21x1_ASAP7_75t_R _27620_ (.A1(_05337_),
    .A2(_07792_),
    .B(_07798_),
    .Y(_07799_));
 OR3x1_ASAP7_75t_R _27621_ (.A(_07786_),
    .B(_07700_),
    .C(_07799_),
    .Y(_07800_));
 OAI21x1_ASAP7_75t_R _27622_ (.A1(_07702_),
    .A2(_07785_),
    .B(_07800_),
    .Y(_02732_));
 NOR2x1_ASAP7_75t_R _27623_ (.A(_01847_),
    .B(_07771_),
    .Y(_07801_));
 AO21x1_ASAP7_75t_R _27624_ (.A1(_06639_),
    .A2(_07770_),
    .B(_07801_),
    .Y(_07802_));
 BUFx4f_ASAP7_75t_R _27625_ (.A(_05329_),
    .Y(_07803_));
 OR4x2_ASAP7_75t_R _27626_ (.A(_07787_),
    .B(_00020_),
    .C(_00023_),
    .D(_02315_),
    .Y(_07804_));
 OR3x2_ASAP7_75t_R _27627_ (.A(_00026_),
    .B(_00028_),
    .C(_07804_),
    .Y(_07805_));
 OR5x2_ASAP7_75t_R _27628_ (.A(_00030_),
    .B(_00033_),
    .C(_00036_),
    .D(_00039_),
    .E(_07805_),
    .Y(_07806_));
 XNOR2x1_ASAP7_75t_R _27629_ (.B(_07806_),
    .Y(_07807_),
    .A(_14806_));
 AND2x2_ASAP7_75t_R _27630_ (.A(_07778_),
    .B(_14231_),
    .Y(_07808_));
 AO21x1_ASAP7_75t_R _27631_ (.A1(_07777_),
    .A2(_00041_),
    .B(_07808_),
    .Y(_07809_));
 OA222x2_ASAP7_75t_R _27632_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01541_),
    .C1(_07809_),
    .C2(_07781_),
    .Y(_07810_));
 INVx1_ASAP7_75t_R _27633_ (.A(_07810_),
    .Y(_07811_));
 AND2x2_ASAP7_75t_R _27634_ (.A(_05455_),
    .B(_07498_),
    .Y(_07812_));
 BUFx3_ASAP7_75t_R _27635_ (.A(_07812_),
    .Y(_07813_));
 OA211x2_ASAP7_75t_R _27636_ (.A1(_07803_),
    .A2(_07807_),
    .B(_07811_),
    .C(_07813_),
    .Y(_07814_));
 AO21x1_ASAP7_75t_R _27637_ (.A1(_07697_),
    .A2(_07802_),
    .B(_07814_),
    .Y(_02733_));
 BUFx4f_ASAP7_75t_R _27638_ (.A(_07700_),
    .Y(_07815_));
 NOR2x1_ASAP7_75t_R _27639_ (.A(_01846_),
    .B(_07771_),
    .Y(_07816_));
 AO21x1_ASAP7_75t_R _27640_ (.A1(_06883_),
    .A2(_07770_),
    .B(_07816_),
    .Y(_07817_));
 OR2x2_ASAP7_75t_R _27641_ (.A(_00039_),
    .B(_07791_),
    .Y(_07818_));
 NOR2x1_ASAP7_75t_R _27642_ (.A(_00042_),
    .B(_07818_),
    .Y(_07819_));
 XNOR2x1_ASAP7_75t_R _27643_ (.B(_07819_),
    .Y(_07820_),
    .A(_00044_));
 AND2x2_ASAP7_75t_R _27644_ (.A(_13561_),
    .B(_13417_),
    .Y(_07821_));
 AO21x1_ASAP7_75t_R _27645_ (.A1(_07776_),
    .A2(_00043_),
    .B(_07821_),
    .Y(_07822_));
 OA222x2_ASAP7_75t_R _27646_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01540_),
    .C1(_07822_),
    .C2(_07781_),
    .Y(_07823_));
 INVx1_ASAP7_75t_R _27647_ (.A(_07823_),
    .Y(_07824_));
 OA211x2_ASAP7_75t_R _27648_ (.A1(_07803_),
    .A2(_07820_),
    .B(_07824_),
    .C(_07813_),
    .Y(_07825_));
 AO21x1_ASAP7_75t_R _27649_ (.A1(_07815_),
    .A2(_07817_),
    .B(_07825_),
    .Y(_02734_));
 BUFx3_ASAP7_75t_R _27650_ (.A(_07812_),
    .Y(_07826_));
 BUFx6f_ASAP7_75t_R _27651_ (.A(_05337_),
    .Y(_07827_));
 OR3x1_ASAP7_75t_R _27652_ (.A(_00042_),
    .B(_00044_),
    .C(_07806_),
    .Y(_07828_));
 XNOR2x1_ASAP7_75t_R _27653_ (.B(_07828_),
    .Y(_07829_),
    .A(_00046_));
 BUFx3_ASAP7_75t_R _27654_ (.A(_04930_),
    .Y(_07830_));
 AND2x2_ASAP7_75t_R _27655_ (.A(_13585_),
    .B(_07778_),
    .Y(_07831_));
 AO21x1_ASAP7_75t_R _27656_ (.A1(_07777_),
    .A2(_00045_),
    .B(_07831_),
    .Y(_07832_));
 OA222x2_ASAP7_75t_R _27657_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01539_),
    .C1(_07832_),
    .C2(_07781_),
    .Y(_07833_));
 AOI21x1_ASAP7_75t_R _27658_ (.A1(_07827_),
    .A2(_07829_),
    .B(_07833_),
    .Y(_07834_));
 BUFx4f_ASAP7_75t_R _27659_ (.A(_07769_),
    .Y(_07835_));
 BUFx6f_ASAP7_75t_R _27660_ (.A(_07769_),
    .Y(_07836_));
 NOR2x1_ASAP7_75t_R _27661_ (.A(_01845_),
    .B(_07836_),
    .Y(_07837_));
 AO21x1_ASAP7_75t_R _27662_ (.A1(_06650_),
    .A2(_07835_),
    .B(_07837_),
    .Y(_07838_));
 BUFx3_ASAP7_75t_R _27663_ (.A(_07546_),
    .Y(_07839_));
 AO22x1_ASAP7_75t_R _27664_ (.A1(_07826_),
    .A2(_07834_),
    .B1(_07838_),
    .B2(_07839_),
    .Y(_02735_));
 AND2x2_ASAP7_75t_R _27665_ (.A(_13595_),
    .B(_07778_),
    .Y(_07840_));
 AO21x1_ASAP7_75t_R _27666_ (.A1(_07777_),
    .A2(_00047_),
    .B(_07840_),
    .Y(_07841_));
 OA222x2_ASAP7_75t_R _27667_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01538_),
    .C1(_07841_),
    .C2(_07781_),
    .Y(_07842_));
 INVx1_ASAP7_75t_R _27668_ (.A(_07842_),
    .Y(_07843_));
 OR4x1_ASAP7_75t_R _27669_ (.A(_00042_),
    .B(_00044_),
    .C(_00046_),
    .D(_07818_),
    .Y(_07844_));
 NAND2x1_ASAP7_75t_R _27670_ (.A(_00048_),
    .B(_07844_),
    .Y(_07845_));
 OR2x4_ASAP7_75t_R _27671_ (.A(_00048_),
    .B(_07844_),
    .Y(_07846_));
 AO21x1_ASAP7_75t_R _27672_ (.A1(_07845_),
    .A2(_07846_),
    .B(_07803_),
    .Y(_07847_));
 BUFx4f_ASAP7_75t_R _27673_ (.A(_07769_),
    .Y(_07848_));
 NOR2x1_ASAP7_75t_R _27674_ (.A(_01844_),
    .B(_07769_),
    .Y(_07849_));
 AO21x1_ASAP7_75t_R _27675_ (.A1(_06065_),
    .A2(_07848_),
    .B(_07849_),
    .Y(_07850_));
 AO32x1_ASAP7_75t_R _27676_ (.A1(_07813_),
    .A2(_07843_),
    .A3(_07847_),
    .B1(_07850_),
    .B2(_07698_),
    .Y(_02736_));
 NOR2x1_ASAP7_75t_R _27677_ (.A(_01843_),
    .B(_07771_),
    .Y(_07851_));
 AO21x1_ASAP7_75t_R _27678_ (.A1(_06660_),
    .A2(_07770_),
    .B(_07851_),
    .Y(_07852_));
 OR5x2_ASAP7_75t_R _27679_ (.A(_00042_),
    .B(_00044_),
    .C(_00046_),
    .D(_00048_),
    .E(_07806_),
    .Y(_07853_));
 XNOR2x1_ASAP7_75t_R _27680_ (.B(_07853_),
    .Y(_07854_),
    .A(_16003_));
 AND2x2_ASAP7_75t_R _27681_ (.A(_14990_),
    .B(_13417_),
    .Y(_07855_));
 AO21x1_ASAP7_75t_R _27682_ (.A1(_07776_),
    .A2(_00049_),
    .B(_07855_),
    .Y(_07856_));
 OA222x2_ASAP7_75t_R _27683_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01537_),
    .C1(_07856_),
    .C2(_05328_),
    .Y(_07857_));
 INVx1_ASAP7_75t_R _27684_ (.A(_07857_),
    .Y(_07858_));
 OA211x2_ASAP7_75t_R _27685_ (.A1(_07803_),
    .A2(_07854_),
    .B(_07858_),
    .C(_07813_),
    .Y(_07859_));
 AO21x1_ASAP7_75t_R _27686_ (.A1(_07815_),
    .A2(_07852_),
    .B(_07859_),
    .Y(_02737_));
 NOR2x1_ASAP7_75t_R _27687_ (.A(_01842_),
    .B(_07771_),
    .Y(_07860_));
 AO21x1_ASAP7_75t_R _27688_ (.A1(_06111_),
    .A2(_07770_),
    .B(_07860_),
    .Y(_07861_));
 NOR2x1_ASAP7_75t_R _27689_ (.A(_00050_),
    .B(_07846_),
    .Y(_07862_));
 XNOR2x1_ASAP7_75t_R _27690_ (.B(_07862_),
    .Y(_07863_),
    .A(_00051_));
 BUFx4f_ASAP7_75t_R _27691_ (.A(_05061_),
    .Y(_07864_));
 BUFx3_ASAP7_75t_R _27692_ (.A(_07493_),
    .Y(_07865_));
 NAND2x2_ASAP7_75t_R _27693_ (.A(_13417_),
    .B(_07492_),
    .Y(_07866_));
 BUFx3_ASAP7_75t_R _27694_ (.A(_07866_),
    .Y(_07867_));
 OA222x2_ASAP7_75t_R _27695_ (.A1(_07864_),
    .A2(_07794_),
    .B1(_07865_),
    .B2(_01536_),
    .C1(_07867_),
    .C2(_14011_),
    .Y(_07868_));
 INVx1_ASAP7_75t_R _27696_ (.A(_07868_),
    .Y(_07869_));
 OA211x2_ASAP7_75t_R _27697_ (.A1(_07803_),
    .A2(_07863_),
    .B(_07869_),
    .C(_07813_),
    .Y(_07870_));
 AO21x1_ASAP7_75t_R _27698_ (.A1(_07815_),
    .A2(_07861_),
    .B(_07870_),
    .Y(_02738_));
 OR3x1_ASAP7_75t_R _27699_ (.A(_00050_),
    .B(_00051_),
    .C(_07853_),
    .Y(_07871_));
 XNOR2x1_ASAP7_75t_R _27700_ (.B(_07871_),
    .Y(_07872_),
    .A(_00052_));
 OA222x2_ASAP7_75t_R _27701_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01535_),
    .C1(_07867_),
    .C2(_15038_),
    .Y(_07873_));
 AOI21x1_ASAP7_75t_R _27702_ (.A1(_07827_),
    .A2(_07872_),
    .B(_07873_),
    .Y(_07874_));
 BUFx6f_ASAP7_75t_R _27703_ (.A(_07769_),
    .Y(_07875_));
 NOR2x1_ASAP7_75t_R _27704_ (.A(_01841_),
    .B(_07875_),
    .Y(_07876_));
 AO21x1_ASAP7_75t_R _27705_ (.A1(_06136_),
    .A2(_07835_),
    .B(_07876_),
    .Y(_07877_));
 AO22x1_ASAP7_75t_R _27706_ (.A1(_07826_),
    .A2(_07874_),
    .B1(_07877_),
    .B2(_07839_),
    .Y(_02739_));
 OR4x1_ASAP7_75t_R _27707_ (.A(_00050_),
    .B(_00051_),
    .C(_00052_),
    .D(_07846_),
    .Y(_07878_));
 XNOR2x1_ASAP7_75t_R _27708_ (.B(_07878_),
    .Y(_07879_),
    .A(_00053_));
 OA222x2_ASAP7_75t_R _27709_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01534_),
    .C1(_07867_),
    .C2(_13903_),
    .Y(_07880_));
 AOI21x1_ASAP7_75t_R _27710_ (.A1(_07827_),
    .A2(_07879_),
    .B(_07880_),
    .Y(_07881_));
 NOR2x1_ASAP7_75t_R _27711_ (.A(_01840_),
    .B(_07875_),
    .Y(_07882_));
 AO21x1_ASAP7_75t_R _27712_ (.A1(_06161_),
    .A2(_07848_),
    .B(_07882_),
    .Y(_07883_));
 AO22x1_ASAP7_75t_R _27713_ (.A1(_07826_),
    .A2(_07881_),
    .B1(_07883_),
    .B2(_07839_),
    .Y(_02740_));
 OR5x1_ASAP7_75t_R _27714_ (.A(_00050_),
    .B(_00051_),
    .C(_00052_),
    .D(_00053_),
    .E(_07853_),
    .Y(_07884_));
 XNOR2x1_ASAP7_75t_R _27715_ (.B(_07884_),
    .Y(_07885_),
    .A(_00054_));
 OA222x2_ASAP7_75t_R _27716_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01533_),
    .C1(_07867_),
    .C2(_15025_),
    .Y(_07886_));
 AOI21x1_ASAP7_75t_R _27717_ (.A1(_07827_),
    .A2(_07885_),
    .B(_07886_),
    .Y(_07887_));
 NOR2x1_ASAP7_75t_R _27718_ (.A(_01839_),
    .B(_07875_),
    .Y(_07888_));
 AO21x1_ASAP7_75t_R _27719_ (.A1(_06180_),
    .A2(_07848_),
    .B(_07888_),
    .Y(_07889_));
 AO22x1_ASAP7_75t_R _27720_ (.A1(_07826_),
    .A2(_07887_),
    .B1(_07889_),
    .B2(_07839_),
    .Y(_02741_));
 NOR2x1_ASAP7_75t_R _27721_ (.A(_01838_),
    .B(_07771_),
    .Y(_07890_));
 AO21x1_ASAP7_75t_R _27722_ (.A1(_06475_),
    .A2(_07770_),
    .B(_07890_),
    .Y(_07891_));
 XOR2x1_ASAP7_75t_R _27723_ (.A(_07787_),
    .Y(_07892_),
    .B(_01544_));
 AND2x2_ASAP7_75t_R _27724_ (.A(_07778_),
    .B(_00013_),
    .Y(_07893_));
 AO21x1_ASAP7_75t_R _27725_ (.A1(_07776_),
    .A2(_00014_),
    .B(_07893_),
    .Y(_07894_));
 OA222x2_ASAP7_75t_R _27726_ (.A1(_07864_),
    .A2(_07794_),
    .B1(_07865_),
    .B2(_01532_),
    .C1(_07894_),
    .C2(_05328_),
    .Y(_07895_));
 INVx1_ASAP7_75t_R _27727_ (.A(_07895_),
    .Y(_07896_));
 OA211x2_ASAP7_75t_R _27728_ (.A1(_07803_),
    .A2(_07892_),
    .B(_07896_),
    .C(_07813_),
    .Y(_07897_));
 AO21x1_ASAP7_75t_R _27729_ (.A1(_07815_),
    .A2(_07891_),
    .B(_07897_),
    .Y(_02742_));
 NOR2x1_ASAP7_75t_R _27730_ (.A(_01837_),
    .B(_07771_),
    .Y(_07898_));
 AO21x1_ASAP7_75t_R _27731_ (.A1(_06218_),
    .A2(_07770_),
    .B(_07898_),
    .Y(_07899_));
 OR5x2_ASAP7_75t_R _27732_ (.A(_00050_),
    .B(_00051_),
    .C(_00052_),
    .D(_00053_),
    .E(_00054_),
    .Y(_07900_));
 NOR2x1_ASAP7_75t_R _27733_ (.A(_07846_),
    .B(_07900_),
    .Y(_07901_));
 XNOR2x1_ASAP7_75t_R _27734_ (.B(_07901_),
    .Y(_07902_),
    .A(_00055_));
 BUFx3_ASAP7_75t_R _27735_ (.A(_04930_),
    .Y(_07903_));
 OA222x2_ASAP7_75t_R _27736_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01531_),
    .C1(_07866_),
    .C2(_15510_),
    .Y(_07904_));
 INVx1_ASAP7_75t_R _27737_ (.A(_07904_),
    .Y(_07905_));
 BUFx3_ASAP7_75t_R _27738_ (.A(_07812_),
    .Y(_07906_));
 OA211x2_ASAP7_75t_R _27739_ (.A1(_07803_),
    .A2(_07902_),
    .B(_07905_),
    .C(_07906_),
    .Y(_07907_));
 AO21x1_ASAP7_75t_R _27740_ (.A1(_07815_),
    .A2(_07899_),
    .B(_07907_),
    .Y(_02743_));
 NOR2x1_ASAP7_75t_R _27741_ (.A(_01836_),
    .B(_07836_),
    .Y(_07908_));
 AO21x1_ASAP7_75t_R _27742_ (.A1(_06695_),
    .A2(_07770_),
    .B(_07908_),
    .Y(_07909_));
 OR3x1_ASAP7_75t_R _27743_ (.A(_00055_),
    .B(_07853_),
    .C(_07900_),
    .Y(_07910_));
 XNOR2x1_ASAP7_75t_R _27744_ (.B(_07910_),
    .Y(_07911_),
    .A(_16752_));
 OA222x2_ASAP7_75t_R _27745_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01530_),
    .C1(_07866_),
    .C2(_16650_),
    .Y(_07912_));
 INVx1_ASAP7_75t_R _27746_ (.A(_07912_),
    .Y(_07913_));
 OA211x2_ASAP7_75t_R _27747_ (.A1(_07774_),
    .A2(_07911_),
    .B(_07913_),
    .C(_07906_),
    .Y(_07914_));
 AO21x1_ASAP7_75t_R _27748_ (.A1(_07815_),
    .A2(_07909_),
    .B(_07914_),
    .Y(_02744_));
 NOR2x1_ASAP7_75t_R _27749_ (.A(_01835_),
    .B(_07836_),
    .Y(_07915_));
 AO21x1_ASAP7_75t_R _27750_ (.A1(_06260_),
    .A2(_07835_),
    .B(_07915_),
    .Y(_07916_));
 OR4x1_ASAP7_75t_R _27751_ (.A(_00055_),
    .B(_00056_),
    .C(_07846_),
    .D(_07900_),
    .Y(_07917_));
 XNOR2x1_ASAP7_75t_R _27752_ (.B(_07917_),
    .Y(_07918_),
    .A(_16883_));
 OA222x2_ASAP7_75t_R _27753_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01529_),
    .C1(_07866_),
    .C2(_15747_),
    .Y(_07919_));
 INVx1_ASAP7_75t_R _27754_ (.A(_07919_),
    .Y(_07920_));
 OA211x2_ASAP7_75t_R _27755_ (.A1(_07774_),
    .A2(_07918_),
    .B(_07920_),
    .C(_07906_),
    .Y(_07921_));
 AO21x1_ASAP7_75t_R _27756_ (.A1(_07815_),
    .A2(_07916_),
    .B(_07921_),
    .Y(_02745_));
 OA222x2_ASAP7_75t_R _27757_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01528_),
    .C1(_07867_),
    .C2(_15568_),
    .Y(_07922_));
 INVx1_ASAP7_75t_R _27758_ (.A(_07922_),
    .Y(_07923_));
 OR4x2_ASAP7_75t_R _27759_ (.A(_00055_),
    .B(_00056_),
    .C(_00057_),
    .D(_07900_),
    .Y(_07924_));
 OAI21x1_ASAP7_75t_R _27760_ (.A1(_07853_),
    .A2(_07924_),
    .B(_00058_),
    .Y(_07925_));
 OR3x2_ASAP7_75t_R _27761_ (.A(_00058_),
    .B(_07853_),
    .C(_07924_),
    .Y(_07926_));
 AO21x1_ASAP7_75t_R _27762_ (.A1(_07925_),
    .A2(_07926_),
    .B(_07803_),
    .Y(_07927_));
 NOR2x1_ASAP7_75t_R _27763_ (.A(_01834_),
    .B(_07769_),
    .Y(_07928_));
 AO21x1_ASAP7_75t_R _27764_ (.A1(_06705_),
    .A2(_07771_),
    .B(_07928_),
    .Y(_07929_));
 AO32x1_ASAP7_75t_R _27765_ (.A1(_07813_),
    .A2(_07923_),
    .A3(_07927_),
    .B1(_07929_),
    .B2(_07700_),
    .Y(_02746_));
 NOR2x1_ASAP7_75t_R _27766_ (.A(_01833_),
    .B(_07836_),
    .Y(_07930_));
 AO21x1_ASAP7_75t_R _27767_ (.A1(_06299_),
    .A2(_07835_),
    .B(_07930_),
    .Y(_07931_));
 OR3x2_ASAP7_75t_R _27768_ (.A(_00058_),
    .B(_07846_),
    .C(_07924_),
    .Y(_07932_));
 XNOR2x1_ASAP7_75t_R _27769_ (.B(_07932_),
    .Y(_07933_),
    .A(_17122_));
 OA222x2_ASAP7_75t_R _27770_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01527_),
    .C1(_07866_),
    .C2(_15555_),
    .Y(_07934_));
 INVx1_ASAP7_75t_R _27771_ (.A(_07934_),
    .Y(_07935_));
 OA211x2_ASAP7_75t_R _27772_ (.A1(_07774_),
    .A2(_07933_),
    .B(_07935_),
    .C(_07906_),
    .Y(_07936_));
 AO21x1_ASAP7_75t_R _27773_ (.A1(_07815_),
    .A2(_07931_),
    .B(_07936_),
    .Y(_02747_));
 NOR2x1_ASAP7_75t_R _27774_ (.A(_01832_),
    .B(_07836_),
    .Y(_07937_));
 AO21x1_ASAP7_75t_R _27775_ (.A1(_06320_),
    .A2(_07835_),
    .B(_07937_),
    .Y(_07938_));
 NOR2x1_ASAP7_75t_R _27776_ (.A(_00059_),
    .B(_07926_),
    .Y(_07939_));
 XNOR2x1_ASAP7_75t_R _27777_ (.B(_07939_),
    .Y(_07940_),
    .A(_00060_));
 OA222x2_ASAP7_75t_R _27778_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01526_),
    .C1(_07866_),
    .C2(_13601_),
    .Y(_07941_));
 INVx1_ASAP7_75t_R _27779_ (.A(_07941_),
    .Y(_07942_));
 OA211x2_ASAP7_75t_R _27780_ (.A1(_07774_),
    .A2(_07940_),
    .B(_07942_),
    .C(_07906_),
    .Y(_07943_));
 AO21x1_ASAP7_75t_R _27781_ (.A1(_07815_),
    .A2(_07938_),
    .B(_07943_),
    .Y(_02748_));
 OR3x1_ASAP7_75t_R _27782_ (.A(_00059_),
    .B(_00060_),
    .C(_07932_),
    .Y(_07944_));
 XNOR2x1_ASAP7_75t_R _27783_ (.B(_07944_),
    .Y(_07945_),
    .A(_00061_));
 OA222x2_ASAP7_75t_R _27784_ (.A1(_07793_),
    .A2(_07830_),
    .B1(_07795_),
    .B2(_01525_),
    .C1(_07867_),
    .C2(_13589_),
    .Y(_07946_));
 AOI21x1_ASAP7_75t_R _27785_ (.A1(_07827_),
    .A2(_07945_),
    .B(_07946_),
    .Y(_07947_));
 NOR2x1_ASAP7_75t_R _27786_ (.A(_01831_),
    .B(_07875_),
    .Y(_07948_));
 AO21x1_ASAP7_75t_R _27787_ (.A1(_06968_),
    .A2(_07848_),
    .B(_07948_),
    .Y(_07949_));
 AO22x1_ASAP7_75t_R _27788_ (.A1(_07826_),
    .A2(_07947_),
    .B1(_07949_),
    .B2(_07839_),
    .Y(_02749_));
 NOR2x1_ASAP7_75t_R _27789_ (.A(_01830_),
    .B(_07836_),
    .Y(_07950_));
 AO21x1_ASAP7_75t_R _27790_ (.A1(_07431_),
    .A2(_07835_),
    .B(_07950_),
    .Y(_07951_));
 OR4x2_ASAP7_75t_R _27791_ (.A(_00059_),
    .B(_00060_),
    .C(_00061_),
    .D(_07926_),
    .Y(_07952_));
 XNOR2x1_ASAP7_75t_R _27792_ (.B(_07952_),
    .Y(_07953_),
    .A(_04389_));
 OA222x2_ASAP7_75t_R _27793_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01524_),
    .C1(_07866_),
    .C2(_13579_),
    .Y(_07954_));
 INVx1_ASAP7_75t_R _27794_ (.A(_07954_),
    .Y(_07955_));
 OA211x2_ASAP7_75t_R _27795_ (.A1(_07774_),
    .A2(_07953_),
    .B(_07955_),
    .C(_07906_),
    .Y(_07956_));
 AO21x1_ASAP7_75t_R _27796_ (.A1(_07815_),
    .A2(_07951_),
    .B(_07956_),
    .Y(_02750_));
 OR2x2_ASAP7_75t_R _27797_ (.A(_00061_),
    .B(_07944_),
    .Y(_07957_));
 NOR2x1_ASAP7_75t_R _27798_ (.A(_00062_),
    .B(_07957_),
    .Y(_07958_));
 XNOR2x1_ASAP7_75t_R _27799_ (.B(_07958_),
    .Y(_07959_),
    .A(_04519_));
 OA222x2_ASAP7_75t_R _27800_ (.A1(_07793_),
    .A2(_07830_),
    .B1(_07795_),
    .B2(_01523_),
    .C1(_07867_),
    .C2(_13578_),
    .Y(_07960_));
 AOI21x1_ASAP7_75t_R _27801_ (.A1(_07827_),
    .A2(_07959_),
    .B(_07960_),
    .Y(_07961_));
 NOR2x1_ASAP7_75t_R _27802_ (.A(_01829_),
    .B(_07875_),
    .Y(_07962_));
 AO21x1_ASAP7_75t_R _27803_ (.A1(_06738_),
    .A2(_07848_),
    .B(_07962_),
    .Y(_07963_));
 AO22x1_ASAP7_75t_R _27804_ (.A1(_07826_),
    .A2(_07961_),
    .B1(_07963_),
    .B2(_07839_),
    .Y(_02751_));
 OR3x1_ASAP7_75t_R _27805_ (.A(_00062_),
    .B(_00063_),
    .C(_07952_),
    .Y(_07964_));
 XNOR2x1_ASAP7_75t_R _27806_ (.B(_07964_),
    .Y(_07965_),
    .A(_00064_));
 OA222x2_ASAP7_75t_R _27807_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01522_),
    .C1(_07867_),
    .C2(_13577_),
    .Y(_07966_));
 AOI21x1_ASAP7_75t_R _27808_ (.A1(_07827_),
    .A2(_07965_),
    .B(_07966_),
    .Y(_07967_));
 NOR2x1_ASAP7_75t_R _27809_ (.A(_01828_),
    .B(_07875_),
    .Y(_07968_));
 AO21x1_ASAP7_75t_R _27810_ (.A1(_06411_),
    .A2(_07848_),
    .B(_07968_),
    .Y(_07969_));
 AO22x1_ASAP7_75t_R _27811_ (.A1(_07826_),
    .A2(_07967_),
    .B1(_07969_),
    .B2(_07698_),
    .Y(_02752_));
 NAND2x1_ASAP7_75t_R _27812_ (.A(\cs_registers_i.pc_id_i[2] ),
    .B(_07787_),
    .Y(_07970_));
 OA211x2_ASAP7_75t_R _27813_ (.A1(_00017_),
    .A2(_07787_),
    .B(_05337_),
    .C(_07970_),
    .Y(_07971_));
 INVx1_ASAP7_75t_R _27814_ (.A(_07971_),
    .Y(_07972_));
 AND2x2_ASAP7_75t_R _27815_ (.A(_07778_),
    .B(net2020),
    .Y(_07973_));
 AO21x1_ASAP7_75t_R _27816_ (.A1(_07777_),
    .A2(_00016_),
    .B(_07973_),
    .Y(_07974_));
 OA222x2_ASAP7_75t_R _27817_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01521_),
    .C1(_07974_),
    .C2(_07781_),
    .Y(_07975_));
 INVx1_ASAP7_75t_R _27818_ (.A(_07975_),
    .Y(_07976_));
 NOR2x1_ASAP7_75t_R _27819_ (.A(_01827_),
    .B(_07769_),
    .Y(_07977_));
 AO21x1_ASAP7_75t_R _27820_ (.A1(_05872_),
    .A2(_07771_),
    .B(_07977_),
    .Y(_07978_));
 AO32x1_ASAP7_75t_R _27821_ (.A1(_07813_),
    .A2(_07972_),
    .A3(_07976_),
    .B1(_07978_),
    .B2(_07700_),
    .Y(_02753_));
 OR4x1_ASAP7_75t_R _27822_ (.A(_00062_),
    .B(_00063_),
    .C(_00064_),
    .D(_07957_),
    .Y(_07979_));
 XNOR2x1_ASAP7_75t_R _27823_ (.B(_07979_),
    .Y(_07980_),
    .A(_00065_));
 OA222x2_ASAP7_75t_R _27824_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01520_),
    .C1(_07867_),
    .C2(_13575_),
    .Y(_07981_));
 AOI21x1_ASAP7_75t_R _27825_ (.A1(_07827_),
    .A2(_07980_),
    .B(_07981_),
    .Y(_07982_));
 NOR2x1_ASAP7_75t_R _27826_ (.A(_01826_),
    .B(_07875_),
    .Y(_07983_));
 AO21x1_ASAP7_75t_R _27827_ (.A1(_06750_),
    .A2(_07848_),
    .B(_07983_),
    .Y(_07984_));
 AO22x1_ASAP7_75t_R _27828_ (.A1(_07826_),
    .A2(_07982_),
    .B1(_07984_),
    .B2(_07698_),
    .Y(_02754_));
 OR5x2_ASAP7_75t_R _27829_ (.A(_00062_),
    .B(_00063_),
    .C(_00064_),
    .D(_00065_),
    .E(_07952_),
    .Y(_07985_));
 XNOR2x1_ASAP7_75t_R _27830_ (.B(_07985_),
    .Y(_07986_),
    .A(_00066_));
 OA222x2_ASAP7_75t_R _27831_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01519_),
    .C1(_07867_),
    .C2(_13576_),
    .Y(_07987_));
 AOI21x1_ASAP7_75t_R _27832_ (.A1(_07827_),
    .A2(_07986_),
    .B(_07987_),
    .Y(_07988_));
 NOR2x1_ASAP7_75t_R _27833_ (.A(_01825_),
    .B(_07875_),
    .Y(_07989_));
 AO21x1_ASAP7_75t_R _27834_ (.A1(_07369_),
    .A2(_07848_),
    .B(_07989_),
    .Y(_07990_));
 AO22x1_ASAP7_75t_R _27835_ (.A1(_07826_),
    .A2(_07988_),
    .B1(_07990_),
    .B2(_07698_),
    .Y(_02755_));
 OR3x1_ASAP7_75t_R _27836_ (.A(_07787_),
    .B(_00020_),
    .C(_02315_),
    .Y(_07991_));
 OAI21x1_ASAP7_75t_R _27837_ (.A1(_07787_),
    .A2(_02315_),
    .B(_00020_),
    .Y(_07992_));
 AO21x1_ASAP7_75t_R _27838_ (.A1(_07991_),
    .A2(_07992_),
    .B(_07803_),
    .Y(_07993_));
 AND2x2_ASAP7_75t_R _27839_ (.A(_07778_),
    .B(_13383_),
    .Y(_07994_));
 AO21x1_ASAP7_75t_R _27840_ (.A1(_07777_),
    .A2(_00019_),
    .B(_07994_),
    .Y(_07995_));
 OA222x2_ASAP7_75t_R _27841_ (.A1(_05062_),
    .A2(_07830_),
    .B1(_07775_),
    .B2(_01518_),
    .C1(_07995_),
    .C2(_07781_),
    .Y(_07996_));
 INVx1_ASAP7_75t_R _27842_ (.A(_07996_),
    .Y(_07997_));
 NOR2x1_ASAP7_75t_R _27843_ (.A(_01824_),
    .B(_07769_),
    .Y(_07998_));
 AO21x1_ASAP7_75t_R _27844_ (.A1(_06500_),
    .A2(_07771_),
    .B(_07998_),
    .Y(_07999_));
 AO32x1_ASAP7_75t_R _27845_ (.A1(_07813_),
    .A2(_07993_),
    .A3(_07997_),
    .B1(_07999_),
    .B2(_07700_),
    .Y(_02756_));
 NOR2x1_ASAP7_75t_R _27846_ (.A(_01823_),
    .B(_07836_),
    .Y(_08000_));
 AO21x1_ASAP7_75t_R _27847_ (.A1(_07042_),
    .A2(_07835_),
    .B(_08000_),
    .Y(_08001_));
 XNOR2x1_ASAP7_75t_R _27848_ (.B(_07788_),
    .Y(_08002_),
    .A(_15054_));
 AND2x2_ASAP7_75t_R _27849_ (.A(_13417_),
    .B(_13569_),
    .Y(_08003_));
 AO21x1_ASAP7_75t_R _27850_ (.A1(_07776_),
    .A2(_00022_),
    .B(_08003_),
    .Y(_08004_));
 OA222x2_ASAP7_75t_R _27851_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01517_),
    .C1(_08004_),
    .C2(_05328_),
    .Y(_08005_));
 INVx1_ASAP7_75t_R _27852_ (.A(_08005_),
    .Y(_08006_));
 OA211x2_ASAP7_75t_R _27853_ (.A1(_07774_),
    .A2(_08002_),
    .B(_08006_),
    .C(_07906_),
    .Y(_08007_));
 AO21x1_ASAP7_75t_R _27854_ (.A1(_07839_),
    .A2(_08001_),
    .B(_08007_),
    .Y(_02757_));
 NOR2x1_ASAP7_75t_R _27855_ (.A(_01822_),
    .B(_07836_),
    .Y(_08008_));
 AO21x1_ASAP7_75t_R _27856_ (.A1(_06534_),
    .A2(_07835_),
    .B(_08008_),
    .Y(_08009_));
 XNOR2x1_ASAP7_75t_R _27857_ (.B(_07804_),
    .Y(_08010_),
    .A(_15116_));
 AND2x2_ASAP7_75t_R _27858_ (.A(_13417_),
    .B(net2013),
    .Y(_08011_));
 AO21x1_ASAP7_75t_R _27859_ (.A1(_07776_),
    .A2(_00025_),
    .B(_08011_),
    .Y(_08012_));
 OA222x2_ASAP7_75t_R _27860_ (.A1(_07864_),
    .A2(_07903_),
    .B1(_07865_),
    .B2(_01516_),
    .C1(_08012_),
    .C2(_05328_),
    .Y(_08013_));
 INVx1_ASAP7_75t_R _27861_ (.A(_08013_),
    .Y(_08014_));
 OA211x2_ASAP7_75t_R _27862_ (.A1(_07774_),
    .A2(_08010_),
    .B(_08014_),
    .C(_07906_),
    .Y(_08015_));
 AO21x1_ASAP7_75t_R _27863_ (.A1(_07839_),
    .A2(_08009_),
    .B(_08015_),
    .Y(_02758_));
 AND2x2_ASAP7_75t_R _27864_ (.A(_13554_),
    .B(_07778_),
    .Y(_08016_));
 AO21x1_ASAP7_75t_R _27865_ (.A1(_07777_),
    .A2(_00027_),
    .B(_08016_),
    .Y(_08017_));
 OAI22x1_ASAP7_75t_R _27866_ (.A1(_01515_),
    .A2(_07775_),
    .B1(_08017_),
    .B2(_07781_),
    .Y(_08018_));
 NAND2x1_ASAP7_75t_R _27867_ (.A(_00028_),
    .B(_07789_),
    .Y(_08019_));
 AND3x1_ASAP7_75t_R _27868_ (.A(_05337_),
    .B(_07790_),
    .C(_08019_),
    .Y(_08020_));
 AO21x1_ASAP7_75t_R _27869_ (.A1(_07803_),
    .A2(_08018_),
    .B(_08020_),
    .Y(_08021_));
 NOR2x1_ASAP7_75t_R _27870_ (.A(_01821_),
    .B(_07875_),
    .Y(_08022_));
 AO21x1_ASAP7_75t_R _27871_ (.A1(_06559_),
    .A2(_07848_),
    .B(_08022_),
    .Y(_08023_));
 AO22x1_ASAP7_75t_R _27872_ (.A1(_07826_),
    .A2(_08021_),
    .B1(_08023_),
    .B2(_07698_),
    .Y(_02759_));
 NOR2x1_ASAP7_75t_R _27873_ (.A(_01820_),
    .B(_07836_),
    .Y(_08024_));
 AO21x1_ASAP7_75t_R _27874_ (.A1(_06584_),
    .A2(_07835_),
    .B(_08024_),
    .Y(_08025_));
 XNOR2x1_ASAP7_75t_R _27875_ (.B(_07805_),
    .Y(_08026_),
    .A(_15235_));
 BUFx6f_ASAP7_75t_R _27876_ (.A(_00446_),
    .Y(_08027_));
 AND2x2_ASAP7_75t_R _27877_ (.A(_08027_),
    .B(_13417_),
    .Y(_08028_));
 AO21x1_ASAP7_75t_R _27878_ (.A1(_07776_),
    .A2(_00029_),
    .B(_08028_),
    .Y(_08029_));
 OA222x2_ASAP7_75t_R _27879_ (.A1(_05061_),
    .A2(_07903_),
    .B1(_07493_),
    .B2(_01514_),
    .C1(_08029_),
    .C2(_05328_),
    .Y(_08030_));
 INVx1_ASAP7_75t_R _27880_ (.A(_08030_),
    .Y(_08031_));
 OA211x2_ASAP7_75t_R _27881_ (.A1(_07774_),
    .A2(_08026_),
    .B(_08031_),
    .C(_07906_),
    .Y(_08032_));
 AO21x1_ASAP7_75t_R _27882_ (.A1(_07839_),
    .A2(_08025_),
    .B(_08032_),
    .Y(_02760_));
 NOR2x1_ASAP7_75t_R _27883_ (.A(_01819_),
    .B(_07836_),
    .Y(_08033_));
 AO21x1_ASAP7_75t_R _27884_ (.A1(_06609_),
    .A2(_07835_),
    .B(_08033_),
    .Y(_08034_));
 NOR2x1_ASAP7_75t_R _27885_ (.A(_00030_),
    .B(_07790_),
    .Y(_08035_));
 XNOR2x1_ASAP7_75t_R _27886_ (.B(_08035_),
    .Y(_08036_),
    .A(_00033_));
 AND2x2_ASAP7_75t_R _27887_ (.A(_13417_),
    .B(_13438_),
    .Y(_08037_));
 AO21x1_ASAP7_75t_R _27888_ (.A1(_07776_),
    .A2(_00032_),
    .B(_08037_),
    .Y(_08038_));
 OA222x2_ASAP7_75t_R _27889_ (.A1(_05061_),
    .A2(_07903_),
    .B1(_07493_),
    .B2(_01513_),
    .C1(_08038_),
    .C2(_05328_),
    .Y(_08039_));
 INVx1_ASAP7_75t_R _27890_ (.A(_08039_),
    .Y(_08040_));
 OA211x2_ASAP7_75t_R _27891_ (.A1(_07774_),
    .A2(_08036_),
    .B(_08040_),
    .C(_07906_),
    .Y(_08041_));
 AO21x1_ASAP7_75t_R _27892_ (.A1(_07839_),
    .A2(_08034_),
    .B(_08041_),
    .Y(_02761_));
 OR3x1_ASAP7_75t_R _27893_ (.A(_00030_),
    .B(_00033_),
    .C(_07805_),
    .Y(_08042_));
 XNOR2x1_ASAP7_75t_R _27894_ (.B(_08042_),
    .Y(_08043_),
    .A(_00036_));
 AND2x2_ASAP7_75t_R _27895_ (.A(_07778_),
    .B(_14049_),
    .Y(_08044_));
 AO21x1_ASAP7_75t_R _27896_ (.A1(_07777_),
    .A2(_00035_),
    .B(_08044_),
    .Y(_08045_));
 OA222x2_ASAP7_75t_R _27897_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_01512_),
    .C1(_08045_),
    .C2(_07781_),
    .Y(_08046_));
 AOI21x1_ASAP7_75t_R _27898_ (.A1(_07827_),
    .A2(_08043_),
    .B(_08046_),
    .Y(_08047_));
 NOR2x1_ASAP7_75t_R _27899_ (.A(_01818_),
    .B(_07875_),
    .Y(_08048_));
 AO21x1_ASAP7_75t_R _27900_ (.A1(_06627_),
    .A2(_07848_),
    .B(_08048_),
    .Y(_08049_));
 AO22x1_ASAP7_75t_R _27901_ (.A1(_07813_),
    .A2(_08047_),
    .B1(_08049_),
    .B2(_07698_),
    .Y(_02762_));
 NAND2x2_ASAP7_75t_R _27902_ (.A(_04932_),
    .B(_05380_),
    .Y(_08050_));
 BUFx4f_ASAP7_75t_R _27903_ (.A(_08050_),
    .Y(_08051_));
 BUFx6f_ASAP7_75t_R _27904_ (.A(_08050_),
    .Y(_08052_));
 AND2x4_ASAP7_75t_R _27905_ (.A(_05877_),
    .B(_05811_),
    .Y(_08053_));
 OR3x4_ASAP7_75t_R _27906_ (.A(_05058_),
    .B(_05765_),
    .C(_05809_),
    .Y(_08054_));
 BUFx4f_ASAP7_75t_R _27907_ (.A(_08054_),
    .Y(_08055_));
 AND2x2_ASAP7_75t_R _27908_ (.A(_01467_),
    .B(_08055_),
    .Y(_08056_));
 AO21x1_ASAP7_75t_R _27909_ (.A1(_05956_),
    .A2(_08053_),
    .B(_08056_),
    .Y(_08057_));
 NAND2x1_ASAP7_75t_R _27910_ (.A(_08052_),
    .B(_08057_),
    .Y(_08058_));
 OA21x2_ASAP7_75t_R _27911_ (.A1(net23),
    .A2(_08051_),
    .B(_08058_),
    .Y(_02763_));
 AND2x2_ASAP7_75t_R _27912_ (.A(_00785_),
    .B(_08055_),
    .Y(_08059_));
 AO21x1_ASAP7_75t_R _27913_ (.A1(_06000_),
    .A2(_08053_),
    .B(_08059_),
    .Y(_08060_));
 NAND2x1_ASAP7_75t_R _27914_ (.A(_08052_),
    .B(_08060_),
    .Y(_08061_));
 OA21x2_ASAP7_75t_R _27915_ (.A1(net24),
    .A2(_08051_),
    .B(_08061_),
    .Y(_02764_));
 AND2x2_ASAP7_75t_R _27916_ (.A(_00784_),
    .B(_08055_),
    .Y(_08062_));
 AO21x1_ASAP7_75t_R _27917_ (.A1(_06017_),
    .A2(_08053_),
    .B(_08062_),
    .Y(_08063_));
 NAND2x1_ASAP7_75t_R _27918_ (.A(_08052_),
    .B(_08063_),
    .Y(_08064_));
 OA21x2_ASAP7_75t_R _27919_ (.A1(net25),
    .A2(_08051_),
    .B(_08064_),
    .Y(_02765_));
 BUFx6f_ASAP7_75t_R _27920_ (.A(_08055_),
    .Y(_08065_));
 NAND2x1_ASAP7_75t_R _27921_ (.A(_01468_),
    .B(_08065_),
    .Y(_08066_));
 BUFx6f_ASAP7_75t_R _27922_ (.A(_08054_),
    .Y(_08067_));
 OR2x2_ASAP7_75t_R _27923_ (.A(_06042_),
    .B(_08067_),
    .Y(_08068_));
 AND3x1_ASAP7_75t_R _27924_ (.A(_04932_),
    .B(_04934_),
    .C(_04935_),
    .Y(_08069_));
 BUFx4f_ASAP7_75t_R _27925_ (.A(_08069_),
    .Y(_08070_));
 BUFx4f_ASAP7_75t_R _27926_ (.A(_08070_),
    .Y(_08071_));
 AO21x1_ASAP7_75t_R _27927_ (.A1(_08066_),
    .A2(_08068_),
    .B(_08071_),
    .Y(_08072_));
 OA21x2_ASAP7_75t_R _27928_ (.A1(net26),
    .A2(_08051_),
    .B(_08072_),
    .Y(_02766_));
 NAND2x1_ASAP7_75t_R _27929_ (.A(_01469_),
    .B(_08065_),
    .Y(_08073_));
 OR2x2_ASAP7_75t_R _27930_ (.A(_06065_),
    .B(_08067_),
    .Y(_08074_));
 AO21x1_ASAP7_75t_R _27931_ (.A1(_08073_),
    .A2(_08074_),
    .B(_08071_),
    .Y(_08075_));
 OA21x2_ASAP7_75t_R _27932_ (.A1(net27),
    .A2(_08051_),
    .B(_08075_),
    .Y(_02767_));
 NAND2x1_ASAP7_75t_R _27933_ (.A(_01470_),
    .B(_08065_),
    .Y(_08076_));
 BUFx3_ASAP7_75t_R _27934_ (.A(_08054_),
    .Y(_08077_));
 OR2x2_ASAP7_75t_R _27935_ (.A(_06088_),
    .B(_08077_),
    .Y(_08078_));
 AO21x1_ASAP7_75t_R _27936_ (.A1(_08076_),
    .A2(_08078_),
    .B(_08071_),
    .Y(_08079_));
 OA21x2_ASAP7_75t_R _27937_ (.A1(net28),
    .A2(_08051_),
    .B(_08079_),
    .Y(_02768_));
 NAND2x1_ASAP7_75t_R _27938_ (.A(_01471_),
    .B(_08065_),
    .Y(_08080_));
 OR2x2_ASAP7_75t_R _27939_ (.A(_06111_),
    .B(_08077_),
    .Y(_08081_));
 AO21x1_ASAP7_75t_R _27940_ (.A1(_08080_),
    .A2(_08081_),
    .B(_08071_),
    .Y(_08082_));
 OA21x2_ASAP7_75t_R _27941_ (.A1(net29),
    .A2(_08051_),
    .B(_08082_),
    .Y(_02769_));
 NAND2x1_ASAP7_75t_R _27942_ (.A(_01472_),
    .B(_08065_),
    .Y(_08083_));
 OR2x2_ASAP7_75t_R _27943_ (.A(_06136_),
    .B(_08077_),
    .Y(_08084_));
 AO21x1_ASAP7_75t_R _27944_ (.A1(_08083_),
    .A2(_08084_),
    .B(_08071_),
    .Y(_08085_));
 OA21x2_ASAP7_75t_R _27945_ (.A1(net30),
    .A2(_08051_),
    .B(_08085_),
    .Y(_02770_));
 NAND2x1_ASAP7_75t_R _27946_ (.A(_01473_),
    .B(_08065_),
    .Y(_08086_));
 OR2x2_ASAP7_75t_R _27947_ (.A(_06160_),
    .B(_08077_),
    .Y(_08087_));
 AO21x1_ASAP7_75t_R _27948_ (.A1(_08086_),
    .A2(_08087_),
    .B(_08071_),
    .Y(_08088_));
 OA21x2_ASAP7_75t_R _27949_ (.A1(net31),
    .A2(_08051_),
    .B(_08088_),
    .Y(_02771_));
 NAND2x1_ASAP7_75t_R _27950_ (.A(_01474_),
    .B(_08065_),
    .Y(_08089_));
 OR2x2_ASAP7_75t_R _27951_ (.A(_06179_),
    .B(_08077_),
    .Y(_08090_));
 AO21x1_ASAP7_75t_R _27952_ (.A1(_08089_),
    .A2(_08090_),
    .B(_08071_),
    .Y(_08091_));
 OA21x2_ASAP7_75t_R _27953_ (.A1(net32),
    .A2(_08051_),
    .B(_08091_),
    .Y(_02772_));
 BUFx4f_ASAP7_75t_R _27954_ (.A(_08050_),
    .Y(_08092_));
 NAND2x1_ASAP7_75t_R _27955_ (.A(_01475_),
    .B(_08065_),
    .Y(_08093_));
 OR2x2_ASAP7_75t_R _27956_ (.A(_06217_),
    .B(_08077_),
    .Y(_08094_));
 AO21x1_ASAP7_75t_R _27957_ (.A1(_08093_),
    .A2(_08094_),
    .B(_08071_),
    .Y(_08095_));
 OA21x2_ASAP7_75t_R _27958_ (.A1(net33),
    .A2(_08092_),
    .B(_08095_),
    .Y(_02773_));
 NAND2x1_ASAP7_75t_R _27959_ (.A(_01476_),
    .B(_08065_),
    .Y(_08096_));
 OR2x2_ASAP7_75t_R _27960_ (.A(_06241_),
    .B(_08077_),
    .Y(_08097_));
 AO21x1_ASAP7_75t_R _27961_ (.A1(_08096_),
    .A2(_08097_),
    .B(_08071_),
    .Y(_08098_));
 OA21x2_ASAP7_75t_R _27962_ (.A1(net34),
    .A2(_08092_),
    .B(_08098_),
    .Y(_02774_));
 NAND2x1_ASAP7_75t_R _27963_ (.A(_01477_),
    .B(_08065_),
    .Y(_08099_));
 OR2x2_ASAP7_75t_R _27964_ (.A(_06259_),
    .B(_08077_),
    .Y(_08100_));
 AO21x1_ASAP7_75t_R _27965_ (.A1(_08099_),
    .A2(_08100_),
    .B(_08071_),
    .Y(_08101_));
 OA21x2_ASAP7_75t_R _27966_ (.A1(net35),
    .A2(_08092_),
    .B(_08101_),
    .Y(_02775_));
 NAND2x1_ASAP7_75t_R _27967_ (.A(_01478_),
    .B(_08067_),
    .Y(_08102_));
 OR2x2_ASAP7_75t_R _27968_ (.A(_06280_),
    .B(_08077_),
    .Y(_08103_));
 AO21x1_ASAP7_75t_R _27969_ (.A1(_08102_),
    .A2(_08103_),
    .B(_08070_),
    .Y(_08104_));
 OA21x2_ASAP7_75t_R _27970_ (.A1(net36),
    .A2(_08092_),
    .B(_08104_),
    .Y(_02776_));
 NAND2x1_ASAP7_75t_R _27971_ (.A(_01479_),
    .B(_08067_),
    .Y(_08105_));
 OR2x2_ASAP7_75t_R _27972_ (.A(_06298_),
    .B(_08077_),
    .Y(_08106_));
 AO21x1_ASAP7_75t_R _27973_ (.A1(_08105_),
    .A2(_08106_),
    .B(_08070_),
    .Y(_08107_));
 OA21x2_ASAP7_75t_R _27974_ (.A1(net37),
    .A2(_08092_),
    .B(_08107_),
    .Y(_02777_));
 NAND2x1_ASAP7_75t_R _27975_ (.A(_01480_),
    .B(_08067_),
    .Y(_08108_));
 OR2x2_ASAP7_75t_R _27976_ (.A(_06319_),
    .B(_08055_),
    .Y(_08109_));
 AO21x1_ASAP7_75t_R _27977_ (.A1(_08108_),
    .A2(_08109_),
    .B(_08070_),
    .Y(_08110_));
 OA21x2_ASAP7_75t_R _27978_ (.A1(net38),
    .A2(_08092_),
    .B(_08110_),
    .Y(_02778_));
 AND2x2_ASAP7_75t_R _27979_ (.A(_01481_),
    .B(_08054_),
    .Y(_08111_));
 AO21x1_ASAP7_75t_R _27980_ (.A1(_06347_),
    .A2(_08053_),
    .B(_08111_),
    .Y(_08112_));
 NAND2x1_ASAP7_75t_R _27981_ (.A(_08052_),
    .B(_08112_),
    .Y(_08113_));
 OA21x2_ASAP7_75t_R _27982_ (.A1(net39),
    .A2(_08092_),
    .B(_08113_),
    .Y(_02779_));
 AND2x2_ASAP7_75t_R _27983_ (.A(_00007_),
    .B(_08054_),
    .Y(_08114_));
 AO21x1_ASAP7_75t_R _27984_ (.A1(_06370_),
    .A2(_08053_),
    .B(_08114_),
    .Y(_08115_));
 NAND2x1_ASAP7_75t_R _27985_ (.A(_08052_),
    .B(_08115_),
    .Y(_08116_));
 OA21x2_ASAP7_75t_R _27986_ (.A1(net40),
    .A2(_08092_),
    .B(_08116_),
    .Y(_02780_));
 NAND2x1_ASAP7_75t_R _27987_ (.A(_00008_),
    .B(_08067_),
    .Y(_08117_));
 OR2x2_ASAP7_75t_R _27988_ (.A(_06392_),
    .B(_08055_),
    .Y(_08118_));
 AO21x1_ASAP7_75t_R _27989_ (.A1(_08117_),
    .A2(_08118_),
    .B(_08070_),
    .Y(_08119_));
 OA21x2_ASAP7_75t_R _27990_ (.A1(net41),
    .A2(_08092_),
    .B(_08119_),
    .Y(_02781_));
 NAND2x1_ASAP7_75t_R _27991_ (.A(_00009_),
    .B(_08067_),
    .Y(_08120_));
 OR2x2_ASAP7_75t_R _27992_ (.A(_06411_),
    .B(_08055_),
    .Y(_08121_));
 AO21x1_ASAP7_75t_R _27993_ (.A1(_08120_),
    .A2(_08121_),
    .B(_08070_),
    .Y(_08122_));
 OA21x2_ASAP7_75t_R _27994_ (.A1(net42),
    .A2(_08092_),
    .B(_08122_),
    .Y(_02782_));
 NAND2x1_ASAP7_75t_R _27995_ (.A(_00010_),
    .B(_08067_),
    .Y(_08123_));
 OR2x2_ASAP7_75t_R _27996_ (.A(_06439_),
    .B(_08055_),
    .Y(_08124_));
 AO21x1_ASAP7_75t_R _27997_ (.A1(_08123_),
    .A2(_08124_),
    .B(_08070_),
    .Y(_08125_));
 OA21x2_ASAP7_75t_R _27998_ (.A1(net43),
    .A2(_08052_),
    .B(_08125_),
    .Y(_02783_));
 AND2x2_ASAP7_75t_R _27999_ (.A(_00011_),
    .B(_08054_),
    .Y(_08126_));
 AO21x1_ASAP7_75t_R _28000_ (.A1(_06455_),
    .A2(_08053_),
    .B(_08126_),
    .Y(_08127_));
 NAND2x1_ASAP7_75t_R _28001_ (.A(_08052_),
    .B(_08127_),
    .Y(_08128_));
 OA21x2_ASAP7_75t_R _28002_ (.A1(net44),
    .A2(_08052_),
    .B(_08128_),
    .Y(_02784_));
 NAND2x1_ASAP7_75t_R _28003_ (.A(_01465_),
    .B(_08067_),
    .Y(_08129_));
 OR2x2_ASAP7_75t_R _28004_ (.A(_06609_),
    .B(_08055_),
    .Y(_08130_));
 AO21x1_ASAP7_75t_R _28005_ (.A1(_08129_),
    .A2(_08130_),
    .B(_08070_),
    .Y(_08131_));
 OA21x2_ASAP7_75t_R _28006_ (.A1(net45),
    .A2(_08052_),
    .B(_08131_),
    .Y(_02785_));
 NAND2x1_ASAP7_75t_R _28007_ (.A(_01466_),
    .B(_08067_),
    .Y(_08132_));
 OR2x2_ASAP7_75t_R _28008_ (.A(_06626_),
    .B(_08055_),
    .Y(_08133_));
 AO21x1_ASAP7_75t_R _28009_ (.A1(_08132_),
    .A2(_08133_),
    .B(_08070_),
    .Y(_08134_));
 OA21x2_ASAP7_75t_R _28010_ (.A1(net46),
    .A2(_08052_),
    .B(_08134_),
    .Y(_02786_));
 OA21x2_ASAP7_75t_R _28011_ (.A1(_13560_),
    .A2(_13589_),
    .B(_13585_),
    .Y(_08135_));
 NAND2x2_ASAP7_75t_R _28012_ (.A(_05096_),
    .B(_08135_),
    .Y(_08136_));
 BUFx6f_ASAP7_75t_R _28013_ (.A(_08136_),
    .Y(_08137_));
 BUFx4f_ASAP7_75t_R _28014_ (.A(_08137_),
    .Y(_08138_));
 OR3x1_ASAP7_75t_R _28015_ (.A(_02211_),
    .B(_05098_),
    .C(_08138_),
    .Y(_08139_));
 NAND2x1_ASAP7_75t_R _28016_ (.A(_01817_),
    .B(_08139_),
    .Y(_08140_));
 OA21x2_ASAP7_75t_R _28017_ (.A1(_05137_),
    .A2(_08139_),
    .B(_08140_),
    .Y(_02787_));
 AND3x4_ASAP7_75t_R _28018_ (.A(_05524_),
    .B(_02211_),
    .C(_02212_),
    .Y(_08141_));
 AND3x1_ASAP7_75t_R _28019_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_05158_),
    .C(_08141_),
    .Y(_08142_));
 AOI21x1_ASAP7_75t_R _28020_ (.A1(_05162_),
    .A2(_05099_),
    .B(_08142_),
    .Y(_02788_));
 BUFx6f_ASAP7_75t_R _28021_ (.A(_02316_),
    .Y(_08143_));
 INVx2_ASAP7_75t_R _28022_ (.A(_08143_),
    .Y(_08144_));
 AND3x1_ASAP7_75t_R _28023_ (.A(_08144_),
    .B(_05132_),
    .C(_08141_),
    .Y(_08145_));
 AOI21x1_ASAP7_75t_R _28024_ (.A1(_18868_),
    .A2(_05099_),
    .B(_08145_),
    .Y(_02789_));
 XNOR2x1_ASAP7_75t_R _28025_ (.B(_02317_),
    .Y(_08146_),
    .A(_00069_));
 AND3x1_ASAP7_75t_R _28026_ (.A(_05158_),
    .B(_08141_),
    .C(_08146_),
    .Y(_08147_));
 AOI21x1_ASAP7_75t_R _28027_ (.A1(_05101_),
    .A2(_05099_),
    .B(_08147_),
    .Y(_02790_));
 BUFx4f_ASAP7_75t_R _28028_ (.A(_05094_),
    .Y(_08148_));
 AND3x1_ASAP7_75t_R _28029_ (.A(_00069_),
    .B(_18867_),
    .C(_18868_),
    .Y(_08149_));
 XNOR2x2_ASAP7_75t_R _28030_ (.A(_05095_),
    .B(_08149_),
    .Y(_08150_));
 AND3x1_ASAP7_75t_R _28031_ (.A(_05158_),
    .B(_08141_),
    .C(_08150_),
    .Y(_08151_));
 AOI21x1_ASAP7_75t_R _28032_ (.A1(_08148_),
    .A2(_05099_),
    .B(_08151_),
    .Y(_02791_));
 INVx1_ASAP7_75t_R _28033_ (.A(_05101_),
    .Y(_08152_));
 OR3x1_ASAP7_75t_R _28034_ (.A(_08152_),
    .B(_05095_),
    .C(_02317_),
    .Y(_08153_));
 AO21x1_ASAP7_75t_R _28035_ (.A1(_08141_),
    .A2(_08153_),
    .B(_05099_),
    .Y(_08154_));
 INVx2_ASAP7_75t_R _28036_ (.A(_05100_),
    .Y(_08155_));
 INVx1_ASAP7_75t_R _28037_ (.A(_02317_),
    .Y(_08156_));
 AND3x1_ASAP7_75t_R _28038_ (.A(_05101_),
    .B(_05094_),
    .C(_08156_),
    .Y(_08157_));
 AND4x1_ASAP7_75t_R _28039_ (.A(_08155_),
    .B(_05132_),
    .C(_08141_),
    .D(_08157_),
    .Y(_08158_));
 AOI21x1_ASAP7_75t_R _28040_ (.A1(_05100_),
    .A2(_08154_),
    .B(_08158_),
    .Y(_02792_));
 NAND2x2_ASAP7_75t_R _28041_ (.A(_05109_),
    .B(_05132_),
    .Y(_08159_));
 BUFx6f_ASAP7_75t_R _28042_ (.A(_08159_),
    .Y(_08160_));
 NAND2x1_ASAP7_75t_R _28043_ (.A(_04861_),
    .B(_05306_),
    .Y(_08161_));
 BUFx4f_ASAP7_75t_R _28044_ (.A(_08161_),
    .Y(_08162_));
 BUFx3_ASAP7_75t_R _28045_ (.A(_08162_),
    .Y(_08163_));
 AND2x2_ASAP7_75t_R _28046_ (.A(_05109_),
    .B(_05132_),
    .Y(_08164_));
 BUFx2_ASAP7_75t_R _28047_ (.A(_08164_),
    .Y(_08165_));
 AND2x2_ASAP7_75t_R _28048_ (.A(_04861_),
    .B(_05306_),
    .Y(_08166_));
 BUFx3_ASAP7_75t_R _28049_ (.A(_08166_),
    .Y(_08167_));
 OR2x2_ASAP7_75t_R _28050_ (.A(_05671_),
    .B(_08167_),
    .Y(_08168_));
 OA211x2_ASAP7_75t_R _28051_ (.A1(_18769_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08168_),
    .Y(_08169_));
 AOI21x1_ASAP7_75t_R _28052_ (.A1(_00106_),
    .A2(_08160_),
    .B(_08169_),
    .Y(_02793_));
 INVx1_ASAP7_75t_R _28053_ (.A(_00116_),
    .Y(_08170_));
 BUFx3_ASAP7_75t_R _28054_ (.A(_08159_),
    .Y(_08171_));
 BUFx3_ASAP7_75t_R _28055_ (.A(_08162_),
    .Y(_08172_));
 BUFx4f_ASAP7_75t_R _28056_ (.A(_08164_),
    .Y(_08173_));
 OR2x2_ASAP7_75t_R _28057_ (.A(_05256_),
    .B(_08167_),
    .Y(_08174_));
 OA211x2_ASAP7_75t_R _28058_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08174_),
    .Y(_08175_));
 AO21x1_ASAP7_75t_R _28059_ (.A1(_08170_),
    .A2(_08171_),
    .B(_08175_),
    .Y(_02794_));
 NAND2x1_ASAP7_75t_R _28060_ (.A(\alu_adder_result_ex[11] ),
    .B(_08167_),
    .Y(_08176_));
 OA211x2_ASAP7_75t_R _28061_ (.A1(_05588_),
    .A2(_08167_),
    .B(_08165_),
    .C(_08176_),
    .Y(_08177_));
 AOI21x1_ASAP7_75t_R _28062_ (.A1(_00115_),
    .A2(_08160_),
    .B(_08177_),
    .Y(_02795_));
 INVx1_ASAP7_75t_R _28063_ (.A(_00118_),
    .Y(_08178_));
 OR2x2_ASAP7_75t_R _28064_ (.A(_05700_),
    .B(_08167_),
    .Y(_08179_));
 OA211x2_ASAP7_75t_R _28065_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08179_),
    .Y(_08180_));
 AO21x1_ASAP7_75t_R _28066_ (.A1(_08178_),
    .A2(_08171_),
    .B(_08180_),
    .Y(_02796_));
 INVx1_ASAP7_75t_R _28067_ (.A(_00117_),
    .Y(_08181_));
 OR2x2_ASAP7_75t_R _28068_ (.A(_05597_),
    .B(_08167_),
    .Y(_08182_));
 OA211x2_ASAP7_75t_R _28069_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08182_),
    .Y(_08183_));
 AO21x1_ASAP7_75t_R _28070_ (.A1(_08181_),
    .A2(_08171_),
    .B(_08183_),
    .Y(_02797_));
 BUFx3_ASAP7_75t_R _28071_ (.A(_08162_),
    .Y(_08184_));
 NAND2x1_ASAP7_75t_R _28072_ (.A(_05603_),
    .B(_08184_),
    .Y(_08185_));
 OA211x2_ASAP7_75t_R _28073_ (.A1(_16028_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08185_),
    .Y(_08186_));
 AOI21x1_ASAP7_75t_R _28074_ (.A1(_00120_),
    .A2(_08160_),
    .B(_08186_),
    .Y(_02798_));
 INVx1_ASAP7_75t_R _28075_ (.A(_00119_),
    .Y(_08187_));
 BUFx3_ASAP7_75t_R _28076_ (.A(_08166_),
    .Y(_08188_));
 OR2x2_ASAP7_75t_R _28077_ (.A(_05300_),
    .B(_08188_),
    .Y(_08189_));
 OA211x2_ASAP7_75t_R _28078_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08189_),
    .Y(_08190_));
 AO21x1_ASAP7_75t_R _28079_ (.A1(_08187_),
    .A2(_08171_),
    .B(_08190_),
    .Y(_02799_));
 INVx1_ASAP7_75t_R _28080_ (.A(_00122_),
    .Y(_08191_));
 OR2x2_ASAP7_75t_R _28081_ (.A(_05169_),
    .B(_08188_),
    .Y(_08192_));
 OA211x2_ASAP7_75t_R _28082_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08192_),
    .Y(_08193_));
 AO21x1_ASAP7_75t_R _28083_ (.A1(_08191_),
    .A2(_08171_),
    .B(_08193_),
    .Y(_02800_));
 AND3x1_ASAP7_75t_R _28084_ (.A(\alu_adder_result_ex[17] ),
    .B(_04861_),
    .C(_05306_),
    .Y(_08194_));
 AO21x1_ASAP7_75t_R _28085_ (.A1(_05189_),
    .A2(_08163_),
    .B(_08194_),
    .Y(_08195_));
 NAND2x1_ASAP7_75t_R _28086_ (.A(_00121_),
    .B(_08159_),
    .Y(_08196_));
 OA21x2_ASAP7_75t_R _28087_ (.A1(_08171_),
    .A2(_08195_),
    .B(_08196_),
    .Y(_02801_));
 NAND2x1_ASAP7_75t_R _28088_ (.A(_05715_),
    .B(_08162_),
    .Y(_08197_));
 OA211x2_ASAP7_75t_R _28089_ (.A1(_16531_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08197_),
    .Y(_08198_));
 AOI21x1_ASAP7_75t_R _28090_ (.A1(_00124_),
    .A2(_08160_),
    .B(_08198_),
    .Y(_02802_));
 INVx1_ASAP7_75t_R _28091_ (.A(_00123_),
    .Y(_08199_));
 OR2x2_ASAP7_75t_R _28092_ (.A(_05621_),
    .B(_08188_),
    .Y(_08200_));
 OA211x2_ASAP7_75t_R _28093_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08200_),
    .Y(_08201_));
 AO21x1_ASAP7_75t_R _28094_ (.A1(_08199_),
    .A2(_08171_),
    .B(_08201_),
    .Y(_02803_));
 INVx1_ASAP7_75t_R _28095_ (.A(_00105_),
    .Y(_08202_));
 OR2x2_ASAP7_75t_R _28096_ (.A(_05531_),
    .B(_08188_),
    .Y(_08203_));
 OA211x2_ASAP7_75t_R _28097_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08203_),
    .Y(_08204_));
 AO21x1_ASAP7_75t_R _28098_ (.A1(_08202_),
    .A2(_08171_),
    .B(_08204_),
    .Y(_02804_));
 INVx1_ASAP7_75t_R _28099_ (.A(_00126_),
    .Y(_08205_));
 BUFx3_ASAP7_75t_R _28100_ (.A(_08159_),
    .Y(_08206_));
 OR2x2_ASAP7_75t_R _28101_ (.A(_05631_),
    .B(_08188_),
    .Y(_08207_));
 OA211x2_ASAP7_75t_R _28102_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_08172_),
    .B(_08173_),
    .C(_08207_),
    .Y(_08208_));
 AO21x1_ASAP7_75t_R _28103_ (.A1(_08205_),
    .A2(_08206_),
    .B(_08208_),
    .Y(_02805_));
 AND2x2_ASAP7_75t_R _28104_ (.A(_05217_),
    .B(_08162_),
    .Y(_08209_));
 AO21x1_ASAP7_75t_R _28105_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_08167_),
    .B(_08209_),
    .Y(_08210_));
 NAND2x1_ASAP7_75t_R _28106_ (.A(_00125_),
    .B(_08159_),
    .Y(_08211_));
 OA21x2_ASAP7_75t_R _28107_ (.A1(_08171_),
    .A2(_08210_),
    .B(_08211_),
    .Y(_02806_));
 INVx1_ASAP7_75t_R _28108_ (.A(_00128_),
    .Y(_08212_));
 BUFx2_ASAP7_75t_R _28109_ (.A(_08164_),
    .Y(_08213_));
 OR2x2_ASAP7_75t_R _28110_ (.A(_05225_),
    .B(_08188_),
    .Y(_08214_));
 OA211x2_ASAP7_75t_R _28111_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_08172_),
    .B(_08213_),
    .C(_08214_),
    .Y(_08215_));
 AO21x1_ASAP7_75t_R _28112_ (.A1(_08212_),
    .A2(_08206_),
    .B(_08215_),
    .Y(_02807_));
 INVx1_ASAP7_75t_R _28113_ (.A(_00127_),
    .Y(_08216_));
 OR2x2_ASAP7_75t_R _28114_ (.A(_05234_),
    .B(_08188_),
    .Y(_08217_));
 OA211x2_ASAP7_75t_R _28115_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08217_),
    .Y(_08218_));
 AO21x1_ASAP7_75t_R _28116_ (.A1(_08216_),
    .A2(_08206_),
    .B(_08218_),
    .Y(_02808_));
 NAND2x1_ASAP7_75t_R _28117_ (.A(_05241_),
    .B(_08162_),
    .Y(_08219_));
 OA211x2_ASAP7_75t_R _28118_ (.A1(_17257_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08219_),
    .Y(_08220_));
 AOI21x1_ASAP7_75t_R _28119_ (.A1(_00130_),
    .A2(_08160_),
    .B(_08220_),
    .Y(_02809_));
 INVx1_ASAP7_75t_R _28120_ (.A(_00129_),
    .Y(_08221_));
 OR2x2_ASAP7_75t_R _28121_ (.A(_05249_),
    .B(_08188_),
    .Y(_08222_));
 OA211x2_ASAP7_75t_R _28122_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08222_),
    .Y(_08223_));
 AO21x1_ASAP7_75t_R _28123_ (.A1(_08221_),
    .A2(_08206_),
    .B(_08223_),
    .Y(_02810_));
 OR2x2_ASAP7_75t_R _28124_ (.A(_05649_),
    .B(_08167_),
    .Y(_08224_));
 OA211x2_ASAP7_75t_R _28125_ (.A1(_04414_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08224_),
    .Y(_08225_));
 AOI21x1_ASAP7_75t_R _28126_ (.A1(_00132_),
    .A2(_08160_),
    .B(_08225_),
    .Y(_02811_));
 INVx1_ASAP7_75t_R _28127_ (.A(_00131_),
    .Y(_08226_));
 OR2x2_ASAP7_75t_R _28128_ (.A(_05265_),
    .B(_08188_),
    .Y(_08227_));
 OA211x2_ASAP7_75t_R _28129_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08227_),
    .Y(_08228_));
 AO21x1_ASAP7_75t_R _28130_ (.A1(_08226_),
    .A2(_08206_),
    .B(_08228_),
    .Y(_02812_));
 INVx1_ASAP7_75t_R _28131_ (.A(_00134_),
    .Y(_08229_));
 OR2x2_ASAP7_75t_R _28132_ (.A(_05273_),
    .B(_08188_),
    .Y(_08230_));
 OA211x2_ASAP7_75t_R _28133_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08230_),
    .Y(_08231_));
 AO21x1_ASAP7_75t_R _28134_ (.A1(_08229_),
    .A2(_08206_),
    .B(_08231_),
    .Y(_02813_));
 INVx1_ASAP7_75t_R _28135_ (.A(_00133_),
    .Y(_08232_));
 OR2x2_ASAP7_75t_R _28136_ (.A(_05281_),
    .B(_08166_),
    .Y(_08233_));
 OA211x2_ASAP7_75t_R _28137_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08233_),
    .Y(_08234_));
 AO21x1_ASAP7_75t_R _28138_ (.A1(_08232_),
    .A2(_08206_),
    .B(_08234_),
    .Y(_02814_));
 INVx1_ASAP7_75t_R _28139_ (.A(_00108_),
    .Y(_08235_));
 OR2x2_ASAP7_75t_R _28140_ (.A(_05196_),
    .B(_08166_),
    .Y(_08236_));
 OA211x2_ASAP7_75t_R _28141_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08236_),
    .Y(_08237_));
 AO21x1_ASAP7_75t_R _28142_ (.A1(_08235_),
    .A2(_08206_),
    .B(_08237_),
    .Y(_02815_));
 NAND2x1_ASAP7_75t_R _28143_ (.A(_05289_),
    .B(_08162_),
    .Y(_08238_));
 OA211x2_ASAP7_75t_R _28144_ (.A1(_04917_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08238_),
    .Y(_08239_));
 AOI21x1_ASAP7_75t_R _28145_ (.A1(_00136_),
    .A2(_08160_),
    .B(_08239_),
    .Y(_02816_));
 INVx1_ASAP7_75t_R _28146_ (.A(_00135_),
    .Y(_08240_));
 OA211x2_ASAP7_75t_R _28147_ (.A1(\alu_adder_result_ex[31] ),
    .A2(_05310_),
    .B(_08213_),
    .C(_04861_),
    .Y(_08241_));
 AO21x1_ASAP7_75t_R _28148_ (.A1(_08240_),
    .A2(_08206_),
    .B(_08241_),
    .Y(_02817_));
 NAND2x1_ASAP7_75t_R _28149_ (.A(_05204_),
    .B(_08162_),
    .Y(_08242_));
 OA211x2_ASAP7_75t_R _28150_ (.A1(_05461_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08242_),
    .Y(_08243_));
 AOI21x1_ASAP7_75t_R _28151_ (.A1(_00107_),
    .A2(_08160_),
    .B(_08243_),
    .Y(_02818_));
 INVx1_ASAP7_75t_R _28152_ (.A(_00110_),
    .Y(_08244_));
 OR2x2_ASAP7_75t_R _28153_ (.A(_05210_),
    .B(_08166_),
    .Y(_08245_));
 OA211x2_ASAP7_75t_R _28154_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08245_),
    .Y(_08246_));
 AO21x1_ASAP7_75t_R _28155_ (.A1(_08244_),
    .A2(_08206_),
    .B(_08246_),
    .Y(_02819_));
 INVx1_ASAP7_75t_R _28156_ (.A(_00109_),
    .Y(_08247_));
 OR2x2_ASAP7_75t_R _28157_ (.A(_05553_),
    .B(_08166_),
    .Y(_08248_));
 OA211x2_ASAP7_75t_R _28158_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_08184_),
    .B(_08213_),
    .C(_08248_),
    .Y(_08249_));
 AO21x1_ASAP7_75t_R _28159_ (.A1(_08247_),
    .A2(_08159_),
    .B(_08249_),
    .Y(_02820_));
 OR2x2_ASAP7_75t_R _28160_ (.A(_05559_),
    .B(_08167_),
    .Y(_08250_));
 OA211x2_ASAP7_75t_R _28161_ (.A1(_15272_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08250_),
    .Y(_08251_));
 AOI21x1_ASAP7_75t_R _28162_ (.A1(_00112_),
    .A2(_08160_),
    .B(_08251_),
    .Y(_02821_));
 NAND2x1_ASAP7_75t_R _28163_ (.A(_05568_),
    .B(_08162_),
    .Y(_08252_));
 OA211x2_ASAP7_75t_R _28164_ (.A1(_15247_),
    .A2(_08163_),
    .B(_08165_),
    .C(_08252_),
    .Y(_08253_));
 AOI21x1_ASAP7_75t_R _28165_ (.A1(_00111_),
    .A2(_08160_),
    .B(_08253_),
    .Y(_02822_));
 OR2x2_ASAP7_75t_R _28166_ (.A(_05692_),
    .B(_08167_),
    .Y(_08254_));
 OA211x2_ASAP7_75t_R _28167_ (.A1(_15417_),
    .A2(_08172_),
    .B(_08173_),
    .C(_08254_),
    .Y(_08255_));
 AOI21x1_ASAP7_75t_R _28168_ (.A1(_00114_),
    .A2(_08171_),
    .B(_08255_),
    .Y(_02823_));
 INVx1_ASAP7_75t_R _28169_ (.A(_00113_),
    .Y(_08256_));
 NAND2x1_ASAP7_75t_R _28170_ (.A(_05577_),
    .B(_08162_),
    .Y(_08257_));
 OA211x2_ASAP7_75t_R _28171_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_08184_),
    .B(_08164_),
    .C(_08257_),
    .Y(_08258_));
 AO21x1_ASAP7_75t_R _28172_ (.A1(_08256_),
    .A2(_08159_),
    .B(_08258_),
    .Y(_02824_));
 BUFx3_ASAP7_75t_R _28173_ (.A(_00068_),
    .Y(_08259_));
 NAND2x2_ASAP7_75t_R _28174_ (.A(_05091_),
    .B(_05132_),
    .Y(_08260_));
 BUFx3_ASAP7_75t_R _28175_ (.A(_08260_),
    .Y(_08261_));
 AO31x2_ASAP7_75t_R _28176_ (.A1(_01751_),
    .A2(_04898_),
    .A3(_04908_),
    .B(_04869_),
    .Y(_08262_));
 AO21x2_ASAP7_75t_R _28177_ (.A1(_04898_),
    .A2(_04908_),
    .B(_01751_),
    .Y(_08263_));
 AND2x4_ASAP7_75t_R _28178_ (.A(_08262_),
    .B(_08263_),
    .Y(_08264_));
 NAND2x2_ASAP7_75t_R _28179_ (.A(_08148_),
    .B(_08264_),
    .Y(_08265_));
 OR4x1_ASAP7_75t_R _28180_ (.A(_08259_),
    .B(_05103_),
    .C(_08261_),
    .D(_08265_),
    .Y(_08266_));
 AND3x1_ASAP7_75t_R _28181_ (.A(_05109_),
    .B(_05159_),
    .C(_05132_),
    .Y(_08267_));
 BUFx6f_ASAP7_75t_R _28182_ (.A(_08267_),
    .Y(_08268_));
 BUFx6f_ASAP7_75t_R _28183_ (.A(_08268_),
    .Y(_08269_));
 AOI21x1_ASAP7_75t_R _28184_ (.A1(_00071_),
    .A2(_08266_),
    .B(_08269_),
    .Y(_02825_));
 BUFx4f_ASAP7_75t_R _28185_ (.A(_00074_),
    .Y(_08270_));
 NAND2x2_ASAP7_75t_R _28186_ (.A(_08262_),
    .B(_08263_),
    .Y(_08271_));
 BUFx4f_ASAP7_75t_R _28187_ (.A(_08271_),
    .Y(_08272_));
 BUFx4f_ASAP7_75t_R _28188_ (.A(_08272_),
    .Y(_08273_));
 OR5x1_ASAP7_75t_R _28189_ (.A(_08148_),
    .B(_08270_),
    .C(_05103_),
    .D(_08260_),
    .E(_08273_),
    .Y(_08274_));
 AOI21x1_ASAP7_75t_R _28190_ (.A1(_00082_),
    .A2(_08274_),
    .B(_08269_),
    .Y(_02826_));
 BUFx4f_ASAP7_75t_R _28191_ (.A(_00067_),
    .Y(_08275_));
 OR5x1_ASAP7_75t_R _28192_ (.A(_08148_),
    .B(_08275_),
    .C(_05103_),
    .D(_08260_),
    .E(_08273_),
    .Y(_08276_));
 AOI21x1_ASAP7_75t_R _28193_ (.A1(_00083_),
    .A2(_08276_),
    .B(_08269_),
    .Y(_02827_));
 BUFx3_ASAP7_75t_R _28194_ (.A(_08260_),
    .Y(_08277_));
 OR4x2_ASAP7_75t_R _28195_ (.A(_08155_),
    .B(_05101_),
    .C(_05094_),
    .D(_08271_),
    .Y(_08278_));
 OR3x1_ASAP7_75t_R _28196_ (.A(_08259_),
    .B(_08277_),
    .C(_08278_),
    .Y(_08279_));
 AOI21x1_ASAP7_75t_R _28197_ (.A1(_00084_),
    .A2(_08279_),
    .B(_08269_),
    .Y(_02828_));
 OR3x1_ASAP7_75t_R _28198_ (.A(_05093_),
    .B(_08277_),
    .C(_08278_),
    .Y(_08280_));
 AOI21x1_ASAP7_75t_R _28199_ (.A1(_00085_),
    .A2(_08280_),
    .B(_08269_),
    .Y(_02829_));
 OR3x1_ASAP7_75t_R _28200_ (.A(_08270_),
    .B(_08277_),
    .C(_08278_),
    .Y(_08281_));
 AOI21x1_ASAP7_75t_R _28201_ (.A1(_00086_),
    .A2(_08281_),
    .B(_08269_),
    .Y(_02830_));
 OR3x1_ASAP7_75t_R _28202_ (.A(_08275_),
    .B(_08277_),
    .C(_08278_),
    .Y(_08282_));
 AOI21x1_ASAP7_75t_R _28203_ (.A1(_00087_),
    .A2(_08282_),
    .B(_08269_),
    .Y(_02831_));
 AND2x2_ASAP7_75t_R _28204_ (.A(_05091_),
    .B(_05132_),
    .Y(_08283_));
 INVx1_ASAP7_75t_R _28205_ (.A(_00068_),
    .Y(_08284_));
 AND3x2_ASAP7_75t_R _28206_ (.A(_05094_),
    .B(_08284_),
    .C(_08264_),
    .Y(_08285_));
 AND2x4_ASAP7_75t_R _28207_ (.A(_08155_),
    .B(_05101_),
    .Y(_08286_));
 NAND2x2_ASAP7_75t_R _28208_ (.A(_08173_),
    .B(_08260_),
    .Y(_08287_));
 INVx1_ASAP7_75t_R _28209_ (.A(_00088_),
    .Y(_08288_));
 AO32x1_ASAP7_75t_R _28210_ (.A1(_08283_),
    .A2(_08285_),
    .A3(_08286_),
    .B1(_08287_),
    .B2(_08288_),
    .Y(_02832_));
 INVx1_ASAP7_75t_R _28211_ (.A(_01458_),
    .Y(_08289_));
 AND3x2_ASAP7_75t_R _28212_ (.A(_08289_),
    .B(_08148_),
    .C(_08264_),
    .Y(_08290_));
 INVx1_ASAP7_75t_R _28213_ (.A(_00089_),
    .Y(_08291_));
 AO32x1_ASAP7_75t_R _28214_ (.A1(_08283_),
    .A2(_08286_),
    .A3(_08290_),
    .B1(_08287_),
    .B2(_08291_),
    .Y(_02833_));
 INVx1_ASAP7_75t_R _28215_ (.A(_00074_),
    .Y(_08292_));
 AND3x4_ASAP7_75t_R _28216_ (.A(_05094_),
    .B(_08292_),
    .C(_08264_),
    .Y(_08293_));
 INVx1_ASAP7_75t_R _28217_ (.A(_00090_),
    .Y(_08294_));
 AO32x1_ASAP7_75t_R _28218_ (.A1(_08283_),
    .A2(_08286_),
    .A3(_08293_),
    .B1(_08287_),
    .B2(_08294_),
    .Y(_02834_));
 INVx1_ASAP7_75t_R _28219_ (.A(_00067_),
    .Y(_08295_));
 AND3x2_ASAP7_75t_R _28220_ (.A(_05094_),
    .B(_08295_),
    .C(_08264_),
    .Y(_08296_));
 INVx1_ASAP7_75t_R _28221_ (.A(_00091_),
    .Y(_08297_));
 AO32x1_ASAP7_75t_R _28222_ (.A1(_08283_),
    .A2(_08286_),
    .A3(_08296_),
    .B1(_08287_),
    .B2(_08297_),
    .Y(_02835_));
 BUFx4f_ASAP7_75t_R _28223_ (.A(_08271_),
    .Y(_08298_));
 OR4x1_ASAP7_75t_R _28224_ (.A(_01458_),
    .B(_05095_),
    .C(_05102_),
    .D(_08298_),
    .Y(_08299_));
 OR2x2_ASAP7_75t_R _28225_ (.A(_08261_),
    .B(_08299_),
    .Y(_08300_));
 AOI21x1_ASAP7_75t_R _28226_ (.A1(_00072_),
    .A2(_08300_),
    .B(_08269_),
    .Y(_02836_));
 OR2x4_ASAP7_75t_R _28227_ (.A(_05100_),
    .B(_05101_),
    .Y(_08301_));
 OR4x1_ASAP7_75t_R _28228_ (.A(_08259_),
    .B(_08261_),
    .C(_08265_),
    .D(_08301_),
    .Y(_08302_));
 AOI21x1_ASAP7_75t_R _28229_ (.A1(_00092_),
    .A2(_08302_),
    .B(_08269_),
    .Y(_02837_));
 OR4x1_ASAP7_75t_R _28230_ (.A(_05093_),
    .B(_08261_),
    .C(_08265_),
    .D(_08301_),
    .Y(_08303_));
 AOI21x1_ASAP7_75t_R _28231_ (.A1(_00093_),
    .A2(_08303_),
    .B(_08269_),
    .Y(_02838_));
 OR4x1_ASAP7_75t_R _28232_ (.A(_08270_),
    .B(_08261_),
    .C(_08265_),
    .D(_08301_),
    .Y(_08304_));
 BUFx6f_ASAP7_75t_R _28233_ (.A(_08268_),
    .Y(_08305_));
 AOI21x1_ASAP7_75t_R _28234_ (.A1(_00094_),
    .A2(_08304_),
    .B(_08305_),
    .Y(_02839_));
 OR4x1_ASAP7_75t_R _28235_ (.A(_08275_),
    .B(_08261_),
    .C(_08265_),
    .D(_08301_),
    .Y(_08306_));
 AOI21x1_ASAP7_75t_R _28236_ (.A1(_00095_),
    .A2(_08306_),
    .B(_08305_),
    .Y(_02840_));
 OR4x2_ASAP7_75t_R _28237_ (.A(_05100_),
    .B(_08152_),
    .C(_05094_),
    .D(_08271_),
    .Y(_08307_));
 OR3x1_ASAP7_75t_R _28238_ (.A(_08259_),
    .B(_08277_),
    .C(_08307_),
    .Y(_08308_));
 AOI21x1_ASAP7_75t_R _28239_ (.A1(_00096_),
    .A2(_08308_),
    .B(_08305_),
    .Y(_02841_));
 OR3x1_ASAP7_75t_R _28240_ (.A(_05093_),
    .B(_08277_),
    .C(_08307_),
    .Y(_08309_));
 AOI21x1_ASAP7_75t_R _28241_ (.A1(_00097_),
    .A2(_08309_),
    .B(_08305_),
    .Y(_02842_));
 OR3x1_ASAP7_75t_R _28242_ (.A(_08270_),
    .B(_08277_),
    .C(_08307_),
    .Y(_08310_));
 AOI21x1_ASAP7_75t_R _28243_ (.A1(_00098_),
    .A2(_08310_),
    .B(_08305_),
    .Y(_02843_));
 OR3x1_ASAP7_75t_R _28244_ (.A(_08275_),
    .B(_08277_),
    .C(_08307_),
    .Y(_08311_));
 AOI21x1_ASAP7_75t_R _28245_ (.A1(_00099_),
    .A2(_08311_),
    .B(_08305_),
    .Y(_02844_));
 OR3x4_ASAP7_75t_R _28246_ (.A(_05094_),
    .B(_08298_),
    .C(_08301_),
    .Y(_08312_));
 OR3x1_ASAP7_75t_R _28247_ (.A(_08259_),
    .B(_08277_),
    .C(_08312_),
    .Y(_08313_));
 AOI21x1_ASAP7_75t_R _28248_ (.A1(_00100_),
    .A2(_08313_),
    .B(_08305_),
    .Y(_02845_));
 OR3x1_ASAP7_75t_R _28249_ (.A(_05093_),
    .B(_08277_),
    .C(_08312_),
    .Y(_08314_));
 AOI21x1_ASAP7_75t_R _28250_ (.A1(_00101_),
    .A2(_08314_),
    .B(_08305_),
    .Y(_02846_));
 OR4x1_ASAP7_75t_R _28251_ (.A(_08270_),
    .B(_05103_),
    .C(_08261_),
    .D(_08265_),
    .Y(_08315_));
 AOI21x1_ASAP7_75t_R _28252_ (.A1(_00073_),
    .A2(_08315_),
    .B(_08305_),
    .Y(_02847_));
 OR3x1_ASAP7_75t_R _28253_ (.A(_08270_),
    .B(_08261_),
    .C(_08312_),
    .Y(_08316_));
 AOI21x1_ASAP7_75t_R _28254_ (.A1(_00102_),
    .A2(_08316_),
    .B(_08305_),
    .Y(_02848_));
 OR3x1_ASAP7_75t_R _28255_ (.A(_08275_),
    .B(_08261_),
    .C(_08312_),
    .Y(_08317_));
 AOI21x1_ASAP7_75t_R _28256_ (.A1(_00103_),
    .A2(_08317_),
    .B(_08268_),
    .Y(_02849_));
 OR4x1_ASAP7_75t_R _28257_ (.A(_08275_),
    .B(_05103_),
    .C(_08260_),
    .D(_08265_),
    .Y(_08318_));
 AOI21x1_ASAP7_75t_R _28258_ (.A1(_00075_),
    .A2(_08318_),
    .B(_08268_),
    .Y(_02850_));
 AND2x2_ASAP7_75t_R _28259_ (.A(_05100_),
    .B(_08152_),
    .Y(_08319_));
 NAND2x1_ASAP7_75t_R _28260_ (.A(_08283_),
    .B(_08319_),
    .Y(_08320_));
 OR3x1_ASAP7_75t_R _28261_ (.A(_08259_),
    .B(_08265_),
    .C(_08320_),
    .Y(_08321_));
 AOI21x1_ASAP7_75t_R _28262_ (.A1(_00076_),
    .A2(_08321_),
    .B(_08268_),
    .Y(_02851_));
 OR3x1_ASAP7_75t_R _28263_ (.A(_05093_),
    .B(_08265_),
    .C(_08320_),
    .Y(_08322_));
 AOI21x1_ASAP7_75t_R _28264_ (.A1(_00077_),
    .A2(_08322_),
    .B(_08268_),
    .Y(_02852_));
 INVx1_ASAP7_75t_R _28265_ (.A(_00078_),
    .Y(_08323_));
 AND3x1_ASAP7_75t_R _28266_ (.A(_08283_),
    .B(_08319_),
    .C(_08293_),
    .Y(_08324_));
 OA21x2_ASAP7_75t_R _28267_ (.A1(_08323_),
    .A2(_08324_),
    .B(_08287_),
    .Y(_02853_));
 OR3x1_ASAP7_75t_R _28268_ (.A(_08275_),
    .B(_08265_),
    .C(_08320_),
    .Y(_08325_));
 AOI21x1_ASAP7_75t_R _28269_ (.A1(_00079_),
    .A2(_08325_),
    .B(_08268_),
    .Y(_02854_));
 OR5x1_ASAP7_75t_R _28270_ (.A(_08148_),
    .B(_08259_),
    .C(_05103_),
    .D(_08260_),
    .E(_08273_),
    .Y(_08326_));
 AOI21x1_ASAP7_75t_R _28271_ (.A1(_00080_),
    .A2(_08326_),
    .B(_08268_),
    .Y(_02855_));
 OR4x1_ASAP7_75t_R _28272_ (.A(_01458_),
    .B(_08148_),
    .C(_05103_),
    .D(_08272_),
    .Y(_08327_));
 OA21x2_ASAP7_75t_R _28273_ (.A1(_08261_),
    .A2(_08327_),
    .B(_00081_),
    .Y(_08328_));
 NOR2x1_ASAP7_75t_R _28274_ (.A(_08268_),
    .B(_08328_),
    .Y(_02856_));
 OR2x2_ASAP7_75t_R _28275_ (.A(_05497_),
    .B(net106),
    .Y(_02857_));
 BUFx4f_ASAP7_75t_R _28276_ (.A(_14726_),
    .Y(_08329_));
 BUFx3_ASAP7_75t_R _28277_ (.A(_13438_),
    .Y(_08330_));
 AND2x2_ASAP7_75t_R _28278_ (.A(_04920_),
    .B(_01508_),
    .Y(_08331_));
 NAND2x2_ASAP7_75t_R _28279_ (.A(_13648_),
    .B(_13774_),
    .Y(_08332_));
 AO33x2_ASAP7_75t_R _28280_ (.A1(_13554_),
    .A2(_13383_),
    .A3(_13377_),
    .B1(_13621_),
    .B2(_13371_),
    .B3(_14880_),
    .Y(_08333_));
 NAND2x1_ASAP7_75t_R _28281_ (.A(_13422_),
    .B(_08333_),
    .Y(_08334_));
 AO21x1_ASAP7_75t_R _28282_ (.A1(_08332_),
    .A2(_08334_),
    .B(_06785_),
    .Y(_08335_));
 INVx1_ASAP7_75t_R _28283_ (.A(_08335_),
    .Y(_08336_));
 AO33x2_ASAP7_75t_R _28284_ (.A1(_01454_),
    .A2(_08331_),
    .A3(_04923_),
    .B1(_05097_),
    .B2(_06833_),
    .B3(_08336_),
    .Y(_08337_));
 BUFx3_ASAP7_75t_R _28285_ (.A(_08337_),
    .Y(_08338_));
 BUFx4f_ASAP7_75t_R _28286_ (.A(_08338_),
    .Y(_08339_));
 AND3x1_ASAP7_75t_R _28287_ (.A(_08329_),
    .B(_08330_),
    .C(_08339_),
    .Y(_08340_));
 BUFx10_ASAP7_75t_R _28288_ (.A(_08340_),
    .Y(_08341_));
 NAND2x2_ASAP7_75t_R _28289_ (.A(_14051_),
    .B(_08341_),
    .Y(_08342_));
 OA21x2_ASAP7_75t_R _28290_ (.A1(_05058_),
    .A2(_06832_),
    .B(_14071_),
    .Y(_08343_));
 OR3x4_ASAP7_75t_R _28291_ (.A(_05143_),
    .B(_08343_),
    .C(_08335_),
    .Y(_08344_));
 BUFx6f_ASAP7_75t_R _28292_ (.A(_08344_),
    .Y(_08345_));
 AO21x1_ASAP7_75t_R _28293_ (.A1(_05078_),
    .A2(_05839_),
    .B(_08345_),
    .Y(_08346_));
 AOI211x1_ASAP7_75t_R _28294_ (.A1(_05135_),
    .A2(_05136_),
    .B(_06811_),
    .C(_14904_),
    .Y(_08347_));
 NOR2x1_ASAP7_75t_R _28295_ (.A(\alu_adder_result_ex[28] ),
    .B(_06824_),
    .Y(_08348_));
 NOR2x1_ASAP7_75t_R _28296_ (.A(_06808_),
    .B(_06822_),
    .Y(_08349_));
 AO21x1_ASAP7_75t_R _28297_ (.A1(_05136_),
    .A2(_08348_),
    .B(_08349_),
    .Y(_08350_));
 NOR2x1_ASAP7_75t_R _28298_ (.A(_08347_),
    .B(_08350_),
    .Y(_08351_));
 BUFx4f_ASAP7_75t_R _28299_ (.A(_06793_),
    .Y(_08352_));
 NOR2x1_ASAP7_75t_R _28300_ (.A(_08352_),
    .B(_06813_),
    .Y(_08353_));
 AO21x1_ASAP7_75t_R _28301_ (.A1(_14904_),
    .A2(_08352_),
    .B(_08353_),
    .Y(_08354_));
 AO221x1_ASAP7_75t_R _28302_ (.A1(_02295_),
    .A2(_14912_),
    .B1(_08354_),
    .B2(net1996),
    .C(_06798_),
    .Y(_08355_));
 OA21x2_ASAP7_75t_R _28303_ (.A1(_08352_),
    .A2(_06812_),
    .B(_08355_),
    .Y(_08356_));
 OR4x2_ASAP7_75t_R _28304_ (.A(_13571_),
    .B(_14915_),
    .C(_14917_),
    .D(_14918_),
    .Y(_08357_));
 NOR2x1_ASAP7_75t_R _28305_ (.A(_14912_),
    .B(_08357_),
    .Y(_08358_));
 OA211x2_ASAP7_75t_R _28306_ (.A1(_15251_),
    .A2(_06810_),
    .B(_06793_),
    .C(_08358_),
    .Y(_08359_));
 BUFx4f_ASAP7_75t_R _28307_ (.A(_08359_),
    .Y(_08360_));
 AND2x2_ASAP7_75t_R _28308_ (.A(net1995),
    .B(_02295_),
    .Y(_08361_));
 NOR3x1_ASAP7_75t_R _28309_ (.A(_08352_),
    .B(_08357_),
    .C(_08361_),
    .Y(_08362_));
 INVx1_ASAP7_75t_R _28310_ (.A(_06794_),
    .Y(_08363_));
 AND3x2_ASAP7_75t_R _28311_ (.A(_08363_),
    .B(_13636_),
    .C(_14912_),
    .Y(_08364_));
 BUFx3_ASAP7_75t_R _28312_ (.A(_08364_),
    .Y(_08365_));
 BUFx4f_ASAP7_75t_R _28313_ (.A(_08365_),
    .Y(_08366_));
 AND2x2_ASAP7_75t_R _28314_ (.A(_13636_),
    .B(_14898_),
    .Y(_08367_));
 OR3x1_ASAP7_75t_R _28315_ (.A(_15251_),
    .B(_06800_),
    .C(_06810_),
    .Y(_08368_));
 AND3x1_ASAP7_75t_R _28316_ (.A(_14912_),
    .B(_08367_),
    .C(_08368_),
    .Y(_08369_));
 OR4x1_ASAP7_75t_R _28317_ (.A(_08360_),
    .B(_08362_),
    .C(_08366_),
    .D(_08369_),
    .Y(_08370_));
 NAND2x1_ASAP7_75t_R _28318_ (.A(_02296_),
    .B(_08352_),
    .Y(_08371_));
 OA21x2_ASAP7_75t_R _28319_ (.A1(_15251_),
    .A2(_08352_),
    .B(_08371_),
    .Y(_08372_));
 OA21x2_ASAP7_75t_R _28320_ (.A1(_08363_),
    .A2(_08372_),
    .B(_08358_),
    .Y(_08373_));
 NOR2x1_ASAP7_75t_R _28321_ (.A(_08370_),
    .B(_08373_),
    .Y(_08374_));
 AOI21x1_ASAP7_75t_R _28322_ (.A1(_08356_),
    .A2(_08374_),
    .B(_05304_),
    .Y(_08375_));
 BUFx4f_ASAP7_75t_R _28323_ (.A(_08375_),
    .Y(_08376_));
 BUFx6f_ASAP7_75t_R _28324_ (.A(_08376_),
    .Y(_08377_));
 NOR2x1_ASAP7_75t_R _28325_ (.A(_06794_),
    .B(_08352_),
    .Y(_08378_));
 AO21x1_ASAP7_75t_R _28326_ (.A1(_08352_),
    .A2(_06814_),
    .B(_08378_),
    .Y(_08379_));
 AND2x6_ASAP7_75t_R _28327_ (.A(_08367_),
    .B(_08379_),
    .Y(_08380_));
 INVx4_ASAP7_75t_R _28328_ (.A(_08380_),
    .Y(_08381_));
 BUFx4f_ASAP7_75t_R _28329_ (.A(_08381_),
    .Y(_08382_));
 OR3x1_ASAP7_75t_R _28330_ (.A(_08352_),
    .B(_08357_),
    .C(_08361_),
    .Y(_08383_));
 BUFx3_ASAP7_75t_R _28331_ (.A(_08383_),
    .Y(_08384_));
 BUFx6f_ASAP7_75t_R _28332_ (.A(_08384_),
    .Y(_08385_));
 OR5x1_ASAP7_75t_R _28333_ (.A(_06794_),
    .B(_15248_),
    .C(_14912_),
    .D(_14913_),
    .E(_06790_),
    .Y(_08386_));
 OA21x2_ASAP7_75t_R _28334_ (.A1(_00406_),
    .A2(_08352_),
    .B(_08386_),
    .Y(_08387_));
 OR3x1_ASAP7_75t_R _28335_ (.A(_08357_),
    .B(_08362_),
    .C(_08387_),
    .Y(_08388_));
 BUFx3_ASAP7_75t_R _28336_ (.A(_08388_),
    .Y(_08389_));
 BUFx6f_ASAP7_75t_R _28337_ (.A(_08389_),
    .Y(_08390_));
 OAI22x1_ASAP7_75t_R _28338_ (.A1(_02252_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_02253_),
    .Y(_08391_));
 AND2x2_ASAP7_75t_R _28339_ (.A(_08382_),
    .B(_08391_),
    .Y(_08392_));
 BUFx4f_ASAP7_75t_R _28340_ (.A(_08360_),
    .Y(_08393_));
 BUFx4f_ASAP7_75t_R _28341_ (.A(_08380_),
    .Y(_08394_));
 BUFx4f_ASAP7_75t_R _28342_ (.A(_08394_),
    .Y(_08395_));
 AO22x1_ASAP7_75t_R _28343_ (.A1(\alu_adder_result_ex[0] ),
    .A2(_08393_),
    .B1(_08395_),
    .B2(_00297_),
    .Y(_08396_));
 AND2x2_ASAP7_75t_R _28344_ (.A(_14149_),
    .B(_14155_),
    .Y(_08397_));
 OR4x2_ASAP7_75t_R _28345_ (.A(_04522_),
    .B(_13553_),
    .C(_13855_),
    .D(_08397_),
    .Y(_08398_));
 OR4x2_ASAP7_75t_R _28346_ (.A(_02251_),
    .B(_14301_),
    .C(_14302_),
    .D(_14305_),
    .Y(_08399_));
 AO21x1_ASAP7_75t_R _28347_ (.A1(_13621_),
    .A2(_08399_),
    .B(_18629_),
    .Y(_08400_));
 BUFx4f_ASAP7_75t_R _28348_ (.A(_08400_),
    .Y(_08401_));
 NAND3x1_ASAP7_75t_R _28349_ (.A(_13621_),
    .B(_18629_),
    .C(_08399_),
    .Y(_08402_));
 BUFx4f_ASAP7_75t_R _28350_ (.A(_08402_),
    .Y(_08403_));
 AO221x2_ASAP7_75t_R _28351_ (.A1(_13621_),
    .A2(_08398_),
    .B1(_08401_),
    .B2(_08403_),
    .C(_18623_),
    .Y(_08404_));
 OR4x2_ASAP7_75t_R _28352_ (.A(_13568_),
    .B(_18625_),
    .C(_06775_),
    .D(_08402_),
    .Y(_08405_));
 OR3x4_ASAP7_75t_R _28353_ (.A(_06794_),
    .B(_13571_),
    .C(_14904_),
    .Y(_08406_));
 BUFx3_ASAP7_75t_R _28354_ (.A(_08406_),
    .Y(_08407_));
 AND3x2_ASAP7_75t_R _28355_ (.A(_06810_),
    .B(_14912_),
    .C(_08367_),
    .Y(_08408_));
 OR3x2_ASAP7_75t_R _28356_ (.A(_04883_),
    .B(_04884_),
    .C(_08364_),
    .Y(_08409_));
 OA211x2_ASAP7_75t_R _28357_ (.A1(_18609_),
    .A2(_08407_),
    .B(_08408_),
    .C(_08409_),
    .Y(_08410_));
 BUFx4f_ASAP7_75t_R _28358_ (.A(_08410_),
    .Y(_08411_));
 AND3x1_ASAP7_75t_R _28359_ (.A(_08404_),
    .B(_08405_),
    .C(_08411_),
    .Y(_08412_));
 AOI221x1_ASAP7_75t_R _28360_ (.A1(_13622_),
    .A2(_08398_),
    .B1(_08401_),
    .B2(_08403_),
    .C(_18623_),
    .Y(_08413_));
 AND3x1_ASAP7_75t_R _28361_ (.A(_13622_),
    .B(_18629_),
    .C(_08399_),
    .Y(_08414_));
 AND4x1_ASAP7_75t_R _28362_ (.A(_13622_),
    .B(_18623_),
    .C(_08398_),
    .D(_08414_),
    .Y(_08415_));
 AND2x2_ASAP7_75t_R _28363_ (.A(_02251_),
    .B(_13621_),
    .Y(_08416_));
 INVx1_ASAP7_75t_R _28364_ (.A(_08416_),
    .Y(_08417_));
 AO31x2_ASAP7_75t_R _28365_ (.A1(_13367_),
    .A2(_04980_),
    .A3(_04981_),
    .B(_08417_),
    .Y(_08418_));
 OR4x2_ASAP7_75t_R _28366_ (.A(_13642_),
    .B(_14301_),
    .C(_14302_),
    .D(_08416_),
    .Y(_08419_));
 AND3x2_ASAP7_75t_R _28367_ (.A(_13361_),
    .B(_13363_),
    .C(_13568_),
    .Y(_08420_));
 NOR2x2_ASAP7_75t_R _28368_ (.A(_00296_),
    .B(_13568_),
    .Y(_08421_));
 AOI221x1_ASAP7_75t_R _28369_ (.A1(_08418_),
    .A2(_08419_),
    .B1(_08420_),
    .B2(_13553_),
    .C(_08421_),
    .Y(_08422_));
 BUFx4f_ASAP7_75t_R _28370_ (.A(_08407_),
    .Y(_08423_));
 OA221x2_ASAP7_75t_R _28371_ (.A1(_18609_),
    .A2(_08423_),
    .B1(_08408_),
    .B2(_18608_),
    .C(_08409_),
    .Y(_08424_));
 AND2x6_ASAP7_75t_R _28372_ (.A(_08418_),
    .B(_08419_),
    .Y(_08425_));
 BUFx4f_ASAP7_75t_R _28373_ (.A(_08425_),
    .Y(_08426_));
 OA22x2_ASAP7_75t_R _28374_ (.A1(_08410_),
    .A2(_08422_),
    .B1(_08424_),
    .B2(_08426_),
    .Y(_08427_));
 OA21x2_ASAP7_75t_R _28375_ (.A1(_08413_),
    .A2(_08415_),
    .B(_08427_),
    .Y(_08428_));
 BUFx4f_ASAP7_75t_R _28376_ (.A(_08366_),
    .Y(_08429_));
 OA21x2_ASAP7_75t_R _28377_ (.A1(_08412_),
    .A2(_08428_),
    .B(_08429_),
    .Y(_08430_));
 OR3x1_ASAP7_75t_R _28378_ (.A(_08392_),
    .B(_08396_),
    .C(_08430_),
    .Y(_08431_));
 AND2x4_ASAP7_75t_R _28379_ (.A(_08401_),
    .B(_08403_),
    .Y(_08432_));
 BUFx4f_ASAP7_75t_R _28380_ (.A(_08432_),
    .Y(_08433_));
 AOI21x1_ASAP7_75t_R _28381_ (.A1(_13553_),
    .A2(_08420_),
    .B(_08421_),
    .Y(_08434_));
 BUFx4f_ASAP7_75t_R _28382_ (.A(_08434_),
    .Y(_08435_));
 AO221x1_ASAP7_75t_R _28383_ (.A1(_15727_),
    .A2(_04522_),
    .B1(_15953_),
    .B2(_15726_),
    .C(_08406_),
    .Y(_08436_));
 OA211x2_ASAP7_75t_R _28384_ (.A1(_18697_),
    .A2(_08365_),
    .B(_08436_),
    .C(_18608_),
    .Y(_08437_));
 AO221x1_ASAP7_75t_R _28385_ (.A1(_16516_),
    .A2(_04522_),
    .B1(_15953_),
    .B2(_16515_),
    .C(_08365_),
    .Y(_08438_));
 OA211x2_ASAP7_75t_R _28386_ (.A1(_18667_),
    .A2(_08407_),
    .B(_08438_),
    .C(_18610_),
    .Y(_08439_));
 OR4x1_ASAP7_75t_R _28387_ (.A(_08425_),
    .B(_08435_),
    .C(_08437_),
    .D(_08439_),
    .Y(_08440_));
 AO221x2_ASAP7_75t_R _28388_ (.A1(_08418_),
    .A2(_08419_),
    .B1(_08420_),
    .B2(_13553_),
    .C(_08421_),
    .Y(_08441_));
 AO221x1_ASAP7_75t_R _28389_ (.A1(_15867_),
    .A2(_04522_),
    .B1(_15953_),
    .B2(_15866_),
    .C(_08406_),
    .Y(_08442_));
 OA211x2_ASAP7_75t_R _28390_ (.A1(_18692_),
    .A2(_08366_),
    .B(_08442_),
    .C(_18610_),
    .Y(_08443_));
 AO221x1_ASAP7_75t_R _28391_ (.A1(_16006_),
    .A2(_04522_),
    .B1(_15953_),
    .B2(_16005_),
    .C(_08406_),
    .Y(_08444_));
 OA211x2_ASAP7_75t_R _28392_ (.A1(_18687_),
    .A2(_08365_),
    .B(_08444_),
    .C(_18608_),
    .Y(_08445_));
 OR3x1_ASAP7_75t_R _28393_ (.A(_08441_),
    .B(_08443_),
    .C(_08445_),
    .Y(_08446_));
 AO21x2_ASAP7_75t_R _28394_ (.A1(_13786_),
    .A2(_13853_),
    .B(_08364_),
    .Y(_08447_));
 NOR3x2_ASAP7_75t_R _28395_ (.B(_13783_),
    .C(_13785_),
    .Y(_08448_),
    .A(_13782_));
 AND3x2_ASAP7_75t_R _28396_ (.A(_13788_),
    .B(_13821_),
    .C(_13852_),
    .Y(_08449_));
 OR3x1_ASAP7_75t_R _28397_ (.A(_08448_),
    .B(_08449_),
    .C(_08364_),
    .Y(_08450_));
 BUFx3_ASAP7_75t_R _28398_ (.A(_08450_),
    .Y(_08451_));
 OA22x2_ASAP7_75t_R _28399_ (.A1(_18725_),
    .A2(_08447_),
    .B1(_08451_),
    .B2(_18717_),
    .Y(_08452_));
 OR3x1_ASAP7_75t_R _28400_ (.A(_08448_),
    .B(_08449_),
    .C(_08406_),
    .Y(_08453_));
 BUFx4f_ASAP7_75t_R _28401_ (.A(_08453_),
    .Y(_08454_));
 AO21x1_ASAP7_75t_R _28402_ (.A1(_13786_),
    .A2(_13853_),
    .B(_08406_),
    .Y(_08455_));
 BUFx4f_ASAP7_75t_R _28403_ (.A(_08455_),
    .Y(_08456_));
 OA22x2_ASAP7_75t_R _28404_ (.A1(_18653_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18647_),
    .Y(_08457_));
 NAND2x2_ASAP7_75t_R _28405_ (.A(_08418_),
    .B(_08419_),
    .Y(_08458_));
 AO211x2_ASAP7_75t_R _28406_ (.A1(_08452_),
    .A2(_08457_),
    .B(_08458_),
    .C(_08435_),
    .Y(_08459_));
 OA22x2_ASAP7_75t_R _28407_ (.A1(_18715_),
    .A2(_08447_),
    .B1(_08451_),
    .B2(_18707_),
    .Y(_08460_));
 OA22x2_ASAP7_75t_R _28408_ (.A1(_18662_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18657_),
    .Y(_08461_));
 AO21x2_ASAP7_75t_R _28409_ (.A1(_13553_),
    .A2(_08420_),
    .B(_08421_),
    .Y(_08462_));
 BUFx4f_ASAP7_75t_R _28410_ (.A(_08462_),
    .Y(_08463_));
 AO211x2_ASAP7_75t_R _28411_ (.A1(_08460_),
    .A2(_08461_),
    .B(_08458_),
    .C(_08463_),
    .Y(_08464_));
 AND4x2_ASAP7_75t_R _28412_ (.A(_08440_),
    .B(_08446_),
    .C(_08459_),
    .D(_08464_),
    .Y(_08465_));
 BUFx4f_ASAP7_75t_R _28413_ (.A(_08434_),
    .Y(_08466_));
 BUFx6f_ASAP7_75t_R _28414_ (.A(_08466_),
    .Y(_08467_));
 BUFx4f_ASAP7_75t_R _28415_ (.A(_08451_),
    .Y(_08468_));
 OR2x2_ASAP7_75t_R _28416_ (.A(_18642_),
    .B(_08447_),
    .Y(_08469_));
 BUFx4f_ASAP7_75t_R _28417_ (.A(_08454_),
    .Y(_08470_));
 OA22x2_ASAP7_75t_R _28418_ (.A1(_18732_),
    .A2(_08470_),
    .B1(_08456_),
    .B2(_18730_),
    .Y(_08471_));
 OA211x2_ASAP7_75t_R _28419_ (.A1(_18637_),
    .A2(_08468_),
    .B(_08469_),
    .C(_08471_),
    .Y(_08472_));
 BUFx4f_ASAP7_75t_R _28420_ (.A(_08447_),
    .Y(_08473_));
 OA22x2_ASAP7_75t_R _28421_ (.A1(_18633_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18630_),
    .Y(_08474_));
 BUFx4f_ASAP7_75t_R _28422_ (.A(_08456_),
    .Y(_08475_));
 OA22x2_ASAP7_75t_R _28423_ (.A1(_18742_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18740_),
    .Y(_08476_));
 BUFx6f_ASAP7_75t_R _28424_ (.A(_08463_),
    .Y(_08477_));
 AO21x1_ASAP7_75t_R _28425_ (.A1(_08474_),
    .A2(_08476_),
    .B(_08477_),
    .Y(_08478_));
 OA21x2_ASAP7_75t_R _28426_ (.A1(_08467_),
    .A2(_08472_),
    .B(_08478_),
    .Y(_08479_));
 NAND2x2_ASAP7_75t_R _28427_ (.A(_08401_),
    .B(_08403_),
    .Y(_08480_));
 BUFx6f_ASAP7_75t_R _28428_ (.A(_08480_),
    .Y(_08481_));
 BUFx4f_ASAP7_75t_R _28429_ (.A(_08425_),
    .Y(_08482_));
 AND2x2_ASAP7_75t_R _28430_ (.A(_08481_),
    .B(_08482_),
    .Y(_08483_));
 AND3x4_ASAP7_75t_R _28431_ (.A(_13786_),
    .B(_13853_),
    .C(_08364_),
    .Y(_08484_));
 OA21x2_ASAP7_75t_R _28432_ (.A1(_08448_),
    .A2(_08449_),
    .B(_08365_),
    .Y(_08485_));
 OA21x2_ASAP7_75t_R _28433_ (.A1(_08448_),
    .A2(_08449_),
    .B(_08407_),
    .Y(_08486_));
 BUFx4f_ASAP7_75t_R _28434_ (.A(_08486_),
    .Y(_08487_));
 AND3x1_ASAP7_75t_R _28435_ (.A(_13786_),
    .B(_13853_),
    .C(_08406_),
    .Y(_08488_));
 BUFx4f_ASAP7_75t_R _28436_ (.A(_08488_),
    .Y(_08489_));
 AO22x1_ASAP7_75t_R _28437_ (.A1(_18622_),
    .A2(_08487_),
    .B1(_08489_),
    .B2(_18618_),
    .Y(_08490_));
 AO221x1_ASAP7_75t_R _28438_ (.A1(_18752_),
    .A2(_08484_),
    .B1(_08485_),
    .B2(_18747_),
    .C(_08490_),
    .Y(_08491_));
 AO22x1_ASAP7_75t_R _28439_ (.A1(_18613_),
    .A2(_08487_),
    .B1(_08485_),
    .B2(_18760_),
    .Y(_08492_));
 OR3x1_ASAP7_75t_R _28440_ (.A(_04883_),
    .B(_04884_),
    .C(_08423_),
    .Y(_08493_));
 OA211x2_ASAP7_75t_R _28441_ (.A1(_18609_),
    .A2(_08366_),
    .B(_08493_),
    .C(_18608_),
    .Y(_08494_));
 OR3x1_ASAP7_75t_R _28442_ (.A(_08477_),
    .B(_08492_),
    .C(_08494_),
    .Y(_08495_));
 AOI21x1_ASAP7_75t_R _28443_ (.A1(_13622_),
    .A2(_08399_),
    .B(_18629_),
    .Y(_08496_));
 BUFx6f_ASAP7_75t_R _28444_ (.A(_08458_),
    .Y(_08497_));
 OA21x2_ASAP7_75t_R _28445_ (.A1(_08496_),
    .A2(_08414_),
    .B(_08497_),
    .Y(_08498_));
 OA211x2_ASAP7_75t_R _28446_ (.A1(_08467_),
    .A2(_08491_),
    .B(_08495_),
    .C(_08498_),
    .Y(_08499_));
 AO221x2_ASAP7_75t_R _28447_ (.A1(_08433_),
    .A2(_08465_),
    .B1(_08479_),
    .B2(_08483_),
    .C(_08499_),
    .Y(_08500_));
 AO21x1_ASAP7_75t_R _28448_ (.A1(_13622_),
    .A2(_08398_),
    .B(_18623_),
    .Y(_08501_));
 BUFx4f_ASAP7_75t_R _28449_ (.A(_08501_),
    .Y(_08502_));
 OR3x1_ASAP7_75t_R _28450_ (.A(_13568_),
    .B(_18625_),
    .C(_06775_),
    .Y(_08503_));
 BUFx4f_ASAP7_75t_R _28451_ (.A(_08503_),
    .Y(_08504_));
 NAND2x1_ASAP7_75t_R _28452_ (.A(_08502_),
    .B(_08504_),
    .Y(_08505_));
 AND2x6_ASAP7_75t_R _28453_ (.A(_06794_),
    .B(_08369_),
    .Y(_08506_));
 AND2x2_ASAP7_75t_R _28454_ (.A(_08505_),
    .B(_08506_),
    .Y(_08507_));
 AND2x6_ASAP7_75t_R _28455_ (.A(_08502_),
    .B(_08504_),
    .Y(_08508_));
 BUFx4f_ASAP7_75t_R _28456_ (.A(_08508_),
    .Y(_08509_));
 OA22x2_ASAP7_75t_R _28457_ (.A1(_18742_),
    .A2(_08447_),
    .B1(_08451_),
    .B2(_18740_),
    .Y(_08510_));
 OA22x2_ASAP7_75t_R _28458_ (.A1(_18633_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18630_),
    .Y(_08511_));
 AO211x2_ASAP7_75t_R _28459_ (.A1(_08510_),
    .A2(_08511_),
    .B(_08425_),
    .C(_08435_),
    .Y(_08512_));
 OA22x2_ASAP7_75t_R _28460_ (.A1(_18732_),
    .A2(_08447_),
    .B1(_08451_),
    .B2(_18730_),
    .Y(_08513_));
 OA22x2_ASAP7_75t_R _28461_ (.A1(_18642_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18637_),
    .Y(_08514_));
 AO21x1_ASAP7_75t_R _28462_ (.A1(_08513_),
    .A2(_08514_),
    .B(_08441_),
    .Y(_08515_));
 AO221x1_ASAP7_75t_R _28463_ (.A1(_04523_),
    .A2(_15119_),
    .B1(_15953_),
    .B2(_04521_),
    .C(_08365_),
    .Y(_08516_));
 OA211x2_ASAP7_75t_R _28464_ (.A1(_18622_),
    .A2(_08407_),
    .B(_08516_),
    .C(_18608_),
    .Y(_08517_));
 AO221x1_ASAP7_75t_R _28465_ (.A1(_04632_),
    .A2(_15119_),
    .B1(_15953_),
    .B2(_04631_),
    .C(_08365_),
    .Y(_08518_));
 OA211x2_ASAP7_75t_R _28466_ (.A1(_18618_),
    .A2(_08407_),
    .B(_08518_),
    .C(_18610_),
    .Y(_08519_));
 OR4x1_ASAP7_75t_R _28467_ (.A(_08458_),
    .B(_08462_),
    .C(_08517_),
    .D(_08519_),
    .Y(_08520_));
 AO22x1_ASAP7_75t_R _28468_ (.A1(_18760_),
    .A2(_08489_),
    .B1(_08484_),
    .B2(_18613_),
    .Y(_08521_));
 OA211x2_ASAP7_75t_R _28469_ (.A1(_18609_),
    .A2(_08407_),
    .B(_08409_),
    .C(_18610_),
    .Y(_08522_));
 OR4x1_ASAP7_75t_R _28470_ (.A(_08458_),
    .B(_08435_),
    .C(_08521_),
    .D(_08522_),
    .Y(_08523_));
 AND4x2_ASAP7_75t_R _28471_ (.A(_08512_),
    .B(_08515_),
    .C(_08520_),
    .D(_08523_),
    .Y(_08524_));
 OAI22x1_ASAP7_75t_R _28472_ (.A1(_18653_),
    .A2(_08473_),
    .B1(_08451_),
    .B2(_18647_),
    .Y(_08525_));
 OAI22x1_ASAP7_75t_R _28473_ (.A1(_18725_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18717_),
    .Y(_08526_));
 BUFx4f_ASAP7_75t_R _28474_ (.A(_08435_),
    .Y(_08527_));
 OAI21x1_ASAP7_75t_R _28475_ (.A1(_08525_),
    .A2(_08526_),
    .B(_08527_),
    .Y(_08528_));
 OAI22x1_ASAP7_75t_R _28476_ (.A1(_18662_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18657_),
    .Y(_08529_));
 OAI22x1_ASAP7_75t_R _28477_ (.A1(_18715_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18707_),
    .Y(_08530_));
 BUFx6f_ASAP7_75t_R _28478_ (.A(_08462_),
    .Y(_08531_));
 OAI21x1_ASAP7_75t_R _28479_ (.A1(_08529_),
    .A2(_08530_),
    .B(_08531_),
    .Y(_08532_));
 AND3x1_ASAP7_75t_R _28480_ (.A(_08528_),
    .B(_08532_),
    .C(_08498_),
    .Y(_08533_));
 OA22x2_ASAP7_75t_R _28481_ (.A1(_18672_),
    .A2(_08447_),
    .B1(_08451_),
    .B2(_18667_),
    .Y(_08534_));
 OA22x2_ASAP7_75t_R _28482_ (.A1(_18702_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18697_),
    .Y(_08535_));
 AO21x1_ASAP7_75t_R _28483_ (.A1(_08534_),
    .A2(_08535_),
    .B(_08463_),
    .Y(_08536_));
 OA22x2_ASAP7_75t_R _28484_ (.A1(_18685_),
    .A2(_08447_),
    .B1(_08451_),
    .B2(_18680_),
    .Y(_08537_));
 OA22x2_ASAP7_75t_R _28485_ (.A1(_18692_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18687_),
    .Y(_08538_));
 AO21x1_ASAP7_75t_R _28486_ (.A1(_08537_),
    .A2(_08538_),
    .B(_08466_),
    .Y(_08539_));
 AND4x1_ASAP7_75t_R _28487_ (.A(_08480_),
    .B(_08426_),
    .C(_08536_),
    .D(_08539_),
    .Y(_08540_));
 AO211x2_ASAP7_75t_R _28488_ (.A1(_08432_),
    .A2(_08524_),
    .B(_08533_),
    .C(_08540_),
    .Y(_08541_));
 BUFx4f_ASAP7_75t_R _28489_ (.A(_08506_),
    .Y(_08542_));
 AND3x1_ASAP7_75t_R _28490_ (.A(_08509_),
    .B(_08541_),
    .C(_08542_),
    .Y(_08543_));
 AOI221x1_ASAP7_75t_R _28491_ (.A1(_08377_),
    .A2(_08431_),
    .B1(_08500_),
    .B2(_08507_),
    .C(_08543_),
    .Y(_08544_));
 OR2x2_ASAP7_75t_R _28492_ (.A(_04867_),
    .B(_05147_),
    .Y(_08545_));
 NAND3x2_ASAP7_75t_R _28493_ (.B(_02216_),
    .C(_08545_),
    .Y(_08546_),
    .A(_05154_));
 NAND2x2_ASAP7_75t_R _28494_ (.A(_13593_),
    .B(_08546_),
    .Y(_08547_));
 BUFx3_ASAP7_75t_R _28495_ (.A(_08547_),
    .Y(_08548_));
 BUFx4f_ASAP7_75t_R _28496_ (.A(_08546_),
    .Y(_08549_));
 BUFx4f_ASAP7_75t_R _28497_ (.A(_08549_),
    .Y(_08550_));
 BUFx6f_ASAP7_75t_R _28498_ (.A(_08550_),
    .Y(_08551_));
 AND3x1_ASAP7_75t_R _28499_ (.A(net2004),
    .B(_00104_),
    .C(_08551_),
    .Y(_08552_));
 AO21x1_ASAP7_75t_R _28500_ (.A1(_00447_),
    .A2(_08548_),
    .B(_08552_),
    .Y(_08553_));
 BUFx4f_ASAP7_75t_R _28501_ (.A(_08332_),
    .Y(_08554_));
 OA21x2_ASAP7_75t_R _28502_ (.A1(_05141_),
    .A2(_08553_),
    .B(_08554_),
    .Y(_08555_));
 OA211x2_ASAP7_75t_R _28503_ (.A1(_08351_),
    .A2(_08356_),
    .B(_08544_),
    .C(_08555_),
    .Y(_08556_));
 BUFx4f_ASAP7_75t_R _28504_ (.A(_01506_),
    .Y(_08557_));
 INVx2_ASAP7_75t_R _28505_ (.A(_08557_),
    .Y(_08558_));
 BUFx4f_ASAP7_75t_R _28506_ (.A(_01507_),
    .Y(_08559_));
 AND2x2_ASAP7_75t_R _28507_ (.A(_08558_),
    .B(_08559_),
    .Y(_08560_));
 INVx1_ASAP7_75t_R _28508_ (.A(_08559_),
    .Y(_08561_));
 BUFx4f_ASAP7_75t_R _28509_ (.A(_08561_),
    .Y(_08562_));
 AND2x4_ASAP7_75t_R _28510_ (.A(_08557_),
    .B(_08562_),
    .Y(_08563_));
 BUFx6f_ASAP7_75t_R _28511_ (.A(_02215_),
    .Y(_08564_));
 AND2x2_ASAP7_75t_R _28512_ (.A(_02210_),
    .B(_08564_),
    .Y(_08565_));
 BUFx4f_ASAP7_75t_R _28513_ (.A(_08565_),
    .Y(_08566_));
 AO221x1_ASAP7_75t_R _28514_ (.A1(net78),
    .A2(_08560_),
    .B1(_08563_),
    .B2(net102),
    .C(_08566_),
    .Y(_08567_));
 INVx1_ASAP7_75t_R _28515_ (.A(_01483_),
    .Y(_08568_));
 INVx1_ASAP7_75t_R _28516_ (.A(_01505_),
    .Y(_08569_));
 NAND2x2_ASAP7_75t_R _28517_ (.A(_05749_),
    .B(_08564_),
    .Y(_08570_));
 AO221x1_ASAP7_75t_R _28518_ (.A1(_08568_),
    .A2(_08560_),
    .B1(_08563_),
    .B2(_08569_),
    .C(_08570_),
    .Y(_08571_));
 BUFx4f_ASAP7_75t_R _28519_ (.A(_08557_),
    .Y(_08572_));
 BUFx4f_ASAP7_75t_R _28520_ (.A(_08559_),
    .Y(_08573_));
 BUFx6f_ASAP7_75t_R _28521_ (.A(_08573_),
    .Y(_08574_));
 NOR2x2_ASAP7_75t_R _28522_ (.A(_08572_),
    .B(_08574_),
    .Y(_08575_));
 AND2x2_ASAP7_75t_R _28523_ (.A(_05749_),
    .B(_05760_),
    .Y(_08576_));
 BUFx6f_ASAP7_75t_R _28524_ (.A(_08576_),
    .Y(_08577_));
 NOR2x1_ASAP7_75t_R _28525_ (.A(_01498_),
    .B(_08577_),
    .Y(_08578_));
 AO21x1_ASAP7_75t_R _28526_ (.A1(net87),
    .A2(_05760_),
    .B(_08578_),
    .Y(_08579_));
 BUFx4f_ASAP7_75t_R _28527_ (.A(_08573_),
    .Y(_08580_));
 AND2x6_ASAP7_75t_R _28528_ (.A(_08572_),
    .B(_08580_),
    .Y(_08581_));
 AO222x2_ASAP7_75t_R _28529_ (.A1(_08567_),
    .A2(_08571_),
    .B1(_08575_),
    .B2(_08579_),
    .C1(_08581_),
    .C2(net48),
    .Y(_08582_));
 NAND2x1_ASAP7_75t_R _28530_ (.A(_08345_),
    .B(_08582_),
    .Y(_08583_));
 OAI21x1_ASAP7_75t_R _28531_ (.A1(_08346_),
    .A2(_08556_),
    .B(_08583_),
    .Y(_08584_));
 BUFx6f_ASAP7_75t_R _28532_ (.A(_08584_),
    .Y(_08585_));
 OR3x1_ASAP7_75t_R _28533_ (.A(_14153_),
    .B(_14303_),
    .C(_14232_),
    .Y(_08586_));
 OA33x2_ASAP7_75t_R _28534_ (.A1(_04924_),
    .A2(_04921_),
    .A3(_06782_),
    .B1(_05143_),
    .B2(_08343_),
    .B3(_08335_),
    .Y(_08587_));
 BUFx3_ASAP7_75t_R _28535_ (.A(_08587_),
    .Y(_08588_));
 NAND2x2_ASAP7_75t_R _28536_ (.A(_14726_),
    .B(_13438_),
    .Y(_08589_));
 OR3x4_ASAP7_75t_R _28537_ (.A(_08586_),
    .B(_08588_),
    .C(_08589_),
    .Y(_08590_));
 BUFx6f_ASAP7_75t_R _28538_ (.A(_08590_),
    .Y(_08591_));
 NAND2x1_ASAP7_75t_R _28539_ (.A(_01814_),
    .B(_08591_),
    .Y(_08592_));
 OA21x2_ASAP7_75t_R _28540_ (.A1(_08342_),
    .A2(_08585_),
    .B(_08592_),
    .Y(_02858_));
 BUFx3_ASAP7_75t_R _28541_ (.A(_08027_),
    .Y(_08593_));
 BUFx3_ASAP7_75t_R _28542_ (.A(_13438_),
    .Y(_08594_));
 BUFx4f_ASAP7_75t_R _28543_ (.A(_08338_),
    .Y(_08595_));
 AND3x2_ASAP7_75t_R _28544_ (.A(_14153_),
    .B(_14050_),
    .C(_14231_),
    .Y(_08596_));
 AND4x2_ASAP7_75t_R _28545_ (.A(_08593_),
    .B(_08594_),
    .C(_08595_),
    .D(_08596_),
    .Y(_08597_));
 BUFx10_ASAP7_75t_R _28546_ (.A(_08597_),
    .Y(_08598_));
 AND3x4_ASAP7_75t_R _28547_ (.A(_05097_),
    .B(_06833_),
    .C(_08336_),
    .Y(_08599_));
 BUFx6f_ASAP7_75t_R _28548_ (.A(_08599_),
    .Y(_08600_));
 AO221x1_ASAP7_75t_R _28549_ (.A1(net83),
    .A2(_08560_),
    .B1(_08563_),
    .B2(net51),
    .C(_08566_),
    .Y(_08601_));
 INVx1_ASAP7_75t_R _28550_ (.A(_01502_),
    .Y(_08602_));
 BUFx3_ASAP7_75t_R _28551_ (.A(_08560_),
    .Y(_08603_));
 BUFx3_ASAP7_75t_R _28552_ (.A(_08563_),
    .Y(_08604_));
 INVx1_ASAP7_75t_R _28553_ (.A(_01487_),
    .Y(_08605_));
 AO221x1_ASAP7_75t_R _28554_ (.A1(_08602_),
    .A2(_08603_),
    .B1(_08604_),
    .B2(_08605_),
    .C(_08570_),
    .Y(_08606_));
 INVx1_ASAP7_75t_R _28555_ (.A(net91),
    .Y(_08607_));
 OAI22x1_ASAP7_75t_R _28556_ (.A1(_08607_),
    .A2(_08564_),
    .B1(_08577_),
    .B2(_01493_),
    .Y(_08608_));
 AO222x2_ASAP7_75t_R _28557_ (.A1(net98),
    .A2(_08581_),
    .B1(_08601_),
    .B2(_08606_),
    .C1(_08608_),
    .C2(_08575_),
    .Y(_08609_));
 INVx1_ASAP7_75t_R _28558_ (.A(_00151_),
    .Y(_08610_));
 AND3x1_ASAP7_75t_R _28559_ (.A(_13593_),
    .B(_08610_),
    .C(_08549_),
    .Y(_08611_));
 AO21x1_ASAP7_75t_R _28560_ (.A1(_05683_),
    .A2(_08547_),
    .B(_08611_),
    .Y(_08612_));
 AO21x1_ASAP7_75t_R _28561_ (.A1(_05304_),
    .A2(_08612_),
    .B(_13776_),
    .Y(_08613_));
 OA22x2_ASAP7_75t_R _28562_ (.A1(_08554_),
    .A2(_06516_),
    .B1(_08377_),
    .B2(_08613_),
    .Y(_08614_));
 OR3x4_ASAP7_75t_R _28563_ (.A(_08496_),
    .B(_08414_),
    .C(_08411_),
    .Y(_08615_));
 AND2x2_ASAP7_75t_R _28564_ (.A(_08366_),
    .B(_08615_),
    .Y(_08616_));
 OA211x2_ASAP7_75t_R _28565_ (.A1(_08411_),
    .A2(_08466_),
    .B(_08424_),
    .C(_08425_),
    .Y(_08617_));
 OA22x2_ASAP7_75t_R _28566_ (.A1(_18760_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18752_),
    .Y(_08618_));
 OA22x2_ASAP7_75t_R _28567_ (.A1(_18618_),
    .A2(_08454_),
    .B1(_08456_),
    .B2(_18613_),
    .Y(_08619_));
 AND4x1_ASAP7_75t_R _28568_ (.A(_08497_),
    .B(_08531_),
    .C(_08618_),
    .D(_08619_),
    .Y(_08620_));
 AO221x1_ASAP7_75t_R _28569_ (.A1(_04392_),
    .A2(_04522_),
    .B1(_15953_),
    .B2(_04391_),
    .C(_08365_),
    .Y(_08621_));
 OA211x2_ASAP7_75t_R _28570_ (.A1(_18630_),
    .A2(_08407_),
    .B(_08621_),
    .C(_18608_),
    .Y(_08622_));
 OA211x2_ASAP7_75t_R _28571_ (.A1(_18622_),
    .A2(_08407_),
    .B(_08516_),
    .C(_18610_),
    .Y(_08623_));
 OA21x2_ASAP7_75t_R _28572_ (.A1(_08622_),
    .A2(_08623_),
    .B(_08422_),
    .Y(_08624_));
 OR3x1_ASAP7_75t_R _28573_ (.A(_08617_),
    .B(_08620_),
    .C(_08624_),
    .Y(_08625_));
 OA21x2_ASAP7_75t_R _28574_ (.A1(_13568_),
    .A2(_06775_),
    .B(_18625_),
    .Y(_08626_));
 AND3x4_ASAP7_75t_R _28575_ (.A(_13622_),
    .B(_18623_),
    .C(_08398_),
    .Y(_08627_));
 OR3x1_ASAP7_75t_R _28576_ (.A(_08626_),
    .B(_08627_),
    .C(_08411_),
    .Y(_08628_));
 OAI21x1_ASAP7_75t_R _28577_ (.A1(_08508_),
    .A2(_08625_),
    .B(_08628_),
    .Y(_08629_));
 NAND2x1_ASAP7_75t_R _28578_ (.A(_08481_),
    .B(_08629_),
    .Y(_08630_));
 NAND2x2_ASAP7_75t_R _28579_ (.A(_08404_),
    .B(_08405_),
    .Y(_08631_));
 BUFx4f_ASAP7_75t_R _28580_ (.A(_08631_),
    .Y(_08632_));
 BUFx4f_ASAP7_75t_R _28581_ (.A(_08497_),
    .Y(_08633_));
 AND3x1_ASAP7_75t_R _28582_ (.A(_08482_),
    .B(_08528_),
    .C(_08532_),
    .Y(_08634_));
 AOI21x1_ASAP7_75t_R _28583_ (.A1(_08633_),
    .A2(_08479_),
    .B(_08634_),
    .Y(_08635_));
 AND3x4_ASAP7_75t_R _28584_ (.A(_08480_),
    .B(_08502_),
    .C(_08504_),
    .Y(_08636_));
 AND2x2_ASAP7_75t_R _28585_ (.A(_08426_),
    .B(_08527_),
    .Y(_08637_));
 NOR2x1_ASAP7_75t_R _28586_ (.A(_08443_),
    .B(_08445_),
    .Y(_08638_));
 NOR2x1_ASAP7_75t_R _28587_ (.A(_08437_),
    .B(_08439_),
    .Y(_08639_));
 AND2x2_ASAP7_75t_R _28588_ (.A(_08425_),
    .B(_08463_),
    .Y(_08640_));
 NAND2x1_ASAP7_75t_R _28589_ (.A(_08534_),
    .B(_08535_),
    .Y(_08641_));
 NAND2x1_ASAP7_75t_R _28590_ (.A(_08537_),
    .B(_08538_),
    .Y(_08642_));
 AND2x4_ASAP7_75t_R _28591_ (.A(_08458_),
    .B(_08463_),
    .Y(_08643_));
 AO22x1_ASAP7_75t_R _28592_ (.A1(_08422_),
    .A2(_08641_),
    .B1(_08642_),
    .B2(_08643_),
    .Y(_08644_));
 AO221x2_ASAP7_75t_R _28593_ (.A1(_08637_),
    .A2(_08638_),
    .B1(_08639_),
    .B2(_08640_),
    .C(_08644_),
    .Y(_08645_));
 BUFx4f_ASAP7_75t_R _28594_ (.A(_08422_),
    .Y(_08646_));
 OR2x2_ASAP7_75t_R _28595_ (.A(_08517_),
    .B(_08519_),
    .Y(_08647_));
 OR2x2_ASAP7_75t_R _28596_ (.A(_08521_),
    .B(_08522_),
    .Y(_08648_));
 OA211x2_ASAP7_75t_R _28597_ (.A1(_18609_),
    .A2(_08423_),
    .B(_08408_),
    .C(_08409_),
    .Y(_08649_));
 AND2x2_ASAP7_75t_R _28598_ (.A(_08426_),
    .B(_08649_),
    .Y(_08650_));
 AO221x1_ASAP7_75t_R _28599_ (.A1(_08646_),
    .A2(_08647_),
    .B1(_08648_),
    .B2(_08643_),
    .C(_08650_),
    .Y(_08651_));
 OR3x4_ASAP7_75t_R _28600_ (.A(_08480_),
    .B(_08626_),
    .C(_08627_),
    .Y(_08652_));
 AO21x2_ASAP7_75t_R _28601_ (.A1(_08502_),
    .A2(_08504_),
    .B(_08480_),
    .Y(_08653_));
 AO211x2_ASAP7_75t_R _28602_ (.A1(_08452_),
    .A2(_08457_),
    .B(_08426_),
    .C(_08527_),
    .Y(_08654_));
 BUFx4f_ASAP7_75t_R _28603_ (.A(_08441_),
    .Y(_08655_));
 AO21x1_ASAP7_75t_R _28604_ (.A1(_08460_),
    .A2(_08461_),
    .B(_08655_),
    .Y(_08656_));
 BUFx4f_ASAP7_75t_R _28605_ (.A(_08458_),
    .Y(_08657_));
 AO211x2_ASAP7_75t_R _28606_ (.A1(_08510_),
    .A2(_08511_),
    .B(_08657_),
    .C(_08527_),
    .Y(_08658_));
 AO211x2_ASAP7_75t_R _28607_ (.A1(_08513_),
    .A2(_08514_),
    .B(_08657_),
    .C(_08531_),
    .Y(_08659_));
 AND4x2_ASAP7_75t_R _28608_ (.A(_08654_),
    .B(_08656_),
    .C(_08658_),
    .D(_08659_),
    .Y(_08660_));
 OAI22x1_ASAP7_75t_R _28609_ (.A1(_08651_),
    .A2(_08652_),
    .B1(_08653_),
    .B2(_08660_),
    .Y(_08661_));
 AOI221x1_ASAP7_75t_R _28610_ (.A1(_08632_),
    .A2(_08635_),
    .B1(_08636_),
    .B2(_08645_),
    .C(_08661_),
    .Y(_08662_));
 BUFx4f_ASAP7_75t_R _28611_ (.A(_08382_),
    .Y(_08663_));
 BUFx6f_ASAP7_75t_R _28612_ (.A(_08384_),
    .Y(_08664_));
 BUFx10_ASAP7_75t_R _28613_ (.A(_08664_),
    .Y(_08665_));
 BUFx6f_ASAP7_75t_R _28614_ (.A(_08389_),
    .Y(_08666_));
 BUFx6f_ASAP7_75t_R _28615_ (.A(_08666_),
    .Y(_08667_));
 OAI22x1_ASAP7_75t_R _28616_ (.A1(_00305_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00304_),
    .Y(_08668_));
 BUFx3_ASAP7_75t_R _28617_ (.A(_08360_),
    .Y(_08669_));
 BUFx3_ASAP7_75t_R _28618_ (.A(_08380_),
    .Y(_08670_));
 AO221x1_ASAP7_75t_R _28619_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_08669_),
    .B1(_08670_),
    .B2(_02257_),
    .C(_08613_),
    .Y(_08671_));
 AO21x1_ASAP7_75t_R _28620_ (.A1(_08663_),
    .A2(_08668_),
    .B(_08671_),
    .Y(_08672_));
 AO221x1_ASAP7_75t_R _28621_ (.A1(_08616_),
    .A2(_08630_),
    .B1(_08662_),
    .B2(_08542_),
    .C(_08672_),
    .Y(_08673_));
 AO21x1_ASAP7_75t_R _28622_ (.A1(_08614_),
    .A2(_08673_),
    .B(_08345_),
    .Y(_08674_));
 OA21x2_ASAP7_75t_R _28623_ (.A1(_08600_),
    .A2(_08609_),
    .B(_08674_),
    .Y(_08675_));
 BUFx4f_ASAP7_75t_R _28624_ (.A(_08675_),
    .Y(_08676_));
 NAND2x2_ASAP7_75t_R _28625_ (.A(_08027_),
    .B(_13438_),
    .Y(_08677_));
 OR3x1_ASAP7_75t_R _28626_ (.A(_14049_),
    .B(_14303_),
    .C(_14232_),
    .Y(_08678_));
 OR3x1_ASAP7_75t_R _28627_ (.A(_08677_),
    .B(_08588_),
    .C(_08678_),
    .Y(_08679_));
 BUFx10_ASAP7_75t_R _28628_ (.A(_08679_),
    .Y(_08680_));
 AND2x2_ASAP7_75t_R _28629_ (.A(_14271_),
    .B(_08680_),
    .Y(_08681_));
 AO21x1_ASAP7_75t_R _28630_ (.A1(_08598_),
    .A2(_08676_),
    .B(_08681_),
    .Y(_02859_));
 BUFx6f_ASAP7_75t_R _28631_ (.A(_08680_),
    .Y(_08682_));
 BUFx4f_ASAP7_75t_R _28632_ (.A(_08344_),
    .Y(_08683_));
 BUFx6f_ASAP7_75t_R _28633_ (.A(_08683_),
    .Y(_08684_));
 BUFx4f_ASAP7_75t_R _28634_ (.A(_08566_),
    .Y(_08685_));
 AO221x1_ASAP7_75t_R _28635_ (.A1(net84),
    .A2(_08603_),
    .B1(_08604_),
    .B2(net75),
    .C(_08685_),
    .Y(_08686_));
 INVx1_ASAP7_75t_R _28636_ (.A(_01501_),
    .Y(_08687_));
 INVx1_ASAP7_75t_R _28637_ (.A(_01486_),
    .Y(_08688_));
 BUFx4f_ASAP7_75t_R _28638_ (.A(_08570_),
    .Y(_08689_));
 AO221x1_ASAP7_75t_R _28639_ (.A1(_08687_),
    .A2(_08603_),
    .B1(_08604_),
    .B2(_08688_),
    .C(_08689_),
    .Y(_08690_));
 INVx1_ASAP7_75t_R _28640_ (.A(net92),
    .Y(_08691_));
 OAI22x1_ASAP7_75t_R _28641_ (.A1(_08691_),
    .A2(_08564_),
    .B1(_08577_),
    .B2(_01492_),
    .Y(_08692_));
 AO222x2_ASAP7_75t_R _28642_ (.A1(net99),
    .A2(_08581_),
    .B1(_08686_),
    .B2(_08690_),
    .C1(_08692_),
    .C2(_08575_),
    .Y(_08693_));
 BUFx4f_ASAP7_75t_R _28643_ (.A(_08599_),
    .Y(_08694_));
 AND2x4_ASAP7_75t_R _28644_ (.A(_08404_),
    .B(_08405_),
    .Y(_08695_));
 OR3x1_ASAP7_75t_R _28645_ (.A(_08463_),
    .B(_08521_),
    .C(_08522_),
    .Y(_08696_));
 OA21x2_ASAP7_75t_R _28646_ (.A1(_08410_),
    .A2(_08466_),
    .B(_08425_),
    .Y(_08697_));
 AND3x1_ASAP7_75t_R _28647_ (.A(_08422_),
    .B(_08510_),
    .C(_08511_),
    .Y(_08698_));
 OA211x2_ASAP7_75t_R _28648_ (.A1(_08517_),
    .A2(_08519_),
    .B(_08458_),
    .C(_08463_),
    .Y(_08699_));
 AO211x2_ASAP7_75t_R _28649_ (.A1(_08696_),
    .A2(_08697_),
    .B(_08698_),
    .C(_08699_),
    .Y(_08700_));
 OR2x2_ASAP7_75t_R _28650_ (.A(_08695_),
    .B(_08700_),
    .Y(_08701_));
 OR3x4_ASAP7_75t_R _28651_ (.A(_08413_),
    .B(_08415_),
    .C(_08411_),
    .Y(_08702_));
 AND2x2_ASAP7_75t_R _28652_ (.A(_08429_),
    .B(_08702_),
    .Y(_08703_));
 OR3x2_ASAP7_75t_R _28653_ (.A(_08432_),
    .B(_08626_),
    .C(_08627_),
    .Y(_08704_));
 OA22x2_ASAP7_75t_R _28654_ (.A1(_18707_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18702_),
    .Y(_08705_));
 AOI22x1_ASAP7_75t_R _28655_ (.A1(_18669_),
    .A2(_08484_),
    .B1(_08485_),
    .B2(_18664_),
    .Y(_08706_));
 NAND2x1_ASAP7_75t_R _28656_ (.A(_08705_),
    .B(_08706_),
    .Y(_08707_));
 AOI22x1_ASAP7_75t_R _28657_ (.A1(_18699_),
    .A2(_08487_),
    .B1(_08489_),
    .B2(_18694_),
    .Y(_08708_));
 OA22x2_ASAP7_75t_R _28658_ (.A1(_18680_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18672_),
    .Y(_08709_));
 AOI21x1_ASAP7_75t_R _28659_ (.A1(_08708_),
    .A2(_08709_),
    .B(_08477_),
    .Y(_08710_));
 AOI21x1_ASAP7_75t_R _28660_ (.A1(_08477_),
    .A2(_08707_),
    .B(_08710_),
    .Y(_08711_));
 OAI22x1_ASAP7_75t_R _28661_ (.A1(_18680_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18672_),
    .Y(_08712_));
 AO22x2_ASAP7_75t_R _28662_ (.A1(_18699_),
    .A2(_08484_),
    .B1(_08485_),
    .B2(_18694_),
    .Y(_08713_));
 NOR3x2_ASAP7_75t_R _28663_ (.B(_08712_),
    .C(_08713_),
    .Y(_08714_),
    .A(_08531_));
 AO21x1_ASAP7_75t_R _28664_ (.A1(_08468_),
    .A2(_08475_),
    .B(_18685_),
    .Y(_08715_));
 OR3x1_ASAP7_75t_R _28665_ (.A(_18687_),
    .B(_08489_),
    .C(_08485_),
    .Y(_08716_));
 AND3x1_ASAP7_75t_R _28666_ (.A(_08531_),
    .B(_08715_),
    .C(_08716_),
    .Y(_08717_));
 OA21x2_ASAP7_75t_R _28667_ (.A1(_08714_),
    .A2(_08717_),
    .B(_08633_),
    .Y(_08718_));
 AO21x1_ASAP7_75t_R _28668_ (.A1(_08482_),
    .A2(_08711_),
    .B(_08718_),
    .Y(_08719_));
 OAI22x1_ASAP7_75t_R _28669_ (.A1(_18637_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18633_),
    .Y(_08720_));
 OAI22x1_ASAP7_75t_R _28670_ (.A1(_18740_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18732_),
    .Y(_08721_));
 OR2x2_ASAP7_75t_R _28671_ (.A(_08720_),
    .B(_08721_),
    .Y(_08722_));
 OA22x2_ASAP7_75t_R _28672_ (.A1(_18647_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18642_),
    .Y(_08723_));
 OA22x2_ASAP7_75t_R _28673_ (.A1(_18730_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18725_),
    .Y(_08724_));
 NAND2x1_ASAP7_75t_R _28674_ (.A(_08723_),
    .B(_08724_),
    .Y(_08725_));
 AO22x1_ASAP7_75t_R _28675_ (.A1(_08646_),
    .A2(_08722_),
    .B1(_08725_),
    .B2(_08643_),
    .Y(_08726_));
 OAI22x1_ASAP7_75t_R _28676_ (.A1(_18717_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18715_),
    .Y(_08727_));
 AO221x2_ASAP7_75t_R _28677_ (.A1(_18659_),
    .A2(_08487_),
    .B1(_08489_),
    .B2(_18655_),
    .C(_08727_),
    .Y(_08728_));
 AOI22x1_ASAP7_75t_R _28678_ (.A1(_18669_),
    .A2(_08487_),
    .B1(_08489_),
    .B2(_18664_),
    .Y(_08729_));
 OA22x2_ASAP7_75t_R _28679_ (.A1(_18707_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18702_),
    .Y(_08730_));
 NAND2x1_ASAP7_75t_R _28680_ (.A(_08729_),
    .B(_08730_),
    .Y(_08731_));
 AO22x1_ASAP7_75t_R _28681_ (.A1(_08637_),
    .A2(_08728_),
    .B1(_08731_),
    .B2(_08640_),
    .Y(_08732_));
 OAI21x1_ASAP7_75t_R _28682_ (.A1(_08726_),
    .A2(_08732_),
    .B(_08631_),
    .Y(_08733_));
 OA22x2_ASAP7_75t_R _28683_ (.A1(_18730_),
    .A2(_08473_),
    .B1(_08451_),
    .B2(_18725_),
    .Y(_08734_));
 OA22x2_ASAP7_75t_R _28684_ (.A1(_18647_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18642_),
    .Y(_08735_));
 AO211x2_ASAP7_75t_R _28685_ (.A1(_08734_),
    .A2(_08735_),
    .B(_08426_),
    .C(_08466_),
    .Y(_08736_));
 OA22x2_ASAP7_75t_R _28686_ (.A1(_18717_),
    .A2(_08473_),
    .B1(_08468_),
    .B2(_18715_),
    .Y(_08737_));
 OA22x2_ASAP7_75t_R _28687_ (.A1(_18657_),
    .A2(_08470_),
    .B1(_08475_),
    .B2(_18653_),
    .Y(_08738_));
 AO21x1_ASAP7_75t_R _28688_ (.A1(_08737_),
    .A2(_08738_),
    .B(_08655_),
    .Y(_08739_));
 AO221x1_ASAP7_75t_R _28689_ (.A1(_17234_),
    .A2(_04522_),
    .B1(_15953_),
    .B2(_17233_),
    .C(_08365_),
    .Y(_08740_));
 OA211x2_ASAP7_75t_R _28690_ (.A1(_18637_),
    .A2(_08423_),
    .B(_08740_),
    .C(_18608_),
    .Y(_08741_));
 AO221x1_ASAP7_75t_R _28691_ (.A1(_04283_),
    .A2(_04522_),
    .B1(_15953_),
    .B2(_04282_),
    .C(_08365_),
    .Y(_08742_));
 OA211x2_ASAP7_75t_R _28692_ (.A1(_18633_),
    .A2(_08407_),
    .B(_08742_),
    .C(_18610_),
    .Y(_08743_));
 OR4x1_ASAP7_75t_R _28693_ (.A(_08497_),
    .B(_08463_),
    .C(_08741_),
    .D(_08743_),
    .Y(_08744_));
 OR4x1_ASAP7_75t_R _28694_ (.A(_08497_),
    .B(_08435_),
    .C(_08622_),
    .D(_08623_),
    .Y(_08745_));
 AND4x2_ASAP7_75t_R _28695_ (.A(_08736_),
    .B(_08739_),
    .C(_08744_),
    .D(_08745_),
    .Y(_08746_));
 AO21x1_ASAP7_75t_R _28696_ (.A1(_13367_),
    .A2(_13553_),
    .B(_13622_),
    .Y(_08747_));
 NAND2x1_ASAP7_75t_R _28697_ (.A(_00296_),
    .B(_13622_),
    .Y(_08748_));
 AO33x2_ASAP7_75t_R _28698_ (.A1(_08747_),
    .A2(_08748_),
    .A3(_08424_),
    .B1(_08618_),
    .B2(_08619_),
    .B3(_08466_),
    .Y(_08749_));
 AO21x1_ASAP7_75t_R _28699_ (.A1(_08633_),
    .A2(_08749_),
    .B(_08650_),
    .Y(_08750_));
 OA22x2_ASAP7_75t_R _28700_ (.A1(_08653_),
    .A2(_08746_),
    .B1(_08750_),
    .B2(_08652_),
    .Y(_08751_));
 OA211x2_ASAP7_75t_R _28701_ (.A1(_08704_),
    .A2(_08719_),
    .B(_08733_),
    .C(_08751_),
    .Y(_08752_));
 BUFx4f_ASAP7_75t_R _28702_ (.A(_13593_),
    .Y(_08753_));
 AO21x1_ASAP7_75t_R _28703_ (.A1(_08753_),
    .A2(_08550_),
    .B(_00801_),
    .Y(_08754_));
 OAI21x1_ASAP7_75t_R _28704_ (.A1(_00158_),
    .A2(_08547_),
    .B(_08754_),
    .Y(_08755_));
 OAI22x1_ASAP7_75t_R _28705_ (.A1(_00307_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00306_),
    .Y(_08756_));
 AO22x1_ASAP7_75t_R _28706_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_08360_),
    .B1(_08380_),
    .B2(_02258_),
    .Y(_08757_));
 AO21x1_ASAP7_75t_R _28707_ (.A1(_08381_),
    .A2(_08756_),
    .B(_08757_),
    .Y(_08758_));
 AO221x1_ASAP7_75t_R _28708_ (.A1(_05514_),
    .A2(_08755_),
    .B1(_08758_),
    .B2(_08376_),
    .C(_05078_),
    .Y(_08759_));
 AO221x1_ASAP7_75t_R _28709_ (.A1(_08701_),
    .A2(_08703_),
    .B1(_08752_),
    .B2(_08542_),
    .C(_08759_),
    .Y(_08760_));
 OA211x2_ASAP7_75t_R _28710_ (.A1(_08554_),
    .A2(_06532_),
    .B(_08694_),
    .C(_08760_),
    .Y(_08761_));
 AO21x2_ASAP7_75t_R _28711_ (.A1(_08684_),
    .A2(_08693_),
    .B(_08761_),
    .Y(_08762_));
 BUFx4f_ASAP7_75t_R _28712_ (.A(_08762_),
    .Y(_08763_));
 BUFx6f_ASAP7_75t_R _28713_ (.A(_08680_),
    .Y(_08764_));
 NAND2x1_ASAP7_75t_R _28714_ (.A(_00575_),
    .B(_08764_),
    .Y(_08765_));
 OA21x2_ASAP7_75t_R _28715_ (.A1(_08682_),
    .A2(_08763_),
    .B(_08765_),
    .Y(_02860_));
 AO221x1_ASAP7_75t_R _28716_ (.A1(net85),
    .A2(_08603_),
    .B1(_08604_),
    .B2(net76),
    .C(_08566_),
    .Y(_08766_));
 INVx1_ASAP7_75t_R _28717_ (.A(_01500_),
    .Y(_08767_));
 INVx1_ASAP7_75t_R _28718_ (.A(_01485_),
    .Y(_08768_));
 AO221x1_ASAP7_75t_R _28719_ (.A1(_08767_),
    .A2(_08603_),
    .B1(_08604_),
    .B2(_08768_),
    .C(_08570_),
    .Y(_08769_));
 INVx1_ASAP7_75t_R _28720_ (.A(net94),
    .Y(_08770_));
 OAI22x1_ASAP7_75t_R _28721_ (.A1(_08770_),
    .A2(_08564_),
    .B1(_08577_),
    .B2(_01491_),
    .Y(_08771_));
 AO222x2_ASAP7_75t_R _28722_ (.A1(net100),
    .A2(_08581_),
    .B1(_08766_),
    .B2(_08769_),
    .C1(_08771_),
    .C2(_08575_),
    .Y(_08772_));
 XOR2x2_ASAP7_75t_R _28723_ (.A(_00167_),
    .B(_00165_),
    .Y(_08773_));
 BUFx4f_ASAP7_75t_R _28724_ (.A(_13595_),
    .Y(_08774_));
 AO21x1_ASAP7_75t_R _28725_ (.A1(_08774_),
    .A2(_08551_),
    .B(_05688_),
    .Y(_08775_));
 OA211x2_ASAP7_75t_R _28726_ (.A1(_08548_),
    .A2(_08773_),
    .B(_08775_),
    .C(_05515_),
    .Y(_08776_));
 BUFx4f_ASAP7_75t_R _28727_ (.A(_08429_),
    .Y(_08777_));
 OR2x2_ASAP7_75t_R _28728_ (.A(_08622_),
    .B(_08623_),
    .Y(_08778_));
 OR2x2_ASAP7_75t_R _28729_ (.A(_08741_),
    .B(_08743_),
    .Y(_08779_));
 AO222x2_ASAP7_75t_R _28730_ (.A1(_08643_),
    .A2(_08778_),
    .B1(_08779_),
    .B2(_08646_),
    .C1(_08482_),
    .C2(_08749_),
    .Y(_08780_));
 OR2x2_ASAP7_75t_R _28731_ (.A(_08695_),
    .B(_08780_),
    .Y(_08781_));
 OAI22x1_ASAP7_75t_R _28732_ (.A1(_00309_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00308_),
    .Y(_08782_));
 AO22x1_ASAP7_75t_R _28733_ (.A1(\alu_adder_result_ex[6] ),
    .A2(_08669_),
    .B1(_08670_),
    .B2(_02259_),
    .Y(_08783_));
 AO21x1_ASAP7_75t_R _28734_ (.A1(_08382_),
    .A2(_08782_),
    .B(_08783_),
    .Y(_08784_));
 AO32x1_ASAP7_75t_R _28735_ (.A1(_08777_),
    .A2(_08702_),
    .A3(_08781_),
    .B1(_08784_),
    .B2(_08376_),
    .Y(_08785_));
 BUFx4f_ASAP7_75t_R _28736_ (.A(_08505_),
    .Y(_08786_));
 AO21x1_ASAP7_75t_R _28737_ (.A1(_08452_),
    .A2(_08457_),
    .B(_08655_),
    .Y(_08787_));
 AO211x2_ASAP7_75t_R _28738_ (.A1(_08510_),
    .A2(_08511_),
    .B(_08657_),
    .C(_08477_),
    .Y(_08788_));
 AO211x2_ASAP7_75t_R _28739_ (.A1(_08513_),
    .A2(_08514_),
    .B(_08426_),
    .C(_08467_),
    .Y(_08789_));
 OR4x1_ASAP7_75t_R _28740_ (.A(_08657_),
    .B(_08527_),
    .C(_08517_),
    .D(_08519_),
    .Y(_08790_));
 AND4x2_ASAP7_75t_R _28741_ (.A(_08787_),
    .B(_08788_),
    .C(_08789_),
    .D(_08790_),
    .Y(_08791_));
 OR2x2_ASAP7_75t_R _28742_ (.A(_08411_),
    .B(_08422_),
    .Y(_08792_));
 OR3x1_ASAP7_75t_R _28743_ (.A(_08655_),
    .B(_08521_),
    .C(_08522_),
    .Y(_08793_));
 AND4x2_ASAP7_75t_R _28744_ (.A(_08502_),
    .B(_08504_),
    .C(_08792_),
    .D(_08793_),
    .Y(_08794_));
 AOI21x1_ASAP7_75t_R _28745_ (.A1(_08786_),
    .A2(_08791_),
    .B(_08794_),
    .Y(_08795_));
 NAND2x1_ASAP7_75t_R _28746_ (.A(_08460_),
    .B(_08461_),
    .Y(_08796_));
 AO22x1_ASAP7_75t_R _28747_ (.A1(_08643_),
    .A2(_08638_),
    .B1(_08639_),
    .B2(_08637_),
    .Y(_08797_));
 AO221x2_ASAP7_75t_R _28748_ (.A1(_08646_),
    .A2(_08642_),
    .B1(_08796_),
    .B2(_08640_),
    .C(_08797_),
    .Y(_08798_));
 NOR2x1_ASAP7_75t_R _28749_ (.A(_08655_),
    .B(_08472_),
    .Y(_08799_));
 OA21x2_ASAP7_75t_R _28750_ (.A1(_08529_),
    .A2(_08530_),
    .B(_08637_),
    .Y(_08800_));
 OR2x2_ASAP7_75t_R _28751_ (.A(_08525_),
    .B(_08526_),
    .Y(_08801_));
 AO22x1_ASAP7_75t_R _28752_ (.A1(_08640_),
    .A2(_08641_),
    .B1(_08801_),
    .B2(_08643_),
    .Y(_08802_));
 OR4x1_ASAP7_75t_R _28753_ (.A(_08508_),
    .B(_08799_),
    .C(_08800_),
    .D(_08802_),
    .Y(_08803_));
 OA211x2_ASAP7_75t_R _28754_ (.A1(_08786_),
    .A2(_08798_),
    .B(_08803_),
    .C(_08481_),
    .Y(_08804_));
 AND4x2_ASAP7_75t_R _28755_ (.A(_06794_),
    .B(_14912_),
    .C(_08367_),
    .D(_08368_),
    .Y(_08805_));
 INVx1_ASAP7_75t_R _28756_ (.A(_08805_),
    .Y(_08806_));
 AOI211x1_ASAP7_75t_R _28757_ (.A1(_08433_),
    .A2(_08795_),
    .B(_08804_),
    .C(_08806_),
    .Y(_08807_));
 OR5x2_ASAP7_75t_R _28758_ (.A(_06557_),
    .B(_08683_),
    .C(_08776_),
    .D(_08785_),
    .E(_08807_),
    .Y(_08808_));
 OA21x2_ASAP7_75t_R _28759_ (.A1(_08600_),
    .A2(_08772_),
    .B(_08808_),
    .Y(_08809_));
 BUFx6f_ASAP7_75t_R _28760_ (.A(_08809_),
    .Y(_08810_));
 NAND2x1_ASAP7_75t_R _28761_ (.A(_00605_),
    .B(_08764_),
    .Y(_08811_));
 OA21x2_ASAP7_75t_R _28762_ (.A1(_08682_),
    .A2(_08810_),
    .B(_08811_),
    .Y(_02861_));
 AO221x1_ASAP7_75t_R _28763_ (.A1(net86),
    .A2(_08560_),
    .B1(_08563_),
    .B2(net77),
    .C(_08566_),
    .Y(_08812_));
 INVx1_ASAP7_75t_R _28764_ (.A(_01499_),
    .Y(_08813_));
 INVx1_ASAP7_75t_R _28765_ (.A(_01484_),
    .Y(_08814_));
 AO221x1_ASAP7_75t_R _28766_ (.A1(_08813_),
    .A2(_08603_),
    .B1(_08604_),
    .B2(_08814_),
    .C(_08570_),
    .Y(_08815_));
 INVx1_ASAP7_75t_R _28767_ (.A(net96),
    .Y(_08816_));
 OAI22x1_ASAP7_75t_R _28768_ (.A1(_08816_),
    .A2(_08564_),
    .B1(_08577_),
    .B2(_01490_),
    .Y(_08817_));
 AO222x2_ASAP7_75t_R _28769_ (.A1(net101),
    .A2(_08581_),
    .B1(_08812_),
    .B2(_08815_),
    .C1(_08817_),
    .C2(_08575_),
    .Y(_08818_));
 AND2x2_ASAP7_75t_R _28770_ (.A(_08632_),
    .B(_08524_),
    .Y(_08819_));
 OA21x2_ASAP7_75t_R _28771_ (.A1(_08412_),
    .A2(_08819_),
    .B(_08777_),
    .Y(_08820_));
 OAI22x1_ASAP7_75t_R _28772_ (.A1(_00311_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00310_),
    .Y(_08821_));
 AO22x1_ASAP7_75t_R _28773_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_08393_),
    .B1(_08670_),
    .B2(_02260_),
    .Y(_08822_));
 AO21x1_ASAP7_75t_R _28774_ (.A1(_08663_),
    .A2(_08821_),
    .B(_08822_),
    .Y(_08823_));
 OA21x2_ASAP7_75t_R _28775_ (.A1(_00157_),
    .A2(_02328_),
    .B(_00166_),
    .Y(_08824_));
 OA21x2_ASAP7_75t_R _28776_ (.A1(_00165_),
    .A2(_08824_),
    .B(_00172_),
    .Y(_08825_));
 XOR2x2_ASAP7_75t_R _28777_ (.A(_00171_),
    .B(_08825_),
    .Y(_08826_));
 BUFx4f_ASAP7_75t_R _28778_ (.A(_08549_),
    .Y(_08827_));
 AO21x1_ASAP7_75t_R _28779_ (.A1(net2004),
    .A2(_08827_),
    .B(_05566_),
    .Y(_08828_));
 OA211x2_ASAP7_75t_R _28780_ (.A1(_08548_),
    .A2(_08826_),
    .B(_08828_),
    .C(_05515_),
    .Y(_08829_));
 AO21x1_ASAP7_75t_R _28781_ (.A1(_08377_),
    .A2(_08823_),
    .B(_08829_),
    .Y(_08830_));
 BUFx4f_ASAP7_75t_R _28782_ (.A(_08805_),
    .Y(_08831_));
 AO21x1_ASAP7_75t_R _28783_ (.A1(_08618_),
    .A2(_08619_),
    .B(_08466_),
    .Y(_08832_));
 OA211x2_ASAP7_75t_R _28784_ (.A1(_08477_),
    .A2(_08778_),
    .B(_08832_),
    .C(_08482_),
    .Y(_08833_));
 AO21x1_ASAP7_75t_R _28785_ (.A1(_08734_),
    .A2(_08735_),
    .B(_08531_),
    .Y(_08834_));
 OA211x2_ASAP7_75t_R _28786_ (.A1(_08467_),
    .A2(_08779_),
    .B(_08834_),
    .C(_08657_),
    .Y(_08835_));
 OR3x1_ASAP7_75t_R _28787_ (.A(_08626_),
    .B(_08627_),
    .C(_08427_),
    .Y(_08836_));
 OA31x2_ASAP7_75t_R _28788_ (.A1(_08508_),
    .A2(_08833_),
    .A3(_08835_),
    .B1(_08836_),
    .Y(_08837_));
 NAND2x1_ASAP7_75t_R _28789_ (.A(_08426_),
    .B(_08527_),
    .Y(_08838_));
 AND2x2_ASAP7_75t_R _28790_ (.A(_08705_),
    .B(_08706_),
    .Y(_08839_));
 AND3x1_ASAP7_75t_R _28791_ (.A(_08531_),
    .B(_08708_),
    .C(_08709_),
    .Y(_08840_));
 AO32x1_ASAP7_75t_R _28792_ (.A1(_08527_),
    .A2(_08715_),
    .A3(_08716_),
    .B1(_08419_),
    .B2(_08418_),
    .Y(_08841_));
 AO211x2_ASAP7_75t_R _28793_ (.A1(_08737_),
    .A2(_08738_),
    .B(_08657_),
    .C(_08467_),
    .Y(_08842_));
 OA221x2_ASAP7_75t_R _28794_ (.A1(_08838_),
    .A2(_08839_),
    .B1(_08840_),
    .B2(_08841_),
    .C(_08842_),
    .Y(_08843_));
 AO22x1_ASAP7_75t_R _28795_ (.A1(_08637_),
    .A2(_08731_),
    .B1(_08725_),
    .B2(_08646_),
    .Y(_08844_));
 OA21x2_ASAP7_75t_R _28796_ (.A1(_08712_),
    .A2(_08713_),
    .B(_08640_),
    .Y(_08845_));
 AOI211x1_ASAP7_75t_R _28797_ (.A1(_08643_),
    .A2(_08728_),
    .B(_08844_),
    .C(_08845_),
    .Y(_08846_));
 AO222x2_ASAP7_75t_R _28798_ (.A1(_08433_),
    .A2(_08837_),
    .B1(_08843_),
    .B2(_08636_),
    .C1(_08846_),
    .C2(_08632_),
    .Y(_08847_));
 AO21x1_ASAP7_75t_R _28799_ (.A1(_08831_),
    .A2(_08847_),
    .B(_06582_),
    .Y(_08848_));
 OR4x2_ASAP7_75t_R _28800_ (.A(_08683_),
    .B(_08820_),
    .C(_08830_),
    .D(_08848_),
    .Y(_08849_));
 OA21x2_ASAP7_75t_R _28801_ (.A1(_08600_),
    .A2(_08818_),
    .B(_08849_),
    .Y(_08850_));
 BUFx6f_ASAP7_75t_R _28802_ (.A(_08850_),
    .Y(_08851_));
 NAND2x1_ASAP7_75t_R _28803_ (.A(_00635_),
    .B(_08764_),
    .Y(_08852_));
 OA21x2_ASAP7_75t_R _28804_ (.A1(_08682_),
    .A2(_08851_),
    .B(_08852_),
    .Y(_02862_));
 OR2x2_ASAP7_75t_R _28805_ (.A(_08432_),
    .B(_08465_),
    .Y(_08853_));
 AND3x1_ASAP7_75t_R _28806_ (.A(_08508_),
    .B(_08506_),
    .C(_08615_),
    .Y(_08854_));
 OAI22x1_ASAP7_75t_R _28807_ (.A1(_00313_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00312_),
    .Y(_08855_));
 AO32x1_ASAP7_75t_R _28808_ (.A1(_15414_),
    .A2(_15416_),
    .A3(_08360_),
    .B1(_08380_),
    .B2(_02261_),
    .Y(_08856_));
 AO21x1_ASAP7_75t_R _28809_ (.A1(_08381_),
    .A2(_08855_),
    .B(_08856_),
    .Y(_08857_));
 AO221x1_ASAP7_75t_R _28810_ (.A1(_08541_),
    .A2(_08507_),
    .B1(_08853_),
    .B2(_08854_),
    .C(_08857_),
    .Y(_08858_));
 NAND2x1_ASAP7_75t_R _28811_ (.A(_08376_),
    .B(_08858_),
    .Y(_08859_));
 NAND2x1_ASAP7_75t_R _28812_ (.A(_08481_),
    .B(_08837_),
    .Y(_08860_));
 AND3x4_ASAP7_75t_R _28813_ (.A(_08401_),
    .B(_08403_),
    .C(_08649_),
    .Y(_08861_));
 INVx1_ASAP7_75t_R _28814_ (.A(_08861_),
    .Y(_08862_));
 AO21x1_ASAP7_75t_R _28815_ (.A1(_08860_),
    .A2(_08862_),
    .B(_08423_),
    .Y(_08863_));
 OA21x2_ASAP7_75t_R _28816_ (.A1(_00167_),
    .A2(_00165_),
    .B(_00172_),
    .Y(_08864_));
 OA21x2_ASAP7_75t_R _28817_ (.A1(_00171_),
    .A2(_08864_),
    .B(_00179_),
    .Y(_08865_));
 XOR2x2_ASAP7_75t_R _28818_ (.A(_00178_),
    .B(_08865_),
    .Y(_08866_));
 AO21x1_ASAP7_75t_R _28819_ (.A1(_08753_),
    .A2(_08550_),
    .B(_05571_),
    .Y(_08867_));
 OA211x2_ASAP7_75t_R _28820_ (.A1(_08547_),
    .A2(_08866_),
    .B(_08867_),
    .C(_05514_),
    .Y(_08868_));
 NOR2x1_ASAP7_75t_R _28821_ (.A(_06607_),
    .B(_08868_),
    .Y(_08869_));
 AND4x2_ASAP7_75t_R _28822_ (.A(_08599_),
    .B(_08859_),
    .C(_08863_),
    .D(_08869_),
    .Y(_08870_));
 AND2x2_ASAP7_75t_R _28823_ (.A(net101),
    .B(_08559_),
    .Y(_08871_));
 AOI21x1_ASAP7_75t_R _28824_ (.A1(net77),
    .A2(_08562_),
    .B(_08871_),
    .Y(_08872_));
 INVx1_ASAP7_75t_R _28825_ (.A(net86),
    .Y(_08873_));
 NAND2x1_ASAP7_75t_R _28826_ (.A(_08873_),
    .B(_08559_),
    .Y(_08874_));
 OA21x2_ASAP7_75t_R _28827_ (.A1(net96),
    .A2(_08559_),
    .B(_08874_),
    .Y(_08875_));
 NOR2x1_ASAP7_75t_R _28828_ (.A(_08557_),
    .B(_08875_),
    .Y(_08876_));
 AO21x1_ASAP7_75t_R _28829_ (.A1(_08557_),
    .A2(_08872_),
    .B(_08876_),
    .Y(_08877_));
 OR3x1_ASAP7_75t_R _28830_ (.A(_01511_),
    .B(_08564_),
    .C(_08877_),
    .Y(_08878_));
 BUFx3_ASAP7_75t_R _28831_ (.A(_08878_),
    .Y(_08879_));
 BUFx4f_ASAP7_75t_R _28832_ (.A(_08572_),
    .Y(_08880_));
 BUFx4f_ASAP7_75t_R _28833_ (.A(_08574_),
    .Y(_08881_));
 NAND2x1_ASAP7_75t_R _28834_ (.A(net102),
    .B(_08573_),
    .Y(_08882_));
 OAI21x1_ASAP7_75t_R _28835_ (.A1(_01483_),
    .A2(_08881_),
    .B(_08882_),
    .Y(_08883_));
 NAND2x1_ASAP7_75t_R _28836_ (.A(_01498_),
    .B(_08573_),
    .Y(_08884_));
 BUFx4f_ASAP7_75t_R _28837_ (.A(_08558_),
    .Y(_08885_));
 OA211x2_ASAP7_75t_R _28838_ (.A1(net48),
    .A2(_08574_),
    .B(_08884_),
    .C(_08885_),
    .Y(_08886_));
 AO21x1_ASAP7_75t_R _28839_ (.A1(_08880_),
    .A2(_08883_),
    .B(_08886_),
    .Y(_08887_));
 AND2x2_ASAP7_75t_R _28840_ (.A(net87),
    .B(_08573_),
    .Y(_08888_));
 AO21x1_ASAP7_75t_R _28841_ (.A1(net48),
    .A2(_08562_),
    .B(_08888_),
    .Y(_08889_));
 INVx1_ASAP7_75t_R _28842_ (.A(net78),
    .Y(_08890_));
 OA21x2_ASAP7_75t_R _28843_ (.A1(_08890_),
    .A2(_08573_),
    .B(_08882_),
    .Y(_08891_));
 NAND2x1_ASAP7_75t_R _28844_ (.A(_08572_),
    .B(_08891_),
    .Y(_08892_));
 OA211x2_ASAP7_75t_R _28845_ (.A1(_08880_),
    .A2(_08889_),
    .B(_08892_),
    .C(_05750_),
    .Y(_08893_));
 AOI21x1_ASAP7_75t_R _28846_ (.A1(_08566_),
    .A2(_08887_),
    .B(_08893_),
    .Y(_08894_));
 AND3x2_ASAP7_75t_R _28847_ (.A(_08344_),
    .B(_08879_),
    .C(_08894_),
    .Y(_08895_));
 OR2x2_ASAP7_75t_R _28848_ (.A(_08870_),
    .B(_08895_),
    .Y(_08896_));
 BUFx2_ASAP7_75t_R _28849_ (.A(_08896_),
    .Y(_08897_));
 BUFx10_ASAP7_75t_R _28850_ (.A(_08897_),
    .Y(_08898_));
 OR2x2_ASAP7_75t_R _28851_ (.A(_00665_),
    .B(_08597_),
    .Y(_08899_));
 OAI21x1_ASAP7_75t_R _28852_ (.A1(_08682_),
    .A2(_08898_),
    .B(_08899_),
    .Y(_02863_));
 INVx1_ASAP7_75t_R _28853_ (.A(net103),
    .Y(_08900_));
 INVx1_ASAP7_75t_R _28854_ (.A(_08581_),
    .Y(_08901_));
 BUFx4f_ASAP7_75t_R _28855_ (.A(_08574_),
    .Y(_08902_));
 AOI22x1_ASAP7_75t_R _28856_ (.A1(net88),
    .A2(_08574_),
    .B1(_08563_),
    .B2(net79),
    .Y(_08903_));
 OR3x1_ASAP7_75t_R _28857_ (.A(_01497_),
    .B(_08557_),
    .C(_08561_),
    .Y(_08904_));
 OA211x2_ASAP7_75t_R _28858_ (.A1(_01482_),
    .A2(_08558_),
    .B(_05749_),
    .C(_08904_),
    .Y(_08905_));
 AO21x1_ASAP7_75t_R _28859_ (.A1(_05750_),
    .A2(_08903_),
    .B(_08905_),
    .Y(_08906_));
 OR2x2_ASAP7_75t_R _28860_ (.A(_08902_),
    .B(_08906_),
    .Y(_08907_));
 BUFx4f_ASAP7_75t_R _28861_ (.A(_08562_),
    .Y(_08908_));
 NAND2x1_ASAP7_75t_R _28862_ (.A(net82),
    .B(_08908_),
    .Y(_08909_));
 BUFx3_ASAP7_75t_R _28863_ (.A(_08572_),
    .Y(_08910_));
 AO21x1_ASAP7_75t_R _28864_ (.A1(_08906_),
    .A2(_08909_),
    .B(_08910_),
    .Y(_08911_));
 OA211x2_ASAP7_75t_R _28865_ (.A1(_08900_),
    .A2(_08901_),
    .B(_08907_),
    .C(_08911_),
    .Y(_08912_));
 OA211x2_ASAP7_75t_R _28866_ (.A1(_08577_),
    .A2(_08912_),
    .B(_08879_),
    .C(_08683_),
    .Y(_08913_));
 NAND2x2_ASAP7_75t_R _28867_ (.A(_08481_),
    .B(_08795_),
    .Y(_08914_));
 OAI22x1_ASAP7_75t_R _28868_ (.A1(_00315_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00314_),
    .Y(_08915_));
 AO22x1_ASAP7_75t_R _28869_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_08393_),
    .B1(_08395_),
    .B2(_02262_),
    .Y(_08916_));
 AO21x1_ASAP7_75t_R _28870_ (.A1(_08663_),
    .A2(_08915_),
    .B(_08916_),
    .Y(_08917_));
 AOI22x1_ASAP7_75t_R _28871_ (.A1(_08616_),
    .A2(_08914_),
    .B1(_08917_),
    .B2(_08377_),
    .Y(_08918_));
 OA21x2_ASAP7_75t_R _28872_ (.A1(_08626_),
    .A2(_08627_),
    .B(_08432_),
    .Y(_08919_));
 OAI21x1_ASAP7_75t_R _28873_ (.A1(_08714_),
    .A2(_08717_),
    .B(_08482_),
    .Y(_08920_));
 AOI21x1_ASAP7_75t_R _28874_ (.A1(_08729_),
    .A2(_08730_),
    .B(_08467_),
    .Y(_08921_));
 AO221x1_ASAP7_75t_R _28875_ (.A1(_08418_),
    .A2(_08419_),
    .B1(_08467_),
    .B2(_08728_),
    .C(_08921_),
    .Y(_08922_));
 NAND2x1_ASAP7_75t_R _28876_ (.A(_08920_),
    .B(_08922_),
    .Y(_08923_));
 AO211x2_ASAP7_75t_R _28877_ (.A1(_08705_),
    .A2(_08706_),
    .B(_08426_),
    .C(_08466_),
    .Y(_08924_));
 AO21x1_ASAP7_75t_R _28878_ (.A1(_08708_),
    .A2(_08709_),
    .B(_08655_),
    .Y(_08925_));
 AO211x2_ASAP7_75t_R _28879_ (.A1(_08734_),
    .A2(_08735_),
    .B(_08497_),
    .C(_08466_),
    .Y(_08926_));
 AO211x2_ASAP7_75t_R _28880_ (.A1(_08737_),
    .A2(_08738_),
    .B(_08497_),
    .C(_08531_),
    .Y(_08927_));
 AND4x2_ASAP7_75t_R _28881_ (.A(_08924_),
    .B(_08925_),
    .C(_08926_),
    .D(_08927_),
    .Y(_08928_));
 AND3x1_ASAP7_75t_R _28882_ (.A(_08502_),
    .B(_08504_),
    .C(_08615_),
    .Y(_08929_));
 OA21x2_ASAP7_75t_R _28883_ (.A1(_08432_),
    .A2(_08928_),
    .B(_08929_),
    .Y(_08930_));
 AO221x2_ASAP7_75t_R _28884_ (.A1(_08919_),
    .A2(_08780_),
    .B1(_08923_),
    .B2(_08632_),
    .C(_08930_),
    .Y(_08931_));
 AND2x2_ASAP7_75t_R _28885_ (.A(_08753_),
    .B(_08549_),
    .Y(_08932_));
 OA21x2_ASAP7_75t_R _28886_ (.A1(_00171_),
    .A2(_08825_),
    .B(_00179_),
    .Y(_08933_));
 OA21x2_ASAP7_75t_R _28887_ (.A1(_00178_),
    .A2(_08933_),
    .B(_00187_),
    .Y(_08934_));
 XNOR2x1_ASAP7_75t_R _28888_ (.B(_08934_),
    .Y(_08935_),
    .A(_00186_));
 OR3x2_ASAP7_75t_R _28889_ (.A(_08753_),
    .B(_13601_),
    .C(_14923_),
    .Y(_08936_));
 NAND2x1_ASAP7_75t_R _28890_ (.A(_08551_),
    .B(_08936_),
    .Y(_08937_));
 AO221x1_ASAP7_75t_R _28891_ (.A1(_08932_),
    .A2(_08935_),
    .B1(_08937_),
    .B2(_00812_),
    .C(_05141_),
    .Y(_08938_));
 INVx2_ASAP7_75t_R _28892_ (.A(_08938_),
    .Y(_08939_));
 AOI211x1_ASAP7_75t_R _28893_ (.A1(_08831_),
    .A2(_08931_),
    .B(_08939_),
    .C(_06625_),
    .Y(_08940_));
 AND3x4_ASAP7_75t_R _28894_ (.A(_08694_),
    .B(_08918_),
    .C(_08940_),
    .Y(_08941_));
 NOR2x2_ASAP7_75t_R _28895_ (.A(_08913_),
    .B(_08941_),
    .Y(_08942_));
 BUFx6f_ASAP7_75t_R _28896_ (.A(_08942_),
    .Y(_08943_));
 NAND2x1_ASAP7_75t_R _28897_ (.A(_00695_),
    .B(_08764_),
    .Y(_08944_));
 OA21x2_ASAP7_75t_R _28898_ (.A1(_08682_),
    .A2(_08943_),
    .B(_08944_),
    .Y(_02864_));
 BUFx4f_ASAP7_75t_R _28899_ (.A(_08880_),
    .Y(_08945_));
 INVx1_ASAP7_75t_R _28900_ (.A(net89),
    .Y(_08946_));
 BUFx3_ASAP7_75t_R _28901_ (.A(_08580_),
    .Y(_08947_));
 NOR2x1_ASAP7_75t_R _28902_ (.A(net93),
    .B(_08902_),
    .Y(_08948_));
 AO21x1_ASAP7_75t_R _28903_ (.A1(_08946_),
    .A2(_08947_),
    .B(_08948_),
    .Y(_08949_));
 BUFx4f_ASAP7_75t_R _28904_ (.A(_08572_),
    .Y(_08950_));
 INVx1_ASAP7_75t_R _28905_ (.A(net49),
    .Y(_08951_));
 NAND2x1_ASAP7_75t_R _28906_ (.A(_08951_),
    .B(_08881_),
    .Y(_08952_));
 OA21x2_ASAP7_75t_R _28907_ (.A1(net80),
    .A2(_08902_),
    .B(_08952_),
    .Y(_08953_));
 NAND2x1_ASAP7_75t_R _28908_ (.A(_08950_),
    .B(_08953_),
    .Y(_08954_));
 OA21x2_ASAP7_75t_R _28909_ (.A1(_08945_),
    .A2(_08949_),
    .B(_08954_),
    .Y(_08955_));
 BUFx4f_ASAP7_75t_R _28910_ (.A(_08881_),
    .Y(_08956_));
 AOI211x1_ASAP7_75t_R _28911_ (.A1(_01496_),
    .A2(_08956_),
    .B(_08948_),
    .C(_08945_),
    .Y(_08957_));
 INVx1_ASAP7_75t_R _28912_ (.A(_01504_),
    .Y(_08958_));
 OA211x2_ASAP7_75t_R _28913_ (.A1(_08958_),
    .A2(_08956_),
    .B(_08952_),
    .C(_08950_),
    .Y(_08959_));
 OAI21x1_ASAP7_75t_R _28914_ (.A1(_08957_),
    .A2(_08959_),
    .B(_08685_),
    .Y(_08960_));
 OA211x2_ASAP7_75t_R _28915_ (.A1(_05749_),
    .A2(_08955_),
    .B(_08960_),
    .C(_08879_),
    .Y(_08961_));
 OAI22x1_ASAP7_75t_R _28916_ (.A1(_00317_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00316_),
    .Y(_08962_));
 AO22x1_ASAP7_75t_R _28917_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_08360_),
    .B1(_08380_),
    .B2(_02263_),
    .Y(_08963_));
 AO21x1_ASAP7_75t_R _28918_ (.A1(_08381_),
    .A2(_08962_),
    .B(_08963_),
    .Y(_08964_));
 AO21x1_ASAP7_75t_R _28919_ (.A1(_08429_),
    .A2(_08861_),
    .B(_08964_),
    .Y(_08965_));
 AND2x4_ASAP7_75t_R _28920_ (.A(_08366_),
    .B(_08480_),
    .Y(_08966_));
 AND3x1_ASAP7_75t_R _28921_ (.A(_08508_),
    .B(_08750_),
    .C(_08966_),
    .Y(_08967_));
 AND3x1_ASAP7_75t_R _28922_ (.A(_08366_),
    .B(_08632_),
    .C(_08746_),
    .Y(_08968_));
 OR3x1_ASAP7_75t_R _28923_ (.A(_08965_),
    .B(_08967_),
    .C(_08968_),
    .Y(_08969_));
 OR4x1_ASAP7_75t_R _28924_ (.A(_08458_),
    .B(_08435_),
    .C(_08443_),
    .D(_08445_),
    .Y(_08970_));
 OAI21x1_ASAP7_75t_R _28925_ (.A1(_08529_),
    .A2(_08530_),
    .B(_08422_),
    .Y(_08971_));
 AO211x2_ASAP7_75t_R _28926_ (.A1(_08537_),
    .A2(_08538_),
    .B(_08497_),
    .C(_08463_),
    .Y(_08972_));
 AO211x2_ASAP7_75t_R _28927_ (.A1(_08534_),
    .A2(_08535_),
    .B(_08425_),
    .C(_08435_),
    .Y(_08973_));
 AND4x1_ASAP7_75t_R _28928_ (.A(_08970_),
    .B(_08971_),
    .C(_08972_),
    .D(_08973_),
    .Y(_08974_));
 OR3x1_ASAP7_75t_R _28929_ (.A(_08441_),
    .B(_08437_),
    .C(_08439_),
    .Y(_08975_));
 AO211x2_ASAP7_75t_R _28930_ (.A1(_08452_),
    .A2(_08457_),
    .B(_08497_),
    .C(_08463_),
    .Y(_08976_));
 AO211x2_ASAP7_75t_R _28931_ (.A1(_08460_),
    .A2(_08461_),
    .B(_08425_),
    .C(_08435_),
    .Y(_08977_));
 AO211x2_ASAP7_75t_R _28932_ (.A1(_08513_),
    .A2(_08514_),
    .B(_08458_),
    .C(_08435_),
    .Y(_08978_));
 AND4x2_ASAP7_75t_R _28933_ (.A(_08975_),
    .B(_08976_),
    .C(_08977_),
    .D(_08978_),
    .Y(_08979_));
 OA21x2_ASAP7_75t_R _28934_ (.A1(_08433_),
    .A2(_08979_),
    .B(_08929_),
    .Y(_08980_));
 AO221x1_ASAP7_75t_R _28935_ (.A1(_08919_),
    .A2(_08700_),
    .B1(_08974_),
    .B2(_08632_),
    .C(_08980_),
    .Y(_08981_));
 AOI22x1_ASAP7_75t_R _28936_ (.A1(_08377_),
    .A2(_08969_),
    .B1(_08981_),
    .B2(_08542_),
    .Y(_08982_));
 OA21x2_ASAP7_75t_R _28937_ (.A1(_00178_),
    .A2(_08865_),
    .B(_00187_),
    .Y(_08983_));
 OA21x2_ASAP7_75t_R _28938_ (.A1(_00186_),
    .A2(_08983_),
    .B(_00193_),
    .Y(_08984_));
 XNOR2x2_ASAP7_75t_R _28939_ (.A(_00192_),
    .B(_08984_),
    .Y(_08985_));
 AO221x2_ASAP7_75t_R _28940_ (.A1(_00815_),
    .A2(_08937_),
    .B1(_08985_),
    .B2(_08932_),
    .C(_05141_),
    .Y(_08986_));
 AND5x2_ASAP7_75t_R _28941_ (.A(_05933_),
    .B(_05953_),
    .C(_08599_),
    .D(_08982_),
    .E(_08986_),
    .Y(_08987_));
 AOI21x1_ASAP7_75t_R _28942_ (.A1(_08684_),
    .A2(_08961_),
    .B(_08987_),
    .Y(_08988_));
 BUFx6f_ASAP7_75t_R _28943_ (.A(_08988_),
    .Y(_08989_));
 BUFx10_ASAP7_75t_R _28944_ (.A(_08680_),
    .Y(_08990_));
 NAND2x1_ASAP7_75t_R _28945_ (.A(_00725_),
    .B(_08990_),
    .Y(_08991_));
 OA21x2_ASAP7_75t_R _28946_ (.A1(_08682_),
    .A2(_08989_),
    .B(_08991_),
    .Y(_02865_));
 INVx1_ASAP7_75t_R _28947_ (.A(net90),
    .Y(_08992_));
 NOR2x1_ASAP7_75t_R _28948_ (.A(net97),
    .B(_08574_),
    .Y(_08993_));
 AO21x1_ASAP7_75t_R _28949_ (.A1(_08992_),
    .A2(_08580_),
    .B(_08993_),
    .Y(_08994_));
 INVx1_ASAP7_75t_R _28950_ (.A(net50),
    .Y(_08995_));
 NAND2x1_ASAP7_75t_R _28951_ (.A(_08995_),
    .B(_08580_),
    .Y(_08996_));
 OA21x2_ASAP7_75t_R _28952_ (.A1(net81),
    .A2(_08881_),
    .B(_08996_),
    .Y(_08997_));
 NAND2x1_ASAP7_75t_R _28953_ (.A(_08950_),
    .B(_08997_),
    .Y(_08998_));
 OA21x2_ASAP7_75t_R _28954_ (.A1(_08945_),
    .A2(_08994_),
    .B(_08998_),
    .Y(_08999_));
 AOI211x1_ASAP7_75t_R _28955_ (.A1(_01495_),
    .A2(_08956_),
    .B(_08993_),
    .C(_08950_),
    .Y(_09000_));
 INVx1_ASAP7_75t_R _28956_ (.A(_01503_),
    .Y(_09001_));
 OA211x2_ASAP7_75t_R _28957_ (.A1(_09001_),
    .A2(_08956_),
    .B(_08996_),
    .C(_08910_),
    .Y(_09002_));
 OAI21x1_ASAP7_75t_R _28958_ (.A1(_09000_),
    .A2(_09002_),
    .B(_08685_),
    .Y(_09003_));
 OA211x2_ASAP7_75t_R _28959_ (.A1(_05749_),
    .A2(_08999_),
    .B(_09003_),
    .C(_08879_),
    .Y(_09004_));
 OR2x2_ASAP7_75t_R _28960_ (.A(_08508_),
    .B(_08660_),
    .Y(_09005_));
 OA21x2_ASAP7_75t_R _28961_ (.A1(_08786_),
    .A2(_08651_),
    .B(_09005_),
    .Y(_09006_));
 AO21x1_ASAP7_75t_R _28962_ (.A1(_08705_),
    .A2(_08706_),
    .B(_08655_),
    .Y(_09007_));
 AO211x2_ASAP7_75t_R _28963_ (.A1(_08734_),
    .A2(_08735_),
    .B(_08657_),
    .C(_08477_),
    .Y(_09008_));
 AO211x2_ASAP7_75t_R _28964_ (.A1(_08737_),
    .A2(_08738_),
    .B(_08426_),
    .C(_08527_),
    .Y(_09009_));
 OR4x1_ASAP7_75t_R _28965_ (.A(_08657_),
    .B(_08527_),
    .C(_08741_),
    .D(_08743_),
    .Y(_09010_));
 AND4x2_ASAP7_75t_R _28966_ (.A(_09007_),
    .B(_09008_),
    .C(_09009_),
    .D(_09010_),
    .Y(_09011_));
 NAND2x1_ASAP7_75t_R _28967_ (.A(_08633_),
    .B(_08477_),
    .Y(_09012_));
 NOR2x1_ASAP7_75t_R _28968_ (.A(_08712_),
    .B(_08713_),
    .Y(_09013_));
 AO31x2_ASAP7_75t_R _28969_ (.A1(_08467_),
    .A2(_08715_),
    .A3(_08716_),
    .B(_08657_),
    .Y(_09014_));
 AO21x1_ASAP7_75t_R _28970_ (.A1(_08729_),
    .A2(_08730_),
    .B(_08655_),
    .Y(_09015_));
 OA221x2_ASAP7_75t_R _28971_ (.A1(_09012_),
    .A2(_09013_),
    .B1(_08840_),
    .B2(_09014_),
    .C(_09015_),
    .Y(_09016_));
 AOI22x1_ASAP7_75t_R _28972_ (.A1(_08636_),
    .A2(_09011_),
    .B1(_09016_),
    .B2(_08632_),
    .Y(_09017_));
 OAI21x1_ASAP7_75t_R _28973_ (.A1(_08481_),
    .A2(_08629_),
    .B(_09017_),
    .Y(_09018_));
 OAI22x1_ASAP7_75t_R _28974_ (.A1(_00319_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00318_),
    .Y(_09019_));
 AO22x1_ASAP7_75t_R _28975_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_08669_),
    .B1(_08670_),
    .B2(_02264_),
    .Y(_09020_));
 AO21x1_ASAP7_75t_R _28976_ (.A1(_08663_),
    .A2(_09019_),
    .B(_09020_),
    .Y(_09021_));
 AO21x1_ASAP7_75t_R _28977_ (.A1(_00178_),
    .A2(_00187_),
    .B(_00186_),
    .Y(_09022_));
 AO21x1_ASAP7_75t_R _28978_ (.A1(_00193_),
    .A2(_09022_),
    .B(_00192_),
    .Y(_09023_));
 AND2x2_ASAP7_75t_R _28979_ (.A(_00198_),
    .B(_09023_),
    .Y(_09024_));
 AND4x1_ASAP7_75t_R _28980_ (.A(_00179_),
    .B(_00187_),
    .C(_00193_),
    .D(_00198_),
    .Y(_09025_));
 OA21x2_ASAP7_75t_R _28981_ (.A1(_00171_),
    .A2(_08825_),
    .B(_09025_),
    .Y(_09026_));
 NOR2x1_ASAP7_75t_R _28982_ (.A(_09024_),
    .B(_09026_),
    .Y(_09027_));
 XNOR2x2_ASAP7_75t_R _28983_ (.A(_00197_),
    .B(_09027_),
    .Y(_09028_));
 NAND2x1_ASAP7_75t_R _28984_ (.A(_05506_),
    .B(_08547_),
    .Y(_09029_));
 OA211x2_ASAP7_75t_R _28985_ (.A1(_08548_),
    .A2(_09028_),
    .B(_09029_),
    .C(_05514_),
    .Y(_09030_));
 AO21x1_ASAP7_75t_R _28986_ (.A1(_08376_),
    .A2(_09021_),
    .B(_09030_),
    .Y(_09031_));
 AOI221x1_ASAP7_75t_R _28987_ (.A1(_09006_),
    .A2(_08966_),
    .B1(_09018_),
    .B2(_08831_),
    .C(_09031_),
    .Y(_09032_));
 AND2x2_ASAP7_75t_R _28988_ (.A(_05999_),
    .B(_09032_),
    .Y(_09033_));
 AND3x4_ASAP7_75t_R _28989_ (.A(_08401_),
    .B(_08403_),
    .C(_08411_),
    .Y(_09034_));
 AOI21x1_ASAP7_75t_R _28990_ (.A1(_08777_),
    .A2(_09034_),
    .B(_08345_),
    .Y(_09035_));
 AOI22x1_ASAP7_75t_R _28991_ (.A1(_08684_),
    .A2(_09004_),
    .B1(_09033_),
    .B2(_09035_),
    .Y(_09036_));
 BUFx6f_ASAP7_75t_R _28992_ (.A(_09036_),
    .Y(_09037_));
 NAND2x1_ASAP7_75t_R _28993_ (.A(_00755_),
    .B(_08990_),
    .Y(_09038_));
 OA21x2_ASAP7_75t_R _28994_ (.A1(_08682_),
    .A2(_09037_),
    .B(_09038_),
    .Y(_02866_));
 NOR2x1_ASAP7_75t_R _28995_ (.A(net98),
    .B(_08574_),
    .Y(_09039_));
 AO21x1_ASAP7_75t_R _28996_ (.A1(_08607_),
    .A2(_08580_),
    .B(_09039_),
    .Y(_09040_));
 OR2x2_ASAP7_75t_R _28997_ (.A(net51),
    .B(_08562_),
    .Y(_09041_));
 OA21x2_ASAP7_75t_R _28998_ (.A1(net83),
    .A2(_08902_),
    .B(_09041_),
    .Y(_09042_));
 NAND2x1_ASAP7_75t_R _28999_ (.A(_08950_),
    .B(_09042_),
    .Y(_09043_));
 OA21x2_ASAP7_75t_R _29000_ (.A1(_08945_),
    .A2(_09040_),
    .B(_09043_),
    .Y(_09044_));
 AOI211x1_ASAP7_75t_R _29001_ (.A1(_01493_),
    .A2(_08956_),
    .B(_09039_),
    .C(_08950_),
    .Y(_09045_));
 OA211x2_ASAP7_75t_R _29002_ (.A1(_08602_),
    .A2(_08956_),
    .B(_09041_),
    .C(_08910_),
    .Y(_09046_));
 OAI21x1_ASAP7_75t_R _29003_ (.A1(_09045_),
    .A2(_09046_),
    .B(_08685_),
    .Y(_09047_));
 OA211x2_ASAP7_75t_R _29004_ (.A1(_05749_),
    .A2(_09044_),
    .B(_09047_),
    .C(_08879_),
    .Y(_09048_));
 OR3x1_ASAP7_75t_R _29005_ (.A(_08531_),
    .B(_08517_),
    .C(_08519_),
    .Y(_09049_));
 OA21x2_ASAP7_75t_R _29006_ (.A1(_08467_),
    .A2(_08648_),
    .B(_09049_),
    .Y(_09050_));
 NAND2x1_ASAP7_75t_R _29007_ (.A(_08633_),
    .B(_09050_),
    .Y(_09051_));
 OAI22x1_ASAP7_75t_R _29008_ (.A1(_08695_),
    .A2(_08645_),
    .B1(_08653_),
    .B2(_09051_),
    .Y(_09052_));
 AO32x1_ASAP7_75t_R _29009_ (.A1(_08502_),
    .A2(_08504_),
    .A3(_08861_),
    .B1(_08650_),
    .B2(_08433_),
    .Y(_09053_));
 AO21x1_ASAP7_75t_R _29010_ (.A1(_08660_),
    .A2(_08636_),
    .B(_09053_),
    .Y(_09054_));
 NOR2x2_ASAP7_75t_R _29011_ (.A(_09052_),
    .B(_09054_),
    .Y(_09055_));
 INVx3_ASAP7_75t_R _29012_ (.A(_08375_),
    .Y(_09056_));
 OA22x2_ASAP7_75t_R _29013_ (.A1(_00321_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00320_),
    .Y(_09057_));
 AOI22x1_ASAP7_75t_R _29014_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_08393_),
    .B1(_08395_),
    .B2(_02265_),
    .Y(_09058_));
 OA21x2_ASAP7_75t_R _29015_ (.A1(_08395_),
    .A2(_09057_),
    .B(_09058_),
    .Y(_09059_));
 OR5x2_ASAP7_75t_R _29016_ (.A(_08626_),
    .B(_08627_),
    .C(_08617_),
    .D(_08620_),
    .E(_08624_),
    .Y(_09060_));
 OAI21x1_ASAP7_75t_R _29017_ (.A1(_08508_),
    .A2(_09011_),
    .B(_09060_),
    .Y(_09061_));
 AO21x1_ASAP7_75t_R _29018_ (.A1(_08401_),
    .A2(_08403_),
    .B(_08423_),
    .Y(_09062_));
 AND3x1_ASAP7_75t_R _29019_ (.A(_00193_),
    .B(_00198_),
    .C(_00206_),
    .Y(_09063_));
 OA21x2_ASAP7_75t_R _29020_ (.A1(_00186_),
    .A2(_08983_),
    .B(_09063_),
    .Y(_09064_));
 AND3x1_ASAP7_75t_R _29021_ (.A(_00192_),
    .B(_00198_),
    .C(_00206_),
    .Y(_09065_));
 AO21x1_ASAP7_75t_R _29022_ (.A1(_00197_),
    .A2(_00206_),
    .B(_09065_),
    .Y(_09066_));
 OR2x2_ASAP7_75t_R _29023_ (.A(_09064_),
    .B(_09066_),
    .Y(_09067_));
 XNOR2x2_ASAP7_75t_R _29024_ (.A(net2022),
    .B(_09067_),
    .Y(_09068_));
 AND3x1_ASAP7_75t_R _29025_ (.A(_13595_),
    .B(_08827_),
    .C(_09068_),
    .Y(_09069_));
 AO21x2_ASAP7_75t_R _29026_ (.A1(_00821_),
    .A2(_08548_),
    .B(_09069_),
    .Y(_09070_));
 OA222x2_ASAP7_75t_R _29027_ (.A1(_09056_),
    .A2(_09059_),
    .B1(_09061_),
    .B2(_09062_),
    .C1(_09070_),
    .C2(_05141_),
    .Y(_09071_));
 OA211x2_ASAP7_75t_R _29028_ (.A1(_08806_),
    .A2(_09055_),
    .B(_09071_),
    .C(_06016_),
    .Y(_09072_));
 AOI22x1_ASAP7_75t_R _29029_ (.A1(_08684_),
    .A2(_09048_),
    .B1(_09072_),
    .B2(_09035_),
    .Y(_09073_));
 BUFx4f_ASAP7_75t_R _29030_ (.A(_09073_),
    .Y(_09074_));
 NAND2x1_ASAP7_75t_R _29031_ (.A(_00451_),
    .B(_08990_),
    .Y(_09075_));
 OA21x2_ASAP7_75t_R _29032_ (.A1(_08682_),
    .A2(_09074_),
    .B(_09075_),
    .Y(_02867_));
 OR2x2_ASAP7_75t_R _29033_ (.A(_08509_),
    .B(_08979_),
    .Y(_09076_));
 OA21x2_ASAP7_75t_R _29034_ (.A1(_08786_),
    .A2(_08700_),
    .B(_09076_),
    .Y(_09077_));
 OAI22x1_ASAP7_75t_R _29035_ (.A1(_00323_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00322_),
    .Y(_09078_));
 AO22x1_ASAP7_75t_R _29036_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_08393_),
    .B1(_08670_),
    .B2(_02266_),
    .Y(_09079_));
 AO21x1_ASAP7_75t_R _29037_ (.A1(_08663_),
    .A2(_09078_),
    .B(_09079_),
    .Y(_09080_));
 OR3x1_ASAP7_75t_R _29038_ (.A(_00197_),
    .B(_09024_),
    .C(_09026_),
    .Y(_09081_));
 AO21x1_ASAP7_75t_R _29039_ (.A1(_00206_),
    .A2(_09081_),
    .B(net2022),
    .Y(_09082_));
 NAND2x1_ASAP7_75t_R _29040_ (.A(_00211_),
    .B(_09082_),
    .Y(_09083_));
 XNOR2x2_ASAP7_75t_R _29041_ (.A(_00210_),
    .B(_09083_),
    .Y(_09084_));
 AO21x1_ASAP7_75t_R _29042_ (.A1(_13595_),
    .A2(_08827_),
    .B(_05598_),
    .Y(_09085_));
 OA211x2_ASAP7_75t_R _29043_ (.A1(_08548_),
    .A2(_09084_),
    .B(_09085_),
    .C(_05515_),
    .Y(_09086_));
 AO21x1_ASAP7_75t_R _29044_ (.A1(_08377_),
    .A2(_09080_),
    .B(_09086_),
    .Y(_09087_));
 AOI211x1_ASAP7_75t_R _29045_ (.A1(_08966_),
    .A2(_09077_),
    .B(_09087_),
    .C(_06041_),
    .Y(_09088_));
 AND3x1_ASAP7_75t_R _29046_ (.A(_08432_),
    .B(_08633_),
    .C(_08749_),
    .Y(_09089_));
 AO221x2_ASAP7_75t_R _29047_ (.A1(_08481_),
    .A2(_08719_),
    .B1(_08861_),
    .B2(_08482_),
    .C(_09089_),
    .Y(_09090_));
 OR2x2_ASAP7_75t_R _29048_ (.A(_08433_),
    .B(_08746_),
    .Y(_09091_));
 AOI22x1_ASAP7_75t_R _29049_ (.A1(_08507_),
    .A2(_09090_),
    .B1(_09091_),
    .B2(_08854_),
    .Y(_09092_));
 AND2x2_ASAP7_75t_R _29050_ (.A(_09088_),
    .B(_09092_),
    .Y(_09093_));
 AOI22x1_ASAP7_75t_R _29051_ (.A1(net92),
    .A2(_08574_),
    .B1(_08563_),
    .B2(net84),
    .Y(_09094_));
 OR3x1_ASAP7_75t_R _29052_ (.A(_01492_),
    .B(_08557_),
    .C(_08562_),
    .Y(_09095_));
 OA211x2_ASAP7_75t_R _29053_ (.A1(_01501_),
    .A2(_08558_),
    .B(_05749_),
    .C(_09095_),
    .Y(_09096_));
 AO21x1_ASAP7_75t_R _29054_ (.A1(_05750_),
    .A2(_09094_),
    .B(_09096_),
    .Y(_09097_));
 NAND2x1_ASAP7_75t_R _29055_ (.A(net75),
    .B(_08581_),
    .Y(_09098_));
 NAND2x1_ASAP7_75t_R _29056_ (.A(net99),
    .B(_08562_),
    .Y(_09099_));
 AO21x1_ASAP7_75t_R _29057_ (.A1(_09097_),
    .A2(_09099_),
    .B(_08910_),
    .Y(_09100_));
 OA211x2_ASAP7_75t_R _29058_ (.A1(_08956_),
    .A2(_09097_),
    .B(_09098_),
    .C(_09100_),
    .Y(_09101_));
 OA211x2_ASAP7_75t_R _29059_ (.A1(_08577_),
    .A2(_09101_),
    .B(_08879_),
    .C(_08683_),
    .Y(_09102_));
 AOI21x1_ASAP7_75t_R _29060_ (.A1(_09035_),
    .A2(_09093_),
    .B(_09102_),
    .Y(_09103_));
 BUFx6f_ASAP7_75t_R _29061_ (.A(_09103_),
    .Y(_09104_));
 NAND2x1_ASAP7_75t_R _29062_ (.A(_00826_),
    .B(_08990_),
    .Y(_09105_));
 OA21x2_ASAP7_75t_R _29063_ (.A1(_08682_),
    .A2(_09104_),
    .B(_09105_),
    .Y(_02868_));
 BUFx10_ASAP7_75t_R _29064_ (.A(_08590_),
    .Y(_09106_));
 BUFx6f_ASAP7_75t_R _29065_ (.A(_09106_),
    .Y(_09107_));
 BUFx6f_ASAP7_75t_R _29066_ (.A(_08988_),
    .Y(_09108_));
 NAND2x1_ASAP7_75t_R _29067_ (.A(_01813_),
    .B(_08591_),
    .Y(_09109_));
 OA21x2_ASAP7_75t_R _29068_ (.A1(_09107_),
    .A2(_09108_),
    .B(_09109_),
    .Y(_02869_));
 AO21x2_ASAP7_75t_R _29069_ (.A1(_08401_),
    .A2(_08403_),
    .B(_08806_),
    .Y(_09110_));
 NOR2x1_ASAP7_75t_R _29070_ (.A(_08798_),
    .B(_09110_),
    .Y(_09111_));
 AO221x1_ASAP7_75t_R _29071_ (.A1(_08502_),
    .A2(_08504_),
    .B1(_08966_),
    .B2(_08928_),
    .C(_09111_),
    .Y(_09112_));
 AO21x1_ASAP7_75t_R _29072_ (.A1(_08780_),
    .A2(_08966_),
    .B(_08786_),
    .Y(_09113_));
 OA211x2_ASAP7_75t_R _29073_ (.A1(_13568_),
    .A2(_06775_),
    .B(_08646_),
    .C(_18625_),
    .Y(_09114_));
 AND4x1_ASAP7_75t_R _29074_ (.A(_13622_),
    .B(_18623_),
    .C(_08398_),
    .D(_08646_),
    .Y(_09115_));
 OAI21x1_ASAP7_75t_R _29075_ (.A1(_09114_),
    .A2(_09115_),
    .B(_08648_),
    .Y(_09116_));
 INVx1_ASAP7_75t_R _29076_ (.A(_08411_),
    .Y(_09117_));
 OR3x1_ASAP7_75t_R _29077_ (.A(_09117_),
    .B(_09114_),
    .C(_09115_),
    .Y(_09118_));
 NAND2x2_ASAP7_75t_R _29078_ (.A(_09116_),
    .B(_09118_),
    .Y(_09119_));
 AND3x1_ASAP7_75t_R _29079_ (.A(_08481_),
    .B(_08509_),
    .C(_08791_),
    .Y(_09120_));
 AO21x1_ASAP7_75t_R _29080_ (.A1(_08433_),
    .A2(_09119_),
    .B(_09120_),
    .Y(_09121_));
 AND2x4_ASAP7_75t_R _29081_ (.A(_04867_),
    .B(_08360_),
    .Y(_09122_));
 OAI22x1_ASAP7_75t_R _29082_ (.A1(_00325_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00324_),
    .Y(_09123_));
 AND2x2_ASAP7_75t_R _29083_ (.A(_02267_),
    .B(_08670_),
    .Y(_09124_));
 AO21x1_ASAP7_75t_R _29084_ (.A1(_08663_),
    .A2(_09123_),
    .B(_09124_),
    .Y(_09125_));
 OA21x2_ASAP7_75t_R _29085_ (.A1(_00205_),
    .A2(_09067_),
    .B(_00211_),
    .Y(_09126_));
 OA21x2_ASAP7_75t_R _29086_ (.A1(_00210_),
    .A2(_09126_),
    .B(_00216_),
    .Y(_09127_));
 XNOR2x2_ASAP7_75t_R _29087_ (.A(_00215_),
    .B(_09127_),
    .Y(_09128_));
 NOR2x1_ASAP7_75t_R _29088_ (.A(_08548_),
    .B(_09128_),
    .Y(_09129_));
 AO21x1_ASAP7_75t_R _29089_ (.A1(_05604_),
    .A2(_08548_),
    .B(_09129_),
    .Y(_09130_));
 AO222x2_ASAP7_75t_R _29090_ (.A1(\alu_adder_result_ex[14] ),
    .A2(_09122_),
    .B1(_09125_),
    .B2(_08376_),
    .C1(_09130_),
    .C2(_05515_),
    .Y(_09131_));
 AO21x1_ASAP7_75t_R _29091_ (.A1(_08831_),
    .A2(_09121_),
    .B(_09131_),
    .Y(_09132_));
 AOI211x1_ASAP7_75t_R _29092_ (.A1(_09112_),
    .A2(_09113_),
    .B(_06063_),
    .C(_09132_),
    .Y(_09133_));
 AO221x1_ASAP7_75t_R _29093_ (.A1(net94),
    .A2(_08574_),
    .B1(_08563_),
    .B2(net85),
    .C(_05749_),
    .Y(_09134_));
 INVx1_ASAP7_75t_R _29094_ (.A(_01491_),
    .Y(_09135_));
 AO221x1_ASAP7_75t_R _29095_ (.A1(_09135_),
    .A2(_08560_),
    .B1(_08563_),
    .B2(_08767_),
    .C(_05750_),
    .Y(_09136_));
 NAND2x1_ASAP7_75t_R _29096_ (.A(_09134_),
    .B(_09136_),
    .Y(_09137_));
 NAND2x1_ASAP7_75t_R _29097_ (.A(net76),
    .B(_08581_),
    .Y(_09138_));
 NAND2x1_ASAP7_75t_R _29098_ (.A(net100),
    .B(_08908_),
    .Y(_09139_));
 AO21x1_ASAP7_75t_R _29099_ (.A1(_09137_),
    .A2(_09139_),
    .B(_08910_),
    .Y(_09140_));
 OA211x2_ASAP7_75t_R _29100_ (.A1(_08956_),
    .A2(_09137_),
    .B(_09138_),
    .C(_09140_),
    .Y(_09141_));
 OA211x2_ASAP7_75t_R _29101_ (.A1(_08577_),
    .A2(_09141_),
    .B(_08879_),
    .C(_08683_),
    .Y(_09142_));
 AOI21x1_ASAP7_75t_R _29102_ (.A1(_09035_),
    .A2(_09133_),
    .B(_09142_),
    .Y(_09143_));
 BUFx6f_ASAP7_75t_R _29103_ (.A(_09143_),
    .Y(_09144_));
 NAND2x1_ASAP7_75t_R _29104_ (.A(_00859_),
    .B(_08990_),
    .Y(_09145_));
 OA21x2_ASAP7_75t_R _29105_ (.A1(_08682_),
    .A2(_09144_),
    .B(_09145_),
    .Y(_02870_));
 BUFx4f_ASAP7_75t_R _29106_ (.A(_08680_),
    .Y(_09146_));
 OR2x2_ASAP7_75t_R _29107_ (.A(_08786_),
    .B(_08524_),
    .Y(_09147_));
 OA211x2_ASAP7_75t_R _29108_ (.A1(_08509_),
    .A2(_08465_),
    .B(_08966_),
    .C(_09147_),
    .Y(_09148_));
 OAI22x1_ASAP7_75t_R _29109_ (.A1(_00327_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00326_),
    .Y(_09149_));
 AO22x1_ASAP7_75t_R _29110_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_08669_),
    .B1(_08394_),
    .B2(_02268_),
    .Y(_09150_));
 AO21x1_ASAP7_75t_R _29111_ (.A1(_08382_),
    .A2(_09149_),
    .B(_09150_),
    .Y(_09151_));
 AO21x1_ASAP7_75t_R _29112_ (.A1(_08429_),
    .A2(_08861_),
    .B(_09151_),
    .Y(_09152_));
 OA21x2_ASAP7_75t_R _29113_ (.A1(_09148_),
    .A2(_09152_),
    .B(_08377_),
    .Y(_09153_));
 AO21x1_ASAP7_75t_R _29114_ (.A1(_00210_),
    .A2(_00216_),
    .B(_00215_),
    .Y(_09154_));
 AND3x1_ASAP7_75t_R _29115_ (.A(_00211_),
    .B(_00216_),
    .C(_00223_),
    .Y(_09155_));
 AO22x1_ASAP7_75t_R _29116_ (.A1(_00223_),
    .A2(_09154_),
    .B1(_09155_),
    .B2(_09082_),
    .Y(_09156_));
 XOR2x2_ASAP7_75t_R _29117_ (.A(_00222_),
    .B(_09156_),
    .Y(_09157_));
 AND2x2_ASAP7_75t_R _29118_ (.A(_08932_),
    .B(_09157_),
    .Y(_09158_));
 AO21x1_ASAP7_75t_R _29119_ (.A1(_05609_),
    .A2(_08548_),
    .B(_09158_),
    .Y(_09159_));
 OA21x2_ASAP7_75t_R _29120_ (.A1(_08833_),
    .A2(_08835_),
    .B(_08480_),
    .Y(_09160_));
 OR3x1_ASAP7_75t_R _29121_ (.A(_08626_),
    .B(_08627_),
    .C(_08861_),
    .Y(_09161_));
 AO32x1_ASAP7_75t_R _29122_ (.A1(_08401_),
    .A2(_08403_),
    .A3(_08427_),
    .B1(_08504_),
    .B2(_08502_),
    .Y(_09162_));
 AO21x1_ASAP7_75t_R _29123_ (.A1(_08481_),
    .A2(_08843_),
    .B(_09162_),
    .Y(_09163_));
 OA21x2_ASAP7_75t_R _29124_ (.A1(_09160_),
    .A2(_09161_),
    .B(_09163_),
    .Y(_09164_));
 AO221x1_ASAP7_75t_R _29125_ (.A1(_05515_),
    .A2(_09159_),
    .B1(_09164_),
    .B2(_08542_),
    .C(_05078_),
    .Y(_09165_));
 OR2x2_ASAP7_75t_R _29126_ (.A(_08554_),
    .B(_06087_),
    .Y(_09166_));
 OA21x2_ASAP7_75t_R _29127_ (.A1(_09153_),
    .A2(_09165_),
    .B(_09166_),
    .Y(_09167_));
 NOR2x1_ASAP7_75t_R _29128_ (.A(net101),
    .B(_08559_),
    .Y(_09168_));
 AO21x1_ASAP7_75t_R _29129_ (.A1(_01490_),
    .A2(_08947_),
    .B(_09168_),
    .Y(_09169_));
 NAND2x1_ASAP7_75t_R _29130_ (.A(net77),
    .B(_08559_),
    .Y(_09170_));
 OA211x2_ASAP7_75t_R _29131_ (.A1(_01499_),
    .A2(_08902_),
    .B(_09170_),
    .C(_08880_),
    .Y(_09171_));
 AO21x1_ASAP7_75t_R _29132_ (.A1(_08885_),
    .A2(_09169_),
    .B(_09171_),
    .Y(_09172_));
 OAI21x1_ASAP7_75t_R _29133_ (.A1(_08873_),
    .A2(_08573_),
    .B(_09170_),
    .Y(_09173_));
 NAND2x1_ASAP7_75t_R _29134_ (.A(_08557_),
    .B(_09173_),
    .Y(_09174_));
 AO21x1_ASAP7_75t_R _29135_ (.A1(_08816_),
    .A2(_08559_),
    .B(_09168_),
    .Y(_09175_));
 OR2x2_ASAP7_75t_R _29136_ (.A(_08557_),
    .B(_09175_),
    .Y(_09176_));
 AO21x1_ASAP7_75t_R _29137_ (.A1(_09174_),
    .A2(_09176_),
    .B(_05749_),
    .Y(_09177_));
 OA211x2_ASAP7_75t_R _29138_ (.A1(_08689_),
    .A2(_09172_),
    .B(_09177_),
    .C(_08879_),
    .Y(_09178_));
 NAND2x1_ASAP7_75t_R _29139_ (.A(_08345_),
    .B(_09178_),
    .Y(_09179_));
 OA21x2_ASAP7_75t_R _29140_ (.A1(_08684_),
    .A2(_09167_),
    .B(_09179_),
    .Y(_09180_));
 BUFx6f_ASAP7_75t_R _29141_ (.A(_09180_),
    .Y(_09181_));
 NAND2x1_ASAP7_75t_R _29142_ (.A(_00892_),
    .B(_08990_),
    .Y(_09182_));
 OA21x2_ASAP7_75t_R _29143_ (.A1(_09146_),
    .A2(_09181_),
    .B(_09182_),
    .Y(_02871_));
 OA21x2_ASAP7_75t_R _29144_ (.A1(_08509_),
    .A2(_08465_),
    .B(_09147_),
    .Y(_09183_));
 INVx2_ASAP7_75t_R _29145_ (.A(_09110_),
    .Y(_09184_));
 AND3x2_ASAP7_75t_R _29146_ (.A(_05154_),
    .B(_02216_),
    .C(_08545_),
    .Y(_09185_));
 BUFx4f_ASAP7_75t_R _29147_ (.A(_09185_),
    .Y(_09186_));
 AO21x1_ASAP7_75t_R _29148_ (.A1(_00223_),
    .A2(_09154_),
    .B(_00222_),
    .Y(_09187_));
 OA31x2_ASAP7_75t_R _29149_ (.A1(net2022),
    .A2(_09064_),
    .A3(_09066_),
    .B1(_09155_),
    .Y(_09188_));
 OR2x2_ASAP7_75t_R _29150_ (.A(_09187_),
    .B(_09188_),
    .Y(_09189_));
 AND2x2_ASAP7_75t_R _29151_ (.A(_00228_),
    .B(_09189_),
    .Y(_09190_));
 XNOR2x1_ASAP7_75t_R _29152_ (.B(_09190_),
    .Y(_09191_),
    .A(net2009));
 OR2x2_ASAP7_75t_R _29153_ (.A(_00104_),
    .B(_08549_),
    .Y(_09192_));
 OAI21x1_ASAP7_75t_R _29154_ (.A1(_09186_),
    .A2(_09191_),
    .B(_09192_),
    .Y(_09193_));
 NAND2x1_ASAP7_75t_R _29155_ (.A(_13566_),
    .B(_05180_),
    .Y(_09194_));
 OA211x2_ASAP7_75t_R _29156_ (.A1(_13566_),
    .A2(_09193_),
    .B(_09194_),
    .C(_05304_),
    .Y(_09195_));
 AO21x1_ASAP7_75t_R _29157_ (.A1(_08831_),
    .A2(_09034_),
    .B(_13776_),
    .Y(_09196_));
 OAI22x1_ASAP7_75t_R _29158_ (.A1(_00329_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00328_),
    .Y(_09197_));
 AND2x2_ASAP7_75t_R _29159_ (.A(_02269_),
    .B(_08380_),
    .Y(_09198_));
 AO221x1_ASAP7_75t_R _29160_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_08669_),
    .B1(_08381_),
    .B2(_09197_),
    .C(_09198_),
    .Y(_09199_));
 OR3x1_ASAP7_75t_R _29161_ (.A(_09195_),
    .B(_09196_),
    .C(_09199_),
    .Y(_09200_));
 AO221x1_ASAP7_75t_R _29162_ (.A1(_08429_),
    .A2(_09164_),
    .B1(_09183_),
    .B2(_09184_),
    .C(_09200_),
    .Y(_09201_));
 OR2x2_ASAP7_75t_R _29163_ (.A(_08376_),
    .B(_09195_),
    .Y(_09202_));
 AO21x1_ASAP7_75t_R _29164_ (.A1(_08554_),
    .A2(_09202_),
    .B(_06109_),
    .Y(_09203_));
 AO21x2_ASAP7_75t_R _29165_ (.A1(_09201_),
    .A2(_09203_),
    .B(_08344_),
    .Y(_09204_));
 OAI21x1_ASAP7_75t_R _29166_ (.A1(_01511_),
    .A2(_09177_),
    .B(_08879_),
    .Y(_09205_));
 AND2x2_ASAP7_75t_R _29167_ (.A(net48),
    .B(_08574_),
    .Y(_09206_));
 AO21x1_ASAP7_75t_R _29168_ (.A1(net102),
    .A2(_08908_),
    .B(_09206_),
    .Y(_09207_));
 OR2x2_ASAP7_75t_R _29169_ (.A(_01498_),
    .B(_08573_),
    .Y(_09208_));
 OA211x2_ASAP7_75t_R _29170_ (.A1(_08890_),
    .A2(_08562_),
    .B(_09208_),
    .C(_08572_),
    .Y(_09209_));
 INVx1_ASAP7_75t_R _29171_ (.A(_09209_),
    .Y(_09210_));
 OA211x2_ASAP7_75t_R _29172_ (.A1(_08910_),
    .A2(_09207_),
    .B(_09210_),
    .C(_08566_),
    .Y(_09211_));
 OR3x4_ASAP7_75t_R _29173_ (.A(_08599_),
    .B(_09205_),
    .C(_09211_),
    .Y(_09212_));
 AND2x6_ASAP7_75t_R _29174_ (.A(_09204_),
    .B(_09212_),
    .Y(_09213_));
 NOR2x1_ASAP7_75t_R _29175_ (.A(_00925_),
    .B(_08598_),
    .Y(_09214_));
 AO21x1_ASAP7_75t_R _29176_ (.A1(_08598_),
    .A2(_09213_),
    .B(_09214_),
    .Y(_02872_));
 OA21x2_ASAP7_75t_R _29177_ (.A1(_01511_),
    .A2(_09177_),
    .B(_08879_),
    .Y(_09215_));
 NAND2x1_ASAP7_75t_R _29178_ (.A(net82),
    .B(_08881_),
    .Y(_09216_));
 OA211x2_ASAP7_75t_R _29179_ (.A1(_08900_),
    .A2(_08947_),
    .B(_09216_),
    .C(_08885_),
    .Y(_09217_));
 NAND2x1_ASAP7_75t_R _29180_ (.A(net79),
    .B(_08881_),
    .Y(_09218_));
 OA211x2_ASAP7_75t_R _29181_ (.A1(_01497_),
    .A2(_08947_),
    .B(_09218_),
    .C(_08880_),
    .Y(_09219_));
 OR3x1_ASAP7_75t_R _29182_ (.A(_08689_),
    .B(_09217_),
    .C(_09219_),
    .Y(_09220_));
 AND3x4_ASAP7_75t_R _29183_ (.A(_08683_),
    .B(_09215_),
    .C(_09220_),
    .Y(_09221_));
 OAI22x1_ASAP7_75t_R _29184_ (.A1(_00331_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00330_),
    .Y(_09222_));
 AO221x1_ASAP7_75t_R _29185_ (.A1(_08636_),
    .A2(_08780_),
    .B1(_08928_),
    .B2(_08632_),
    .C(_09034_),
    .Y(_09223_));
 AO22x1_ASAP7_75t_R _29186_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_08393_),
    .B1(_08395_),
    .B2(_02270_),
    .Y(_09224_));
 AO221x1_ASAP7_75t_R _29187_ (.A1(_08663_),
    .A2(_09222_),
    .B1(_09223_),
    .B2(_08831_),
    .C(_09224_),
    .Y(_09225_));
 NAND2x1_ASAP7_75t_R _29188_ (.A(_08377_),
    .B(_09225_),
    .Y(_09226_));
 NAND2x1_ASAP7_75t_R _29189_ (.A(_08509_),
    .B(_08791_),
    .Y(_09227_));
 OA21x2_ASAP7_75t_R _29190_ (.A1(_08509_),
    .A2(_08798_),
    .B(_09227_),
    .Y(_09228_));
 AND3x2_ASAP7_75t_R _29191_ (.A(_08366_),
    .B(_08401_),
    .C(_08403_),
    .Y(_09229_));
 OR4x1_ASAP7_75t_R _29192_ (.A(_00197_),
    .B(net2022),
    .C(net2008),
    .D(_09187_),
    .Y(_09230_));
 OR3x1_ASAP7_75t_R _29193_ (.A(_09024_),
    .B(_09026_),
    .C(_09230_),
    .Y(_09231_));
 OA21x2_ASAP7_75t_R _29194_ (.A1(_00206_),
    .A2(net2022),
    .B(_09155_),
    .Y(_09232_));
 OA21x2_ASAP7_75t_R _29195_ (.A1(_00228_),
    .A2(_00227_),
    .B(_00231_),
    .Y(_09233_));
 OA31x2_ASAP7_75t_R _29196_ (.A1(net2008),
    .A2(_09187_),
    .A3(_09232_),
    .B1(_09233_),
    .Y(_09234_));
 AND2x2_ASAP7_75t_R _29197_ (.A(_09231_),
    .B(_09234_),
    .Y(_09235_));
 XNOR2x1_ASAP7_75t_R _29198_ (.B(_09235_),
    .Y(_09236_),
    .A(_00230_));
 AND2x2_ASAP7_75t_R _29199_ (.A(_08549_),
    .B(_09236_),
    .Y(_09237_));
 AO21x1_ASAP7_75t_R _29200_ (.A1(_00137_),
    .A2(_09186_),
    .B(_09237_),
    .Y(_09238_));
 NAND2x1_ASAP7_75t_R _29201_ (.A(_13595_),
    .B(_09238_),
    .Y(_09239_));
 OA211x2_ASAP7_75t_R _29202_ (.A1(net2004),
    .A2(_05710_),
    .B(_05514_),
    .C(_09239_),
    .Y(_09240_));
 AOI21x1_ASAP7_75t_R _29203_ (.A1(_09119_),
    .A2(_09229_),
    .B(_09240_),
    .Y(_09241_));
 OA21x2_ASAP7_75t_R _29204_ (.A1(_09062_),
    .A2(_09228_),
    .B(_09241_),
    .Y(_09242_));
 AND4x2_ASAP7_75t_R _29205_ (.A(_06135_),
    .B(_08694_),
    .C(_09226_),
    .D(_09242_),
    .Y(_09243_));
 NOR2x2_ASAP7_75t_R _29206_ (.A(_09221_),
    .B(_09243_),
    .Y(_09244_));
 BUFx4f_ASAP7_75t_R _29207_ (.A(_09244_),
    .Y(_09245_));
 NAND2x1_ASAP7_75t_R _29208_ (.A(_00958_),
    .B(_08990_),
    .Y(_09246_));
 OA21x2_ASAP7_75t_R _29209_ (.A1(_09146_),
    .A2(_09245_),
    .B(_09246_),
    .Y(_02873_));
 NAND2x1_ASAP7_75t_R _29210_ (.A(net80),
    .B(_08881_),
    .Y(_09247_));
 OA211x2_ASAP7_75t_R _29211_ (.A1(_01496_),
    .A2(_08947_),
    .B(_09247_),
    .C(_08880_),
    .Y(_09248_));
 NAND2x1_ASAP7_75t_R _29212_ (.A(net93),
    .B(_08881_),
    .Y(_09249_));
 OA211x2_ASAP7_75t_R _29213_ (.A1(_08951_),
    .A2(_08947_),
    .B(_09249_),
    .C(_08885_),
    .Y(_09250_));
 OR3x2_ASAP7_75t_R _29214_ (.A(_08689_),
    .B(_09248_),
    .C(_09250_),
    .Y(_09251_));
 NAND2x2_ASAP7_75t_R _29215_ (.A(_09215_),
    .B(_09251_),
    .Y(_09252_));
 AND2x2_ASAP7_75t_R _29216_ (.A(_08429_),
    .B(_08786_),
    .Y(_09253_));
 AND2x2_ASAP7_75t_R _29217_ (.A(_08509_),
    .B(_08616_),
    .Y(_09254_));
 OAI22x1_ASAP7_75t_R _29218_ (.A1(_00333_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00332_),
    .Y(_09255_));
 AND2x2_ASAP7_75t_R _29219_ (.A(_02271_),
    .B(_08394_),
    .Y(_09256_));
 AO221x1_ASAP7_75t_R _29220_ (.A1(\alu_adder_result_ex[18] ),
    .A2(_08669_),
    .B1(_08381_),
    .B2(_09255_),
    .C(_09256_),
    .Y(_09257_));
 AO21x1_ASAP7_75t_R _29221_ (.A1(_08831_),
    .A2(_09034_),
    .B(_09257_),
    .Y(_09258_));
 AO221x1_ASAP7_75t_R _29222_ (.A1(_09090_),
    .A2(_09253_),
    .B1(_09254_),
    .B2(_09091_),
    .C(_09258_),
    .Y(_09259_));
 AO21x1_ASAP7_75t_R _29223_ (.A1(_09077_),
    .A2(_09184_),
    .B(_09259_),
    .Y(_09260_));
 AND2x2_ASAP7_75t_R _29224_ (.A(_08599_),
    .B(_08377_),
    .Y(_09261_));
 OA21x2_ASAP7_75t_R _29225_ (.A1(net2008),
    .A2(_09189_),
    .B(_09233_),
    .Y(_09262_));
 OA21x2_ASAP7_75t_R _29226_ (.A1(_00230_),
    .A2(_09262_),
    .B(_00235_),
    .Y(_09263_));
 XNOR2x1_ASAP7_75t_R _29227_ (.B(_09263_),
    .Y(_09264_),
    .A(_00234_));
 AND2x2_ASAP7_75t_R _29228_ (.A(_00140_),
    .B(_09186_),
    .Y(_09265_));
 AO21x1_ASAP7_75t_R _29229_ (.A1(_08827_),
    .A2(_09264_),
    .B(_09265_),
    .Y(_09266_));
 NAND2x1_ASAP7_75t_R _29230_ (.A(_08774_),
    .B(_09266_),
    .Y(_09267_));
 OA211x2_ASAP7_75t_R _29231_ (.A1(_13595_),
    .A2(_05716_),
    .B(_05515_),
    .C(_09267_),
    .Y(_09268_));
 OA21x2_ASAP7_75t_R _29232_ (.A1(_06159_),
    .A2(_09268_),
    .B(_08694_),
    .Y(_09269_));
 AO221x2_ASAP7_75t_R _29233_ (.A1(_08345_),
    .A2(_09252_),
    .B1(_09260_),
    .B2(_09261_),
    .C(_09269_),
    .Y(_09270_));
 BUFx6f_ASAP7_75t_R _29234_ (.A(_09270_),
    .Y(_09271_));
 NAND2x1_ASAP7_75t_R _29235_ (.A(_00991_),
    .B(_08990_),
    .Y(_09272_));
 OA21x2_ASAP7_75t_R _29236_ (.A1(_09146_),
    .A2(_09271_),
    .B(_09272_),
    .Y(_02874_));
 AND2x2_ASAP7_75t_R _29237_ (.A(_00235_),
    .B(_00238_),
    .Y(_09273_));
 AND2x2_ASAP7_75t_R _29238_ (.A(_09234_),
    .B(_09273_),
    .Y(_09274_));
 AO21x1_ASAP7_75t_R _29239_ (.A1(_00230_),
    .A2(_00235_),
    .B(_00234_),
    .Y(_09275_));
 AND2x2_ASAP7_75t_R _29240_ (.A(_00238_),
    .B(_09275_),
    .Y(_09276_));
 AO21x1_ASAP7_75t_R _29241_ (.A1(_09231_),
    .A2(_09274_),
    .B(_09276_),
    .Y(_09277_));
 XNOR2x1_ASAP7_75t_R _29242_ (.B(_09277_),
    .Y(_09278_),
    .A(_00237_));
 AND2x2_ASAP7_75t_R _29243_ (.A(_08550_),
    .B(_09278_),
    .Y(_09279_));
 AO21x1_ASAP7_75t_R _29244_ (.A1(_00146_),
    .A2(_09186_),
    .B(_09279_),
    .Y(_09280_));
 NAND2x1_ASAP7_75t_R _29245_ (.A(_08774_),
    .B(_09280_),
    .Y(_09281_));
 OA211x2_ASAP7_75t_R _29246_ (.A1(_08774_),
    .A2(_05623_),
    .B(_05515_),
    .C(_09281_),
    .Y(_09282_));
 AOI21x1_ASAP7_75t_R _29247_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_09122_),
    .B(_09282_),
    .Y(_09283_));
 NAND2x1_ASAP7_75t_R _29248_ (.A(_06178_),
    .B(_09283_),
    .Y(_09284_));
 INVx2_ASAP7_75t_R _29249_ (.A(_08506_),
    .Y(_09285_));
 OA22x2_ASAP7_75t_R _29250_ (.A1(_00335_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00334_),
    .Y(_09286_));
 NAND2x1_ASAP7_75t_R _29251_ (.A(_02272_),
    .B(_08395_),
    .Y(_09287_));
 OA21x2_ASAP7_75t_R _29252_ (.A1(_08395_),
    .A2(_09286_),
    .B(_09287_),
    .Y(_09288_));
 OA21x2_ASAP7_75t_R _29253_ (.A1(_09285_),
    .A2(_08862_),
    .B(_09288_),
    .Y(_09289_));
 OA21x2_ASAP7_75t_R _29254_ (.A1(_09061_),
    .A2(_09110_),
    .B(_09289_),
    .Y(_09290_));
 OAI21x1_ASAP7_75t_R _29255_ (.A1(_08423_),
    .A2(_09055_),
    .B(_09290_),
    .Y(_09291_));
 NAND2x1_ASAP7_75t_R _29256_ (.A(net81),
    .B(_08902_),
    .Y(_09292_));
 OA211x2_ASAP7_75t_R _29257_ (.A1(_01495_),
    .A2(_08947_),
    .B(_09292_),
    .C(_08910_),
    .Y(_09293_));
 NAND2x1_ASAP7_75t_R _29258_ (.A(net97),
    .B(_08902_),
    .Y(_09294_));
 OA211x2_ASAP7_75t_R _29259_ (.A1(_08995_),
    .A2(_08947_),
    .B(_09294_),
    .C(_08885_),
    .Y(_09295_));
 OR3x1_ASAP7_75t_R _29260_ (.A(_08689_),
    .B(_09293_),
    .C(_09295_),
    .Y(_09296_));
 AOI21x1_ASAP7_75t_R _29261_ (.A1(_09215_),
    .A2(_09296_),
    .B(_08600_),
    .Y(_09297_));
 AO221x2_ASAP7_75t_R _29262_ (.A1(_08600_),
    .A2(_09284_),
    .B1(_09291_),
    .B2(_09261_),
    .C(_09297_),
    .Y(_09298_));
 BUFx6f_ASAP7_75t_R _29263_ (.A(_09298_),
    .Y(_09299_));
 NAND2x1_ASAP7_75t_R _29264_ (.A(_01024_),
    .B(_08990_),
    .Y(_09300_));
 OA21x2_ASAP7_75t_R _29265_ (.A1(_09146_),
    .A2(_09299_),
    .B(_09300_),
    .Y(_02875_));
 OAI22x1_ASAP7_75t_R _29266_ (.A1(_00337_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00336_),
    .Y(_09301_));
 AND2x2_ASAP7_75t_R _29267_ (.A(_02273_),
    .B(_08394_),
    .Y(_09302_));
 AO21x1_ASAP7_75t_R _29268_ (.A1(_08382_),
    .A2(_09301_),
    .B(_09302_),
    .Y(_09303_));
 AO21x1_ASAP7_75t_R _29269_ (.A1(_08542_),
    .A2(_08861_),
    .B(_09303_),
    .Y(_09304_));
 AO221x1_ASAP7_75t_R _29270_ (.A1(_08777_),
    .A2(_09018_),
    .B1(_09184_),
    .B2(_09006_),
    .C(_09304_),
    .Y(_09305_));
 AO21x1_ASAP7_75t_R _29271_ (.A1(_00227_),
    .A2(_00231_),
    .B(_00230_),
    .Y(_09306_));
 OR2x2_ASAP7_75t_R _29272_ (.A(_09187_),
    .B(_09306_),
    .Y(_09307_));
 OA211x2_ASAP7_75t_R _29273_ (.A1(_00230_),
    .A2(_09233_),
    .B(_09273_),
    .C(_00241_),
    .Y(_09308_));
 OA21x2_ASAP7_75t_R _29274_ (.A1(_09188_),
    .A2(_09307_),
    .B(_09308_),
    .Y(_09309_));
 AO21x1_ASAP7_75t_R _29275_ (.A1(_00234_),
    .A2(_00238_),
    .B(_00237_),
    .Y(_09310_));
 AND2x2_ASAP7_75t_R _29276_ (.A(_00241_),
    .B(_09310_),
    .Y(_09311_));
 NOR2x1_ASAP7_75t_R _29277_ (.A(_09309_),
    .B(_09311_),
    .Y(_09312_));
 XNOR2x1_ASAP7_75t_R _29278_ (.B(_09312_),
    .Y(_09313_),
    .A(_00240_));
 AND2x2_ASAP7_75t_R _29279_ (.A(_08610_),
    .B(_09186_),
    .Y(_09314_));
 AO21x1_ASAP7_75t_R _29280_ (.A1(_08827_),
    .A2(_09313_),
    .B(_09314_),
    .Y(_09315_));
 NOR2x1_ASAP7_75t_R _29281_ (.A(_08774_),
    .B(_05315_),
    .Y(_09316_));
 AO21x1_ASAP7_75t_R _29282_ (.A1(_08774_),
    .A2(_09315_),
    .B(_09316_),
    .Y(_09317_));
 AO221x1_ASAP7_75t_R _29283_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_09122_),
    .B1(_09317_),
    .B2(_05516_),
    .C(_06216_),
    .Y(_09318_));
 AO21x1_ASAP7_75t_R _29284_ (.A1(_08377_),
    .A2(_09305_),
    .B(_09318_),
    .Y(_09319_));
 AND2x2_ASAP7_75t_R _29285_ (.A(net98),
    .B(_08580_),
    .Y(_09320_));
 AO21x1_ASAP7_75t_R _29286_ (.A1(net51),
    .A2(_08908_),
    .B(_09320_),
    .Y(_09321_));
 NAND2x1_ASAP7_75t_R _29287_ (.A(net83),
    .B(_08580_),
    .Y(_09322_));
 OA211x2_ASAP7_75t_R _29288_ (.A1(_01493_),
    .A2(_08881_),
    .B(_09322_),
    .C(_08572_),
    .Y(_09323_));
 INVx1_ASAP7_75t_R _29289_ (.A(_09323_),
    .Y(_09324_));
 OA211x2_ASAP7_75t_R _29290_ (.A1(_08945_),
    .A2(_09321_),
    .B(_09324_),
    .C(_08685_),
    .Y(_09325_));
 OR3x1_ASAP7_75t_R _29291_ (.A(_08694_),
    .B(_09205_),
    .C(_09325_),
    .Y(_09326_));
 OA21x2_ASAP7_75t_R _29292_ (.A1(_08684_),
    .A2(_09319_),
    .B(_09326_),
    .Y(_09327_));
 BUFx4f_ASAP7_75t_R _29293_ (.A(_09327_),
    .Y(_09328_));
 NAND2x1_ASAP7_75t_R _29294_ (.A(_01057_),
    .B(_08990_),
    .Y(_09329_));
 OA21x2_ASAP7_75t_R _29295_ (.A1(_09146_),
    .A2(_09328_),
    .B(_09329_),
    .Y(_02876_));
 OAI22x1_ASAP7_75t_R _29296_ (.A1(_00339_),
    .A2(_08384_),
    .B1(_08389_),
    .B2(_00338_),
    .Y(_09330_));
 AO22x1_ASAP7_75t_R _29297_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_08360_),
    .B1(_08380_),
    .B2(_02274_),
    .Y(_09331_));
 AO21x1_ASAP7_75t_R _29298_ (.A1(_08381_),
    .A2(_09330_),
    .B(_09331_),
    .Y(_09332_));
 AO21x1_ASAP7_75t_R _29299_ (.A1(_08506_),
    .A2(_08861_),
    .B(_09332_),
    .Y(_09333_));
 AND4x1_ASAP7_75t_R _29300_ (.A(_08481_),
    .B(_08508_),
    .C(_08506_),
    .D(_08750_),
    .Y(_09334_));
 AND3x1_ASAP7_75t_R _29301_ (.A(_08631_),
    .B(_08506_),
    .C(_08746_),
    .Y(_09335_));
 OR3x1_ASAP7_75t_R _29302_ (.A(_09333_),
    .B(_09334_),
    .C(_09335_),
    .Y(_09336_));
 OR2x2_ASAP7_75t_R _29303_ (.A(_00237_),
    .B(_00240_),
    .Y(_09337_));
 AO211x2_ASAP7_75t_R _29304_ (.A1(_09231_),
    .A2(_09274_),
    .B(_09337_),
    .C(_09276_),
    .Y(_09338_));
 OA21x2_ASAP7_75t_R _29305_ (.A1(_00241_),
    .A2(_00240_),
    .B(_00244_),
    .Y(_09339_));
 AND2x2_ASAP7_75t_R _29306_ (.A(_09338_),
    .B(_09339_),
    .Y(_09340_));
 XNOR2x1_ASAP7_75t_R _29307_ (.B(_09340_),
    .Y(_09341_),
    .A(_00243_));
 AND2x2_ASAP7_75t_R _29308_ (.A(_00158_),
    .B(_09185_),
    .Y(_09342_));
 AO21x1_ASAP7_75t_R _29309_ (.A1(_08550_),
    .A2(_09341_),
    .B(_09342_),
    .Y(_09343_));
 NAND2x1_ASAP7_75t_R _29310_ (.A(net2004),
    .B(_09343_),
    .Y(_09344_));
 OA211x2_ASAP7_75t_R _29311_ (.A1(_08774_),
    .A2(_05722_),
    .B(_05514_),
    .C(_09344_),
    .Y(_09345_));
 AO221x1_ASAP7_75t_R _29312_ (.A1(_08777_),
    .A2(_08981_),
    .B1(_09336_),
    .B2(_08376_),
    .C(_09345_),
    .Y(_09346_));
 OR2x2_ASAP7_75t_R _29313_ (.A(_08554_),
    .B(_06240_),
    .Y(_09347_));
 OA21x2_ASAP7_75t_R _29314_ (.A1(_05078_),
    .A2(_09346_),
    .B(_09347_),
    .Y(_09348_));
 AND2x2_ASAP7_75t_R _29315_ (.A(net99),
    .B(_08580_),
    .Y(_09349_));
 AO21x1_ASAP7_75t_R _29316_ (.A1(net75),
    .A2(_08908_),
    .B(_09349_),
    .Y(_09350_));
 NAND2x1_ASAP7_75t_R _29317_ (.A(net84),
    .B(_08580_),
    .Y(_09351_));
 OA211x2_ASAP7_75t_R _29318_ (.A1(_01492_),
    .A2(_08881_),
    .B(_09351_),
    .C(_08572_),
    .Y(_09352_));
 INVx1_ASAP7_75t_R _29319_ (.A(_09352_),
    .Y(_09353_));
 OA211x2_ASAP7_75t_R _29320_ (.A1(_08945_),
    .A2(_09350_),
    .B(_09353_),
    .C(_08685_),
    .Y(_09354_));
 OR3x1_ASAP7_75t_R _29321_ (.A(_08694_),
    .B(_09205_),
    .C(_09354_),
    .Y(_09355_));
 OA21x2_ASAP7_75t_R _29322_ (.A1(_08345_),
    .A2(_09348_),
    .B(_09355_),
    .Y(_09356_));
 BUFx6f_ASAP7_75t_R _29323_ (.A(_09356_),
    .Y(_09357_));
 BUFx10_ASAP7_75t_R _29324_ (.A(_08680_),
    .Y(_09358_));
 NAND2x1_ASAP7_75t_R _29325_ (.A(_01090_),
    .B(_09358_),
    .Y(_09359_));
 OA21x2_ASAP7_75t_R _29326_ (.A1(_09146_),
    .A2(_09357_),
    .B(_09359_),
    .Y(_02877_));
 OR2x2_ASAP7_75t_R _29327_ (.A(_08753_),
    .B(_04867_),
    .Y(_09360_));
 BUFx4f_ASAP7_75t_R _29328_ (.A(_09360_),
    .Y(_09361_));
 OR2x2_ASAP7_75t_R _29329_ (.A(_13566_),
    .B(_04867_),
    .Y(_09362_));
 OR2x2_ASAP7_75t_R _29330_ (.A(_00240_),
    .B(_00243_),
    .Y(_09363_));
 OR2x2_ASAP7_75t_R _29331_ (.A(_00244_),
    .B(_00243_),
    .Y(_09364_));
 OA31x2_ASAP7_75t_R _29332_ (.A1(_09309_),
    .A2(_09311_),
    .A3(_09363_),
    .B1(_09364_),
    .Y(_09365_));
 AND2x2_ASAP7_75t_R _29333_ (.A(_00247_),
    .B(_09365_),
    .Y(_09366_));
 XNOR2x1_ASAP7_75t_R _29334_ (.B(_09366_),
    .Y(_09367_),
    .A(_00246_));
 NOR2x1_ASAP7_75t_R _29335_ (.A(_08550_),
    .B(_08773_),
    .Y(_09368_));
 AO21x1_ASAP7_75t_R _29336_ (.A1(_08827_),
    .A2(_09367_),
    .B(_09368_),
    .Y(_09369_));
 OAI22x1_ASAP7_75t_R _29337_ (.A1(_05316_),
    .A2(_09361_),
    .B1(_09362_),
    .B2(_09369_),
    .Y(_09370_));
 AND2x2_ASAP7_75t_R _29338_ (.A(_08831_),
    .B(_08615_),
    .Y(_09371_));
 OAI22x1_ASAP7_75t_R _29339_ (.A1(_00341_),
    .A2(_08384_),
    .B1(_08389_),
    .B2(_00340_),
    .Y(_09372_));
 AND2x2_ASAP7_75t_R _29340_ (.A(_02275_),
    .B(_08380_),
    .Y(_09373_));
 AO221x1_ASAP7_75t_R _29341_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_08669_),
    .B1(_08381_),
    .B2(_09372_),
    .C(_09373_),
    .Y(_09374_));
 OR2x2_ASAP7_75t_R _29342_ (.A(_05078_),
    .B(_09374_),
    .Y(_09375_));
 AO221x1_ASAP7_75t_R _29343_ (.A1(_08429_),
    .A2(_08931_),
    .B1(_09371_),
    .B2(_08914_),
    .C(_09375_),
    .Y(_09376_));
 OR2x2_ASAP7_75t_R _29344_ (.A(_13776_),
    .B(_08375_),
    .Y(_09377_));
 OR2x2_ASAP7_75t_R _29345_ (.A(_09377_),
    .B(_09370_),
    .Y(_09378_));
 NAND2x1_ASAP7_75t_R _29346_ (.A(_05078_),
    .B(_06258_),
    .Y(_09379_));
 OA211x2_ASAP7_75t_R _29347_ (.A1(_09370_),
    .A2(_09376_),
    .B(_09378_),
    .C(_09379_),
    .Y(_09380_));
 AND2x2_ASAP7_75t_R _29348_ (.A(net100),
    .B(_08580_),
    .Y(_09381_));
 AO21x1_ASAP7_75t_R _29349_ (.A1(net76),
    .A2(_08908_),
    .B(_09381_),
    .Y(_09382_));
 INVx1_ASAP7_75t_R _29350_ (.A(net85),
    .Y(_09383_));
 OR2x2_ASAP7_75t_R _29351_ (.A(_01491_),
    .B(_08573_),
    .Y(_09384_));
 OA211x2_ASAP7_75t_R _29352_ (.A1(_09383_),
    .A2(_08908_),
    .B(_09384_),
    .C(_08572_),
    .Y(_09385_));
 INVx1_ASAP7_75t_R _29353_ (.A(_09385_),
    .Y(_09386_));
 OA211x2_ASAP7_75t_R _29354_ (.A1(_08945_),
    .A2(_09382_),
    .B(_09386_),
    .C(_08685_),
    .Y(_09387_));
 OR3x1_ASAP7_75t_R _29355_ (.A(_08694_),
    .B(_09205_),
    .C(_09387_),
    .Y(_09388_));
 OA21x2_ASAP7_75t_R _29356_ (.A1(_08684_),
    .A2(_09380_),
    .B(_09388_),
    .Y(_09389_));
 BUFx6f_ASAP7_75t_R _29357_ (.A(_09389_),
    .Y(_09390_));
 NAND2x1_ASAP7_75t_R _29358_ (.A(_01123_),
    .B(_09358_),
    .Y(_09391_));
 OA21x2_ASAP7_75t_R _29359_ (.A1(_09146_),
    .A2(_09390_),
    .B(_09391_),
    .Y(_02878_));
 OR2x2_ASAP7_75t_R _29360_ (.A(_00243_),
    .B(_00246_),
    .Y(_09392_));
 AO21x1_ASAP7_75t_R _29361_ (.A1(_09338_),
    .A2(_09339_),
    .B(_09392_),
    .Y(_09393_));
 OA211x2_ASAP7_75t_R _29362_ (.A1(_00247_),
    .A2(_00246_),
    .B(_00250_),
    .C(_09393_),
    .Y(_09394_));
 XNOR2x1_ASAP7_75t_R _29363_ (.B(_09394_),
    .Y(_09395_),
    .A(_00249_));
 NOR2x1_ASAP7_75t_R _29364_ (.A(_08827_),
    .B(_08826_),
    .Y(_09396_));
 AO21x1_ASAP7_75t_R _29365_ (.A1(_08827_),
    .A2(_09395_),
    .B(_09396_),
    .Y(_09397_));
 NAND2x1_ASAP7_75t_R _29366_ (.A(_08774_),
    .B(_09397_),
    .Y(_09398_));
 OA211x2_ASAP7_75t_R _29367_ (.A1(_13595_),
    .A2(_05642_),
    .B(_05515_),
    .C(_09398_),
    .Y(_09399_));
 INVx1_ASAP7_75t_R _29368_ (.A(_09399_),
    .Y(_09400_));
 OA211x2_ASAP7_75t_R _29369_ (.A1(_08433_),
    .A2(_08465_),
    .B(_08615_),
    .C(_08509_),
    .Y(_09401_));
 AO21x1_ASAP7_75t_R _29370_ (.A1(_08786_),
    .A2(_08541_),
    .B(_09401_),
    .Y(_09402_));
 OAI22x1_ASAP7_75t_R _29371_ (.A1(_00343_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00342_),
    .Y(_09403_));
 AO22x1_ASAP7_75t_R _29372_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_08669_),
    .B1(_08670_),
    .B2(_02276_),
    .Y(_09404_));
 AO21x1_ASAP7_75t_R _29373_ (.A1(_08663_),
    .A2(_09403_),
    .B(_09404_),
    .Y(_09405_));
 AO221x1_ASAP7_75t_R _29374_ (.A1(_13648_),
    .A2(_13774_),
    .B1(_08831_),
    .B2(_09034_),
    .C(_09405_),
    .Y(_09406_));
 AOI221x1_ASAP7_75t_R _29375_ (.A1(_08777_),
    .A2(_09402_),
    .B1(_09184_),
    .B2(_08837_),
    .C(_09406_),
    .Y(_09407_));
 OAI22x1_ASAP7_75t_R _29376_ (.A1(_08554_),
    .A2(_06279_),
    .B1(_09377_),
    .B2(_09399_),
    .Y(_09408_));
 AO21x1_ASAP7_75t_R _29377_ (.A1(_09400_),
    .A2(_09407_),
    .B(_09408_),
    .Y(_09409_));
 INVx1_ASAP7_75t_R _29378_ (.A(_01490_),
    .Y(_09410_));
 OA211x2_ASAP7_75t_R _29379_ (.A1(_09410_),
    .A2(_08902_),
    .B(_08874_),
    .C(_08880_),
    .Y(_09411_));
 INVx1_ASAP7_75t_R _29380_ (.A(_09411_),
    .Y(_09412_));
 OA21x2_ASAP7_75t_R _29381_ (.A1(_08945_),
    .A2(_08872_),
    .B(_09412_),
    .Y(_09413_));
 OA211x2_ASAP7_75t_R _29382_ (.A1(_08689_),
    .A2(_09413_),
    .B(_09215_),
    .C(_08683_),
    .Y(_09414_));
 AOI21x1_ASAP7_75t_R _29383_ (.A1(_08600_),
    .A2(_09409_),
    .B(_09414_),
    .Y(_09415_));
 BUFx6f_ASAP7_75t_R _29384_ (.A(_09415_),
    .Y(_09416_));
 NAND2x1_ASAP7_75t_R _29385_ (.A(_01156_),
    .B(_09358_),
    .Y(_09417_));
 OA21x2_ASAP7_75t_R _29386_ (.A1(_09146_),
    .A2(_09416_),
    .B(_09417_),
    .Y(_02879_));
 NAND2x1_ASAP7_75t_R _29387_ (.A(_01812_),
    .B(_08591_),
    .Y(_09418_));
 OA21x2_ASAP7_75t_R _29388_ (.A1(_09107_),
    .A2(_09037_),
    .B(_09418_),
    .Y(_02880_));
 AO21x1_ASAP7_75t_R _29389_ (.A1(_00247_),
    .A2(_09365_),
    .B(_00246_),
    .Y(_09419_));
 AND2x2_ASAP7_75t_R _29390_ (.A(_00250_),
    .B(_00253_),
    .Y(_09420_));
 AO22x1_ASAP7_75t_R _29391_ (.A1(_00249_),
    .A2(_00253_),
    .B1(_09419_),
    .B2(_09420_),
    .Y(_09421_));
 XOR2x1_ASAP7_75t_R _29392_ (.A(_00252_),
    .Y(_09422_),
    .B(_09421_));
 AND2x2_ASAP7_75t_R _29393_ (.A(_09185_),
    .B(_08866_),
    .Y(_09423_));
 AO21x1_ASAP7_75t_R _29394_ (.A1(_08550_),
    .A2(_09422_),
    .B(_09423_),
    .Y(_09424_));
 NAND2x1_ASAP7_75t_R _29395_ (.A(_13566_),
    .B(_05317_),
    .Y(_09425_));
 OA211x2_ASAP7_75t_R _29396_ (.A1(_13567_),
    .A2(_09424_),
    .B(_09425_),
    .C(_05514_),
    .Y(_09426_));
 AO21x1_ASAP7_75t_R _29397_ (.A1(\alu_adder_result_ex[24] ),
    .A2(_09122_),
    .B(_09426_),
    .Y(_09427_));
 OAI22x1_ASAP7_75t_R _29398_ (.A1(_00345_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00344_),
    .Y(_09428_));
 AND2x2_ASAP7_75t_R _29399_ (.A(_02277_),
    .B(_08394_),
    .Y(_09429_));
 AO21x1_ASAP7_75t_R _29400_ (.A1(_08382_),
    .A2(_09428_),
    .B(_09429_),
    .Y(_09430_));
 AND3x1_ASAP7_75t_R _29401_ (.A(_08631_),
    .B(_08524_),
    .C(_08506_),
    .Y(_09431_));
 AND3x1_ASAP7_75t_R _29402_ (.A(_08695_),
    .B(_08649_),
    .C(_08506_),
    .Y(_09432_));
 OR4x1_ASAP7_75t_R _29403_ (.A(_05078_),
    .B(_09430_),
    .C(_09431_),
    .D(_09432_),
    .Y(_09433_));
 AO21x1_ASAP7_75t_R _29404_ (.A1(_08777_),
    .A2(_08847_),
    .B(_09433_),
    .Y(_09434_));
 OR2x2_ASAP7_75t_R _29405_ (.A(_08554_),
    .B(_06297_),
    .Y(_09435_));
 OR2x2_ASAP7_75t_R _29406_ (.A(_09377_),
    .B(_09426_),
    .Y(_09436_));
 OA211x2_ASAP7_75t_R _29407_ (.A1(_09427_),
    .A2(_09434_),
    .B(_09435_),
    .C(_09436_),
    .Y(_09437_));
 NAND2x1_ASAP7_75t_R _29408_ (.A(_08885_),
    .B(_08891_),
    .Y(_09438_));
 OA211x2_ASAP7_75t_R _29409_ (.A1(_08885_),
    .A2(_08889_),
    .B(_09438_),
    .C(_08685_),
    .Y(_09439_));
 OA21x2_ASAP7_75t_R _29410_ (.A1(_09205_),
    .A2(_09439_),
    .B(_08345_),
    .Y(_09440_));
 AO21x2_ASAP7_75t_R _29411_ (.A1(_08600_),
    .A2(_09437_),
    .B(_09440_),
    .Y(_09441_));
 BUFx4f_ASAP7_75t_R _29412_ (.A(_09441_),
    .Y(_09442_));
 NAND2x1_ASAP7_75t_R _29413_ (.A(_01189_),
    .B(_09358_),
    .Y(_09443_));
 OA21x2_ASAP7_75t_R _29414_ (.A1(_09146_),
    .A2(_09442_),
    .B(_09443_),
    .Y(_02881_));
 NOR2x1_ASAP7_75t_R _29415_ (.A(net79),
    .B(_08947_),
    .Y(_09444_));
 AO21x1_ASAP7_75t_R _29416_ (.A1(_08900_),
    .A2(_08956_),
    .B(_09444_),
    .Y(_09445_));
 INVx1_ASAP7_75t_R _29417_ (.A(net88),
    .Y(_09446_));
 OA211x2_ASAP7_75t_R _29418_ (.A1(_09446_),
    .A2(_08908_),
    .B(_08909_),
    .C(_08910_),
    .Y(_09447_));
 AO21x1_ASAP7_75t_R _29419_ (.A1(_08885_),
    .A2(_09445_),
    .B(_09447_),
    .Y(_09448_));
 OA21x2_ASAP7_75t_R _29420_ (.A1(_08689_),
    .A2(_09448_),
    .B(_09215_),
    .Y(_09449_));
 OR3x1_ASAP7_75t_R _29421_ (.A(_08799_),
    .B(_08800_),
    .C(_08802_),
    .Y(_09450_));
 OR3x1_ASAP7_75t_R _29422_ (.A(_08423_),
    .B(_08695_),
    .C(_09450_),
    .Y(_09451_));
 OR3x1_ASAP7_75t_R _29423_ (.A(_08786_),
    .B(_08798_),
    .C(_09062_),
    .Y(_09452_));
 AND3x1_ASAP7_75t_R _29424_ (.A(_08786_),
    .B(_08791_),
    .C(_09229_),
    .Y(_09453_));
 AOI21x1_ASAP7_75t_R _29425_ (.A1(_08794_),
    .A2(_09229_),
    .B(_09453_),
    .Y(_09454_));
 AND3x1_ASAP7_75t_R _29426_ (.A(_09451_),
    .B(_09452_),
    .C(_09454_),
    .Y(_09455_));
 OAI22x1_ASAP7_75t_R _29427_ (.A1(_00347_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00346_),
    .Y(_09456_));
 AND2x2_ASAP7_75t_R _29428_ (.A(_02278_),
    .B(_08395_),
    .Y(_09457_));
 AO221x1_ASAP7_75t_R _29429_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_08393_),
    .B1(_08663_),
    .B2(_09456_),
    .C(_09457_),
    .Y(_09458_));
 AND3x1_ASAP7_75t_R _29430_ (.A(_08542_),
    .B(_08702_),
    .C(_08781_),
    .Y(_09459_));
 NOR2x1_ASAP7_75t_R _29431_ (.A(_09458_),
    .B(_09459_),
    .Y(_09460_));
 AO21x1_ASAP7_75t_R _29432_ (.A1(_09455_),
    .A2(_09460_),
    .B(_09056_),
    .Y(_09461_));
 OR2x2_ASAP7_75t_R _29433_ (.A(_05645_),
    .B(_08936_),
    .Y(_09462_));
 OR2x2_ASAP7_75t_R _29434_ (.A(_00249_),
    .B(_00252_),
    .Y(_09463_));
 OA21x2_ASAP7_75t_R _29435_ (.A1(_00253_),
    .A2(_00252_),
    .B(_00256_),
    .Y(_09464_));
 OA21x2_ASAP7_75t_R _29436_ (.A1(_09394_),
    .A2(_09463_),
    .B(_09464_),
    .Y(_09465_));
 XNOR2x2_ASAP7_75t_R _29437_ (.A(_00255_),
    .B(_09465_),
    .Y(_09466_));
 AND3x1_ASAP7_75t_R _29438_ (.A(_08774_),
    .B(_09186_),
    .C(_08935_),
    .Y(_09467_));
 OR2x2_ASAP7_75t_R _29439_ (.A(_05141_),
    .B(_09467_),
    .Y(_09468_));
 AOI21x1_ASAP7_75t_R _29440_ (.A1(_08932_),
    .A2(_09466_),
    .B(_09468_),
    .Y(_09469_));
 AOI211x1_ASAP7_75t_R _29441_ (.A1(_09462_),
    .A2(_09469_),
    .B(_06318_),
    .C(_08345_),
    .Y(_09470_));
 AOI22x1_ASAP7_75t_R _29442_ (.A1(_08684_),
    .A2(_09449_),
    .B1(_09461_),
    .B2(_09470_),
    .Y(_09471_));
 BUFx6f_ASAP7_75t_R _29443_ (.A(_09471_),
    .Y(_09472_));
 NAND2x1_ASAP7_75t_R _29444_ (.A(_01222_),
    .B(_09358_),
    .Y(_09473_));
 OA21x2_ASAP7_75t_R _29445_ (.A1(_09146_),
    .A2(_09472_),
    .B(_09473_),
    .Y(_02882_));
 OAI22x1_ASAP7_75t_R _29446_ (.A1(_00349_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00348_),
    .Y(_09474_));
 AND2x2_ASAP7_75t_R _29447_ (.A(_08382_),
    .B(_09474_),
    .Y(_09475_));
 AO221x1_ASAP7_75t_R _29448_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_08393_),
    .B1(_08395_),
    .B2(_02279_),
    .C(_09475_),
    .Y(_09476_));
 AND3x1_ASAP7_75t_R _29449_ (.A(_08542_),
    .B(_08701_),
    .C(_08702_),
    .Y(_09477_));
 AOI211x1_ASAP7_75t_R _29450_ (.A1(_08777_),
    .A2(_08752_),
    .B(_09476_),
    .C(_09477_),
    .Y(_09478_));
 OR2x2_ASAP7_75t_R _29451_ (.A(_09056_),
    .B(_09478_),
    .Y(_09479_));
 AND4x1_ASAP7_75t_R _29452_ (.A(_00250_),
    .B(_00253_),
    .C(_00256_),
    .D(_00259_),
    .Y(_09480_));
 AO21x1_ASAP7_75t_R _29453_ (.A1(_00249_),
    .A2(_00253_),
    .B(_00252_),
    .Y(_09481_));
 AO21x1_ASAP7_75t_R _29454_ (.A1(_00256_),
    .A2(_09481_),
    .B(_00255_),
    .Y(_09482_));
 AO22x1_ASAP7_75t_R _29455_ (.A1(_09419_),
    .A2(_09480_),
    .B1(_09482_),
    .B2(_00259_),
    .Y(_09483_));
 XOR2x1_ASAP7_75t_R _29456_ (.A(_00258_),
    .Y(_09484_),
    .B(_09483_));
 NOR2x1_ASAP7_75t_R _29457_ (.A(_08551_),
    .B(_08985_),
    .Y(_09485_));
 AO21x1_ASAP7_75t_R _29458_ (.A1(_08551_),
    .A2(_09484_),
    .B(_09485_),
    .Y(_09486_));
 INVx1_ASAP7_75t_R _29459_ (.A(_09486_),
    .Y(_09487_));
 AO21x1_ASAP7_75t_R _29460_ (.A1(_13567_),
    .A2(_05318_),
    .B(_05141_),
    .Y(_09488_));
 AO21x1_ASAP7_75t_R _29461_ (.A1(_13595_),
    .A2(_09487_),
    .B(_09488_),
    .Y(_09489_));
 AND3x1_ASAP7_75t_R _29462_ (.A(_06346_),
    .B(_08600_),
    .C(_09489_),
    .Y(_09490_));
 NOR2x1_ASAP7_75t_R _29463_ (.A(_08950_),
    .B(_08953_),
    .Y(_09491_));
 AO21x1_ASAP7_75t_R _29464_ (.A1(_08945_),
    .A2(_08949_),
    .B(_09491_),
    .Y(_09492_));
 OA211x2_ASAP7_75t_R _29465_ (.A1(_08689_),
    .A2(_09492_),
    .B(_09215_),
    .C(_08683_),
    .Y(_09493_));
 AOI21x1_ASAP7_75t_R _29466_ (.A1(_09479_),
    .A2(_09490_),
    .B(_09493_),
    .Y(_09494_));
 BUFx6f_ASAP7_75t_R _29467_ (.A(_09494_),
    .Y(_09495_));
 NAND2x1_ASAP7_75t_R _29468_ (.A(_01255_),
    .B(_09358_),
    .Y(_09496_));
 OA21x2_ASAP7_75t_R _29469_ (.A1(_08764_),
    .A2(_09495_),
    .B(_09496_),
    .Y(_02883_));
 OA21x2_ASAP7_75t_R _29470_ (.A1(_00255_),
    .A2(_09465_),
    .B(_00259_),
    .Y(_09497_));
 OA21x2_ASAP7_75t_R _29471_ (.A1(_00258_),
    .A2(_09497_),
    .B(_00262_),
    .Y(_09498_));
 XNOR2x1_ASAP7_75t_R _29472_ (.B(_09498_),
    .Y(_09499_),
    .A(_00261_));
 NAND2x1_ASAP7_75t_R _29473_ (.A(_08827_),
    .B(_09499_),
    .Y(_09500_));
 OR2x2_ASAP7_75t_R _29474_ (.A(_08550_),
    .B(_09028_),
    .Y(_09501_));
 AND4x2_ASAP7_75t_R _29475_ (.A(_08774_),
    .B(_05515_),
    .C(_09500_),
    .D(_09501_),
    .Y(_09502_));
 AND2x2_ASAP7_75t_R _29476_ (.A(_08429_),
    .B(_08662_),
    .Y(_09503_));
 OAI22x1_ASAP7_75t_R _29477_ (.A1(_00351_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00350_),
    .Y(_09504_));
 AO22x1_ASAP7_75t_R _29478_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_08360_),
    .B1(_08394_),
    .B2(_02280_),
    .Y(_09505_));
 AO21x1_ASAP7_75t_R _29479_ (.A1(_08382_),
    .A2(_09504_),
    .B(_09505_),
    .Y(_09506_));
 AO222x2_ASAP7_75t_R _29480_ (.A1(_05738_),
    .A2(_05096_),
    .B1(_08630_),
    .B2(_09371_),
    .C1(_09506_),
    .C2(_08376_),
    .Y(_09507_));
 OR5x2_ASAP7_75t_R _29481_ (.A(_06369_),
    .B(_08344_),
    .C(_09502_),
    .D(_09503_),
    .E(_09507_),
    .Y(_09508_));
 NAND2x1_ASAP7_75t_R _29482_ (.A(_08880_),
    .B(_08994_),
    .Y(_09509_));
 OA211x2_ASAP7_75t_R _29483_ (.A1(_08950_),
    .A2(_08997_),
    .B(_09509_),
    .C(_08566_),
    .Y(_09510_));
 OR3x4_ASAP7_75t_R _29484_ (.A(_08599_),
    .B(_09205_),
    .C(_09510_),
    .Y(_09511_));
 AND2x6_ASAP7_75t_R _29485_ (.A(_09508_),
    .B(_09511_),
    .Y(_09512_));
 NOR2x1_ASAP7_75t_R _29486_ (.A(_01288_),
    .B(_08598_),
    .Y(_09513_));
 AO21x1_ASAP7_75t_R _29487_ (.A1(_08598_),
    .A2(_09512_),
    .B(_09513_),
    .Y(_02884_));
 AO21x1_ASAP7_75t_R _29488_ (.A1(_00259_),
    .A2(_09482_),
    .B(_00258_),
    .Y(_09514_));
 AO21x1_ASAP7_75t_R _29489_ (.A1(_00262_),
    .A2(_09514_),
    .B(_00261_),
    .Y(_09515_));
 OA211x2_ASAP7_75t_R _29490_ (.A1(_00262_),
    .A2(_00261_),
    .B(_00265_),
    .C(_09480_),
    .Y(_09516_));
 AO22x1_ASAP7_75t_R _29491_ (.A1(_00265_),
    .A2(_09515_),
    .B1(_09516_),
    .B2(_09419_),
    .Y(_09517_));
 XOR2x1_ASAP7_75t_R _29492_ (.A(_00264_),
    .Y(_09518_),
    .B(_09517_));
 NOR2x1_ASAP7_75t_R _29493_ (.A(_08550_),
    .B(_09068_),
    .Y(_09519_));
 AO21x1_ASAP7_75t_R _29494_ (.A1(_08827_),
    .A2(_09518_),
    .B(_09519_),
    .Y(_09520_));
 NAND2x1_ASAP7_75t_R _29495_ (.A(_13567_),
    .B(_05319_),
    .Y(_09521_));
 OA211x2_ASAP7_75t_R _29496_ (.A1(_13567_),
    .A2(_09520_),
    .B(_09521_),
    .C(_05514_),
    .Y(_09522_));
 AO21x1_ASAP7_75t_R _29497_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_09122_),
    .B(_09522_),
    .Y(_09523_));
 AOI22x1_ASAP7_75t_R _29498_ (.A1(_18630_),
    .A2(_08487_),
    .B1(_08489_),
    .B2(_18622_),
    .Y(_09524_));
 AOI22x1_ASAP7_75t_R _29499_ (.A1(_18747_),
    .A2(_08484_),
    .B1(_08485_),
    .B2(_18742_),
    .Y(_09525_));
 AO32x1_ASAP7_75t_R _29500_ (.A1(_08646_),
    .A2(_09524_),
    .A3(_09525_),
    .B1(_08637_),
    .B2(_08725_),
    .Y(_09526_));
 AO22x1_ASAP7_75t_R _29501_ (.A1(_08640_),
    .A2(_08728_),
    .B1(_08722_),
    .B2(_08643_),
    .Y(_09527_));
 OA21x2_ASAP7_75t_R _29502_ (.A1(_09526_),
    .A2(_09527_),
    .B(_08631_),
    .Y(_09528_));
 NOR2x1_ASAP7_75t_R _29503_ (.A(_08704_),
    .B(_09016_),
    .Y(_09529_));
 AOI211x1_ASAP7_75t_R _29504_ (.A1(_08433_),
    .A2(_09061_),
    .B(_09528_),
    .C(_09529_),
    .Y(_09530_));
 AND2x2_ASAP7_75t_R _29505_ (.A(_08429_),
    .B(_09530_),
    .Y(_09531_));
 OAI22x1_ASAP7_75t_R _29506_ (.A1(_00353_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_00352_),
    .Y(_09532_));
 AND2x2_ASAP7_75t_R _29507_ (.A(_02281_),
    .B(_08394_),
    .Y(_09533_));
 AO21x1_ASAP7_75t_R _29508_ (.A1(_08382_),
    .A2(_09532_),
    .B(_09533_),
    .Y(_09534_));
 OA21x2_ASAP7_75t_R _29509_ (.A1(_08695_),
    .A2(_08482_),
    .B(_08411_),
    .Y(_09535_));
 AND3x1_ASAP7_75t_R _29510_ (.A(_08631_),
    .B(_08633_),
    .C(_09050_),
    .Y(_09536_));
 OA21x2_ASAP7_75t_R _29511_ (.A1(_09535_),
    .A2(_09536_),
    .B(_08831_),
    .Y(_09537_));
 OA21x2_ASAP7_75t_R _29512_ (.A1(_09534_),
    .A2(_09537_),
    .B(_08376_),
    .Y(_09538_));
 OR5x2_ASAP7_75t_R _29513_ (.A(_06391_),
    .B(_08344_),
    .C(_09523_),
    .D(_09531_),
    .E(_09538_),
    .Y(_09539_));
 NAND2x1_ASAP7_75t_R _29514_ (.A(_08910_),
    .B(_09040_),
    .Y(_09540_));
 OA211x2_ASAP7_75t_R _29515_ (.A1(_08950_),
    .A2(_09042_),
    .B(_09540_),
    .C(_08685_),
    .Y(_09541_));
 OR3x2_ASAP7_75t_R _29516_ (.A(_08694_),
    .B(_09205_),
    .C(_09541_),
    .Y(_09542_));
 AND2x6_ASAP7_75t_R _29517_ (.A(_09542_),
    .B(_09539_),
    .Y(_09543_));
 BUFx3_ASAP7_75t_R _29518_ (.A(_09543_),
    .Y(_09544_));
 NOR2x1_ASAP7_75t_R _29519_ (.A(_01321_),
    .B(_08598_),
    .Y(_09545_));
 AO21x1_ASAP7_75t_R _29520_ (.A1(_08598_),
    .A2(net95),
    .B(_09545_),
    .Y(_02885_));
 OAI22x1_ASAP7_75t_R _29521_ (.A1(_08838_),
    .A2(_08472_),
    .B1(_08491_),
    .B2(_08655_),
    .Y(_09546_));
 NAND2x1_ASAP7_75t_R _29522_ (.A(_08474_),
    .B(_08476_),
    .Y(_09547_));
 AO22x1_ASAP7_75t_R _29523_ (.A1(_08640_),
    .A2(_08801_),
    .B1(_09547_),
    .B2(_08643_),
    .Y(_09548_));
 OA21x2_ASAP7_75t_R _29524_ (.A1(_09546_),
    .A2(_09548_),
    .B(_08631_),
    .Y(_09549_));
 NOR2x1_ASAP7_75t_R _29525_ (.A(_08653_),
    .B(_08979_),
    .Y(_09550_));
 OAI22x1_ASAP7_75t_R _29526_ (.A1(_08652_),
    .A2(_08700_),
    .B1(_08974_),
    .B2(_08704_),
    .Y(_09551_));
 OR4x1_ASAP7_75t_R _29527_ (.A(_08423_),
    .B(_09549_),
    .C(_09550_),
    .D(_09551_),
    .Y(_09552_));
 OA22x2_ASAP7_75t_R _29528_ (.A1(_00355_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00354_),
    .Y(_09553_));
 NAND2x1_ASAP7_75t_R _29529_ (.A(_02282_),
    .B(_08394_),
    .Y(_09554_));
 OA21x2_ASAP7_75t_R _29530_ (.A1(_08670_),
    .A2(_09553_),
    .B(_09554_),
    .Y(_09555_));
 AOI21x1_ASAP7_75t_R _29531_ (.A1(_09552_),
    .A2(_09555_),
    .B(_09056_),
    .Y(_09556_));
 AO21x1_ASAP7_75t_R _29532_ (.A1(_00265_),
    .A2(_09515_),
    .B(_00264_),
    .Y(_09557_));
 AND3x1_ASAP7_75t_R _29533_ (.A(_00247_),
    .B(_00268_),
    .C(_09516_),
    .Y(_09558_));
 AO21x1_ASAP7_75t_R _29534_ (.A1(_09338_),
    .A2(_09339_),
    .B(_00243_),
    .Y(_09559_));
 AND3x1_ASAP7_75t_R _29535_ (.A(_00246_),
    .B(_00268_),
    .C(_09516_),
    .Y(_09560_));
 AO221x1_ASAP7_75t_R _29536_ (.A1(_00268_),
    .A2(_09557_),
    .B1(_09558_),
    .B2(_09559_),
    .C(_09560_),
    .Y(_09561_));
 XNOR2x1_ASAP7_75t_R _29537_ (.B(_00267_),
    .Y(_09562_),
    .A(_09561_));
 NOR2x1_ASAP7_75t_R _29538_ (.A(_08546_),
    .B(_09084_),
    .Y(_09563_));
 AO21x2_ASAP7_75t_R _29539_ (.A1(_08549_),
    .A2(_09562_),
    .B(_09563_),
    .Y(_09564_));
 NAND2x1_ASAP7_75t_R _29540_ (.A(_08753_),
    .B(_09564_),
    .Y(_09565_));
 OA211x2_ASAP7_75t_R _29541_ (.A1(_08753_),
    .A2(_05741_),
    .B(_09565_),
    .C(_05304_),
    .Y(_09566_));
 AND3x1_ASAP7_75t_R _29542_ (.A(_08631_),
    .B(_08633_),
    .C(_08749_),
    .Y(_09567_));
 OA21x2_ASAP7_75t_R _29543_ (.A1(_09535_),
    .A2(_09567_),
    .B(_08805_),
    .Y(_09568_));
 AO21x1_ASAP7_75t_R _29544_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_09122_),
    .B(_13776_),
    .Y(_09569_));
 OR3x1_ASAP7_75t_R _29545_ (.A(_09568_),
    .B(_09566_),
    .C(_09569_),
    .Y(_09570_));
 OR2x2_ASAP7_75t_R _29546_ (.A(_08554_),
    .B(_06409_),
    .Y(_09571_));
 OA211x2_ASAP7_75t_R _29547_ (.A1(_09570_),
    .A2(_09556_),
    .B(_09571_),
    .C(_08599_),
    .Y(_09572_));
 AND2x2_ASAP7_75t_R _29548_ (.A(net75),
    .B(_08573_),
    .Y(_09573_));
 AO21x1_ASAP7_75t_R _29549_ (.A1(net84),
    .A2(_08562_),
    .B(_09573_),
    .Y(_09574_));
 OA211x2_ASAP7_75t_R _29550_ (.A1(_08691_),
    .A2(_08562_),
    .B(_09099_),
    .C(_08557_),
    .Y(_09575_));
 INVx1_ASAP7_75t_R _29551_ (.A(_09575_),
    .Y(_09576_));
 OA211x2_ASAP7_75t_R _29552_ (.A1(_08880_),
    .A2(_09574_),
    .B(_09576_),
    .C(_08565_),
    .Y(_09577_));
 OA21x2_ASAP7_75t_R _29553_ (.A1(_09205_),
    .A2(_09577_),
    .B(_08344_),
    .Y(_09578_));
 OR2x2_ASAP7_75t_R _29554_ (.A(_09578_),
    .B(_09572_),
    .Y(_09579_));
 BUFx6f_ASAP7_75t_R _29555_ (.A(_09579_),
    .Y(_09580_));
 NAND2x1_ASAP7_75t_R _29556_ (.A(_01354_),
    .B(_09358_),
    .Y(_09581_));
 OA21x2_ASAP7_75t_R _29557_ (.A1(_08764_),
    .A2(_09580_),
    .B(_09581_),
    .Y(_02886_));
 INVx1_ASAP7_75t_R _29558_ (.A(_06438_),
    .Y(_09582_));
 INVx1_ASAP7_75t_R _29559_ (.A(_00270_),
    .Y(_09583_));
 OA21x2_ASAP7_75t_R _29560_ (.A1(_00264_),
    .A2(_09517_),
    .B(_00268_),
    .Y(_09584_));
 OAI21x1_ASAP7_75t_R _29561_ (.A1(_00267_),
    .A2(_09584_),
    .B(_00271_),
    .Y(_09585_));
 XNOR2x1_ASAP7_75t_R _29562_ (.B(_09585_),
    .Y(_09586_),
    .A(_09583_));
 AND2x2_ASAP7_75t_R _29563_ (.A(_09186_),
    .B(_09128_),
    .Y(_09587_));
 AO211x2_ASAP7_75t_R _29564_ (.A1(_08551_),
    .A2(_09586_),
    .B(_09587_),
    .C(_09362_),
    .Y(_09588_));
 AOI21x1_ASAP7_75t_R _29565_ (.A1(_08737_),
    .A2(_08738_),
    .B(_08477_),
    .Y(_09589_));
 AOI21x1_ASAP7_75t_R _29566_ (.A1(_08734_),
    .A2(_08735_),
    .B(_08467_),
    .Y(_09590_));
 OR3x1_ASAP7_75t_R _29567_ (.A(_08633_),
    .B(_09589_),
    .C(_09590_),
    .Y(_09591_));
 AO221x1_ASAP7_75t_R _29568_ (.A1(_08418_),
    .A2(_08419_),
    .B1(_08477_),
    .B2(_08707_),
    .C(_08710_),
    .Y(_09592_));
 AOI22x1_ASAP7_75t_R _29569_ (.A1(_18618_),
    .A2(_08487_),
    .B1(_08489_),
    .B2(_18613_),
    .Y(_09593_));
 AOI22x1_ASAP7_75t_R _29570_ (.A1(_18760_),
    .A2(_08484_),
    .B1(_08485_),
    .B2(_18752_),
    .Y(_09594_));
 AND3x1_ASAP7_75t_R _29571_ (.A(_08422_),
    .B(_09593_),
    .C(_09594_),
    .Y(_09595_));
 AND4x1_ASAP7_75t_R _29572_ (.A(_08497_),
    .B(_08531_),
    .C(_09524_),
    .D(_09525_),
    .Y(_09596_));
 AOI211x1_ASAP7_75t_R _29573_ (.A1(_08723_),
    .A2(_08724_),
    .B(_08657_),
    .C(_08527_),
    .Y(_09597_));
 OA211x2_ASAP7_75t_R _29574_ (.A1(_08720_),
    .A2(_08721_),
    .B(_08425_),
    .C(_08466_),
    .Y(_09598_));
 OR4x1_ASAP7_75t_R _29575_ (.A(_09595_),
    .B(_09596_),
    .C(_09597_),
    .D(_09598_),
    .Y(_09599_));
 AO32x2_ASAP7_75t_R _29576_ (.A1(_08919_),
    .A2(_09591_),
    .A3(_09592_),
    .B1(_09599_),
    .B2(_08631_),
    .Y(_09600_));
 AND3x1_ASAP7_75t_R _29577_ (.A(_08432_),
    .B(_08502_),
    .C(_08504_),
    .Y(_09601_));
 NAND2x1_ASAP7_75t_R _29578_ (.A(_08482_),
    .B(_08749_),
    .Y(_09602_));
 AOI22x1_ASAP7_75t_R _29579_ (.A1(_08643_),
    .A2(_08778_),
    .B1(_08779_),
    .B2(_08646_),
    .Y(_09603_));
 AO33x2_ASAP7_75t_R _29580_ (.A1(_09601_),
    .A2(_09602_),
    .A3(_09603_),
    .B1(_08920_),
    .B2(_08922_),
    .B3(_08636_),
    .Y(_09604_));
 OR3x1_ASAP7_75t_R _29581_ (.A(_08423_),
    .B(_09600_),
    .C(_09604_),
    .Y(_09605_));
 OA21x2_ASAP7_75t_R _29582_ (.A1(_08695_),
    .A2(_08655_),
    .B(_09117_),
    .Y(_09606_));
 INVx1_ASAP7_75t_R _29583_ (.A(_08648_),
    .Y(_09607_));
 AND3x1_ASAP7_75t_R _29584_ (.A(_08631_),
    .B(_08646_),
    .C(_09607_),
    .Y(_09608_));
 OAI22x1_ASAP7_75t_R _29585_ (.A1(_00357_),
    .A2(_08384_),
    .B1(_08389_),
    .B2(_00356_),
    .Y(_09609_));
 AND2x2_ASAP7_75t_R _29586_ (.A(_08381_),
    .B(_09609_),
    .Y(_09610_));
 AOI221x1_ASAP7_75t_R _29587_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_08669_),
    .B1(_08670_),
    .B2(_02283_),
    .C(_09610_),
    .Y(_09611_));
 OA31x2_ASAP7_75t_R _29588_ (.A1(_09285_),
    .A2(_09606_),
    .A3(_09608_),
    .B1(_09611_),
    .Y(_09612_));
 AO21x1_ASAP7_75t_R _29589_ (.A1(_09605_),
    .A2(_09612_),
    .B(_09056_),
    .Y(_09613_));
 OR3x1_ASAP7_75t_R _29590_ (.A(_13595_),
    .B(_05320_),
    .C(_05141_),
    .Y(_09614_));
 AND5x2_ASAP7_75t_R _29591_ (.A(_09582_),
    .B(_08599_),
    .C(_09588_),
    .D(_09613_),
    .E(_09614_),
    .Y(_09615_));
 OA211x2_ASAP7_75t_R _29592_ (.A1(_08770_),
    .A2(_08908_),
    .B(_09139_),
    .C(_08880_),
    .Y(_09616_));
 NAND2x1_ASAP7_75t_R _29593_ (.A(net76),
    .B(_08902_),
    .Y(_09617_));
 OA211x2_ASAP7_75t_R _29594_ (.A1(_09383_),
    .A2(_08947_),
    .B(_09617_),
    .C(_08885_),
    .Y(_09618_));
 OR3x2_ASAP7_75t_R _29595_ (.A(_08689_),
    .B(_09616_),
    .C(_09618_),
    .Y(_09619_));
 AND3x2_ASAP7_75t_R _29596_ (.A(_08345_),
    .B(_09215_),
    .C(_09619_),
    .Y(_09620_));
 NOR2x2_ASAP7_75t_R _29597_ (.A(_09615_),
    .B(_09620_),
    .Y(_09621_));
 BUFx3_ASAP7_75t_R _29598_ (.A(_09621_),
    .Y(_09622_));
 NOR2x1_ASAP7_75t_R _29599_ (.A(_01387_),
    .B(_08598_),
    .Y(_09623_));
 AO21x1_ASAP7_75t_R _29600_ (.A1(_08598_),
    .A2(net151),
    .B(_09623_),
    .Y(_02887_));
 AND3x1_ASAP7_75t_R _29601_ (.A(_08777_),
    .B(_08509_),
    .C(_08541_),
    .Y(_09624_));
 OAI22x1_ASAP7_75t_R _29602_ (.A1(_00358_),
    .A2(_08385_),
    .B1(_08390_),
    .B2(_01451_),
    .Y(_09625_));
 AND2x2_ASAP7_75t_R _29603_ (.A(_02299_),
    .B(_08394_),
    .Y(_09626_));
 AO21x1_ASAP7_75t_R _29604_ (.A1(_08382_),
    .A2(_09625_),
    .B(_09626_),
    .Y(_09627_));
 OR2x2_ASAP7_75t_R _29605_ (.A(_00267_),
    .B(_00270_),
    .Y(_09628_));
 OA21x2_ASAP7_75t_R _29606_ (.A1(_00271_),
    .A2(_00270_),
    .B(_00275_),
    .Y(_09629_));
 OA21x2_ASAP7_75t_R _29607_ (.A1(_09561_),
    .A2(_09628_),
    .B(_09629_),
    .Y(_09630_));
 OR4x1_ASAP7_75t_R _29608_ (.A(_13566_),
    .B(_00274_),
    .C(_09185_),
    .D(_09630_),
    .Y(_09631_));
 AND4x1_ASAP7_75t_R _29609_ (.A(_13593_),
    .B(_00274_),
    .C(_08549_),
    .D(_09630_),
    .Y(_09632_));
 INVx1_ASAP7_75t_R _29610_ (.A(_09632_),
    .Y(_09633_));
 OR3x1_ASAP7_75t_R _29611_ (.A(_13566_),
    .B(_08549_),
    .C(_09157_),
    .Y(_09634_));
 OA21x2_ASAP7_75t_R _29612_ (.A1(_08753_),
    .A2(_04869_),
    .B(_09634_),
    .Y(_09635_));
 AND4x2_ASAP7_75t_R _29613_ (.A(_05514_),
    .B(_09631_),
    .C(_09633_),
    .D(_09635_),
    .Y(_09636_));
 AND3x1_ASAP7_75t_R _29614_ (.A(_08632_),
    .B(_08427_),
    .C(_08542_),
    .Y(_09637_));
 AO21x1_ASAP7_75t_R _29615_ (.A1(\alu_adder_result_ex[31] ),
    .A2(_08393_),
    .B(_05078_),
    .Y(_09638_));
 OR5x1_ASAP7_75t_R _29616_ (.A(_09432_),
    .B(_09636_),
    .C(_09627_),
    .D(_09637_),
    .E(_09638_),
    .Y(_09639_));
 AOI211x1_ASAP7_75t_R _29617_ (.A1(_08500_),
    .A2(_09253_),
    .B(_09624_),
    .C(_09639_),
    .Y(_09640_));
 NOR2x1_ASAP7_75t_R _29618_ (.A(_09377_),
    .B(_09636_),
    .Y(_09641_));
 AO21x1_ASAP7_75t_R _29619_ (.A1(_05078_),
    .A2(_06453_),
    .B(_09641_),
    .Y(_09642_));
 OA21x2_ASAP7_75t_R _29620_ (.A1(_09642_),
    .A2(_09640_),
    .B(_08600_),
    .Y(_09643_));
 NOR2x1_ASAP7_75t_R _29621_ (.A(_08950_),
    .B(_09173_),
    .Y(_09644_));
 AO21x1_ASAP7_75t_R _29622_ (.A1(_08945_),
    .A2(_09175_),
    .B(_09644_),
    .Y(_09645_));
 OA211x2_ASAP7_75t_R _29623_ (.A1(_08689_),
    .A2(_09645_),
    .B(_09215_),
    .C(_08683_),
    .Y(_09646_));
 NOR2x2_ASAP7_75t_R _29624_ (.A(_09646_),
    .B(_09643_),
    .Y(_09647_));
 BUFx3_ASAP7_75t_R _29625_ (.A(_09647_),
    .Y(_09648_));
 AND2x2_ASAP7_75t_R _29626_ (.A(_04799_),
    .B(_08680_),
    .Y(_09649_));
 AO21x1_ASAP7_75t_R _29627_ (.A1(_08598_),
    .A2(net7),
    .B(_09649_),
    .Y(_02888_));
 BUFx6f_ASAP7_75t_R _29628_ (.A(_08584_),
    .Y(_09650_));
 AND2x2_ASAP7_75t_R _29629_ (.A(_14726_),
    .B(_13438_),
    .Y(_09651_));
 AND2x4_ASAP7_75t_R _29630_ (.A(_09651_),
    .B(_08596_),
    .Y(_09652_));
 NAND2x2_ASAP7_75t_R _29631_ (.A(_08339_),
    .B(_09652_),
    .Y(_09653_));
 BUFx10_ASAP7_75t_R _29632_ (.A(_09653_),
    .Y(_09654_));
 BUFx6f_ASAP7_75t_R _29633_ (.A(_09654_),
    .Y(_09655_));
 BUFx6f_ASAP7_75t_R _29634_ (.A(_09653_),
    .Y(_09656_));
 NAND2x1_ASAP7_75t_R _29635_ (.A(_00419_),
    .B(_09656_),
    .Y(_09657_));
 OA21x2_ASAP7_75t_R _29636_ (.A1(_09650_),
    .A2(_09655_),
    .B(_09657_),
    .Y(_02889_));
 OA21x2_ASAP7_75t_R _29637_ (.A1(_08433_),
    .A2(_09119_),
    .B(_08616_),
    .Y(_09658_));
 OAI22x1_ASAP7_75t_R _29638_ (.A1(_00299_),
    .A2(_08665_),
    .B1(_08667_),
    .B2(_00298_),
    .Y(_09659_));
 AO22x1_ASAP7_75t_R _29639_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_08393_),
    .B1(_08395_),
    .B2(_02254_),
    .Y(_09660_));
 AO21x1_ASAP7_75t_R _29640_ (.A1(_08663_),
    .A2(_09659_),
    .B(_09660_),
    .Y(_09661_));
 NOR3x1_ASAP7_75t_R _29641_ (.A(_09285_),
    .B(_09600_),
    .C(_09604_),
    .Y(_09662_));
 OR3x1_ASAP7_75t_R _29642_ (.A(_09658_),
    .B(_09661_),
    .C(_09662_),
    .Y(_09663_));
 AND3x1_ASAP7_75t_R _29643_ (.A(_13595_),
    .B(_00137_),
    .C(_08551_),
    .Y(_09664_));
 AO21x1_ASAP7_75t_R _29644_ (.A1(_00414_),
    .A2(_08548_),
    .B(_09664_),
    .Y(_09665_));
 OAI21x1_ASAP7_75t_R _29645_ (.A1(_05142_),
    .A2(_09665_),
    .B(_06194_),
    .Y(_09666_));
 INVx1_ASAP7_75t_R _29646_ (.A(_01494_),
    .Y(_09667_));
 AO21x1_ASAP7_75t_R _29647_ (.A1(_09667_),
    .A2(_08566_),
    .B(_08902_),
    .Y(_09668_));
 NOR2x1_ASAP7_75t_R _29648_ (.A(_01482_),
    .B(_08570_),
    .Y(_09669_));
 AO21x1_ASAP7_75t_R _29649_ (.A1(net79),
    .A2(_08570_),
    .B(_09669_),
    .Y(_09670_));
 OAI22x1_ASAP7_75t_R _29650_ (.A1(_09446_),
    .A2(_08564_),
    .B1(_08576_),
    .B2(_01497_),
    .Y(_09671_));
 AO32x1_ASAP7_75t_R _29651_ (.A1(net103),
    .A2(_08563_),
    .A3(_08570_),
    .B1(_08575_),
    .B2(_09671_),
    .Y(_09672_));
 AO221x1_ASAP7_75t_R _29652_ (.A1(_08910_),
    .A2(_09668_),
    .B1(_09670_),
    .B2(_08956_),
    .C(_09672_),
    .Y(_09673_));
 OA211x2_ASAP7_75t_R _29653_ (.A1(net82),
    .A2(_08901_),
    .B(_09673_),
    .C(_08344_),
    .Y(_09674_));
 AO221x2_ASAP7_75t_R _29654_ (.A1(_09261_),
    .A2(_09663_),
    .B1(_09666_),
    .B2(_08600_),
    .C(_09674_),
    .Y(_09675_));
 BUFx6f_ASAP7_75t_R _29655_ (.A(_09675_),
    .Y(_09676_));
 BUFx10_ASAP7_75t_R _29656_ (.A(_09654_),
    .Y(_09677_));
 NAND2x1_ASAP7_75t_R _29657_ (.A(_00372_),
    .B(_09677_),
    .Y(_09678_));
 OA21x2_ASAP7_75t_R _29658_ (.A1(_09655_),
    .A2(_09676_),
    .B(_09678_),
    .Y(_02890_));
 NAND2x1_ASAP7_75t_R _29659_ (.A(_01811_),
    .B(_08591_),
    .Y(_09679_));
 OA21x2_ASAP7_75t_R _29660_ (.A1(_09107_),
    .A2(_09074_),
    .B(_09679_),
    .Y(_02891_));
 AO221x1_ASAP7_75t_R _29661_ (.A1(net80),
    .A2(_08603_),
    .B1(_08604_),
    .B2(net49),
    .C(_08685_),
    .Y(_09680_));
 INVx1_ASAP7_75t_R _29662_ (.A(_01489_),
    .Y(_09681_));
 AO221x1_ASAP7_75t_R _29663_ (.A1(_08958_),
    .A2(_08603_),
    .B1(_08604_),
    .B2(_09681_),
    .C(_08570_),
    .Y(_09682_));
 OAI22x1_ASAP7_75t_R _29664_ (.A1(_08946_),
    .A2(_08564_),
    .B1(_08577_),
    .B2(_01496_),
    .Y(_09683_));
 AO222x2_ASAP7_75t_R _29665_ (.A1(net93),
    .A2(_08581_),
    .B1(_09680_),
    .B2(_09682_),
    .C1(_09683_),
    .C2(_08575_),
    .Y(_09684_));
 OAI21x1_ASAP7_75t_R _29666_ (.A1(_09535_),
    .A2(_09567_),
    .B(_08777_),
    .Y(_09685_));
 AND3x1_ASAP7_75t_R _29667_ (.A(_08753_),
    .B(_00140_),
    .C(_08550_),
    .Y(_09686_));
 AO21x1_ASAP7_75t_R _29668_ (.A1(_00792_),
    .A2(_08547_),
    .B(_09686_),
    .Y(_09687_));
 OA22x2_ASAP7_75t_R _29669_ (.A1(_00301_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00300_),
    .Y(_09688_));
 AOI22x1_ASAP7_75t_R _29670_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_08669_),
    .B1(_08394_),
    .B2(_02255_),
    .Y(_09689_));
 OA21x2_ASAP7_75t_R _29671_ (.A1(_08670_),
    .A2(_09688_),
    .B(_09689_),
    .Y(_09690_));
 OA222x2_ASAP7_75t_R _29672_ (.A1(_13603_),
    .A2(_14730_),
    .B1(_05141_),
    .B2(_09687_),
    .C1(_09690_),
    .C2(_09056_),
    .Y(_09691_));
 OR4x1_ASAP7_75t_R _29673_ (.A(_09285_),
    .B(_09549_),
    .C(_09550_),
    .D(_09551_),
    .Y(_09692_));
 NAND3x1_ASAP7_75t_R _29674_ (.A(_09685_),
    .B(_09691_),
    .C(_09692_),
    .Y(_09693_));
 OA211x2_ASAP7_75t_R _29675_ (.A1(_08554_),
    .A2(_05870_),
    .B(_08694_),
    .C(_09693_),
    .Y(_09694_));
 AO21x2_ASAP7_75t_R _29676_ (.A1(_08684_),
    .A2(_09684_),
    .B(_09694_),
    .Y(_09695_));
 BUFx6f_ASAP7_75t_R _29677_ (.A(_09695_),
    .Y(_09696_));
 NAND2x1_ASAP7_75t_R _29678_ (.A(_00483_),
    .B(_09677_),
    .Y(_09697_));
 OA21x2_ASAP7_75t_R _29679_ (.A1(_09655_),
    .A2(_09696_),
    .B(_09697_),
    .Y(_02892_));
 AO221x1_ASAP7_75t_R _29680_ (.A1(net81),
    .A2(_08603_),
    .B1(_08604_),
    .B2(net50),
    .C(_08566_),
    .Y(_09698_));
 INVx1_ASAP7_75t_R _29681_ (.A(_01488_),
    .Y(_09699_));
 AO221x1_ASAP7_75t_R _29682_ (.A1(_09001_),
    .A2(_08603_),
    .B1(_08604_),
    .B2(_09699_),
    .C(_08570_),
    .Y(_09700_));
 OAI22x1_ASAP7_75t_R _29683_ (.A1(_08992_),
    .A2(_08564_),
    .B1(_08577_),
    .B2(_01495_),
    .Y(_09701_));
 AO222x2_ASAP7_75t_R _29684_ (.A1(net97),
    .A2(_08581_),
    .B1(_09698_),
    .B2(_09700_),
    .C1(_09701_),
    .C2(_08575_),
    .Y(_09702_));
 AND4x1_ASAP7_75t_R _29685_ (.A(_08366_),
    .B(_08632_),
    .C(_08633_),
    .D(_09050_),
    .Y(_09703_));
 OA211x2_ASAP7_75t_R _29686_ (.A1(_08695_),
    .A2(_08482_),
    .B(_08411_),
    .C(_08366_),
    .Y(_09704_));
 OAI22x1_ASAP7_75t_R _29687_ (.A1(_00303_),
    .A2(_08664_),
    .B1(_08666_),
    .B2(_00302_),
    .Y(_09705_));
 AO22x1_ASAP7_75t_R _29688_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_08360_),
    .B1(_08380_),
    .B2(_02256_),
    .Y(_09706_));
 AO21x1_ASAP7_75t_R _29689_ (.A1(_08381_),
    .A2(_09705_),
    .B(_09706_),
    .Y(_09707_));
 INVx1_ASAP7_75t_R _29690_ (.A(_00146_),
    .Y(_09708_));
 AO21x1_ASAP7_75t_R _29691_ (.A1(_08753_),
    .A2(_08549_),
    .B(_05545_),
    .Y(_09709_));
 OA211x2_ASAP7_75t_R _29692_ (.A1(_09708_),
    .A2(_08547_),
    .B(_09709_),
    .C(_05304_),
    .Y(_09710_));
 AO21x1_ASAP7_75t_R _29693_ (.A1(_08375_),
    .A2(_09707_),
    .B(_09710_),
    .Y(_09711_));
 OR3x1_ASAP7_75t_R _29694_ (.A(_09703_),
    .B(_09704_),
    .C(_09711_),
    .Y(_09712_));
 AO21x1_ASAP7_75t_R _29695_ (.A1(_08542_),
    .A2(_09530_),
    .B(_09712_),
    .Y(_09713_));
 OA21x2_ASAP7_75t_R _29696_ (.A1(_06499_),
    .A2(_09713_),
    .B(_08694_),
    .Y(_09714_));
 AO21x2_ASAP7_75t_R _29697_ (.A1(_08684_),
    .A2(_09702_),
    .B(_09714_),
    .Y(_09715_));
 BUFx6f_ASAP7_75t_R _29698_ (.A(_09715_),
    .Y(_09716_));
 NAND2x1_ASAP7_75t_R _29699_ (.A(_00514_),
    .B(_09677_),
    .Y(_09717_));
 OA21x2_ASAP7_75t_R _29700_ (.A1(_09655_),
    .A2(_09716_),
    .B(_09717_),
    .Y(_02893_));
 BUFx6f_ASAP7_75t_R _29701_ (.A(_08675_),
    .Y(_09718_));
 AND2x6_ASAP7_75t_R _29702_ (.A(_08595_),
    .B(_09652_),
    .Y(_09719_));
 NOR2x1_ASAP7_75t_R _29703_ (.A(_00544_),
    .B(_09719_),
    .Y(_09720_));
 AO21x1_ASAP7_75t_R _29704_ (.A1(_09718_),
    .A2(_09719_),
    .B(_09720_),
    .Y(_02894_));
 BUFx6f_ASAP7_75t_R _29705_ (.A(_08762_),
    .Y(_09721_));
 NAND2x1_ASAP7_75t_R _29706_ (.A(_00576_),
    .B(_09677_),
    .Y(_09722_));
 OA21x2_ASAP7_75t_R _29707_ (.A1(_09721_),
    .A2(_09655_),
    .B(_09722_),
    .Y(_02895_));
 NAND2x1_ASAP7_75t_R _29708_ (.A(_00606_),
    .B(_09677_),
    .Y(_09723_));
 OA21x2_ASAP7_75t_R _29709_ (.A1(_08810_),
    .A2(_09655_),
    .B(_09723_),
    .Y(_02896_));
 NAND2x1_ASAP7_75t_R _29710_ (.A(_00636_),
    .B(_09677_),
    .Y(_09724_));
 OA21x2_ASAP7_75t_R _29711_ (.A1(_08851_),
    .A2(_09655_),
    .B(_09724_),
    .Y(_02897_));
 AO21x1_ASAP7_75t_R _29712_ (.A1(_08595_),
    .A2(_09652_),
    .B(_00666_),
    .Y(_09725_));
 OAI21x1_ASAP7_75t_R _29713_ (.A1(_08898_),
    .A2(_09655_),
    .B(_09725_),
    .Y(_02898_));
 NAND2x1_ASAP7_75t_R _29714_ (.A(_00696_),
    .B(_09677_),
    .Y(_09726_));
 OA21x2_ASAP7_75t_R _29715_ (.A1(_08943_),
    .A2(_09655_),
    .B(_09726_),
    .Y(_02899_));
 NAND2x1_ASAP7_75t_R _29716_ (.A(_00726_),
    .B(_09677_),
    .Y(_09727_));
 OA21x2_ASAP7_75t_R _29717_ (.A1(_08989_),
    .A2(_09655_),
    .B(_09727_),
    .Y(_02900_));
 BUFx10_ASAP7_75t_R _29718_ (.A(_09036_),
    .Y(_09728_));
 BUFx4f_ASAP7_75t_R _29719_ (.A(_09654_),
    .Y(_09729_));
 NAND2x1_ASAP7_75t_R _29720_ (.A(_00756_),
    .B(_09677_),
    .Y(_09730_));
 OA21x2_ASAP7_75t_R _29721_ (.A1(_09728_),
    .A2(_09729_),
    .B(_09730_),
    .Y(_02901_));
 BUFx6f_ASAP7_75t_R _29722_ (.A(_09103_),
    .Y(_09731_));
 NAND2x1_ASAP7_75t_R _29723_ (.A(_01810_),
    .B(_08591_),
    .Y(_09732_));
 OA21x2_ASAP7_75t_R _29724_ (.A1(_09107_),
    .A2(_09731_),
    .B(_09732_),
    .Y(_02902_));
 NAND2x1_ASAP7_75t_R _29725_ (.A(_00452_),
    .B(_09677_),
    .Y(_09733_));
 OA21x2_ASAP7_75t_R _29726_ (.A1(_09074_),
    .A2(_09729_),
    .B(_09733_),
    .Y(_02903_));
 BUFx6f_ASAP7_75t_R _29727_ (.A(_09653_),
    .Y(_09734_));
 NAND2x1_ASAP7_75t_R _29728_ (.A(_00827_),
    .B(_09734_),
    .Y(_09735_));
 OA21x2_ASAP7_75t_R _29729_ (.A1(_09104_),
    .A2(_09729_),
    .B(_09735_),
    .Y(_02904_));
 NAND2x1_ASAP7_75t_R _29730_ (.A(_00860_),
    .B(_09734_),
    .Y(_09736_));
 OA21x2_ASAP7_75t_R _29731_ (.A1(_09144_),
    .A2(_09729_),
    .B(_09736_),
    .Y(_02905_));
 NAND2x1_ASAP7_75t_R _29732_ (.A(_00893_),
    .B(_09734_),
    .Y(_09737_));
 OA21x2_ASAP7_75t_R _29733_ (.A1(_09181_),
    .A2(_09729_),
    .B(_09737_),
    .Y(_02906_));
 BUFx4f_ASAP7_75t_R _29734_ (.A(_09213_),
    .Y(_09738_));
 NAND2x1_ASAP7_75t_R _29735_ (.A(_00926_),
    .B(_09734_),
    .Y(_09739_));
 OA21x2_ASAP7_75t_R _29736_ (.A1(_09738_),
    .A2(_09729_),
    .B(_09739_),
    .Y(_02907_));
 NAND2x1_ASAP7_75t_R _29737_ (.A(_00959_),
    .B(_09734_),
    .Y(_09740_));
 OA21x2_ASAP7_75t_R _29738_ (.A1(_09245_),
    .A2(_09729_),
    .B(_09740_),
    .Y(_02908_));
 NAND2x1_ASAP7_75t_R _29739_ (.A(_00992_),
    .B(_09734_),
    .Y(_09741_));
 OA21x2_ASAP7_75t_R _29740_ (.A1(_09271_),
    .A2(_09729_),
    .B(_09741_),
    .Y(_02909_));
 NAND2x1_ASAP7_75t_R _29741_ (.A(_01025_),
    .B(_09734_),
    .Y(_09742_));
 OA21x2_ASAP7_75t_R _29742_ (.A1(_09299_),
    .A2(_09729_),
    .B(_09742_),
    .Y(_02910_));
 NAND2x1_ASAP7_75t_R _29743_ (.A(_01058_),
    .B(_09734_),
    .Y(_09743_));
 OA21x2_ASAP7_75t_R _29744_ (.A1(_09328_),
    .A2(_09729_),
    .B(_09743_),
    .Y(_02911_));
 NAND2x1_ASAP7_75t_R _29745_ (.A(_01091_),
    .B(_09734_),
    .Y(_09744_));
 OA21x2_ASAP7_75t_R _29746_ (.A1(_09357_),
    .A2(_09656_),
    .B(_09744_),
    .Y(_02912_));
 BUFx4f_ASAP7_75t_R _29747_ (.A(_09143_),
    .Y(_09745_));
 NAND2x1_ASAP7_75t_R _29748_ (.A(_01809_),
    .B(_08591_),
    .Y(_09746_));
 OA21x2_ASAP7_75t_R _29749_ (.A1(_09107_),
    .A2(_09745_),
    .B(_09746_),
    .Y(_02913_));
 NAND2x1_ASAP7_75t_R _29750_ (.A(_01124_),
    .B(_09734_),
    .Y(_09747_));
 OA21x2_ASAP7_75t_R _29751_ (.A1(_09390_),
    .A2(_09656_),
    .B(_09747_),
    .Y(_02914_));
 NAND2x1_ASAP7_75t_R _29752_ (.A(_01157_),
    .B(_09654_),
    .Y(_09748_));
 OA21x2_ASAP7_75t_R _29753_ (.A1(_09416_),
    .A2(_09656_),
    .B(_09748_),
    .Y(_02915_));
 BUFx4f_ASAP7_75t_R _29754_ (.A(_09441_),
    .Y(_09749_));
 NAND2x1_ASAP7_75t_R _29755_ (.A(_01190_),
    .B(_09654_),
    .Y(_09750_));
 OA21x2_ASAP7_75t_R _29756_ (.A1(_09749_),
    .A2(_09656_),
    .B(_09750_),
    .Y(_02916_));
 NAND2x1_ASAP7_75t_R _29757_ (.A(_01223_),
    .B(_09654_),
    .Y(_09751_));
 OA21x2_ASAP7_75t_R _29758_ (.A1(_09472_),
    .A2(_09656_),
    .B(_09751_),
    .Y(_02917_));
 NAND2x1_ASAP7_75t_R _29759_ (.A(_01256_),
    .B(_09654_),
    .Y(_09752_));
 OA21x2_ASAP7_75t_R _29760_ (.A1(_09495_),
    .A2(_09656_),
    .B(_09752_),
    .Y(_02918_));
 BUFx3_ASAP7_75t_R _29761_ (.A(_09512_),
    .Y(_09753_));
 NAND2x1_ASAP7_75t_R _29762_ (.A(_01289_),
    .B(_09654_),
    .Y(_09754_));
 OA21x2_ASAP7_75t_R _29763_ (.A1(_09753_),
    .A2(_09656_),
    .B(_09754_),
    .Y(_02919_));
 BUFx6f_ASAP7_75t_R _29764_ (.A(_09543_),
    .Y(_09755_));
 NAND2x1_ASAP7_75t_R _29765_ (.A(_01322_),
    .B(_09654_),
    .Y(_09756_));
 OA21x2_ASAP7_75t_R _29766_ (.A1(_09755_),
    .A2(_09656_),
    .B(_09756_),
    .Y(_02920_));
 BUFx3_ASAP7_75t_R _29767_ (.A(_09580_),
    .Y(_09757_));
 NAND2x1_ASAP7_75t_R _29768_ (.A(_01355_),
    .B(_09654_),
    .Y(_09758_));
 OA21x2_ASAP7_75t_R _29769_ (.A1(net13),
    .A2(_09656_),
    .B(_09758_),
    .Y(_02921_));
 BUFx3_ASAP7_75t_R _29770_ (.A(_09621_),
    .Y(_09759_));
 NOR2x1_ASAP7_75t_R _29771_ (.A(_01388_),
    .B(_09719_),
    .Y(_09760_));
 AO21x1_ASAP7_75t_R _29772_ (.A1(net152),
    .A2(_09719_),
    .B(_09760_),
    .Y(_02922_));
 BUFx3_ASAP7_75t_R _29773_ (.A(_09647_),
    .Y(_09761_));
 NOR2x1_ASAP7_75t_R _29774_ (.A(_01421_),
    .B(_09719_),
    .Y(_09762_));
 AO21x1_ASAP7_75t_R _29775_ (.A1(net8),
    .A2(_09719_),
    .B(_09762_),
    .Y(_02923_));
 BUFx6f_ASAP7_75t_R _29776_ (.A(_09180_),
    .Y(_09763_));
 BUFx10_ASAP7_75t_R _29777_ (.A(_08590_),
    .Y(_09764_));
 NAND2x1_ASAP7_75t_R _29778_ (.A(_01808_),
    .B(_09764_),
    .Y(_09765_));
 OA21x2_ASAP7_75t_R _29779_ (.A1(_09107_),
    .A2(_09763_),
    .B(_09765_),
    .Y(_02924_));
 BUFx3_ASAP7_75t_R _29780_ (.A(_08587_),
    .Y(_09766_));
 NAND2x2_ASAP7_75t_R _29781_ (.A(_08027_),
    .B(_13439_),
    .Y(_09767_));
 OR3x1_ASAP7_75t_R _29782_ (.A(_09766_),
    .B(_08678_),
    .C(_09767_),
    .Y(_09768_));
 BUFx10_ASAP7_75t_R _29783_ (.A(_09768_),
    .Y(_09769_));
 BUFx6f_ASAP7_75t_R _29784_ (.A(_09769_),
    .Y(_09770_));
 NAND2x1_ASAP7_75t_R _29785_ (.A(_00420_),
    .B(_09770_),
    .Y(_09771_));
 OA21x2_ASAP7_75t_R _29786_ (.A1(_09650_),
    .A2(_09770_),
    .B(_09771_),
    .Y(_02925_));
 BUFx3_ASAP7_75t_R _29787_ (.A(_09675_),
    .Y(_09772_));
 BUFx4f_ASAP7_75t_R _29788_ (.A(_13439_),
    .Y(_09773_));
 AND2x4_ASAP7_75t_R _29789_ (.A(_08027_),
    .B(_09773_),
    .Y(_09774_));
 AND3x1_ASAP7_75t_R _29790_ (.A(_08339_),
    .B(_08596_),
    .C(_09774_),
    .Y(_09775_));
 BUFx6f_ASAP7_75t_R _29791_ (.A(_09775_),
    .Y(_09776_));
 BUFx4f_ASAP7_75t_R _29792_ (.A(_09776_),
    .Y(_09777_));
 BUFx4f_ASAP7_75t_R _29793_ (.A(_09769_),
    .Y(_09778_));
 AND2x2_ASAP7_75t_R _29794_ (.A(_13474_),
    .B(_09778_),
    .Y(_09779_));
 AO21x1_ASAP7_75t_R _29795_ (.A1(_09772_),
    .A2(_09777_),
    .B(_09779_),
    .Y(_02926_));
 BUFx6f_ASAP7_75t_R _29796_ (.A(_09695_),
    .Y(_09780_));
 NAND2x1_ASAP7_75t_R _29797_ (.A(_00484_),
    .B(_09770_),
    .Y(_09781_));
 OA21x2_ASAP7_75t_R _29798_ (.A1(_09780_),
    .A2(_09770_),
    .B(_09781_),
    .Y(_02927_));
 BUFx4f_ASAP7_75t_R _29799_ (.A(_09715_),
    .Y(_09782_));
 AND2x2_ASAP7_75t_R _29800_ (.A(_14218_),
    .B(_09778_),
    .Y(_09783_));
 AO21x1_ASAP7_75t_R _29801_ (.A1(_09782_),
    .A2(_09777_),
    .B(_09783_),
    .Y(_02928_));
 AND2x2_ASAP7_75t_R _29802_ (.A(_15007_),
    .B(_09778_),
    .Y(_09784_));
 AO21x1_ASAP7_75t_R _29803_ (.A1(_09718_),
    .A2(_09777_),
    .B(_09784_),
    .Y(_02929_));
 NAND2x1_ASAP7_75t_R _29804_ (.A(_00577_),
    .B(_09770_),
    .Y(_09785_));
 OA21x2_ASAP7_75t_R _29805_ (.A1(_09721_),
    .A2(_09770_),
    .B(_09785_),
    .Y(_02930_));
 BUFx4f_ASAP7_75t_R _29806_ (.A(_08809_),
    .Y(_09786_));
 AND2x2_ASAP7_75t_R _29807_ (.A(_15144_),
    .B(_09778_),
    .Y(_09787_));
 AO21x1_ASAP7_75t_R _29808_ (.A1(_09786_),
    .A2(_09777_),
    .B(_09787_),
    .Y(_02931_));
 BUFx6f_ASAP7_75t_R _29809_ (.A(_08850_),
    .Y(_09788_));
 AND2x2_ASAP7_75t_R _29810_ (.A(_14450_),
    .B(_09778_),
    .Y(_09789_));
 AO21x1_ASAP7_75t_R _29811_ (.A1(_09788_),
    .A2(_09777_),
    .B(_09789_),
    .Y(_02932_));
 BUFx6f_ASAP7_75t_R _29812_ (.A(_08870_),
    .Y(_09790_));
 BUFx6f_ASAP7_75t_R _29813_ (.A(_08895_),
    .Y(_09791_));
 OR3x1_ASAP7_75t_R _29814_ (.A(_09790_),
    .B(_09791_),
    .C(_09778_),
    .Y(_09792_));
 OAI21x1_ASAP7_75t_R _29815_ (.A1(_00667_),
    .A2(_09777_),
    .B(_09792_),
    .Y(_02933_));
 AND2x2_ASAP7_75t_R _29816_ (.A(_14590_),
    .B(_09778_),
    .Y(_09793_));
 AO21x1_ASAP7_75t_R _29817_ (.A1(_08943_),
    .A2(_09777_),
    .B(_09793_),
    .Y(_02934_));
 AND2x4_ASAP7_75t_R _29818_ (.A(_14051_),
    .B(_08341_),
    .Y(_09794_));
 AND3x1_ASAP7_75t_R _29819_ (.A(_14051_),
    .B(_08595_),
    .C(_09651_),
    .Y(_09795_));
 BUFx4f_ASAP7_75t_R _29820_ (.A(_09795_),
    .Y(_09796_));
 NOR2x1_ASAP7_75t_R _29821_ (.A(_01807_),
    .B(_09796_),
    .Y(_09797_));
 AO21x1_ASAP7_75t_R _29822_ (.A1(_09794_),
    .A2(_09213_),
    .B(_09797_),
    .Y(_02935_));
 AND2x2_ASAP7_75t_R _29823_ (.A(_14609_),
    .B(_09778_),
    .Y(_09798_));
 AO21x1_ASAP7_75t_R _29824_ (.A1(_09108_),
    .A2(_09777_),
    .B(_09798_),
    .Y(_02936_));
 AND2x2_ASAP7_75t_R _29825_ (.A(_14669_),
    .B(_09778_),
    .Y(_09799_));
 AO21x1_ASAP7_75t_R _29826_ (.A1(_09037_),
    .A2(_09777_),
    .B(_09799_),
    .Y(_02937_));
 BUFx4f_ASAP7_75t_R _29827_ (.A(_09073_),
    .Y(_09800_));
 AND2x2_ASAP7_75t_R _29828_ (.A(_13967_),
    .B(_09778_),
    .Y(_09801_));
 AO21x1_ASAP7_75t_R _29829_ (.A1(_09800_),
    .A2(_09777_),
    .B(_09801_),
    .Y(_02938_));
 BUFx4f_ASAP7_75t_R _29830_ (.A(_09776_),
    .Y(_09802_));
 BUFx4f_ASAP7_75t_R _29831_ (.A(_09769_),
    .Y(_09803_));
 AND2x2_ASAP7_75t_R _29832_ (.A(_15616_),
    .B(_09803_),
    .Y(_09804_));
 AO21x1_ASAP7_75t_R _29833_ (.A1(_09731_),
    .A2(_09802_),
    .B(_09804_),
    .Y(_02939_));
 AND2x2_ASAP7_75t_R _29834_ (.A(_15770_),
    .B(_09803_),
    .Y(_09805_));
 AO21x1_ASAP7_75t_R _29835_ (.A1(_09745_),
    .A2(_09802_),
    .B(_09805_),
    .Y(_02940_));
 AND2x2_ASAP7_75t_R _29836_ (.A(_15896_),
    .B(_09803_),
    .Y(_09806_));
 AO21x1_ASAP7_75t_R _29837_ (.A1(_09763_),
    .A2(_09802_),
    .B(_09806_),
    .Y(_02941_));
 AND2x2_ASAP7_75t_R _29838_ (.A(_16047_),
    .B(_09803_),
    .Y(_09807_));
 AO21x1_ASAP7_75t_R _29839_ (.A1(_09738_),
    .A2(_09802_),
    .B(_09807_),
    .Y(_02942_));
 BUFx6f_ASAP7_75t_R _29840_ (.A(_09244_),
    .Y(_09808_));
 AND2x2_ASAP7_75t_R _29841_ (.A(_16165_),
    .B(_09803_),
    .Y(_09809_));
 AO21x1_ASAP7_75t_R _29842_ (.A1(_09808_),
    .A2(_09802_),
    .B(_09809_),
    .Y(_02943_));
 BUFx6f_ASAP7_75t_R _29843_ (.A(_09270_),
    .Y(_09810_));
 AND2x2_ASAP7_75t_R _29844_ (.A(_16307_),
    .B(_09803_),
    .Y(_09811_));
 AO21x1_ASAP7_75t_R _29845_ (.A1(_09810_),
    .A2(_09802_),
    .B(_09811_),
    .Y(_02944_));
 BUFx6f_ASAP7_75t_R _29846_ (.A(_09298_),
    .Y(_09812_));
 AND2x2_ASAP7_75t_R _29847_ (.A(_16421_),
    .B(_09803_),
    .Y(_09813_));
 AO21x1_ASAP7_75t_R _29848_ (.A1(_09812_),
    .A2(_09802_),
    .B(_09813_),
    .Y(_02945_));
 NAND2x1_ASAP7_75t_R _29849_ (.A(_01806_),
    .B(_09764_),
    .Y(_09814_));
 OA21x2_ASAP7_75t_R _29850_ (.A1(_09107_),
    .A2(_09808_),
    .B(_09814_),
    .Y(_02946_));
 BUFx6f_ASAP7_75t_R _29851_ (.A(_09327_),
    .Y(_09815_));
 AND2x2_ASAP7_75t_R _29852_ (.A(_16548_),
    .B(_09803_),
    .Y(_09816_));
 AO21x1_ASAP7_75t_R _29853_ (.A1(_09815_),
    .A2(_09802_),
    .B(_09816_),
    .Y(_02947_));
 BUFx6f_ASAP7_75t_R _29854_ (.A(_09356_),
    .Y(_09817_));
 AND2x2_ASAP7_75t_R _29855_ (.A(_16662_),
    .B(_09803_),
    .Y(_09818_));
 AO21x1_ASAP7_75t_R _29856_ (.A1(_09817_),
    .A2(_09802_),
    .B(_09818_),
    .Y(_02948_));
 BUFx6f_ASAP7_75t_R _29857_ (.A(_09389_),
    .Y(_09819_));
 AND2x2_ASAP7_75t_R _29858_ (.A(_16792_),
    .B(_09803_),
    .Y(_09820_));
 AO21x1_ASAP7_75t_R _29859_ (.A1(_09819_),
    .A2(_09802_),
    .B(_09820_),
    .Y(_02949_));
 BUFx4f_ASAP7_75t_R _29860_ (.A(_09415_),
    .Y(_09821_));
 AND2x2_ASAP7_75t_R _29861_ (.A(_16902_),
    .B(_09769_),
    .Y(_09822_));
 AO21x1_ASAP7_75t_R _29862_ (.A1(_09821_),
    .A2(_09776_),
    .B(_09822_),
    .Y(_02950_));
 NAND2x1_ASAP7_75t_R _29863_ (.A(_01191_),
    .B(_09770_),
    .Y(_09823_));
 OA21x2_ASAP7_75t_R _29864_ (.A1(_09749_),
    .A2(_09770_),
    .B(_09823_),
    .Y(_02951_));
 BUFx6f_ASAP7_75t_R _29865_ (.A(_09471_),
    .Y(_09824_));
 AND2x2_ASAP7_75t_R _29866_ (.A(_17141_),
    .B(_09769_),
    .Y(_09825_));
 AO21x1_ASAP7_75t_R _29867_ (.A1(_09824_),
    .A2(_09776_),
    .B(_09825_),
    .Y(_02952_));
 BUFx6f_ASAP7_75t_R _29868_ (.A(_09494_),
    .Y(_09826_));
 AND2x2_ASAP7_75t_R _29869_ (.A(_17272_),
    .B(_09769_),
    .Y(_09827_));
 AO21x1_ASAP7_75t_R _29870_ (.A1(_09826_),
    .A2(_09776_),
    .B(_09827_),
    .Y(_02953_));
 AND2x2_ASAP7_75t_R _29871_ (.A(_04299_),
    .B(_09769_),
    .Y(_09828_));
 AO21x1_ASAP7_75t_R _29872_ (.A1(_09753_),
    .A2(_09776_),
    .B(_09828_),
    .Y(_02954_));
 AND2x2_ASAP7_75t_R _29873_ (.A(_04429_),
    .B(_09769_),
    .Y(_09829_));
 AO21x1_ASAP7_75t_R _29874_ (.A1(_09755_),
    .A2(_09776_),
    .B(_09829_),
    .Y(_02955_));
 NAND2x1_ASAP7_75t_R _29875_ (.A(_01356_),
    .B(_09770_),
    .Y(_09830_));
 OA21x2_ASAP7_75t_R _29876_ (.A1(_09757_),
    .A2(_09770_),
    .B(_09830_),
    .Y(_02956_));
 NAND2x1_ASAP7_75t_R _29877_ (.A(_01805_),
    .B(_09764_),
    .Y(_09831_));
 OA21x2_ASAP7_75t_R _29878_ (.A1(_09107_),
    .A2(_09810_),
    .B(_09831_),
    .Y(_02957_));
 AND2x2_ASAP7_75t_R _29879_ (.A(_04653_),
    .B(_09769_),
    .Y(_09832_));
 AO21x1_ASAP7_75t_R _29880_ (.A1(net152),
    .A2(_09776_),
    .B(_09832_),
    .Y(_02958_));
 AND2x2_ASAP7_75t_R _29881_ (.A(_04847_),
    .B(_09769_),
    .Y(_09833_));
 AO21x1_ASAP7_75t_R _29882_ (.A1(net8),
    .A2(_09776_),
    .B(_09833_),
    .Y(_02959_));
 BUFx3_ASAP7_75t_R _29883_ (.A(_08338_),
    .Y(_09834_));
 AND4x2_ASAP7_75t_R _29884_ (.A(_08329_),
    .B(_09773_),
    .C(_09834_),
    .D(_08596_),
    .Y(_09835_));
 BUFx10_ASAP7_75t_R _29885_ (.A(_09835_),
    .Y(_09836_));
 INVx1_ASAP7_75t_R _29886_ (.A(_09836_),
    .Y(_09837_));
 BUFx3_ASAP7_75t_R _29887_ (.A(_08587_),
    .Y(_09838_));
 OR4x2_ASAP7_75t_R _29888_ (.A(_08593_),
    .B(_08594_),
    .C(_09838_),
    .D(_08678_),
    .Y(_09839_));
 BUFx6f_ASAP7_75t_R _29889_ (.A(_09839_),
    .Y(_09840_));
 NAND2x1_ASAP7_75t_R _29890_ (.A(_00421_),
    .B(_09840_),
    .Y(_09841_));
 OA21x2_ASAP7_75t_R _29891_ (.A1(_09650_),
    .A2(_09837_),
    .B(_09841_),
    .Y(_02960_));
 BUFx6f_ASAP7_75t_R _29892_ (.A(_09835_),
    .Y(_09842_));
 BUFx4f_ASAP7_75t_R _29893_ (.A(_09842_),
    .Y(_09843_));
 NOR2x1_ASAP7_75t_R _29894_ (.A(_00374_),
    .B(_09836_),
    .Y(_09844_));
 AO21x1_ASAP7_75t_R _29895_ (.A1(_09772_),
    .A2(_09843_),
    .B(_09844_),
    .Y(_02961_));
 NAND2x1_ASAP7_75t_R _29896_ (.A(_00485_),
    .B(_09840_),
    .Y(_09845_));
 OA21x2_ASAP7_75t_R _29897_ (.A1(_09780_),
    .A2(_09840_),
    .B(_09845_),
    .Y(_02962_));
 NOR2x1_ASAP7_75t_R _29898_ (.A(_00516_),
    .B(_09836_),
    .Y(_09846_));
 AO21x1_ASAP7_75t_R _29899_ (.A1(_09782_),
    .A2(_09843_),
    .B(_09846_),
    .Y(_02963_));
 AND2x2_ASAP7_75t_R _29900_ (.A(_14274_),
    .B(_09839_),
    .Y(_09847_));
 AO21x1_ASAP7_75t_R _29901_ (.A1(_09718_),
    .A2(_09843_),
    .B(_09847_),
    .Y(_02964_));
 NAND2x1_ASAP7_75t_R _29902_ (.A(_00578_),
    .B(_09840_),
    .Y(_09848_));
 OA21x2_ASAP7_75t_R _29903_ (.A1(_09721_),
    .A2(_09840_),
    .B(_09848_),
    .Y(_02965_));
 NOR2x1_ASAP7_75t_R _29904_ (.A(_00608_),
    .B(_09836_),
    .Y(_09849_));
 AO21x1_ASAP7_75t_R _29905_ (.A1(_09786_),
    .A2(_09843_),
    .B(_09849_),
    .Y(_02966_));
 BUFx10_ASAP7_75t_R _29906_ (.A(_09835_),
    .Y(_09850_));
 NOR2x1_ASAP7_75t_R _29907_ (.A(_00638_),
    .B(_09850_),
    .Y(_09851_));
 AO21x1_ASAP7_75t_R _29908_ (.A1(_09788_),
    .A2(_09843_),
    .B(_09851_),
    .Y(_02967_));
 NAND2x1_ASAP7_75t_R _29909_ (.A(_01804_),
    .B(_09764_),
    .Y(_09852_));
 OA21x2_ASAP7_75t_R _29910_ (.A1(_09107_),
    .A2(_09812_),
    .B(_09852_),
    .Y(_02968_));
 NAND2x1_ASAP7_75t_R _29911_ (.A(_01803_),
    .B(_09764_),
    .Y(_09853_));
 OA21x2_ASAP7_75t_R _29912_ (.A1(_09107_),
    .A2(_09676_),
    .B(_09853_),
    .Y(_02969_));
 OR3x1_ASAP7_75t_R _29913_ (.A(_09790_),
    .B(_09791_),
    .C(_09840_),
    .Y(_09854_));
 OAI21x1_ASAP7_75t_R _29914_ (.A1(_00668_),
    .A2(_09843_),
    .B(_09854_),
    .Y(_02970_));
 BUFx6f_ASAP7_75t_R _29915_ (.A(_08942_),
    .Y(_09855_));
 NOR2x1_ASAP7_75t_R _29916_ (.A(_00698_),
    .B(_09850_),
    .Y(_09856_));
 AO21x1_ASAP7_75t_R _29917_ (.A1(_09855_),
    .A2(_09843_),
    .B(_09856_),
    .Y(_02971_));
 NOR2x1_ASAP7_75t_R _29918_ (.A(_00728_),
    .B(_09850_),
    .Y(_09857_));
 AO21x1_ASAP7_75t_R _29919_ (.A1(_09108_),
    .A2(_09843_),
    .B(_09857_),
    .Y(_02972_));
 NOR2x1_ASAP7_75t_R _29920_ (.A(_00758_),
    .B(_09850_),
    .Y(_09858_));
 AO21x1_ASAP7_75t_R _29921_ (.A1(_09037_),
    .A2(_09843_),
    .B(_09858_),
    .Y(_02973_));
 NOR2x1_ASAP7_75t_R _29922_ (.A(_00454_),
    .B(_09850_),
    .Y(_09859_));
 AO21x1_ASAP7_75t_R _29923_ (.A1(_09800_),
    .A2(_09843_),
    .B(_09859_),
    .Y(_02974_));
 BUFx4f_ASAP7_75t_R _29924_ (.A(_09842_),
    .Y(_09860_));
 NOR2x1_ASAP7_75t_R _29925_ (.A(_00829_),
    .B(_09850_),
    .Y(_09861_));
 AO21x1_ASAP7_75t_R _29926_ (.A1(_09731_),
    .A2(_09860_),
    .B(_09861_),
    .Y(_02975_));
 NOR2x1_ASAP7_75t_R _29927_ (.A(_00862_),
    .B(_09850_),
    .Y(_09862_));
 AO21x1_ASAP7_75t_R _29928_ (.A1(_09745_),
    .A2(_09860_),
    .B(_09862_),
    .Y(_02976_));
 NOR2x1_ASAP7_75t_R _29929_ (.A(_00895_),
    .B(_09850_),
    .Y(_09863_));
 AO21x1_ASAP7_75t_R _29930_ (.A1(_09763_),
    .A2(_09860_),
    .B(_09863_),
    .Y(_02977_));
 AND3x1_ASAP7_75t_R _29931_ (.A(_09204_),
    .B(_09212_),
    .C(_09842_),
    .Y(_09864_));
 AO21x1_ASAP7_75t_R _29932_ (.A1(_16042_),
    .A2(_09840_),
    .B(_09864_),
    .Y(_02978_));
 NOR2x1_ASAP7_75t_R _29933_ (.A(_00961_),
    .B(_09850_),
    .Y(_09865_));
 AO21x1_ASAP7_75t_R _29934_ (.A1(_09808_),
    .A2(_09860_),
    .B(_09865_),
    .Y(_02979_));
 BUFx6f_ASAP7_75t_R _29935_ (.A(_08590_),
    .Y(_09866_));
 NAND2x1_ASAP7_75t_R _29936_ (.A(_01802_),
    .B(_09764_),
    .Y(_09867_));
 OA21x2_ASAP7_75t_R _29937_ (.A1(_09866_),
    .A2(_09815_),
    .B(_09867_),
    .Y(_02980_));
 NOR2x1_ASAP7_75t_R _29938_ (.A(_00994_),
    .B(_09850_),
    .Y(_09868_));
 AO21x1_ASAP7_75t_R _29939_ (.A1(_09810_),
    .A2(_09860_),
    .B(_09868_),
    .Y(_02981_));
 NOR2x1_ASAP7_75t_R _29940_ (.A(_01027_),
    .B(_09842_),
    .Y(_09869_));
 AO21x1_ASAP7_75t_R _29941_ (.A1(_09812_),
    .A2(_09860_),
    .B(_09869_),
    .Y(_02982_));
 NOR2x1_ASAP7_75t_R _29942_ (.A(_01060_),
    .B(_09842_),
    .Y(_09870_));
 AO21x1_ASAP7_75t_R _29943_ (.A1(_09815_),
    .A2(_09860_),
    .B(_09870_),
    .Y(_02983_));
 NOR2x1_ASAP7_75t_R _29944_ (.A(_01093_),
    .B(_09842_),
    .Y(_09871_));
 AO21x1_ASAP7_75t_R _29945_ (.A1(_09817_),
    .A2(_09860_),
    .B(_09871_),
    .Y(_02984_));
 NOR2x1_ASAP7_75t_R _29946_ (.A(_01126_),
    .B(_09842_),
    .Y(_09872_));
 AO21x1_ASAP7_75t_R _29947_ (.A1(_09819_),
    .A2(_09860_),
    .B(_09872_),
    .Y(_02985_));
 NOR2x1_ASAP7_75t_R _29948_ (.A(_01159_),
    .B(_09842_),
    .Y(_09873_));
 AO21x1_ASAP7_75t_R _29949_ (.A1(_09821_),
    .A2(_09860_),
    .B(_09873_),
    .Y(_02986_));
 NAND2x1_ASAP7_75t_R _29950_ (.A(_01192_),
    .B(_09840_),
    .Y(_09874_));
 OA21x2_ASAP7_75t_R _29951_ (.A1(_09749_),
    .A2(_09837_),
    .B(_09874_),
    .Y(_02987_));
 NOR2x1_ASAP7_75t_R _29952_ (.A(_01225_),
    .B(_09842_),
    .Y(_09875_));
 AO21x1_ASAP7_75t_R _29953_ (.A1(_09824_),
    .A2(_09836_),
    .B(_09875_),
    .Y(_02988_));
 NOR2x1_ASAP7_75t_R _29954_ (.A(_01258_),
    .B(_09842_),
    .Y(_09876_));
 AO21x1_ASAP7_75t_R _29955_ (.A1(_09826_),
    .A2(_09836_),
    .B(_09876_),
    .Y(_02989_));
 AND2x2_ASAP7_75t_R _29956_ (.A(_04296_),
    .B(_09839_),
    .Y(_09877_));
 AO21x1_ASAP7_75t_R _29957_ (.A1(_09753_),
    .A2(_09836_),
    .B(_09877_),
    .Y(_02990_));
 NAND2x1_ASAP7_75t_R _29958_ (.A(_01801_),
    .B(_09764_),
    .Y(_09878_));
 OA21x2_ASAP7_75t_R _29959_ (.A1(_09866_),
    .A2(_09817_),
    .B(_09878_),
    .Y(_02991_));
 AND2x2_ASAP7_75t_R _29960_ (.A(_04426_),
    .B(_09839_),
    .Y(_09879_));
 AO21x1_ASAP7_75t_R _29961_ (.A1(_09755_),
    .A2(_09836_),
    .B(_09879_),
    .Y(_02992_));
 NAND2x1_ASAP7_75t_R _29962_ (.A(_01357_),
    .B(_09840_),
    .Y(_09880_));
 OA21x2_ASAP7_75t_R _29963_ (.A1(net13),
    .A2(_09840_),
    .B(_09880_),
    .Y(_02993_));
 AND2x2_ASAP7_75t_R _29964_ (.A(_04650_),
    .B(_09839_),
    .Y(_09881_));
 AO21x1_ASAP7_75t_R _29965_ (.A1(_09759_),
    .A2(_09836_),
    .B(_09881_),
    .Y(_02994_));
 AND2x2_ASAP7_75t_R _29966_ (.A(_04802_),
    .B(_09839_),
    .Y(_09882_));
 AO21x1_ASAP7_75t_R _29967_ (.A1(_09761_),
    .A2(_09836_),
    .B(_09882_),
    .Y(_02995_));
 OR3x2_ASAP7_75t_R _29968_ (.A(_14153_),
    .B(_14050_),
    .C(_14232_),
    .Y(_09883_));
 OR3x4_ASAP7_75t_R _29969_ (.A(_08677_),
    .B(_09838_),
    .C(_09883_),
    .Y(_09884_));
 BUFx4f_ASAP7_75t_R _29970_ (.A(_09884_),
    .Y(_09885_));
 NAND2x1_ASAP7_75t_R _29971_ (.A(_00422_),
    .B(_09885_),
    .Y(_09886_));
 OA21x2_ASAP7_75t_R _29972_ (.A1(_09650_),
    .A2(_09885_),
    .B(_09886_),
    .Y(_02996_));
 AND3x4_ASAP7_75t_R _29973_ (.A(_14049_),
    .B(_14303_),
    .C(_14231_),
    .Y(_09887_));
 AND4x2_ASAP7_75t_R _29974_ (.A(_08027_),
    .B(_08330_),
    .C(_09834_),
    .D(_09887_),
    .Y(_09888_));
 BUFx4f_ASAP7_75t_R _29975_ (.A(_09888_),
    .Y(_09889_));
 BUFx6f_ASAP7_75t_R _29976_ (.A(_09888_),
    .Y(_09890_));
 NOR2x1_ASAP7_75t_R _29977_ (.A(_00375_),
    .B(_09890_),
    .Y(_09891_));
 AO21x1_ASAP7_75t_R _29978_ (.A1(_09772_),
    .A2(_09889_),
    .B(_09891_),
    .Y(_02997_));
 NAND2x1_ASAP7_75t_R _29979_ (.A(_00486_),
    .B(_09885_),
    .Y(_09892_));
 OA21x2_ASAP7_75t_R _29980_ (.A1(_09780_),
    .A2(_09885_),
    .B(_09892_),
    .Y(_02998_));
 NOR2x1_ASAP7_75t_R _29981_ (.A(_00517_),
    .B(_09890_),
    .Y(_09893_));
 AO21x1_ASAP7_75t_R _29982_ (.A1(_09782_),
    .A2(_09889_),
    .B(_09893_),
    .Y(_02999_));
 AND2x2_ASAP7_75t_R _29983_ (.A(_14263_),
    .B(_09884_),
    .Y(_09894_));
 AO21x1_ASAP7_75t_R _29984_ (.A1(_09718_),
    .A2(_09889_),
    .B(_09894_),
    .Y(_03000_));
 NAND2x1_ASAP7_75t_R _29985_ (.A(_00579_),
    .B(_09885_),
    .Y(_09895_));
 OA21x2_ASAP7_75t_R _29986_ (.A1(_09721_),
    .A2(_09885_),
    .B(_09895_),
    .Y(_03001_));
 NAND2x1_ASAP7_75t_R _29987_ (.A(_01800_),
    .B(_09764_),
    .Y(_09896_));
 OA21x2_ASAP7_75t_R _29988_ (.A1(_09866_),
    .A2(_09390_),
    .B(_09896_),
    .Y(_03002_));
 NOR2x1_ASAP7_75t_R _29989_ (.A(_00609_),
    .B(_09890_),
    .Y(_09897_));
 AO21x1_ASAP7_75t_R _29990_ (.A1(_09786_),
    .A2(_09889_),
    .B(_09897_),
    .Y(_03003_));
 NOR2x1_ASAP7_75t_R _29991_ (.A(_00639_),
    .B(_09890_),
    .Y(_09898_));
 AO21x1_ASAP7_75t_R _29992_ (.A1(_09788_),
    .A2(_09889_),
    .B(_09898_),
    .Y(_03004_));
 OR3x1_ASAP7_75t_R _29993_ (.A(_09790_),
    .B(_09791_),
    .C(_09884_),
    .Y(_09899_));
 OAI21x1_ASAP7_75t_R _29994_ (.A1(_00669_),
    .A2(_09889_),
    .B(_09899_),
    .Y(_03005_));
 BUFx10_ASAP7_75t_R _29995_ (.A(_09888_),
    .Y(_09900_));
 NOR2x1_ASAP7_75t_R _29996_ (.A(_00699_),
    .B(_09900_),
    .Y(_09901_));
 AO21x1_ASAP7_75t_R _29997_ (.A1(_09855_),
    .A2(_09889_),
    .B(_09901_),
    .Y(_03006_));
 NOR2x1_ASAP7_75t_R _29998_ (.A(_00729_),
    .B(_09900_),
    .Y(_09902_));
 AO21x1_ASAP7_75t_R _29999_ (.A1(_09108_),
    .A2(_09889_),
    .B(_09902_),
    .Y(_03007_));
 NAND2x1_ASAP7_75t_R _30000_ (.A(_00759_),
    .B(_09885_),
    .Y(_09903_));
 OA21x2_ASAP7_75t_R _30001_ (.A1(_09728_),
    .A2(_09885_),
    .B(_09903_),
    .Y(_03008_));
 NOR2x1_ASAP7_75t_R _30002_ (.A(_00455_),
    .B(_09900_),
    .Y(_09904_));
 AO21x1_ASAP7_75t_R _30003_ (.A1(_09800_),
    .A2(_09889_),
    .B(_09904_),
    .Y(_03009_));
 NOR2x1_ASAP7_75t_R _30004_ (.A(_00830_),
    .B(_09900_),
    .Y(_09905_));
 AO21x1_ASAP7_75t_R _30005_ (.A1(_09731_),
    .A2(_09889_),
    .B(_09905_),
    .Y(_03010_));
 BUFx4f_ASAP7_75t_R _30006_ (.A(_09888_),
    .Y(_09906_));
 NOR2x1_ASAP7_75t_R _30007_ (.A(_00863_),
    .B(_09900_),
    .Y(_09907_));
 AO21x1_ASAP7_75t_R _30008_ (.A1(_09745_),
    .A2(_09906_),
    .B(_09907_),
    .Y(_03011_));
 NOR2x1_ASAP7_75t_R _30009_ (.A(_00896_),
    .B(_09900_),
    .Y(_09908_));
 AO21x1_ASAP7_75t_R _30010_ (.A1(_09763_),
    .A2(_09906_),
    .B(_09908_),
    .Y(_03012_));
 NAND2x1_ASAP7_75t_R _30011_ (.A(_01799_),
    .B(_09764_),
    .Y(_09909_));
 OA21x2_ASAP7_75t_R _30012_ (.A1(_09866_),
    .A2(_09416_),
    .B(_09909_),
    .Y(_03013_));
 NOR2x1_ASAP7_75t_R _30013_ (.A(_00929_),
    .B(_09900_),
    .Y(_09910_));
 AO21x1_ASAP7_75t_R _30014_ (.A1(_09738_),
    .A2(_09906_),
    .B(_09910_),
    .Y(_03014_));
 NOR2x1_ASAP7_75t_R _30015_ (.A(_00962_),
    .B(_09900_),
    .Y(_09911_));
 AO21x1_ASAP7_75t_R _30016_ (.A1(_09808_),
    .A2(_09906_),
    .B(_09911_),
    .Y(_03015_));
 NOR2x1_ASAP7_75t_R _30017_ (.A(_00995_),
    .B(_09900_),
    .Y(_09912_));
 AO21x1_ASAP7_75t_R _30018_ (.A1(_09810_),
    .A2(_09906_),
    .B(_09912_),
    .Y(_03016_));
 NOR2x1_ASAP7_75t_R _30019_ (.A(_01028_),
    .B(_09900_),
    .Y(_09913_));
 AO21x1_ASAP7_75t_R _30020_ (.A1(_09812_),
    .A2(_09906_),
    .B(_09913_),
    .Y(_03017_));
 BUFx10_ASAP7_75t_R _30021_ (.A(_09888_),
    .Y(_09914_));
 NOR2x1_ASAP7_75t_R _30022_ (.A(_01061_),
    .B(_09914_),
    .Y(_09915_));
 AO21x1_ASAP7_75t_R _30023_ (.A1(_09815_),
    .A2(_09906_),
    .B(_09915_),
    .Y(_03018_));
 NOR2x1_ASAP7_75t_R _30024_ (.A(_01094_),
    .B(_09914_),
    .Y(_09916_));
 AO21x1_ASAP7_75t_R _30025_ (.A1(_09817_),
    .A2(_09906_),
    .B(_09916_),
    .Y(_03019_));
 NOR2x1_ASAP7_75t_R _30026_ (.A(_01127_),
    .B(_09914_),
    .Y(_09917_));
 AO21x1_ASAP7_75t_R _30027_ (.A1(_09819_),
    .A2(_09906_),
    .B(_09917_),
    .Y(_03020_));
 NOR2x1_ASAP7_75t_R _30028_ (.A(_01160_),
    .B(_09914_),
    .Y(_09918_));
 AO21x1_ASAP7_75t_R _30029_ (.A1(_09821_),
    .A2(_09906_),
    .B(_09918_),
    .Y(_03021_));
 NAND2x1_ASAP7_75t_R _30030_ (.A(_01193_),
    .B(_09884_),
    .Y(_09919_));
 OA21x2_ASAP7_75t_R _30031_ (.A1(_09749_),
    .A2(_09885_),
    .B(_09919_),
    .Y(_03022_));
 NOR2x1_ASAP7_75t_R _30032_ (.A(_01226_),
    .B(_09914_),
    .Y(_09920_));
 AO21x1_ASAP7_75t_R _30033_ (.A1(_09824_),
    .A2(_09890_),
    .B(_09920_),
    .Y(_03023_));
 NAND2x1_ASAP7_75t_R _30034_ (.A(_01798_),
    .B(_09764_),
    .Y(_09921_));
 OA21x2_ASAP7_75t_R _30035_ (.A1(_09866_),
    .A2(_09441_),
    .B(_09921_),
    .Y(_03024_));
 NOR2x1_ASAP7_75t_R _30036_ (.A(_01259_),
    .B(_09914_),
    .Y(_09922_));
 AO21x1_ASAP7_75t_R _30037_ (.A1(_09826_),
    .A2(_09890_),
    .B(_09922_),
    .Y(_03025_));
 NOR2x1_ASAP7_75t_R _30038_ (.A(_01292_),
    .B(_09914_),
    .Y(_09923_));
 AO21x1_ASAP7_75t_R _30039_ (.A1(_09753_),
    .A2(_09890_),
    .B(_09923_),
    .Y(_03026_));
 NOR2x1_ASAP7_75t_R _30040_ (.A(_01325_),
    .B(_09914_),
    .Y(_09924_));
 AO21x1_ASAP7_75t_R _30041_ (.A1(_09755_),
    .A2(_09890_),
    .B(_09924_),
    .Y(_03027_));
 NAND2x1_ASAP7_75t_R _30042_ (.A(_01358_),
    .B(_09884_),
    .Y(_09925_));
 OA21x2_ASAP7_75t_R _30043_ (.A1(net13),
    .A2(_09885_),
    .B(_09925_),
    .Y(_03028_));
 NOR2x1_ASAP7_75t_R _30044_ (.A(_01391_),
    .B(_09914_),
    .Y(_09926_));
 AO21x1_ASAP7_75t_R _30045_ (.A1(_09759_),
    .A2(_09890_),
    .B(_09926_),
    .Y(_03029_));
 NOR2x1_ASAP7_75t_R _30046_ (.A(_01424_),
    .B(_09914_),
    .Y(_09927_));
 AO21x1_ASAP7_75t_R _30047_ (.A1(_09761_),
    .A2(_09890_),
    .B(_09927_),
    .Y(_03030_));
 NAND2x2_ASAP7_75t_R _30048_ (.A(_08341_),
    .B(_09887_),
    .Y(_09928_));
 OR3x1_ASAP7_75t_R _30049_ (.A(_09838_),
    .B(_08589_),
    .C(_09883_),
    .Y(_09929_));
 BUFx6f_ASAP7_75t_R _30050_ (.A(_09929_),
    .Y(_09930_));
 NAND2x1_ASAP7_75t_R _30051_ (.A(_00423_),
    .B(_09930_),
    .Y(_09931_));
 OA21x2_ASAP7_75t_R _30052_ (.A1(_09650_),
    .A2(_09928_),
    .B(_09931_),
    .Y(_03031_));
 AND4x1_ASAP7_75t_R _30053_ (.A(_14726_),
    .B(_08330_),
    .C(_08338_),
    .D(_09887_),
    .Y(_09932_));
 BUFx10_ASAP7_75t_R _30054_ (.A(_09932_),
    .Y(_09933_));
 BUFx4f_ASAP7_75t_R _30055_ (.A(_09933_),
    .Y(_09934_));
 BUFx10_ASAP7_75t_R _30056_ (.A(_09933_),
    .Y(_09935_));
 NOR2x1_ASAP7_75t_R _30057_ (.A(_00376_),
    .B(_09935_),
    .Y(_09936_));
 AO21x1_ASAP7_75t_R _30058_ (.A1(_09772_),
    .A2(_09934_),
    .B(_09936_),
    .Y(_03032_));
 NAND2x1_ASAP7_75t_R _30059_ (.A(_00487_),
    .B(_09930_),
    .Y(_09937_));
 OA21x2_ASAP7_75t_R _30060_ (.A1(_09780_),
    .A2(_09930_),
    .B(_09937_),
    .Y(_03033_));
 NOR2x1_ASAP7_75t_R _30061_ (.A(_00518_),
    .B(_09935_),
    .Y(_09938_));
 AO21x1_ASAP7_75t_R _30062_ (.A1(_09782_),
    .A2(_09934_),
    .B(_09938_),
    .Y(_03034_));
 NAND2x1_ASAP7_75t_R _30063_ (.A(_01797_),
    .B(_09106_),
    .Y(_09939_));
 OA21x2_ASAP7_75t_R _30064_ (.A1(_09866_),
    .A2(_09824_),
    .B(_09939_),
    .Y(_03035_));
 NOR2x1_ASAP7_75t_R _30065_ (.A(_00548_),
    .B(_09935_),
    .Y(_09940_));
 AO21x1_ASAP7_75t_R _30066_ (.A1(_09718_),
    .A2(_09934_),
    .B(_09940_),
    .Y(_03036_));
 NAND2x1_ASAP7_75t_R _30067_ (.A(_00580_),
    .B(_09930_),
    .Y(_09941_));
 OA21x2_ASAP7_75t_R _30068_ (.A1(_09721_),
    .A2(_09930_),
    .B(_09941_),
    .Y(_03037_));
 NOR2x1_ASAP7_75t_R _30069_ (.A(_00610_),
    .B(_09935_),
    .Y(_09942_));
 AO21x1_ASAP7_75t_R _30070_ (.A1(_09786_),
    .A2(_09934_),
    .B(_09942_),
    .Y(_03038_));
 BUFx10_ASAP7_75t_R _30071_ (.A(_09933_),
    .Y(_09943_));
 NOR2x1_ASAP7_75t_R _30072_ (.A(_00640_),
    .B(_09943_),
    .Y(_09944_));
 AO21x1_ASAP7_75t_R _30073_ (.A1(_09788_),
    .A2(_09934_),
    .B(_09944_),
    .Y(_03039_));
 OR2x2_ASAP7_75t_R _30074_ (.A(_00670_),
    .B(_09933_),
    .Y(_09945_));
 OAI21x1_ASAP7_75t_R _30075_ (.A1(_08898_),
    .A2(_09928_),
    .B(_09945_),
    .Y(_03040_));
 NOR2x1_ASAP7_75t_R _30076_ (.A(_00700_),
    .B(_09943_),
    .Y(_09946_));
 AO21x1_ASAP7_75t_R _30077_ (.A1(_09855_),
    .A2(_09934_),
    .B(_09946_),
    .Y(_03041_));
 NOR2x1_ASAP7_75t_R _30078_ (.A(_00730_),
    .B(_09943_),
    .Y(_09947_));
 AO21x1_ASAP7_75t_R _30079_ (.A1(_09108_),
    .A2(_09934_),
    .B(_09947_),
    .Y(_03042_));
 NOR2x1_ASAP7_75t_R _30080_ (.A(_00760_),
    .B(_09943_),
    .Y(_09948_));
 AO21x1_ASAP7_75t_R _30081_ (.A1(_09037_),
    .A2(_09934_),
    .B(_09948_),
    .Y(_03043_));
 NOR2x1_ASAP7_75t_R _30082_ (.A(_00456_),
    .B(_09943_),
    .Y(_09949_));
 AO21x1_ASAP7_75t_R _30083_ (.A1(_09800_),
    .A2(_09934_),
    .B(_09949_),
    .Y(_03044_));
 NOR2x1_ASAP7_75t_R _30084_ (.A(_00831_),
    .B(_09943_),
    .Y(_09950_));
 AO21x1_ASAP7_75t_R _30085_ (.A1(_09731_),
    .A2(_09934_),
    .B(_09950_),
    .Y(_03045_));
 NAND2x1_ASAP7_75t_R _30086_ (.A(_01796_),
    .B(_09106_),
    .Y(_09951_));
 OA21x2_ASAP7_75t_R _30087_ (.A1(_09866_),
    .A2(_09826_),
    .B(_09951_),
    .Y(_03046_));
 BUFx4f_ASAP7_75t_R _30088_ (.A(_09933_),
    .Y(_09952_));
 NOR2x1_ASAP7_75t_R _30089_ (.A(_00864_),
    .B(_09943_),
    .Y(_09953_));
 AO21x1_ASAP7_75t_R _30090_ (.A1(_09745_),
    .A2(_09952_),
    .B(_09953_),
    .Y(_03047_));
 NOR2x1_ASAP7_75t_R _30091_ (.A(_00897_),
    .B(_09943_),
    .Y(_09954_));
 AO21x1_ASAP7_75t_R _30092_ (.A1(_09763_),
    .A2(_09952_),
    .B(_09954_),
    .Y(_03048_));
 NOR2x1_ASAP7_75t_R _30093_ (.A(_00930_),
    .B(_09943_),
    .Y(_09955_));
 AO21x1_ASAP7_75t_R _30094_ (.A1(_09738_),
    .A2(_09952_),
    .B(_09955_),
    .Y(_03049_));
 NOR2x1_ASAP7_75t_R _30095_ (.A(_00963_),
    .B(_09943_),
    .Y(_09956_));
 AO21x1_ASAP7_75t_R _30096_ (.A1(_09808_),
    .A2(_09952_),
    .B(_09956_),
    .Y(_03050_));
 BUFx6f_ASAP7_75t_R _30097_ (.A(_09933_),
    .Y(_09957_));
 NOR2x1_ASAP7_75t_R _30098_ (.A(_00996_),
    .B(_09957_),
    .Y(_09958_));
 AO21x1_ASAP7_75t_R _30099_ (.A1(_09810_),
    .A2(_09952_),
    .B(_09958_),
    .Y(_03051_));
 NOR2x1_ASAP7_75t_R _30100_ (.A(_01029_),
    .B(_09957_),
    .Y(_09959_));
 AO21x1_ASAP7_75t_R _30101_ (.A1(_09812_),
    .A2(_09952_),
    .B(_09959_),
    .Y(_03052_));
 NOR2x1_ASAP7_75t_R _30102_ (.A(_01062_),
    .B(_09957_),
    .Y(_09960_));
 AO21x1_ASAP7_75t_R _30103_ (.A1(_09815_),
    .A2(_09952_),
    .B(_09960_),
    .Y(_03053_));
 NOR2x1_ASAP7_75t_R _30104_ (.A(_01095_),
    .B(_09957_),
    .Y(_09961_));
 AO21x1_ASAP7_75t_R _30105_ (.A1(_09817_),
    .A2(_09952_),
    .B(_09961_),
    .Y(_03054_));
 NOR2x1_ASAP7_75t_R _30106_ (.A(_01128_),
    .B(_09957_),
    .Y(_09962_));
 AO21x1_ASAP7_75t_R _30107_ (.A1(_09819_),
    .A2(_09952_),
    .B(_09962_),
    .Y(_03055_));
 NOR2x1_ASAP7_75t_R _30108_ (.A(_01161_),
    .B(_09957_),
    .Y(_09963_));
 AO21x1_ASAP7_75t_R _30109_ (.A1(_09821_),
    .A2(_09952_),
    .B(_09963_),
    .Y(_03056_));
 NOR2x1_ASAP7_75t_R _30110_ (.A(_01795_),
    .B(_09796_),
    .Y(_09964_));
 AO21x1_ASAP7_75t_R _30111_ (.A1(_09794_),
    .A2(_09512_),
    .B(_09964_),
    .Y(_03057_));
 NAND2x1_ASAP7_75t_R _30112_ (.A(_01194_),
    .B(_09930_),
    .Y(_09965_));
 OA21x2_ASAP7_75t_R _30113_ (.A1(_09749_),
    .A2(_09930_),
    .B(_09965_),
    .Y(_03058_));
 NOR2x1_ASAP7_75t_R _30114_ (.A(_01227_),
    .B(_09957_),
    .Y(_09966_));
 AO21x1_ASAP7_75t_R _30115_ (.A1(_09824_),
    .A2(_09935_),
    .B(_09966_),
    .Y(_03059_));
 NOR2x1_ASAP7_75t_R _30116_ (.A(_01260_),
    .B(_09957_),
    .Y(_09967_));
 AO21x1_ASAP7_75t_R _30117_ (.A1(_09826_),
    .A2(_09935_),
    .B(_09967_),
    .Y(_03060_));
 NOR2x1_ASAP7_75t_R _30118_ (.A(_01293_),
    .B(_09957_),
    .Y(_09968_));
 AO21x1_ASAP7_75t_R _30119_ (.A1(_09753_),
    .A2(_09935_),
    .B(_09968_),
    .Y(_03061_));
 NOR2x1_ASAP7_75t_R _30120_ (.A(_01326_),
    .B(_09957_),
    .Y(_09969_));
 AO21x1_ASAP7_75t_R _30121_ (.A1(_09755_),
    .A2(_09935_),
    .B(_09969_),
    .Y(_03062_));
 NAND2x1_ASAP7_75t_R _30122_ (.A(_01359_),
    .B(_09930_),
    .Y(_09970_));
 OA21x2_ASAP7_75t_R _30123_ (.A1(net13),
    .A2(_09930_),
    .B(_09970_),
    .Y(_03063_));
 NOR2x1_ASAP7_75t_R _30124_ (.A(_01392_),
    .B(_09933_),
    .Y(_09971_));
 AO21x1_ASAP7_75t_R _30125_ (.A1(_09759_),
    .A2(_09935_),
    .B(_09971_),
    .Y(_03064_));
 NOR2x1_ASAP7_75t_R _30126_ (.A(_01425_),
    .B(_09933_),
    .Y(_09972_));
 AO21x1_ASAP7_75t_R _30127_ (.A1(_09761_),
    .A2(_09935_),
    .B(_09972_),
    .Y(_03065_));
 OR3x1_ASAP7_75t_R _30128_ (.A(_09766_),
    .B(_09767_),
    .C(_09883_),
    .Y(_09973_));
 BUFx10_ASAP7_75t_R _30129_ (.A(_09973_),
    .Y(_09974_));
 BUFx6f_ASAP7_75t_R _30130_ (.A(_09974_),
    .Y(_09975_));
 NAND2x1_ASAP7_75t_R _30131_ (.A(_00424_),
    .B(_09975_),
    .Y(_09976_));
 OA21x2_ASAP7_75t_R _30132_ (.A1(_09650_),
    .A2(_09975_),
    .B(_09976_),
    .Y(_03066_));
 AND3x1_ASAP7_75t_R _30133_ (.A(_08339_),
    .B(_09774_),
    .C(_09887_),
    .Y(_09977_));
 BUFx6f_ASAP7_75t_R _30134_ (.A(_09977_),
    .Y(_09978_));
 BUFx6f_ASAP7_75t_R _30135_ (.A(_09978_),
    .Y(_09979_));
 BUFx4f_ASAP7_75t_R _30136_ (.A(_09974_),
    .Y(_09980_));
 AND2x2_ASAP7_75t_R _30137_ (.A(_13505_),
    .B(_09980_),
    .Y(_09981_));
 AO21x1_ASAP7_75t_R _30138_ (.A1(_09772_),
    .A2(_09979_),
    .B(_09981_),
    .Y(_03067_));
 NOR2x1_ASAP7_75t_R _30139_ (.A(_01794_),
    .B(_09796_),
    .Y(_09982_));
 AO21x1_ASAP7_75t_R _30140_ (.A1(_09794_),
    .A2(net95),
    .B(_09982_),
    .Y(_03068_));
 NAND2x1_ASAP7_75t_R _30141_ (.A(_00488_),
    .B(_09975_),
    .Y(_09983_));
 OA21x2_ASAP7_75t_R _30142_ (.A1(_09780_),
    .A2(_09975_),
    .B(_09983_),
    .Y(_03069_));
 AND2x2_ASAP7_75t_R _30143_ (.A(_14933_),
    .B(_09980_),
    .Y(_09984_));
 AO21x1_ASAP7_75t_R _30144_ (.A1(_09782_),
    .A2(_09979_),
    .B(_09984_),
    .Y(_03070_));
 AND2x2_ASAP7_75t_R _30145_ (.A(_14997_),
    .B(_09980_),
    .Y(_09985_));
 AO21x1_ASAP7_75t_R _30146_ (.A1(_09718_),
    .A2(_09979_),
    .B(_09985_),
    .Y(_03071_));
 NAND2x1_ASAP7_75t_R _30147_ (.A(_00581_),
    .B(_09975_),
    .Y(_09986_));
 OA21x2_ASAP7_75t_R _30148_ (.A1(_09721_),
    .A2(_09975_),
    .B(_09986_),
    .Y(_03072_));
 AND2x2_ASAP7_75t_R _30149_ (.A(_15132_),
    .B(_09980_),
    .Y(_09987_));
 AO21x1_ASAP7_75t_R _30150_ (.A1(_09786_),
    .A2(_09979_),
    .B(_09987_),
    .Y(_03073_));
 AND2x2_ASAP7_75t_R _30151_ (.A(_14458_),
    .B(_09980_),
    .Y(_09988_));
 AO21x1_ASAP7_75t_R _30152_ (.A1(_09788_),
    .A2(_09979_),
    .B(_09988_),
    .Y(_03074_));
 OR3x1_ASAP7_75t_R _30153_ (.A(_09790_),
    .B(_09791_),
    .C(_09980_),
    .Y(_09989_));
 OAI21x1_ASAP7_75t_R _30154_ (.A1(_00671_),
    .A2(_09979_),
    .B(_09989_),
    .Y(_03075_));
 AND2x2_ASAP7_75t_R _30155_ (.A(_15346_),
    .B(_09980_),
    .Y(_09990_));
 AO21x1_ASAP7_75t_R _30156_ (.A1(_09855_),
    .A2(_09979_),
    .B(_09990_),
    .Y(_03076_));
 AND2x2_ASAP7_75t_R _30157_ (.A(_14616_),
    .B(_09980_),
    .Y(_09991_));
 AO21x1_ASAP7_75t_R _30158_ (.A1(_09108_),
    .A2(_09979_),
    .B(_09991_),
    .Y(_03077_));
 AND2x2_ASAP7_75t_R _30159_ (.A(_14685_),
    .B(_09980_),
    .Y(_09992_));
 AO21x1_ASAP7_75t_R _30160_ (.A1(_09037_),
    .A2(_09979_),
    .B(_09992_),
    .Y(_03078_));
 NAND2x1_ASAP7_75t_R _30161_ (.A(_01793_),
    .B(_09106_),
    .Y(_09993_));
 OA21x2_ASAP7_75t_R _30162_ (.A1(_09866_),
    .A2(_09580_),
    .B(_09993_),
    .Y(_03079_));
 NAND2x1_ASAP7_75t_R _30163_ (.A(_01792_),
    .B(_09106_),
    .Y(_09994_));
 OA21x2_ASAP7_75t_R _30164_ (.A1(_09866_),
    .A2(_09696_),
    .B(_09994_),
    .Y(_03080_));
 AND2x2_ASAP7_75t_R _30165_ (.A(_15521_),
    .B(_09980_),
    .Y(_09995_));
 AO21x1_ASAP7_75t_R _30166_ (.A1(_09800_),
    .A2(_09979_),
    .B(_09995_),
    .Y(_03081_));
 BUFx4f_ASAP7_75t_R _30167_ (.A(_09978_),
    .Y(_09996_));
 BUFx4f_ASAP7_75t_R _30168_ (.A(_09974_),
    .Y(_09997_));
 AND2x2_ASAP7_75t_R _30169_ (.A(_15601_),
    .B(_09997_),
    .Y(_09998_));
 AO21x1_ASAP7_75t_R _30170_ (.A1(_09731_),
    .A2(_09996_),
    .B(_09998_),
    .Y(_03082_));
 AND2x2_ASAP7_75t_R _30171_ (.A(_15760_),
    .B(_09997_),
    .Y(_09999_));
 AO21x1_ASAP7_75t_R _30172_ (.A1(_09745_),
    .A2(_09996_),
    .B(_09999_),
    .Y(_03083_));
 AND2x2_ASAP7_75t_R _30173_ (.A(_15881_),
    .B(_09997_),
    .Y(_10000_));
 AO21x1_ASAP7_75t_R _30174_ (.A1(_09763_),
    .A2(_09996_),
    .B(_10000_),
    .Y(_03084_));
 AND2x2_ASAP7_75t_R _30175_ (.A(_16037_),
    .B(_09997_),
    .Y(_10001_));
 AO21x1_ASAP7_75t_R _30176_ (.A1(_09738_),
    .A2(_09996_),
    .B(_10001_),
    .Y(_03085_));
 AND2x2_ASAP7_75t_R _30177_ (.A(_16155_),
    .B(_09997_),
    .Y(_10002_));
 AO21x1_ASAP7_75t_R _30178_ (.A1(_09808_),
    .A2(_09996_),
    .B(_10002_),
    .Y(_03086_));
 AND2x2_ASAP7_75t_R _30179_ (.A(_16297_),
    .B(_09997_),
    .Y(_10003_));
 AO21x1_ASAP7_75t_R _30180_ (.A1(_09810_),
    .A2(_09996_),
    .B(_10003_),
    .Y(_03087_));
 AND2x2_ASAP7_75t_R _30181_ (.A(_16412_),
    .B(_09997_),
    .Y(_10004_));
 AO21x1_ASAP7_75t_R _30182_ (.A1(_09812_),
    .A2(_09996_),
    .B(_10004_),
    .Y(_03088_));
 AND2x2_ASAP7_75t_R _30183_ (.A(_16539_),
    .B(_09997_),
    .Y(_10005_));
 AO21x1_ASAP7_75t_R _30184_ (.A1(_09815_),
    .A2(_09996_),
    .B(_10005_),
    .Y(_03089_));
 AND2x2_ASAP7_75t_R _30185_ (.A(_16654_),
    .B(_09997_),
    .Y(_10006_));
 AO21x1_ASAP7_75t_R _30186_ (.A1(_09817_),
    .A2(_09996_),
    .B(_10006_),
    .Y(_03090_));
 NOR2x1_ASAP7_75t_R _30187_ (.A(_01791_),
    .B(_09796_),
    .Y(_10007_));
 AO21x1_ASAP7_75t_R _30188_ (.A1(_09794_),
    .A2(_09621_),
    .B(_10007_),
    .Y(_03091_));
 AND2x2_ASAP7_75t_R _30189_ (.A(_16784_),
    .B(_09997_),
    .Y(_10008_));
 AO21x1_ASAP7_75t_R _30190_ (.A1(_09819_),
    .A2(_09996_),
    .B(_10008_),
    .Y(_03092_));
 AND2x2_ASAP7_75t_R _30191_ (.A(_16894_),
    .B(_09974_),
    .Y(_10009_));
 AO21x1_ASAP7_75t_R _30192_ (.A1(_09821_),
    .A2(_09978_),
    .B(_10009_),
    .Y(_03093_));
 NAND2x1_ASAP7_75t_R _30193_ (.A(_01195_),
    .B(_09975_),
    .Y(_10010_));
 OA21x2_ASAP7_75t_R _30194_ (.A1(_09749_),
    .A2(_09975_),
    .B(_10010_),
    .Y(_03094_));
 AND2x2_ASAP7_75t_R _30195_ (.A(_17133_),
    .B(_09974_),
    .Y(_10011_));
 AO21x1_ASAP7_75t_R _30196_ (.A1(_09824_),
    .A2(_09978_),
    .B(_10011_),
    .Y(_03095_));
 AND2x2_ASAP7_75t_R _30197_ (.A(_17264_),
    .B(_09974_),
    .Y(_10012_));
 AO21x1_ASAP7_75t_R _30198_ (.A1(_09826_),
    .A2(_09978_),
    .B(_10012_),
    .Y(_03096_));
 AND2x2_ASAP7_75t_R _30199_ (.A(_04291_),
    .B(_09974_),
    .Y(_10013_));
 AO21x1_ASAP7_75t_R _30200_ (.A1(_09753_),
    .A2(_09978_),
    .B(_10013_),
    .Y(_03097_));
 AND2x2_ASAP7_75t_R _30201_ (.A(_04421_),
    .B(_09974_),
    .Y(_10014_));
 AO21x1_ASAP7_75t_R _30202_ (.A1(_09755_),
    .A2(_09978_),
    .B(_10014_),
    .Y(_03098_));
 NAND2x1_ASAP7_75t_R _30203_ (.A(_01360_),
    .B(_09975_),
    .Y(_10015_));
 OA21x2_ASAP7_75t_R _30204_ (.A1(_09757_),
    .A2(_09975_),
    .B(_10015_),
    .Y(_03099_));
 AND2x2_ASAP7_75t_R _30205_ (.A(_04645_),
    .B(_09974_),
    .Y(_10016_));
 AO21x1_ASAP7_75t_R _30206_ (.A1(net152),
    .A2(_09978_),
    .B(_10016_),
    .Y(_03100_));
 AND2x2_ASAP7_75t_R _30207_ (.A(_04764_),
    .B(_09974_),
    .Y(_10017_));
 AO21x1_ASAP7_75t_R _30208_ (.A1(net8),
    .A2(_09978_),
    .B(_10017_),
    .Y(_03101_));
 NOR2x1_ASAP7_75t_R _30209_ (.A(_01790_),
    .B(_09796_),
    .Y(_10018_));
 AO21x1_ASAP7_75t_R _30210_ (.A1(_09794_),
    .A2(_09647_),
    .B(_10018_),
    .Y(_03102_));
 AND4x2_ASAP7_75t_R _30211_ (.A(_08329_),
    .B(_09773_),
    .C(_09834_),
    .D(_09887_),
    .Y(_10019_));
 BUFx12f_ASAP7_75t_R _30212_ (.A(_10019_),
    .Y(_10020_));
 INVx2_ASAP7_75t_R _30213_ (.A(_10020_),
    .Y(_10021_));
 OR4x2_ASAP7_75t_R _30214_ (.A(_08593_),
    .B(_08594_),
    .C(_09838_),
    .D(_09883_),
    .Y(_10022_));
 BUFx6f_ASAP7_75t_R _30215_ (.A(_10022_),
    .Y(_10023_));
 NAND2x1_ASAP7_75t_R _30216_ (.A(_00425_),
    .B(_10023_),
    .Y(_10024_));
 OA21x2_ASAP7_75t_R _30217_ (.A1(_09650_),
    .A2(_10021_),
    .B(_10024_),
    .Y(_03103_));
 BUFx4f_ASAP7_75t_R _30218_ (.A(_10020_),
    .Y(_10025_));
 BUFx12_ASAP7_75t_R _30219_ (.A(_10019_),
    .Y(_10026_));
 NOR2x1_ASAP7_75t_R _30220_ (.A(_00378_),
    .B(_10026_),
    .Y(_10027_));
 AO21x1_ASAP7_75t_R _30221_ (.A1(_09772_),
    .A2(_10025_),
    .B(_10027_),
    .Y(_03104_));
 NAND2x1_ASAP7_75t_R _30222_ (.A(_00489_),
    .B(_10023_),
    .Y(_10028_));
 OA21x2_ASAP7_75t_R _30223_ (.A1(_09780_),
    .A2(_10023_),
    .B(_10028_),
    .Y(_03105_));
 NOR2x1_ASAP7_75t_R _30224_ (.A(_00520_),
    .B(_10026_),
    .Y(_10029_));
 AO21x1_ASAP7_75t_R _30225_ (.A1(_09782_),
    .A2(_10025_),
    .B(_10029_),
    .Y(_03106_));
 AND2x2_ASAP7_75t_R _30226_ (.A(_14266_),
    .B(_10022_),
    .Y(_10030_));
 AO21x1_ASAP7_75t_R _30227_ (.A1(_09718_),
    .A2(_10025_),
    .B(_10030_),
    .Y(_03107_));
 NAND2x1_ASAP7_75t_R _30228_ (.A(_00582_),
    .B(_10023_),
    .Y(_10031_));
 OA21x2_ASAP7_75t_R _30229_ (.A1(_09721_),
    .A2(_10023_),
    .B(_10031_),
    .Y(_03108_));
 NOR2x1_ASAP7_75t_R _30230_ (.A(_00612_),
    .B(_10026_),
    .Y(_10032_));
 AO21x1_ASAP7_75t_R _30231_ (.A1(_09786_),
    .A2(_10025_),
    .B(_10032_),
    .Y(_03109_));
 NOR2x1_ASAP7_75t_R _30232_ (.A(_00642_),
    .B(_10026_),
    .Y(_10033_));
 AO21x1_ASAP7_75t_R _30233_ (.A1(_09788_),
    .A2(_10025_),
    .B(_10033_),
    .Y(_03110_));
 NAND2x1_ASAP7_75t_R _30234_ (.A(_15279_),
    .B(_10023_),
    .Y(_10034_));
 OAI21x1_ASAP7_75t_R _30235_ (.A1(_08898_),
    .A2(_10021_),
    .B(_10034_),
    .Y(_03111_));
 NOR2x1_ASAP7_75t_R _30236_ (.A(_00702_),
    .B(_10026_),
    .Y(_10035_));
 AO21x1_ASAP7_75t_R _30237_ (.A1(_09855_),
    .A2(_10025_),
    .B(_10035_),
    .Y(_03112_));
 OR3x1_ASAP7_75t_R _30238_ (.A(_08586_),
    .B(_08588_),
    .C(_09767_),
    .Y(_10036_));
 BUFx4f_ASAP7_75t_R _30239_ (.A(_10036_),
    .Y(_10037_));
 BUFx4f_ASAP7_75t_R _30240_ (.A(_10037_),
    .Y(_10038_));
 BUFx6f_ASAP7_75t_R _30241_ (.A(_10037_),
    .Y(_10039_));
 NAND2x1_ASAP7_75t_R _30242_ (.A(_00416_),
    .B(_10039_),
    .Y(_10040_));
 OA21x2_ASAP7_75t_R _30243_ (.A1(_09650_),
    .A2(_10038_),
    .B(_10040_),
    .Y(_03113_));
 BUFx10_ASAP7_75t_R _30244_ (.A(_10020_),
    .Y(_10041_));
 NOR2x1_ASAP7_75t_R _30245_ (.A(_00732_),
    .B(_10041_),
    .Y(_10042_));
 AO21x1_ASAP7_75t_R _30246_ (.A1(_09108_),
    .A2(_10025_),
    .B(_10042_),
    .Y(_03114_));
 NOR2x1_ASAP7_75t_R _30247_ (.A(_00762_),
    .B(_10041_),
    .Y(_10043_));
 AO21x1_ASAP7_75t_R _30248_ (.A1(_09037_),
    .A2(_10025_),
    .B(_10043_),
    .Y(_03115_));
 NOR2x1_ASAP7_75t_R _30249_ (.A(_00458_),
    .B(_10041_),
    .Y(_10044_));
 AO21x1_ASAP7_75t_R _30250_ (.A1(_09800_),
    .A2(_10025_),
    .B(_10044_),
    .Y(_03116_));
 NOR2x1_ASAP7_75t_R _30251_ (.A(_00833_),
    .B(_10041_),
    .Y(_10045_));
 AO21x1_ASAP7_75t_R _30252_ (.A1(_09731_),
    .A2(_10025_),
    .B(_10045_),
    .Y(_03117_));
 BUFx4f_ASAP7_75t_R _30253_ (.A(_10020_),
    .Y(_10046_));
 NOR2x1_ASAP7_75t_R _30254_ (.A(_00866_),
    .B(_10041_),
    .Y(_10047_));
 AO21x1_ASAP7_75t_R _30255_ (.A1(_09745_),
    .A2(_10046_),
    .B(_10047_),
    .Y(_03118_));
 NOR2x1_ASAP7_75t_R _30256_ (.A(_00899_),
    .B(_10041_),
    .Y(_10048_));
 AO21x1_ASAP7_75t_R _30257_ (.A1(_09763_),
    .A2(_10046_),
    .B(_10048_),
    .Y(_03119_));
 AND2x2_ASAP7_75t_R _30258_ (.A(_16033_),
    .B(_10022_),
    .Y(_10049_));
 AO21x1_ASAP7_75t_R _30259_ (.A1(_09738_),
    .A2(_10046_),
    .B(_10049_),
    .Y(_03120_));
 NOR2x1_ASAP7_75t_R _30260_ (.A(_00965_),
    .B(_10041_),
    .Y(_10050_));
 AO21x1_ASAP7_75t_R _30261_ (.A1(_09808_),
    .A2(_10046_),
    .B(_10050_),
    .Y(_03121_));
 NOR2x1_ASAP7_75t_R _30262_ (.A(_00998_),
    .B(_10041_),
    .Y(_10051_));
 AO21x1_ASAP7_75t_R _30263_ (.A1(_09810_),
    .A2(_10046_),
    .B(_10051_),
    .Y(_03122_));
 NOR2x1_ASAP7_75t_R _30264_ (.A(_01031_),
    .B(_10041_),
    .Y(_10052_));
 AO21x1_ASAP7_75t_R _30265_ (.A1(_09812_),
    .A2(_10046_),
    .B(_10052_),
    .Y(_03123_));
 NAND2x1_ASAP7_75t_R _30266_ (.A(_00369_),
    .B(_10039_),
    .Y(_10053_));
 OA21x2_ASAP7_75t_R _30267_ (.A1(_09676_),
    .A2(_10038_),
    .B(_10053_),
    .Y(_03124_));
 NOR2x1_ASAP7_75t_R _30268_ (.A(_01064_),
    .B(_10041_),
    .Y(_10054_));
 AO21x1_ASAP7_75t_R _30269_ (.A1(_09815_),
    .A2(_10046_),
    .B(_10054_),
    .Y(_03125_));
 NOR2x1_ASAP7_75t_R _30270_ (.A(_01097_),
    .B(_10020_),
    .Y(_10055_));
 AO21x1_ASAP7_75t_R _30271_ (.A1(_09817_),
    .A2(_10046_),
    .B(_10055_),
    .Y(_03126_));
 NOR2x1_ASAP7_75t_R _30272_ (.A(_01130_),
    .B(_10020_),
    .Y(_10056_));
 AO21x1_ASAP7_75t_R _30273_ (.A1(_09819_),
    .A2(_10046_),
    .B(_10056_),
    .Y(_03127_));
 NOR2x1_ASAP7_75t_R _30274_ (.A(_01163_),
    .B(_10020_),
    .Y(_10057_));
 AO21x1_ASAP7_75t_R _30275_ (.A1(_09821_),
    .A2(_10046_),
    .B(_10057_),
    .Y(_03128_));
 NAND2x1_ASAP7_75t_R _30276_ (.A(_01196_),
    .B(_10023_),
    .Y(_10058_));
 OA21x2_ASAP7_75t_R _30277_ (.A1(_09749_),
    .A2(_10023_),
    .B(_10058_),
    .Y(_03129_));
 NOR2x1_ASAP7_75t_R _30278_ (.A(_01229_),
    .B(_10020_),
    .Y(_10059_));
 AO21x1_ASAP7_75t_R _30279_ (.A1(_09824_),
    .A2(_10026_),
    .B(_10059_),
    .Y(_03130_));
 NOR2x1_ASAP7_75t_R _30280_ (.A(_01262_),
    .B(_10020_),
    .Y(_10060_));
 AO21x1_ASAP7_75t_R _30281_ (.A1(_09826_),
    .A2(_10026_),
    .B(_10060_),
    .Y(_03131_));
 AND3x2_ASAP7_75t_R _30282_ (.A(_09508_),
    .B(_09511_),
    .C(_10020_),
    .Y(_10061_));
 AO21x1_ASAP7_75t_R _30283_ (.A1(_04288_),
    .A2(_10021_),
    .B(_10061_),
    .Y(_03132_));
 AND2x2_ASAP7_75t_R _30284_ (.A(_04418_),
    .B(_10022_),
    .Y(_10062_));
 AO21x1_ASAP7_75t_R _30285_ (.A1(_09755_),
    .A2(_10026_),
    .B(_10062_),
    .Y(_03133_));
 NAND2x1_ASAP7_75t_R _30286_ (.A(_01361_),
    .B(_10023_),
    .Y(_10063_));
 OA21x2_ASAP7_75t_R _30287_ (.A1(_09757_),
    .A2(_10023_),
    .B(_10063_),
    .Y(_03134_));
 NAND2x1_ASAP7_75t_R _30288_ (.A(_00480_),
    .B(_10039_),
    .Y(_10064_));
 OA21x2_ASAP7_75t_R _30289_ (.A1(_09780_),
    .A2(_10038_),
    .B(_10064_),
    .Y(_03135_));
 AND2x2_ASAP7_75t_R _30290_ (.A(_04642_),
    .B(_10022_),
    .Y(_10065_));
 AO21x1_ASAP7_75t_R _30291_ (.A1(_09759_),
    .A2(_10026_),
    .B(_10065_),
    .Y(_03136_));
 AND2x2_ASAP7_75t_R _30292_ (.A(_04761_),
    .B(_10022_),
    .Y(_10066_));
 AO21x1_ASAP7_75t_R _30293_ (.A1(_09761_),
    .A2(_10026_),
    .B(_10066_),
    .Y(_03137_));
 OR3x2_ASAP7_75t_R _30294_ (.A(_14049_),
    .B(_14050_),
    .C(_14232_),
    .Y(_10067_));
 OR3x4_ASAP7_75t_R _30295_ (.A(_08677_),
    .B(_09766_),
    .C(_10067_),
    .Y(_10068_));
 BUFx6f_ASAP7_75t_R _30296_ (.A(_10068_),
    .Y(_10069_));
 BUFx6f_ASAP7_75t_R _30297_ (.A(_10068_),
    .Y(_10070_));
 NAND2x1_ASAP7_75t_R _30298_ (.A(_00426_),
    .B(_10070_),
    .Y(_10071_));
 OA21x2_ASAP7_75t_R _30299_ (.A1(_09650_),
    .A2(_10069_),
    .B(_10071_),
    .Y(_03138_));
 NAND2x1_ASAP7_75t_R _30300_ (.A(_00379_),
    .B(_10070_),
    .Y(_10072_));
 OA21x2_ASAP7_75t_R _30301_ (.A1(_09676_),
    .A2(_10069_),
    .B(_10072_),
    .Y(_03139_));
 NAND2x1_ASAP7_75t_R _30302_ (.A(_00490_),
    .B(_10070_),
    .Y(_10073_));
 OA21x2_ASAP7_75t_R _30303_ (.A1(_09780_),
    .A2(_10069_),
    .B(_10073_),
    .Y(_03140_));
 NAND2x1_ASAP7_75t_R _30304_ (.A(_00521_),
    .B(_10070_),
    .Y(_10074_));
 OA21x2_ASAP7_75t_R _30305_ (.A1(_09716_),
    .A2(_10069_),
    .B(_10074_),
    .Y(_03141_));
 AND3x4_ASAP7_75t_R _30306_ (.A(_14153_),
    .B(_14303_),
    .C(_14231_),
    .Y(_10075_));
 AND4x2_ASAP7_75t_R _30307_ (.A(_08027_),
    .B(_08330_),
    .C(_09834_),
    .D(_10075_),
    .Y(_10076_));
 BUFx4f_ASAP7_75t_R _30308_ (.A(_10076_),
    .Y(_10077_));
 BUFx6f_ASAP7_75t_R _30309_ (.A(_10077_),
    .Y(_10078_));
 BUFx10_ASAP7_75t_R _30310_ (.A(_10068_),
    .Y(_10079_));
 AND2x2_ASAP7_75t_R _30311_ (.A(_14234_),
    .B(_10079_),
    .Y(_10080_));
 AO21x1_ASAP7_75t_R _30312_ (.A1(_09718_),
    .A2(_10078_),
    .B(_10080_),
    .Y(_03142_));
 NAND2x1_ASAP7_75t_R _30313_ (.A(_00583_),
    .B(_10070_),
    .Y(_10081_));
 OA21x2_ASAP7_75t_R _30314_ (.A1(_09721_),
    .A2(_10069_),
    .B(_10081_),
    .Y(_03143_));
 AND2x2_ASAP7_75t_R _30315_ (.A(_14421_),
    .B(_10079_),
    .Y(_10082_));
 AO21x1_ASAP7_75t_R _30316_ (.A1(_09786_),
    .A2(_10078_),
    .B(_10082_),
    .Y(_03144_));
 NAND2x1_ASAP7_75t_R _30317_ (.A(_00643_),
    .B(_10070_),
    .Y(_10083_));
 OA21x2_ASAP7_75t_R _30318_ (.A1(_08851_),
    .A2(_10069_),
    .B(_10083_),
    .Y(_03145_));
 NAND2x1_ASAP7_75t_R _30319_ (.A(_00511_),
    .B(_10039_),
    .Y(_10084_));
 OA21x2_ASAP7_75t_R _30320_ (.A1(_09716_),
    .A2(_10038_),
    .B(_10084_),
    .Y(_03146_));
 NAND2x1_ASAP7_75t_R _30321_ (.A(_14511_),
    .B(_10070_),
    .Y(_10085_));
 OAI21x1_ASAP7_75t_R _30322_ (.A1(_08898_),
    .A2(_10069_),
    .B(_10085_),
    .Y(_03147_));
 AND2x2_ASAP7_75t_R _30323_ (.A(_14583_),
    .B(_10079_),
    .Y(_10086_));
 AO21x1_ASAP7_75t_R _30324_ (.A1(_09855_),
    .A2(_10078_),
    .B(_10086_),
    .Y(_03148_));
 NAND2x1_ASAP7_75t_R _30325_ (.A(_00733_),
    .B(_10070_),
    .Y(_10087_));
 OA21x2_ASAP7_75t_R _30326_ (.A1(_08989_),
    .A2(_10069_),
    .B(_10087_),
    .Y(_03149_));
 BUFx10_ASAP7_75t_R _30327_ (.A(_10068_),
    .Y(_10088_));
 NAND2x1_ASAP7_75t_R _30328_ (.A(_00763_),
    .B(_10088_),
    .Y(_10089_));
 OA21x2_ASAP7_75t_R _30329_ (.A1(_09728_),
    .A2(_10069_),
    .B(_10089_),
    .Y(_03150_));
 AND2x2_ASAP7_75t_R _30330_ (.A(_14007_),
    .B(_10079_),
    .Y(_10090_));
 AO21x1_ASAP7_75t_R _30331_ (.A1(_09800_),
    .A2(_10078_),
    .B(_10090_),
    .Y(_03151_));
 NAND2x1_ASAP7_75t_R _30332_ (.A(_00834_),
    .B(_10088_),
    .Y(_10091_));
 OA21x2_ASAP7_75t_R _30333_ (.A1(_09104_),
    .A2(_10069_),
    .B(_10091_),
    .Y(_03152_));
 BUFx4f_ASAP7_75t_R _30334_ (.A(_10079_),
    .Y(_10092_));
 NAND2x1_ASAP7_75t_R _30335_ (.A(_00867_),
    .B(_10088_),
    .Y(_10093_));
 OA21x2_ASAP7_75t_R _30336_ (.A1(_09144_),
    .A2(_10092_),
    .B(_10093_),
    .Y(_03153_));
 NAND2x1_ASAP7_75t_R _30337_ (.A(_00900_),
    .B(_10088_),
    .Y(_10094_));
 OA21x2_ASAP7_75t_R _30338_ (.A1(_09181_),
    .A2(_10092_),
    .B(_10094_),
    .Y(_03154_));
 NOR2x1_ASAP7_75t_R _30339_ (.A(_00933_),
    .B(_10077_),
    .Y(_10095_));
 AO21x1_ASAP7_75t_R _30340_ (.A1(_09738_),
    .A2(_10078_),
    .B(_10095_),
    .Y(_03155_));
 NAND2x1_ASAP7_75t_R _30341_ (.A(_00966_),
    .B(_10088_),
    .Y(_10096_));
 OA21x2_ASAP7_75t_R _30342_ (.A1(_09245_),
    .A2(_10092_),
    .B(_10096_),
    .Y(_03156_));
 AND3x4_ASAP7_75t_R _30343_ (.A(_14051_),
    .B(_08595_),
    .C(_09774_),
    .Y(_10097_));
 BUFx6f_ASAP7_75t_R _30344_ (.A(_10097_),
    .Y(_10098_));
 NOR2x1_ASAP7_75t_R _30345_ (.A(_00541_),
    .B(_10098_),
    .Y(_10099_));
 AO21x1_ASAP7_75t_R _30346_ (.A1(_09718_),
    .A2(_10098_),
    .B(_10099_),
    .Y(_03157_));
 NAND2x1_ASAP7_75t_R _30347_ (.A(_00999_),
    .B(_10088_),
    .Y(_10100_));
 OA21x2_ASAP7_75t_R _30348_ (.A1(_09271_),
    .A2(_10092_),
    .B(_10100_),
    .Y(_03158_));
 NAND2x1_ASAP7_75t_R _30349_ (.A(_01032_),
    .B(_10088_),
    .Y(_10101_));
 OA21x2_ASAP7_75t_R _30350_ (.A1(_09299_),
    .A2(_10092_),
    .B(_10101_),
    .Y(_03159_));
 NAND2x1_ASAP7_75t_R _30351_ (.A(_01065_),
    .B(_10088_),
    .Y(_10102_));
 OA21x2_ASAP7_75t_R _30352_ (.A1(_09328_),
    .A2(_10092_),
    .B(_10102_),
    .Y(_03160_));
 NAND2x1_ASAP7_75t_R _30353_ (.A(_01098_),
    .B(_10088_),
    .Y(_10103_));
 OA21x2_ASAP7_75t_R _30354_ (.A1(_09357_),
    .A2(_10092_),
    .B(_10103_),
    .Y(_03161_));
 NAND2x1_ASAP7_75t_R _30355_ (.A(_01131_),
    .B(_10088_),
    .Y(_10104_));
 OA21x2_ASAP7_75t_R _30356_ (.A1(_09390_),
    .A2(_10092_),
    .B(_10104_),
    .Y(_03162_));
 NOR2x1_ASAP7_75t_R _30357_ (.A(_01164_),
    .B(_10077_),
    .Y(_10105_));
 AO21x1_ASAP7_75t_R _30358_ (.A1(_09821_),
    .A2(_10078_),
    .B(_10105_),
    .Y(_03163_));
 NAND2x1_ASAP7_75t_R _30359_ (.A(_01197_),
    .B(_10079_),
    .Y(_10106_));
 OA21x2_ASAP7_75t_R _30360_ (.A1(_09749_),
    .A2(_10092_),
    .B(_10106_),
    .Y(_03164_));
 NAND2x1_ASAP7_75t_R _30361_ (.A(_01230_),
    .B(_10079_),
    .Y(_10107_));
 OA21x2_ASAP7_75t_R _30362_ (.A1(_09472_),
    .A2(_10092_),
    .B(_10107_),
    .Y(_03165_));
 NAND2x1_ASAP7_75t_R _30363_ (.A(_01263_),
    .B(_10079_),
    .Y(_10108_));
 OA21x2_ASAP7_75t_R _30364_ (.A1(_09495_),
    .A2(_10070_),
    .B(_10108_),
    .Y(_03166_));
 NOR2x1_ASAP7_75t_R _30365_ (.A(_01296_),
    .B(_10077_),
    .Y(_10109_));
 AO21x1_ASAP7_75t_R _30366_ (.A1(_09753_),
    .A2(_10078_),
    .B(_10109_),
    .Y(_03167_));
 BUFx10_ASAP7_75t_R _30367_ (.A(_10037_),
    .Y(_10110_));
 NAND2x1_ASAP7_75t_R _30368_ (.A(_00573_),
    .B(_10110_),
    .Y(_10111_));
 OA21x2_ASAP7_75t_R _30369_ (.A1(_09721_),
    .A2(_10038_),
    .B(_10111_),
    .Y(_03168_));
 NOR2x1_ASAP7_75t_R _30370_ (.A(_01329_),
    .B(_10077_),
    .Y(_10112_));
 AO21x1_ASAP7_75t_R _30371_ (.A1(_09755_),
    .A2(_10078_),
    .B(_10112_),
    .Y(_03169_));
 NAND2x1_ASAP7_75t_R _30372_ (.A(_01362_),
    .B(_10079_),
    .Y(_10113_));
 OA21x2_ASAP7_75t_R _30373_ (.A1(_09757_),
    .A2(_10070_),
    .B(_10113_),
    .Y(_03170_));
 NOR2x1_ASAP7_75t_R _30374_ (.A(_01395_),
    .B(_10077_),
    .Y(_10114_));
 AO21x1_ASAP7_75t_R _30375_ (.A1(net152),
    .A2(_10078_),
    .B(_10114_),
    .Y(_03171_));
 AND2x2_ASAP7_75t_R _30376_ (.A(_04810_),
    .B(_10079_),
    .Y(_10115_));
 AO21x1_ASAP7_75t_R _30377_ (.A1(net8),
    .A2(_10078_),
    .B(_10115_),
    .Y(_03172_));
 NAND2x2_ASAP7_75t_R _30378_ (.A(_08341_),
    .B(_10075_),
    .Y(_10116_));
 OR3x1_ASAP7_75t_R _30379_ (.A(_09838_),
    .B(_08589_),
    .C(_10067_),
    .Y(_10117_));
 BUFx6f_ASAP7_75t_R _30380_ (.A(_10117_),
    .Y(_10118_));
 NAND2x1_ASAP7_75t_R _30381_ (.A(_00427_),
    .B(_10118_),
    .Y(_10119_));
 OA21x2_ASAP7_75t_R _30382_ (.A1(_09650_),
    .A2(_10116_),
    .B(_10119_),
    .Y(_03173_));
 AND4x1_ASAP7_75t_R _30383_ (.A(_14726_),
    .B(_08330_),
    .C(_08338_),
    .D(_10075_),
    .Y(_10120_));
 BUFx6f_ASAP7_75t_R _30384_ (.A(_10120_),
    .Y(_10121_));
 BUFx4f_ASAP7_75t_R _30385_ (.A(_10121_),
    .Y(_10122_));
 BUFx10_ASAP7_75t_R _30386_ (.A(_10121_),
    .Y(_10123_));
 NOR2x1_ASAP7_75t_R _30387_ (.A(_00380_),
    .B(_10123_),
    .Y(_10124_));
 AO21x1_ASAP7_75t_R _30388_ (.A1(_09772_),
    .A2(_10122_),
    .B(_10124_),
    .Y(_03174_));
 NAND2x1_ASAP7_75t_R _30389_ (.A(_00491_),
    .B(_10118_),
    .Y(_10125_));
 OA21x2_ASAP7_75t_R _30390_ (.A1(_09780_),
    .A2(_10118_),
    .B(_10125_),
    .Y(_03175_));
 NOR2x1_ASAP7_75t_R _30391_ (.A(_00522_),
    .B(_10123_),
    .Y(_10126_));
 AO21x1_ASAP7_75t_R _30392_ (.A1(_09782_),
    .A2(_10122_),
    .B(_10126_),
    .Y(_03176_));
 NOR2x1_ASAP7_75t_R _30393_ (.A(_00552_),
    .B(_10123_),
    .Y(_10127_));
 AO21x1_ASAP7_75t_R _30394_ (.A1(_09718_),
    .A2(_10122_),
    .B(_10127_),
    .Y(_03177_));
 NAND2x1_ASAP7_75t_R _30395_ (.A(_00584_),
    .B(_10118_),
    .Y(_10128_));
 OA21x2_ASAP7_75t_R _30396_ (.A1(_09721_),
    .A2(_10118_),
    .B(_10128_),
    .Y(_03178_));
 NAND2x1_ASAP7_75t_R _30397_ (.A(_00603_),
    .B(_10110_),
    .Y(_10129_));
 OA21x2_ASAP7_75t_R _30398_ (.A1(_08810_),
    .A2(_10038_),
    .B(_10129_),
    .Y(_03179_));
 NOR2x1_ASAP7_75t_R _30399_ (.A(_00614_),
    .B(_10123_),
    .Y(_10130_));
 AO21x1_ASAP7_75t_R _30400_ (.A1(_09786_),
    .A2(_10122_),
    .B(_10130_),
    .Y(_03180_));
 BUFx10_ASAP7_75t_R _30401_ (.A(_10121_),
    .Y(_10131_));
 NOR2x1_ASAP7_75t_R _30402_ (.A(_00644_),
    .B(_10131_),
    .Y(_10132_));
 AO21x1_ASAP7_75t_R _30403_ (.A1(_09788_),
    .A2(_10122_),
    .B(_10132_),
    .Y(_03181_));
 OR2x2_ASAP7_75t_R _30404_ (.A(_00674_),
    .B(_10121_),
    .Y(_10133_));
 OAI21x1_ASAP7_75t_R _30405_ (.A1(_08898_),
    .A2(_10116_),
    .B(_10133_),
    .Y(_03182_));
 NOR2x1_ASAP7_75t_R _30406_ (.A(_00704_),
    .B(_10131_),
    .Y(_10134_));
 AO21x1_ASAP7_75t_R _30407_ (.A1(_09855_),
    .A2(_10122_),
    .B(_10134_),
    .Y(_03183_));
 NOR2x1_ASAP7_75t_R _30408_ (.A(_00734_),
    .B(_10131_),
    .Y(_10135_));
 AO21x1_ASAP7_75t_R _30409_ (.A1(_09108_),
    .A2(_10122_),
    .B(_10135_),
    .Y(_03184_));
 NOR2x1_ASAP7_75t_R _30410_ (.A(_00764_),
    .B(_10131_),
    .Y(_10136_));
 AO21x1_ASAP7_75t_R _30411_ (.A1(_09037_),
    .A2(_10122_),
    .B(_10136_),
    .Y(_03185_));
 NOR2x1_ASAP7_75t_R _30412_ (.A(_00460_),
    .B(_10131_),
    .Y(_10137_));
 AO21x1_ASAP7_75t_R _30413_ (.A1(_09800_),
    .A2(_10122_),
    .B(_10137_),
    .Y(_03186_));
 NOR2x1_ASAP7_75t_R _30414_ (.A(_00835_),
    .B(_10131_),
    .Y(_10138_));
 AO21x1_ASAP7_75t_R _30415_ (.A1(_09731_),
    .A2(_10122_),
    .B(_10138_),
    .Y(_03187_));
 BUFx4f_ASAP7_75t_R _30416_ (.A(_10121_),
    .Y(_10139_));
 NOR2x1_ASAP7_75t_R _30417_ (.A(_00868_),
    .B(_10131_),
    .Y(_10140_));
 AO21x1_ASAP7_75t_R _30418_ (.A1(_09745_),
    .A2(_10139_),
    .B(_10140_),
    .Y(_03188_));
 NOR2x1_ASAP7_75t_R _30419_ (.A(_00901_),
    .B(_10131_),
    .Y(_10141_));
 AO21x1_ASAP7_75t_R _30420_ (.A1(_09763_),
    .A2(_10139_),
    .B(_10141_),
    .Y(_03189_));
 NAND2x1_ASAP7_75t_R _30421_ (.A(_00633_),
    .B(_10110_),
    .Y(_10142_));
 OA21x2_ASAP7_75t_R _30422_ (.A1(_08851_),
    .A2(_10038_),
    .B(_10142_),
    .Y(_03190_));
 NAND2x1_ASAP7_75t_R _30423_ (.A(_01789_),
    .B(_09106_),
    .Y(_10143_));
 OA21x2_ASAP7_75t_R _30424_ (.A1(_09866_),
    .A2(_09716_),
    .B(_10143_),
    .Y(_03191_));
 NOR2x1_ASAP7_75t_R _30425_ (.A(_00934_),
    .B(_10131_),
    .Y(_10144_));
 AO21x1_ASAP7_75t_R _30426_ (.A1(_09738_),
    .A2(_10139_),
    .B(_10144_),
    .Y(_03192_));
 NOR2x1_ASAP7_75t_R _30427_ (.A(_00967_),
    .B(_10131_),
    .Y(_10145_));
 AO21x1_ASAP7_75t_R _30428_ (.A1(_09808_),
    .A2(_10139_),
    .B(_10145_),
    .Y(_03193_));
 BUFx6f_ASAP7_75t_R _30429_ (.A(_10121_),
    .Y(_10146_));
 NOR2x1_ASAP7_75t_R _30430_ (.A(_01000_),
    .B(_10146_),
    .Y(_10147_));
 AO21x1_ASAP7_75t_R _30431_ (.A1(_09810_),
    .A2(_10139_),
    .B(_10147_),
    .Y(_03194_));
 NOR2x1_ASAP7_75t_R _30432_ (.A(_01033_),
    .B(_10146_),
    .Y(_10148_));
 AO21x1_ASAP7_75t_R _30433_ (.A1(_09812_),
    .A2(_10139_),
    .B(_10148_),
    .Y(_03195_));
 NOR2x1_ASAP7_75t_R _30434_ (.A(_01066_),
    .B(_10146_),
    .Y(_10149_));
 AO21x1_ASAP7_75t_R _30435_ (.A1(_09815_),
    .A2(_10139_),
    .B(_10149_),
    .Y(_03196_));
 NOR2x1_ASAP7_75t_R _30436_ (.A(_01099_),
    .B(_10146_),
    .Y(_10150_));
 AO21x1_ASAP7_75t_R _30437_ (.A1(_09817_),
    .A2(_10139_),
    .B(_10150_),
    .Y(_03197_));
 NOR2x1_ASAP7_75t_R _30438_ (.A(_01132_),
    .B(_10146_),
    .Y(_10151_));
 AO21x1_ASAP7_75t_R _30439_ (.A1(_09819_),
    .A2(_10139_),
    .B(_10151_),
    .Y(_03198_));
 NOR2x1_ASAP7_75t_R _30440_ (.A(_01165_),
    .B(_10146_),
    .Y(_10152_));
 AO21x1_ASAP7_75t_R _30441_ (.A1(_09821_),
    .A2(_10139_),
    .B(_10152_),
    .Y(_03199_));
 NAND2x1_ASAP7_75t_R _30442_ (.A(_01198_),
    .B(_10118_),
    .Y(_10153_));
 OA21x2_ASAP7_75t_R _30443_ (.A1(_09749_),
    .A2(_10118_),
    .B(_10153_),
    .Y(_03200_));
 NOR2x1_ASAP7_75t_R _30444_ (.A(_01231_),
    .B(_10146_),
    .Y(_10154_));
 AO21x1_ASAP7_75t_R _30445_ (.A1(_09824_),
    .A2(_10123_),
    .B(_10154_),
    .Y(_03201_));
 OR2x2_ASAP7_75t_R _30446_ (.A(_00663_),
    .B(_10097_),
    .Y(_10155_));
 OAI21x1_ASAP7_75t_R _30447_ (.A1(_08898_),
    .A2(_10038_),
    .B(_10155_),
    .Y(_03202_));
 NOR2x1_ASAP7_75t_R _30448_ (.A(_01264_),
    .B(_10146_),
    .Y(_10156_));
 AO21x1_ASAP7_75t_R _30449_ (.A1(_09826_),
    .A2(_10123_),
    .B(_10156_),
    .Y(_03203_));
 NOR2x1_ASAP7_75t_R _30450_ (.A(_01297_),
    .B(_10146_),
    .Y(_10157_));
 AO21x1_ASAP7_75t_R _30451_ (.A1(_09753_),
    .A2(_10123_),
    .B(_10157_),
    .Y(_03204_));
 NOR2x1_ASAP7_75t_R _30452_ (.A(_01330_),
    .B(_10146_),
    .Y(_10158_));
 AO21x1_ASAP7_75t_R _30453_ (.A1(_09755_),
    .A2(_10123_),
    .B(_10158_),
    .Y(_03205_));
 NAND2x1_ASAP7_75t_R _30454_ (.A(_01363_),
    .B(_10118_),
    .Y(_10159_));
 OA21x2_ASAP7_75t_R _30455_ (.A1(net13),
    .A2(_10118_),
    .B(_10159_),
    .Y(_03206_));
 NOR2x1_ASAP7_75t_R _30456_ (.A(_01396_),
    .B(_10121_),
    .Y(_10160_));
 AO21x1_ASAP7_75t_R _30457_ (.A1(_09759_),
    .A2(_10123_),
    .B(_10160_),
    .Y(_03207_));
 AND2x2_ASAP7_75t_R _30458_ (.A(_04816_),
    .B(_10118_),
    .Y(_10161_));
 AO21x1_ASAP7_75t_R _30459_ (.A1(_09761_),
    .A2(_10123_),
    .B(_10161_),
    .Y(_03208_));
 BUFx4f_ASAP7_75t_R _30460_ (.A(_08584_),
    .Y(_10162_));
 OR3x4_ASAP7_75t_R _30461_ (.A(_09766_),
    .B(_09767_),
    .C(_10067_),
    .Y(_10163_));
 BUFx10_ASAP7_75t_R _30462_ (.A(_10163_),
    .Y(_10164_));
 BUFx6f_ASAP7_75t_R _30463_ (.A(_10164_),
    .Y(_10165_));
 NAND2x1_ASAP7_75t_R _30464_ (.A(_00428_),
    .B(_10165_),
    .Y(_10166_));
 OA21x2_ASAP7_75t_R _30465_ (.A1(_10162_),
    .A2(_10165_),
    .B(_10166_),
    .Y(_03209_));
 AND3x1_ASAP7_75t_R _30466_ (.A(_08339_),
    .B(_09774_),
    .C(_10075_),
    .Y(_10167_));
 BUFx6f_ASAP7_75t_R _30467_ (.A(_10167_),
    .Y(_10168_));
 BUFx4f_ASAP7_75t_R _30468_ (.A(_10168_),
    .Y(_10169_));
 BUFx6f_ASAP7_75t_R _30469_ (.A(_10163_),
    .Y(_10170_));
 AND2x2_ASAP7_75t_R _30470_ (.A(_13488_),
    .B(_10170_),
    .Y(_10171_));
 AO21x1_ASAP7_75t_R _30471_ (.A1(_09772_),
    .A2(_10169_),
    .B(_10171_),
    .Y(_03210_));
 NAND2x1_ASAP7_75t_R _30472_ (.A(_00492_),
    .B(_10165_),
    .Y(_10172_));
 OA21x2_ASAP7_75t_R _30473_ (.A1(_09780_),
    .A2(_10165_),
    .B(_10172_),
    .Y(_03211_));
 AND2x2_ASAP7_75t_R _30474_ (.A(_14183_),
    .B(_10170_),
    .Y(_10173_));
 AO21x1_ASAP7_75t_R _30475_ (.A1(_09782_),
    .A2(_10169_),
    .B(_10173_),
    .Y(_03212_));
 NAND2x1_ASAP7_75t_R _30476_ (.A(_00693_),
    .B(_10110_),
    .Y(_10174_));
 OA21x2_ASAP7_75t_R _30477_ (.A1(_08943_),
    .A2(_10038_),
    .B(_10174_),
    .Y(_03213_));
 BUFx6f_ASAP7_75t_R _30478_ (.A(_08675_),
    .Y(_10175_));
 AND2x2_ASAP7_75t_R _30479_ (.A(_15018_),
    .B(_10170_),
    .Y(_10176_));
 AO21x1_ASAP7_75t_R _30480_ (.A1(_10175_),
    .A2(_10169_),
    .B(_10176_),
    .Y(_03214_));
 BUFx6f_ASAP7_75t_R _30481_ (.A(_08762_),
    .Y(_10177_));
 NAND2x1_ASAP7_75t_R _30482_ (.A(_00585_),
    .B(_10165_),
    .Y(_10178_));
 OA21x2_ASAP7_75t_R _30483_ (.A1(_10177_),
    .A2(_10165_),
    .B(_10178_),
    .Y(_03215_));
 AND2x2_ASAP7_75t_R _30484_ (.A(_14418_),
    .B(_10170_),
    .Y(_10179_));
 AO21x1_ASAP7_75t_R _30485_ (.A1(_09786_),
    .A2(_10169_),
    .B(_10179_),
    .Y(_03216_));
 AND2x2_ASAP7_75t_R _30486_ (.A(_14455_),
    .B(_10170_),
    .Y(_10180_));
 AO21x1_ASAP7_75t_R _30487_ (.A1(_09788_),
    .A2(_10169_),
    .B(_10180_),
    .Y(_03217_));
 NAND2x1_ASAP7_75t_R _30488_ (.A(_14508_),
    .B(_10165_),
    .Y(_10181_));
 OAI21x1_ASAP7_75t_R _30489_ (.A1(_08898_),
    .A2(_10165_),
    .B(_10181_),
    .Y(_03218_));
 AND2x2_ASAP7_75t_R _30490_ (.A(_14580_),
    .B(_10170_),
    .Y(_10182_));
 AO21x1_ASAP7_75t_R _30491_ (.A1(_09855_),
    .A2(_10169_),
    .B(_10182_),
    .Y(_03219_));
 AND2x2_ASAP7_75t_R _30492_ (.A(_14649_),
    .B(_10170_),
    .Y(_10183_));
 AO21x1_ASAP7_75t_R _30493_ (.A1(_09108_),
    .A2(_10169_),
    .B(_10183_),
    .Y(_03220_));
 AND2x2_ASAP7_75t_R _30494_ (.A(_14700_),
    .B(_10170_),
    .Y(_10184_));
 AO21x1_ASAP7_75t_R _30495_ (.A1(_09037_),
    .A2(_10169_),
    .B(_10184_),
    .Y(_03221_));
 BUFx4f_ASAP7_75t_R _30496_ (.A(_10164_),
    .Y(_10185_));
 AND2x2_ASAP7_75t_R _30497_ (.A(_13985_),
    .B(_10185_),
    .Y(_10186_));
 AO21x1_ASAP7_75t_R _30498_ (.A1(_09800_),
    .A2(_10169_),
    .B(_10186_),
    .Y(_03222_));
 AND2x2_ASAP7_75t_R _30499_ (.A(_15626_),
    .B(_10185_),
    .Y(_10187_));
 AO21x1_ASAP7_75t_R _30500_ (.A1(_09731_),
    .A2(_10169_),
    .B(_10187_),
    .Y(_03223_));
 NAND2x1_ASAP7_75t_R _30501_ (.A(_00723_),
    .B(_10110_),
    .Y(_10188_));
 OA21x2_ASAP7_75t_R _30502_ (.A1(_08989_),
    .A2(_10038_),
    .B(_10188_),
    .Y(_03224_));
 BUFx4f_ASAP7_75t_R _30503_ (.A(_10168_),
    .Y(_10189_));
 AND2x2_ASAP7_75t_R _30504_ (.A(_15777_),
    .B(_10185_),
    .Y(_10190_));
 AO21x1_ASAP7_75t_R _30505_ (.A1(_09745_),
    .A2(_10189_),
    .B(_10190_),
    .Y(_03225_));
 AND2x2_ASAP7_75t_R _30506_ (.A(_15906_),
    .B(_10185_),
    .Y(_10191_));
 AO21x1_ASAP7_75t_R _30507_ (.A1(_09763_),
    .A2(_10189_),
    .B(_10191_),
    .Y(_03226_));
 AND2x2_ASAP7_75t_R _30508_ (.A(_16055_),
    .B(_10185_),
    .Y(_10192_));
 AO21x1_ASAP7_75t_R _30509_ (.A1(_09738_),
    .A2(_10189_),
    .B(_10192_),
    .Y(_03227_));
 AND2x2_ASAP7_75t_R _30510_ (.A(_16172_),
    .B(_10185_),
    .Y(_10193_));
 AO21x1_ASAP7_75t_R _30511_ (.A1(_09808_),
    .A2(_10189_),
    .B(_10193_),
    .Y(_03228_));
 AND2x2_ASAP7_75t_R _30512_ (.A(_16315_),
    .B(_10185_),
    .Y(_10194_));
 AO21x1_ASAP7_75t_R _30513_ (.A1(_09810_),
    .A2(_10189_),
    .B(_10194_),
    .Y(_03229_));
 AND2x2_ASAP7_75t_R _30514_ (.A(_16429_),
    .B(_10185_),
    .Y(_10195_));
 AO21x1_ASAP7_75t_R _30515_ (.A1(_09812_),
    .A2(_10189_),
    .B(_10195_),
    .Y(_03230_));
 AND2x2_ASAP7_75t_R _30516_ (.A(_16555_),
    .B(_10185_),
    .Y(_10196_));
 AO21x1_ASAP7_75t_R _30517_ (.A1(_09815_),
    .A2(_10189_),
    .B(_10196_),
    .Y(_03231_));
 AND2x2_ASAP7_75t_R _30518_ (.A(_16669_),
    .B(_10185_),
    .Y(_10197_));
 AO21x1_ASAP7_75t_R _30519_ (.A1(_09817_),
    .A2(_10189_),
    .B(_10197_),
    .Y(_03232_));
 AND2x2_ASAP7_75t_R _30520_ (.A(_16799_),
    .B(_10164_),
    .Y(_10198_));
 AO21x1_ASAP7_75t_R _30521_ (.A1(_09819_),
    .A2(_10189_),
    .B(_10198_),
    .Y(_03233_));
 AND2x2_ASAP7_75t_R _30522_ (.A(_16909_),
    .B(_10164_),
    .Y(_10199_));
 AO21x1_ASAP7_75t_R _30523_ (.A1(_09821_),
    .A2(_10189_),
    .B(_10199_),
    .Y(_03234_));
 BUFx6f_ASAP7_75t_R _30524_ (.A(_10037_),
    .Y(_10200_));
 NAND2x1_ASAP7_75t_R _30525_ (.A(_00753_),
    .B(_10110_),
    .Y(_10201_));
 OA21x2_ASAP7_75t_R _30526_ (.A1(_09728_),
    .A2(_10200_),
    .B(_10201_),
    .Y(_03235_));
 NAND2x1_ASAP7_75t_R _30527_ (.A(_01199_),
    .B(_10170_),
    .Y(_10202_));
 OA21x2_ASAP7_75t_R _30528_ (.A1(_09749_),
    .A2(_10165_),
    .B(_10202_),
    .Y(_03236_));
 AND2x2_ASAP7_75t_R _30529_ (.A(_17148_),
    .B(_10164_),
    .Y(_10203_));
 AO21x1_ASAP7_75t_R _30530_ (.A1(_09824_),
    .A2(_10168_),
    .B(_10203_),
    .Y(_03237_));
 AND2x2_ASAP7_75t_R _30531_ (.A(_17279_),
    .B(_10164_),
    .Y(_10204_));
 AO21x1_ASAP7_75t_R _30532_ (.A1(_09826_),
    .A2(_10168_),
    .B(_10204_),
    .Y(_03238_));
 AND2x2_ASAP7_75t_R _30533_ (.A(_04306_),
    .B(_10164_),
    .Y(_10205_));
 AO21x1_ASAP7_75t_R _30534_ (.A1(_09753_),
    .A2(_10168_),
    .B(_10205_),
    .Y(_03239_));
 AND2x2_ASAP7_75t_R _30535_ (.A(_04436_),
    .B(_10164_),
    .Y(_10206_));
 AO21x1_ASAP7_75t_R _30536_ (.A1(_09755_),
    .A2(_10168_),
    .B(_10206_),
    .Y(_03240_));
 NAND2x1_ASAP7_75t_R _30537_ (.A(_01364_),
    .B(_10170_),
    .Y(_10207_));
 OA21x2_ASAP7_75t_R _30538_ (.A1(_09757_),
    .A2(_10165_),
    .B(_10207_),
    .Y(_03241_));
 AND2x2_ASAP7_75t_R _30539_ (.A(_04660_),
    .B(_10164_),
    .Y(_10208_));
 AO21x1_ASAP7_75t_R _30540_ (.A1(net152),
    .A2(_10168_),
    .B(_10208_),
    .Y(_03242_));
 AND2x2_ASAP7_75t_R _30541_ (.A(_04787_),
    .B(_10164_),
    .Y(_10209_));
 AO21x1_ASAP7_75t_R _30542_ (.A1(net8),
    .A2(_10168_),
    .B(_10209_),
    .Y(_03243_));
 AND4x2_ASAP7_75t_R _30543_ (.A(_08329_),
    .B(_09773_),
    .C(_09834_),
    .D(_10075_),
    .Y(_10210_));
 BUFx10_ASAP7_75t_R _30544_ (.A(_10210_),
    .Y(_10211_));
 INVx1_ASAP7_75t_R _30545_ (.A(_10211_),
    .Y(_10212_));
 OR4x2_ASAP7_75t_R _30546_ (.A(_08593_),
    .B(_08594_),
    .C(_09838_),
    .D(_10067_),
    .Y(_10213_));
 BUFx6f_ASAP7_75t_R _30547_ (.A(_10213_),
    .Y(_10214_));
 NAND2x1_ASAP7_75t_R _30548_ (.A(_00429_),
    .B(_10214_),
    .Y(_10215_));
 OA21x2_ASAP7_75t_R _30549_ (.A1(_10162_),
    .A2(_10212_),
    .B(_10215_),
    .Y(_03244_));
 BUFx4f_ASAP7_75t_R _30550_ (.A(_10211_),
    .Y(_10216_));
 BUFx10_ASAP7_75t_R _30551_ (.A(_10210_),
    .Y(_10217_));
 NOR2x1_ASAP7_75t_R _30552_ (.A(_00382_),
    .B(_10217_),
    .Y(_10218_));
 AO21x1_ASAP7_75t_R _30553_ (.A1(_09772_),
    .A2(_10216_),
    .B(_10218_),
    .Y(_03245_));
 NAND2x1_ASAP7_75t_R _30554_ (.A(_00449_),
    .B(_10110_),
    .Y(_10219_));
 OA21x2_ASAP7_75t_R _30555_ (.A1(_09074_),
    .A2(_10200_),
    .B(_10219_),
    .Y(_03246_));
 BUFx6f_ASAP7_75t_R _30556_ (.A(_09695_),
    .Y(_10220_));
 NAND2x1_ASAP7_75t_R _30557_ (.A(_00493_),
    .B(_10214_),
    .Y(_10221_));
 OA21x2_ASAP7_75t_R _30558_ (.A1(_10220_),
    .A2(_10214_),
    .B(_10221_),
    .Y(_03247_));
 NOR2x1_ASAP7_75t_R _30559_ (.A(_00524_),
    .B(_10217_),
    .Y(_10222_));
 AO21x1_ASAP7_75t_R _30560_ (.A1(_09782_),
    .A2(_10216_),
    .B(_10222_),
    .Y(_03248_));
 AND2x2_ASAP7_75t_R _30561_ (.A(_15014_),
    .B(_10213_),
    .Y(_10223_));
 AO21x1_ASAP7_75t_R _30562_ (.A1(_10175_),
    .A2(_10216_),
    .B(_10223_),
    .Y(_03249_));
 NAND2x1_ASAP7_75t_R _30563_ (.A(_00586_),
    .B(_10214_),
    .Y(_10224_));
 OA21x2_ASAP7_75t_R _30564_ (.A1(_10177_),
    .A2(_10214_),
    .B(_10224_),
    .Y(_03250_));
 NOR2x1_ASAP7_75t_R _30565_ (.A(_00616_),
    .B(_10217_),
    .Y(_10225_));
 AO21x1_ASAP7_75t_R _30566_ (.A1(_09786_),
    .A2(_10216_),
    .B(_10225_),
    .Y(_03251_));
 NOR2x1_ASAP7_75t_R _30567_ (.A(_00646_),
    .B(_10217_),
    .Y(_10226_));
 AO21x1_ASAP7_75t_R _30568_ (.A1(_09788_),
    .A2(_10216_),
    .B(_10226_),
    .Y(_03252_));
 NAND2x1_ASAP7_75t_R _30569_ (.A(_15296_),
    .B(_10214_),
    .Y(_10227_));
 OAI21x1_ASAP7_75t_R _30570_ (.A1(_08898_),
    .A2(_10212_),
    .B(_10227_),
    .Y(_03253_));
 BUFx10_ASAP7_75t_R _30571_ (.A(_10211_),
    .Y(_10228_));
 NOR2x1_ASAP7_75t_R _30572_ (.A(_00706_),
    .B(_10228_),
    .Y(_10229_));
 AO21x1_ASAP7_75t_R _30573_ (.A1(_09855_),
    .A2(_10216_),
    .B(_10229_),
    .Y(_03254_));
 NOR2x1_ASAP7_75t_R _30574_ (.A(_00736_),
    .B(_10228_),
    .Y(_10230_));
 AO21x1_ASAP7_75t_R _30575_ (.A1(_09108_),
    .A2(_10216_),
    .B(_10230_),
    .Y(_03255_));
 NOR2x1_ASAP7_75t_R _30576_ (.A(_00766_),
    .B(_10228_),
    .Y(_10231_));
 AO21x1_ASAP7_75t_R _30577_ (.A1(_09037_),
    .A2(_10216_),
    .B(_10231_),
    .Y(_03256_));
 NAND2x1_ASAP7_75t_R _30578_ (.A(_00824_),
    .B(_10110_),
    .Y(_10232_));
 OA21x2_ASAP7_75t_R _30579_ (.A1(_09104_),
    .A2(_10200_),
    .B(_10232_),
    .Y(_03257_));
 NOR2x1_ASAP7_75t_R _30580_ (.A(_00462_),
    .B(_10228_),
    .Y(_10233_));
 AO21x1_ASAP7_75t_R _30581_ (.A1(_09800_),
    .A2(_10216_),
    .B(_10233_),
    .Y(_03258_));
 NOR2x1_ASAP7_75t_R _30582_ (.A(_00837_),
    .B(_10228_),
    .Y(_10234_));
 AO21x1_ASAP7_75t_R _30583_ (.A1(_09731_),
    .A2(_10216_),
    .B(_10234_),
    .Y(_03259_));
 BUFx4f_ASAP7_75t_R _30584_ (.A(_10211_),
    .Y(_10235_));
 NOR2x1_ASAP7_75t_R _30585_ (.A(_00870_),
    .B(_10228_),
    .Y(_10236_));
 AO21x1_ASAP7_75t_R _30586_ (.A1(_09745_),
    .A2(_10235_),
    .B(_10236_),
    .Y(_03260_));
 NOR2x1_ASAP7_75t_R _30587_ (.A(_00903_),
    .B(_10228_),
    .Y(_10237_));
 AO21x1_ASAP7_75t_R _30588_ (.A1(_09763_),
    .A2(_10235_),
    .B(_10237_),
    .Y(_03261_));
 BUFx6f_ASAP7_75t_R _30589_ (.A(_09213_),
    .Y(_10238_));
 AND2x2_ASAP7_75t_R _30590_ (.A(_16052_),
    .B(_10213_),
    .Y(_10239_));
 AO21x1_ASAP7_75t_R _30591_ (.A1(_10238_),
    .A2(_10235_),
    .B(_10239_),
    .Y(_03262_));
 NOR2x1_ASAP7_75t_R _30592_ (.A(_00969_),
    .B(_10228_),
    .Y(_10240_));
 AO21x1_ASAP7_75t_R _30593_ (.A1(_09808_),
    .A2(_10235_),
    .B(_10240_),
    .Y(_03263_));
 NOR2x1_ASAP7_75t_R _30594_ (.A(_01002_),
    .B(_10228_),
    .Y(_10241_));
 AO21x1_ASAP7_75t_R _30595_ (.A1(_09810_),
    .A2(_10235_),
    .B(_10241_),
    .Y(_03264_));
 NOR2x1_ASAP7_75t_R _30596_ (.A(_01035_),
    .B(_10228_),
    .Y(_10242_));
 AO21x1_ASAP7_75t_R _30597_ (.A1(_09812_),
    .A2(_10235_),
    .B(_10242_),
    .Y(_03265_));
 NOR2x1_ASAP7_75t_R _30598_ (.A(_01068_),
    .B(_10211_),
    .Y(_10243_));
 AO21x1_ASAP7_75t_R _30599_ (.A1(_09815_),
    .A2(_10235_),
    .B(_10243_),
    .Y(_03266_));
 NOR2x1_ASAP7_75t_R _30600_ (.A(_01101_),
    .B(_10211_),
    .Y(_10244_));
 AO21x1_ASAP7_75t_R _30601_ (.A1(_09817_),
    .A2(_10235_),
    .B(_10244_),
    .Y(_03267_));
 NAND2x1_ASAP7_75t_R _30602_ (.A(_00857_),
    .B(_10110_),
    .Y(_10245_));
 OA21x2_ASAP7_75t_R _30603_ (.A1(_09144_),
    .A2(_10200_),
    .B(_10245_),
    .Y(_03268_));
 NOR2x1_ASAP7_75t_R _30604_ (.A(_01134_),
    .B(_10211_),
    .Y(_10246_));
 AO21x1_ASAP7_75t_R _30605_ (.A1(_09819_),
    .A2(_10235_),
    .B(_10246_),
    .Y(_03269_));
 NOR2x1_ASAP7_75t_R _30606_ (.A(_01167_),
    .B(_10211_),
    .Y(_10247_));
 AO21x1_ASAP7_75t_R _30607_ (.A1(_09821_),
    .A2(_10235_),
    .B(_10247_),
    .Y(_03270_));
 BUFx6f_ASAP7_75t_R _30608_ (.A(_09441_),
    .Y(_10248_));
 NAND2x1_ASAP7_75t_R _30609_ (.A(_01200_),
    .B(_10214_),
    .Y(_10249_));
 OA21x2_ASAP7_75t_R _30610_ (.A1(_10248_),
    .A2(_10214_),
    .B(_10249_),
    .Y(_03271_));
 NOR2x1_ASAP7_75t_R _30611_ (.A(_01233_),
    .B(_10211_),
    .Y(_10250_));
 AO21x1_ASAP7_75t_R _30612_ (.A1(_09824_),
    .A2(_10217_),
    .B(_10250_),
    .Y(_03272_));
 NOR2x1_ASAP7_75t_R _30613_ (.A(_01266_),
    .B(_10211_),
    .Y(_10251_));
 AO21x1_ASAP7_75t_R _30614_ (.A1(_09826_),
    .A2(_10217_),
    .B(_10251_),
    .Y(_03273_));
 AND2x2_ASAP7_75t_R _30615_ (.A(_04303_),
    .B(_10213_),
    .Y(_10252_));
 AO21x1_ASAP7_75t_R _30616_ (.A1(_09753_),
    .A2(_10217_),
    .B(_10252_),
    .Y(_03274_));
 BUFx6f_ASAP7_75t_R _30617_ (.A(_09543_),
    .Y(_10253_));
 AND2x2_ASAP7_75t_R _30618_ (.A(_04433_),
    .B(_10213_),
    .Y(_10254_));
 AO21x1_ASAP7_75t_R _30619_ (.A1(_10253_),
    .A2(_10217_),
    .B(_10254_),
    .Y(_03275_));
 BUFx4f_ASAP7_75t_R _30620_ (.A(_09579_),
    .Y(_10255_));
 NAND2x1_ASAP7_75t_R _30621_ (.A(_01365_),
    .B(_10214_),
    .Y(_10256_));
 OA21x2_ASAP7_75t_R _30622_ (.A1(_10255_),
    .A2(_10214_),
    .B(_10256_),
    .Y(_03276_));
 BUFx3_ASAP7_75t_R _30623_ (.A(_09621_),
    .Y(_10257_));
 AND2x2_ASAP7_75t_R _30624_ (.A(_04657_),
    .B(_10213_),
    .Y(_10258_));
 AO21x1_ASAP7_75t_R _30625_ (.A1(net153),
    .A2(_10217_),
    .B(_10258_),
    .Y(_03277_));
 BUFx3_ASAP7_75t_R _30626_ (.A(_09647_),
    .Y(_10259_));
 AND2x2_ASAP7_75t_R _30627_ (.A(_04784_),
    .B(_10213_),
    .Y(_10260_));
 AO21x1_ASAP7_75t_R _30628_ (.A1(net9),
    .A2(_10217_),
    .B(_10260_),
    .Y(_03278_));
 NAND2x1_ASAP7_75t_R _30629_ (.A(_00890_),
    .B(_10110_),
    .Y(_10261_));
 OA21x2_ASAP7_75t_R _30630_ (.A1(_09181_),
    .A2(_10200_),
    .B(_10261_),
    .Y(_03279_));
 OR3x2_ASAP7_75t_R _30631_ (.A(_14153_),
    .B(_14303_),
    .C(_14231_),
    .Y(_10262_));
 OR3x4_ASAP7_75t_R _30632_ (.A(_08677_),
    .B(_08588_),
    .C(_10262_),
    .Y(_10263_));
 BUFx6f_ASAP7_75t_R _30633_ (.A(_10263_),
    .Y(_10264_));
 BUFx6f_ASAP7_75t_R _30634_ (.A(_10264_),
    .Y(_10265_));
 BUFx6f_ASAP7_75t_R _30635_ (.A(_10264_),
    .Y(_10266_));
 NAND2x1_ASAP7_75t_R _30636_ (.A(_00430_),
    .B(_10266_),
    .Y(_10267_));
 OA21x2_ASAP7_75t_R _30637_ (.A1(_10162_),
    .A2(_10265_),
    .B(_10267_),
    .Y(_03280_));
 NAND2x1_ASAP7_75t_R _30638_ (.A(_00383_),
    .B(_10266_),
    .Y(_10268_));
 OA21x2_ASAP7_75t_R _30639_ (.A1(_09676_),
    .A2(_10265_),
    .B(_10268_),
    .Y(_03281_));
 NAND2x1_ASAP7_75t_R _30640_ (.A(_00494_),
    .B(_10266_),
    .Y(_10269_));
 OA21x2_ASAP7_75t_R _30641_ (.A1(_10220_),
    .A2(_10265_),
    .B(_10269_),
    .Y(_03282_));
 NAND2x1_ASAP7_75t_R _30642_ (.A(_00525_),
    .B(_10266_),
    .Y(_10270_));
 OA21x2_ASAP7_75t_R _30643_ (.A1(_09716_),
    .A2(_10265_),
    .B(_10270_),
    .Y(_03283_));
 AND3x4_ASAP7_75t_R _30644_ (.A(_14049_),
    .B(_14050_),
    .C(_14232_),
    .Y(_10271_));
 AND4x2_ASAP7_75t_R _30645_ (.A(_08593_),
    .B(_08594_),
    .C(_08339_),
    .D(_10271_),
    .Y(_10272_));
 BUFx6f_ASAP7_75t_R _30646_ (.A(_10272_),
    .Y(_10273_));
 NOR2x1_ASAP7_75t_R _30647_ (.A(_00555_),
    .B(_10273_),
    .Y(_10274_));
 AO21x1_ASAP7_75t_R _30648_ (.A1(_10175_),
    .A2(_10273_),
    .B(_10274_),
    .Y(_03284_));
 BUFx12f_ASAP7_75t_R _30649_ (.A(_10264_),
    .Y(_10275_));
 NAND2x1_ASAP7_75t_R _30650_ (.A(_00587_),
    .B(_10275_),
    .Y(_10276_));
 OA21x2_ASAP7_75t_R _30651_ (.A1(_10177_),
    .A2(_10265_),
    .B(_10276_),
    .Y(_03285_));
 NAND2x1_ASAP7_75t_R _30652_ (.A(_00617_),
    .B(_10275_),
    .Y(_10277_));
 OA21x2_ASAP7_75t_R _30653_ (.A1(_08810_),
    .A2(_10265_),
    .B(_10277_),
    .Y(_03286_));
 NAND2x1_ASAP7_75t_R _30654_ (.A(_00647_),
    .B(_10275_),
    .Y(_10278_));
 OA21x2_ASAP7_75t_R _30655_ (.A1(_08851_),
    .A2(_10265_),
    .B(_10278_),
    .Y(_03287_));
 BUFx10_ASAP7_75t_R _30656_ (.A(_08897_),
    .Y(_10279_));
 OR2x2_ASAP7_75t_R _30657_ (.A(_00677_),
    .B(_10272_),
    .Y(_10280_));
 OAI21x1_ASAP7_75t_R _30658_ (.A1(_10279_),
    .A2(_10265_),
    .B(_10280_),
    .Y(_03288_));
 NAND2x1_ASAP7_75t_R _30659_ (.A(_00707_),
    .B(_10275_),
    .Y(_10281_));
 OA21x2_ASAP7_75t_R _30660_ (.A1(_08943_),
    .A2(_10265_),
    .B(_10281_),
    .Y(_03289_));
 NOR2x1_ASAP7_75t_R _30661_ (.A(_00923_),
    .B(_10098_),
    .Y(_10282_));
 AO21x1_ASAP7_75t_R _30662_ (.A1(_10238_),
    .A2(_10098_),
    .B(_10282_),
    .Y(_03290_));
 NAND2x1_ASAP7_75t_R _30663_ (.A(_00737_),
    .B(_10275_),
    .Y(_10283_));
 OA21x2_ASAP7_75t_R _30664_ (.A1(_08989_),
    .A2(_10265_),
    .B(_10283_),
    .Y(_03291_));
 BUFx6f_ASAP7_75t_R _30665_ (.A(_10264_),
    .Y(_10284_));
 NAND2x1_ASAP7_75t_R _30666_ (.A(_00767_),
    .B(_10275_),
    .Y(_10285_));
 OA21x2_ASAP7_75t_R _30667_ (.A1(_09728_),
    .A2(_10284_),
    .B(_10285_),
    .Y(_03292_));
 NAND2x1_ASAP7_75t_R _30668_ (.A(_00463_),
    .B(_10275_),
    .Y(_10286_));
 OA21x2_ASAP7_75t_R _30669_ (.A1(_09074_),
    .A2(_10284_),
    .B(_10286_),
    .Y(_03293_));
 NAND2x1_ASAP7_75t_R _30670_ (.A(_00838_),
    .B(_10275_),
    .Y(_10287_));
 OA21x2_ASAP7_75t_R _30671_ (.A1(_09104_),
    .A2(_10284_),
    .B(_10287_),
    .Y(_03294_));
 NAND2x1_ASAP7_75t_R _30672_ (.A(_00871_),
    .B(_10275_),
    .Y(_10288_));
 OA21x2_ASAP7_75t_R _30673_ (.A1(_09144_),
    .A2(_10284_),
    .B(_10288_),
    .Y(_03295_));
 NAND2x1_ASAP7_75t_R _30674_ (.A(_00904_),
    .B(_10275_),
    .Y(_10289_));
 OA21x2_ASAP7_75t_R _30675_ (.A1(_09181_),
    .A2(_10284_),
    .B(_10289_),
    .Y(_03296_));
 NOR2x1_ASAP7_75t_R _30676_ (.A(_00937_),
    .B(_10273_),
    .Y(_10290_));
 AO21x1_ASAP7_75t_R _30677_ (.A1(_10238_),
    .A2(_10273_),
    .B(_10290_),
    .Y(_03297_));
 BUFx6f_ASAP7_75t_R _30678_ (.A(_10264_),
    .Y(_10291_));
 NAND2x1_ASAP7_75t_R _30679_ (.A(_00970_),
    .B(_10291_),
    .Y(_10292_));
 OA21x2_ASAP7_75t_R _30680_ (.A1(_09245_),
    .A2(_10284_),
    .B(_10292_),
    .Y(_03298_));
 NAND2x1_ASAP7_75t_R _30681_ (.A(_01003_),
    .B(_10291_),
    .Y(_10293_));
 OA21x2_ASAP7_75t_R _30682_ (.A1(_09271_),
    .A2(_10284_),
    .B(_10293_),
    .Y(_03299_));
 NAND2x1_ASAP7_75t_R _30683_ (.A(_01036_),
    .B(_10291_),
    .Y(_10294_));
 OA21x2_ASAP7_75t_R _30684_ (.A1(_09299_),
    .A2(_10284_),
    .B(_10294_),
    .Y(_03300_));
 BUFx6f_ASAP7_75t_R _30685_ (.A(_10037_),
    .Y(_10295_));
 NAND2x1_ASAP7_75t_R _30686_ (.A(_00956_),
    .B(_10295_),
    .Y(_10296_));
 OA21x2_ASAP7_75t_R _30687_ (.A1(_09245_),
    .A2(_10200_),
    .B(_10296_),
    .Y(_03301_));
 NOR2x1_ASAP7_75t_R _30688_ (.A(_01788_),
    .B(_09796_),
    .Y(_10297_));
 AO21x1_ASAP7_75t_R _30689_ (.A1(_09794_),
    .A2(_08675_),
    .B(_10297_),
    .Y(_03302_));
 NAND2x1_ASAP7_75t_R _30690_ (.A(_01069_),
    .B(_10291_),
    .Y(_10298_));
 OA21x2_ASAP7_75t_R _30691_ (.A1(_09328_),
    .A2(_10284_),
    .B(_10298_),
    .Y(_03303_));
 NAND2x1_ASAP7_75t_R _30692_ (.A(_01102_),
    .B(_10291_),
    .Y(_10299_));
 OA21x2_ASAP7_75t_R _30693_ (.A1(_09357_),
    .A2(_10284_),
    .B(_10299_),
    .Y(_03304_));
 NAND2x1_ASAP7_75t_R _30694_ (.A(_01135_),
    .B(_10291_),
    .Y(_10300_));
 OA21x2_ASAP7_75t_R _30695_ (.A1(_09390_),
    .A2(_10266_),
    .B(_10300_),
    .Y(_03305_));
 NAND2x1_ASAP7_75t_R _30696_ (.A(_01168_),
    .B(_10291_),
    .Y(_10301_));
 OA21x2_ASAP7_75t_R _30697_ (.A1(_09416_),
    .A2(_10266_),
    .B(_10301_),
    .Y(_03306_));
 NAND2x1_ASAP7_75t_R _30698_ (.A(_01201_),
    .B(_10291_),
    .Y(_10302_));
 OA21x2_ASAP7_75t_R _30699_ (.A1(_10248_),
    .A2(_10266_),
    .B(_10302_),
    .Y(_03307_));
 NAND2x1_ASAP7_75t_R _30700_ (.A(_01234_),
    .B(_10291_),
    .Y(_10303_));
 OA21x2_ASAP7_75t_R _30701_ (.A1(_09472_),
    .A2(_10266_),
    .B(_10303_),
    .Y(_03308_));
 NAND2x1_ASAP7_75t_R _30702_ (.A(_01267_),
    .B(_10291_),
    .Y(_10304_));
 OA21x2_ASAP7_75t_R _30703_ (.A1(_09495_),
    .A2(_10266_),
    .B(_10304_),
    .Y(_03309_));
 BUFx3_ASAP7_75t_R _30704_ (.A(_09512_),
    .Y(_10305_));
 NOR2x1_ASAP7_75t_R _30705_ (.A(_01300_),
    .B(_10273_),
    .Y(_10306_));
 AO21x1_ASAP7_75t_R _30706_ (.A1(_10305_),
    .A2(_10273_),
    .B(_10306_),
    .Y(_03310_));
 NOR2x1_ASAP7_75t_R _30707_ (.A(_01333_),
    .B(_10273_),
    .Y(_10307_));
 AO21x1_ASAP7_75t_R _30708_ (.A1(_10253_),
    .A2(_10273_),
    .B(_10307_),
    .Y(_03311_));
 NAND2x1_ASAP7_75t_R _30709_ (.A(_01366_),
    .B(_10264_),
    .Y(_10308_));
 OA21x2_ASAP7_75t_R _30710_ (.A1(_10255_),
    .A2(_10266_),
    .B(_10308_),
    .Y(_03312_));
 NAND2x1_ASAP7_75t_R _30711_ (.A(_00989_),
    .B(_10295_),
    .Y(_10309_));
 OA21x2_ASAP7_75t_R _30712_ (.A1(_09271_),
    .A2(_10200_),
    .B(_10309_),
    .Y(_03313_));
 NOR2x1_ASAP7_75t_R _30713_ (.A(_01399_),
    .B(_10272_),
    .Y(_10310_));
 AO21x1_ASAP7_75t_R _30714_ (.A1(_10257_),
    .A2(_10273_),
    .B(_10310_),
    .Y(_03314_));
 NOR2x1_ASAP7_75t_R _30715_ (.A(_01432_),
    .B(_10272_),
    .Y(_10311_));
 AO21x1_ASAP7_75t_R _30716_ (.A1(_10259_),
    .A2(_10273_),
    .B(_10311_),
    .Y(_03315_));
 NAND2x2_ASAP7_75t_R _30717_ (.A(_08341_),
    .B(_10271_),
    .Y(_10312_));
 OR3x4_ASAP7_75t_R _30718_ (.A(_08588_),
    .B(_08589_),
    .C(_10262_),
    .Y(_10313_));
 BUFx12_ASAP7_75t_R _30719_ (.A(_10313_),
    .Y(_10314_));
 NAND2x1_ASAP7_75t_R _30720_ (.A(_00431_),
    .B(_10314_),
    .Y(_10315_));
 OA21x2_ASAP7_75t_R _30721_ (.A1(_10162_),
    .A2(_10312_),
    .B(_10315_),
    .Y(_03316_));
 BUFx12f_ASAP7_75t_R _30722_ (.A(_10313_),
    .Y(_10316_));
 BUFx6f_ASAP7_75t_R _30723_ (.A(_10316_),
    .Y(_10317_));
 NAND2x1_ASAP7_75t_R _30724_ (.A(_00384_),
    .B(_10314_),
    .Y(_10318_));
 OA21x2_ASAP7_75t_R _30725_ (.A1(_09676_),
    .A2(_10317_),
    .B(_10318_),
    .Y(_03317_));
 NAND2x1_ASAP7_75t_R _30726_ (.A(_00495_),
    .B(_10314_),
    .Y(_10319_));
 OA21x2_ASAP7_75t_R _30727_ (.A1(_10220_),
    .A2(_10317_),
    .B(_10319_),
    .Y(_03318_));
 NAND2x1_ASAP7_75t_R _30728_ (.A(_00526_),
    .B(_10314_),
    .Y(_10320_));
 OA21x2_ASAP7_75t_R _30729_ (.A1(_09716_),
    .A2(_10317_),
    .B(_10320_),
    .Y(_03319_));
 AND2x4_ASAP7_75t_R _30730_ (.A(_08341_),
    .B(_10271_),
    .Y(_10321_));
 AND3x1_ASAP7_75t_R _30731_ (.A(_08595_),
    .B(_09651_),
    .C(_10271_),
    .Y(_10322_));
 BUFx6f_ASAP7_75t_R _30732_ (.A(_10322_),
    .Y(_10323_));
 NOR2x1_ASAP7_75t_R _30733_ (.A(_00556_),
    .B(_10323_),
    .Y(_10324_));
 AO21x1_ASAP7_75t_R _30734_ (.A1(_10175_),
    .A2(_10321_),
    .B(_10324_),
    .Y(_03320_));
 NAND2x1_ASAP7_75t_R _30735_ (.A(_00588_),
    .B(_10314_),
    .Y(_10325_));
 OA21x2_ASAP7_75t_R _30736_ (.A1(_10177_),
    .A2(_10317_),
    .B(_10325_),
    .Y(_03321_));
 NAND2x1_ASAP7_75t_R _30737_ (.A(_00618_),
    .B(_10314_),
    .Y(_10326_));
 OA21x2_ASAP7_75t_R _30738_ (.A1(_08810_),
    .A2(_10317_),
    .B(_10326_),
    .Y(_03322_));
 BUFx12f_ASAP7_75t_R _30739_ (.A(_10313_),
    .Y(_10327_));
 NAND2x1_ASAP7_75t_R _30740_ (.A(_00648_),
    .B(_10327_),
    .Y(_10328_));
 OA21x2_ASAP7_75t_R _30741_ (.A1(_08851_),
    .A2(_10317_),
    .B(_10328_),
    .Y(_03323_));
 NAND2x1_ASAP7_75t_R _30742_ (.A(_01022_),
    .B(_10295_),
    .Y(_10329_));
 OA21x2_ASAP7_75t_R _30743_ (.A1(_09299_),
    .A2(_10200_),
    .B(_10329_),
    .Y(_03324_));
 OR2x2_ASAP7_75t_R _30744_ (.A(_00678_),
    .B(_10323_),
    .Y(_10330_));
 OAI21x1_ASAP7_75t_R _30745_ (.A1(_10279_),
    .A2(_10312_),
    .B(_10330_),
    .Y(_03325_));
 NAND2x1_ASAP7_75t_R _30746_ (.A(_00708_),
    .B(_10327_),
    .Y(_10331_));
 OA21x2_ASAP7_75t_R _30747_ (.A1(_08943_),
    .A2(_10317_),
    .B(_10331_),
    .Y(_03326_));
 NAND2x1_ASAP7_75t_R _30748_ (.A(_00738_),
    .B(_10327_),
    .Y(_10332_));
 OA21x2_ASAP7_75t_R _30749_ (.A1(_08989_),
    .A2(_10317_),
    .B(_10332_),
    .Y(_03327_));
 NAND2x1_ASAP7_75t_R _30750_ (.A(_00768_),
    .B(_10327_),
    .Y(_10333_));
 OA21x2_ASAP7_75t_R _30751_ (.A1(_09728_),
    .A2(_10317_),
    .B(_10333_),
    .Y(_03328_));
 NAND2x1_ASAP7_75t_R _30752_ (.A(_00464_),
    .B(_10327_),
    .Y(_10334_));
 OA21x2_ASAP7_75t_R _30753_ (.A1(_09074_),
    .A2(_10317_),
    .B(_10334_),
    .Y(_03329_));
 BUFx6f_ASAP7_75t_R _30754_ (.A(_10313_),
    .Y(_10335_));
 NAND2x1_ASAP7_75t_R _30755_ (.A(_00839_),
    .B(_10327_),
    .Y(_10336_));
 OA21x2_ASAP7_75t_R _30756_ (.A1(_09104_),
    .A2(_10335_),
    .B(_10336_),
    .Y(_03330_));
 NAND2x1_ASAP7_75t_R _30757_ (.A(_00872_),
    .B(_10327_),
    .Y(_10337_));
 OA21x2_ASAP7_75t_R _30758_ (.A1(_09144_),
    .A2(_10335_),
    .B(_10337_),
    .Y(_03331_));
 NAND2x1_ASAP7_75t_R _30759_ (.A(_00905_),
    .B(_10327_),
    .Y(_10338_));
 OA21x2_ASAP7_75t_R _30760_ (.A1(_09181_),
    .A2(_10335_),
    .B(_10338_),
    .Y(_03332_));
 NOR2x1_ASAP7_75t_R _30761_ (.A(_00938_),
    .B(_10323_),
    .Y(_10339_));
 AO21x1_ASAP7_75t_R _30762_ (.A1(_10238_),
    .A2(_10321_),
    .B(_10339_),
    .Y(_03333_));
 NAND2x1_ASAP7_75t_R _30763_ (.A(_00971_),
    .B(_10327_),
    .Y(_10340_));
 OA21x2_ASAP7_75t_R _30764_ (.A1(_09245_),
    .A2(_10335_),
    .B(_10340_),
    .Y(_03334_));
 NAND2x1_ASAP7_75t_R _30765_ (.A(_01055_),
    .B(_10295_),
    .Y(_10341_));
 OA21x2_ASAP7_75t_R _30766_ (.A1(_09328_),
    .A2(_10200_),
    .B(_10341_),
    .Y(_03335_));
 NAND2x1_ASAP7_75t_R _30767_ (.A(_01004_),
    .B(_10327_),
    .Y(_10342_));
 OA21x2_ASAP7_75t_R _30768_ (.A1(_09271_),
    .A2(_10335_),
    .B(_10342_),
    .Y(_03336_));
 NAND2x1_ASAP7_75t_R _30769_ (.A(_01037_),
    .B(_10316_),
    .Y(_10343_));
 OA21x2_ASAP7_75t_R _30770_ (.A1(_09299_),
    .A2(_10335_),
    .B(_10343_),
    .Y(_03337_));
 NAND2x1_ASAP7_75t_R _30771_ (.A(_01070_),
    .B(_10316_),
    .Y(_10344_));
 OA21x2_ASAP7_75t_R _30772_ (.A1(_09328_),
    .A2(_10335_),
    .B(_10344_),
    .Y(_03338_));
 NAND2x1_ASAP7_75t_R _30773_ (.A(_01103_),
    .B(_10316_),
    .Y(_10345_));
 OA21x2_ASAP7_75t_R _30774_ (.A1(_09357_),
    .A2(_10335_),
    .B(_10345_),
    .Y(_03339_));
 NAND2x1_ASAP7_75t_R _30775_ (.A(_01136_),
    .B(_10316_),
    .Y(_10346_));
 OA21x2_ASAP7_75t_R _30776_ (.A1(_09390_),
    .A2(_10335_),
    .B(_10346_),
    .Y(_03340_));
 NAND2x1_ASAP7_75t_R _30777_ (.A(_01169_),
    .B(_10316_),
    .Y(_10347_));
 OA21x2_ASAP7_75t_R _30778_ (.A1(_09416_),
    .A2(_10335_),
    .B(_10347_),
    .Y(_03341_));
 NAND2x1_ASAP7_75t_R _30779_ (.A(_01202_),
    .B(_10316_),
    .Y(_10348_));
 OA21x2_ASAP7_75t_R _30780_ (.A1(_10248_),
    .A2(_10314_),
    .B(_10348_),
    .Y(_03342_));
 NAND2x1_ASAP7_75t_R _30781_ (.A(_01235_),
    .B(_10316_),
    .Y(_10349_));
 OA21x2_ASAP7_75t_R _30782_ (.A1(_09472_),
    .A2(_10314_),
    .B(_10349_),
    .Y(_03343_));
 NAND2x1_ASAP7_75t_R _30783_ (.A(_01268_),
    .B(_10316_),
    .Y(_10350_));
 OA21x2_ASAP7_75t_R _30784_ (.A1(_09495_),
    .A2(_10314_),
    .B(_10350_),
    .Y(_03344_));
 NOR2x1_ASAP7_75t_R _30785_ (.A(_01301_),
    .B(_10323_),
    .Y(_10351_));
 AO21x1_ASAP7_75t_R _30786_ (.A1(_10305_),
    .A2(_10321_),
    .B(_10351_),
    .Y(_03345_));
 NAND2x1_ASAP7_75t_R _30787_ (.A(_01088_),
    .B(_10295_),
    .Y(_10352_));
 OA21x2_ASAP7_75t_R _30788_ (.A1(_09357_),
    .A2(_10200_),
    .B(_10352_),
    .Y(_03346_));
 NOR2x1_ASAP7_75t_R _30789_ (.A(_01334_),
    .B(_10323_),
    .Y(_10353_));
 AO21x1_ASAP7_75t_R _30790_ (.A1(_10253_),
    .A2(_10321_),
    .B(_10353_),
    .Y(_03347_));
 NAND2x1_ASAP7_75t_R _30791_ (.A(_01367_),
    .B(_10316_),
    .Y(_10354_));
 OA21x2_ASAP7_75t_R _30792_ (.A1(_10255_),
    .A2(_10314_),
    .B(_10354_),
    .Y(_03348_));
 NOR2x1_ASAP7_75t_R _30793_ (.A(_01400_),
    .B(_10323_),
    .Y(_10355_));
 AO21x1_ASAP7_75t_R _30794_ (.A1(net153),
    .A2(_10321_),
    .B(_10355_),
    .Y(_03349_));
 NOR2x1_ASAP7_75t_R _30795_ (.A(_01433_),
    .B(_10323_),
    .Y(_10356_));
 AO21x1_ASAP7_75t_R _30796_ (.A1(net9),
    .A2(_10321_),
    .B(_10356_),
    .Y(_03350_));
 OR3x1_ASAP7_75t_R _30797_ (.A(_09766_),
    .B(_09767_),
    .C(_10262_),
    .Y(_10357_));
 BUFx10_ASAP7_75t_R _30798_ (.A(_10357_),
    .Y(_10358_));
 BUFx6f_ASAP7_75t_R _30799_ (.A(_10358_),
    .Y(_10359_));
 NAND2x1_ASAP7_75t_R _30800_ (.A(_00432_),
    .B(_10359_),
    .Y(_10360_));
 OA21x2_ASAP7_75t_R _30801_ (.A1(_10162_),
    .A2(_10359_),
    .B(_10360_),
    .Y(_03351_));
 BUFx6f_ASAP7_75t_R _30802_ (.A(_09675_),
    .Y(_10361_));
 AND3x1_ASAP7_75t_R _30803_ (.A(_08339_),
    .B(_09774_),
    .C(_10271_),
    .Y(_10362_));
 BUFx6f_ASAP7_75t_R _30804_ (.A(_10362_),
    .Y(_10363_));
 BUFx6f_ASAP7_75t_R _30805_ (.A(_10363_),
    .Y(_10364_));
 BUFx6f_ASAP7_75t_R _30806_ (.A(_10358_),
    .Y(_10365_));
 AND2x2_ASAP7_75t_R _30807_ (.A(_13544_),
    .B(_10365_),
    .Y(_10366_));
 AO21x1_ASAP7_75t_R _30808_ (.A1(_10361_),
    .A2(_10364_),
    .B(_10366_),
    .Y(_03352_));
 NAND2x1_ASAP7_75t_R _30809_ (.A(_00496_),
    .B(_10359_),
    .Y(_10367_));
 OA21x2_ASAP7_75t_R _30810_ (.A1(_10220_),
    .A2(_10359_),
    .B(_10367_),
    .Y(_03353_));
 BUFx4f_ASAP7_75t_R _30811_ (.A(_09715_),
    .Y(_10368_));
 AND2x2_ASAP7_75t_R _30812_ (.A(_14165_),
    .B(_10365_),
    .Y(_10369_));
 AO21x1_ASAP7_75t_R _30813_ (.A1(_10368_),
    .A2(_10364_),
    .B(_10369_),
    .Y(_03354_));
 AND2x2_ASAP7_75t_R _30814_ (.A(_14256_),
    .B(_10365_),
    .Y(_10370_));
 AO21x1_ASAP7_75t_R _30815_ (.A1(_10175_),
    .A2(_10364_),
    .B(_10370_),
    .Y(_03355_));
 NAND2x1_ASAP7_75t_R _30816_ (.A(_00589_),
    .B(_10359_),
    .Y(_10371_));
 OA21x2_ASAP7_75t_R _30817_ (.A1(_10177_),
    .A2(_10359_),
    .B(_10371_),
    .Y(_03356_));
 NAND2x1_ASAP7_75t_R _30818_ (.A(_01121_),
    .B(_10295_),
    .Y(_10372_));
 OA21x2_ASAP7_75t_R _30819_ (.A1(_09390_),
    .A2(_10039_),
    .B(_10372_),
    .Y(_03357_));
 BUFx4f_ASAP7_75t_R _30820_ (.A(_08809_),
    .Y(_10373_));
 AND2x2_ASAP7_75t_R _30821_ (.A(_14381_),
    .B(_10365_),
    .Y(_10374_));
 AO21x1_ASAP7_75t_R _30822_ (.A1(_10373_),
    .A2(_10364_),
    .B(_10374_),
    .Y(_03358_));
 BUFx4f_ASAP7_75t_R _30823_ (.A(_08850_),
    .Y(_10375_));
 AND2x2_ASAP7_75t_R _30824_ (.A(_14437_),
    .B(_10365_),
    .Y(_10376_));
 AO21x1_ASAP7_75t_R _30825_ (.A1(_10375_),
    .A2(_10364_),
    .B(_10376_),
    .Y(_03359_));
 OR3x1_ASAP7_75t_R _30826_ (.A(_09790_),
    .B(_09791_),
    .C(_10365_),
    .Y(_10377_));
 OAI21x1_ASAP7_75t_R _30827_ (.A1(_00679_),
    .A2(_10364_),
    .B(_10377_),
    .Y(_03360_));
 AND2x2_ASAP7_75t_R _30828_ (.A(_14555_),
    .B(_10365_),
    .Y(_10378_));
 AO21x1_ASAP7_75t_R _30829_ (.A1(_09855_),
    .A2(_10364_),
    .B(_10378_),
    .Y(_03361_));
 BUFx4f_ASAP7_75t_R _30830_ (.A(_08988_),
    .Y(_10379_));
 AND2x2_ASAP7_75t_R _30831_ (.A(_14661_),
    .B(_10365_),
    .Y(_10380_));
 AO21x1_ASAP7_75t_R _30832_ (.A1(_10379_),
    .A2(_10364_),
    .B(_10380_),
    .Y(_03362_));
 BUFx6f_ASAP7_75t_R _30833_ (.A(_09036_),
    .Y(_10381_));
 BUFx6f_ASAP7_75t_R _30834_ (.A(_10358_),
    .Y(_10382_));
 AND2x2_ASAP7_75t_R _30835_ (.A(_14714_),
    .B(_10382_),
    .Y(_10383_));
 AO21x1_ASAP7_75t_R _30836_ (.A1(_10381_),
    .A2(_10364_),
    .B(_10383_),
    .Y(_03363_));
 BUFx4f_ASAP7_75t_R _30837_ (.A(_09073_),
    .Y(_10384_));
 BUFx6f_ASAP7_75t_R _30838_ (.A(_10363_),
    .Y(_10385_));
 AND2x2_ASAP7_75t_R _30839_ (.A(_13957_),
    .B(_10382_),
    .Y(_10386_));
 AO21x1_ASAP7_75t_R _30840_ (.A1(_10384_),
    .A2(_10385_),
    .B(_10386_),
    .Y(_03364_));
 BUFx6f_ASAP7_75t_R _30841_ (.A(_09103_),
    .Y(_10387_));
 AND2x2_ASAP7_75t_R _30842_ (.A(_15664_),
    .B(_10382_),
    .Y(_10388_));
 AO21x1_ASAP7_75t_R _30843_ (.A1(_10387_),
    .A2(_10385_),
    .B(_10388_),
    .Y(_03365_));
 BUFx4f_ASAP7_75t_R _30844_ (.A(_09143_),
    .Y(_10389_));
 AND2x2_ASAP7_75t_R _30845_ (.A(_15809_),
    .B(_10382_),
    .Y(_10390_));
 AO21x1_ASAP7_75t_R _30846_ (.A1(_10389_),
    .A2(_10385_),
    .B(_10390_),
    .Y(_03366_));
 BUFx4f_ASAP7_75t_R _30847_ (.A(_09180_),
    .Y(_10391_));
 AND2x2_ASAP7_75t_R _30848_ (.A(_15943_),
    .B(_10382_),
    .Y(_10392_));
 AO21x1_ASAP7_75t_R _30849_ (.A1(_10391_),
    .A2(_10385_),
    .B(_10392_),
    .Y(_03367_));
 NAND2x1_ASAP7_75t_R _30850_ (.A(_01154_),
    .B(_10295_),
    .Y(_10393_));
 OA21x2_ASAP7_75t_R _30851_ (.A1(_09416_),
    .A2(_10039_),
    .B(_10393_),
    .Y(_03368_));
 AND3x1_ASAP7_75t_R _30852_ (.A(_09204_),
    .B(_09212_),
    .C(_10363_),
    .Y(_10394_));
 AO21x1_ASAP7_75t_R _30853_ (.A1(_16088_),
    .A2(_10359_),
    .B(_10394_),
    .Y(_03369_));
 BUFx4f_ASAP7_75t_R _30854_ (.A(_09244_),
    .Y(_10395_));
 AND2x2_ASAP7_75t_R _30855_ (.A(_16203_),
    .B(_10382_),
    .Y(_10396_));
 AO21x1_ASAP7_75t_R _30856_ (.A1(_10395_),
    .A2(_10385_),
    .B(_10396_),
    .Y(_03370_));
 BUFx4f_ASAP7_75t_R _30857_ (.A(_09270_),
    .Y(_10397_));
 AND2x2_ASAP7_75t_R _30858_ (.A(_16348_),
    .B(_10382_),
    .Y(_10398_));
 AO21x1_ASAP7_75t_R _30859_ (.A1(_10397_),
    .A2(_10385_),
    .B(_10398_),
    .Y(_03371_));
 BUFx4f_ASAP7_75t_R _30860_ (.A(_09298_),
    .Y(_10399_));
 AND2x2_ASAP7_75t_R _30861_ (.A(_16460_),
    .B(_10382_),
    .Y(_10400_));
 AO21x1_ASAP7_75t_R _30862_ (.A1(_10399_),
    .A2(_10385_),
    .B(_10400_),
    .Y(_03372_));
 BUFx4f_ASAP7_75t_R _30863_ (.A(_09327_),
    .Y(_10401_));
 AND2x2_ASAP7_75t_R _30864_ (.A(_16586_),
    .B(_10382_),
    .Y(_10402_));
 AO21x1_ASAP7_75t_R _30865_ (.A1(_10401_),
    .A2(_10385_),
    .B(_10402_),
    .Y(_03373_));
 BUFx4f_ASAP7_75t_R _30866_ (.A(_09356_),
    .Y(_10403_));
 AND2x2_ASAP7_75t_R _30867_ (.A(_16700_),
    .B(_10382_),
    .Y(_10404_));
 AO21x1_ASAP7_75t_R _30868_ (.A1(_10403_),
    .A2(_10385_),
    .B(_10404_),
    .Y(_03374_));
 AND2x2_ASAP7_75t_R _30869_ (.A(_16830_),
    .B(_10358_),
    .Y(_10405_));
 AO21x1_ASAP7_75t_R _30870_ (.A1(_09819_),
    .A2(_10385_),
    .B(_10405_),
    .Y(_03375_));
 BUFx4f_ASAP7_75t_R _30871_ (.A(_09415_),
    .Y(_10406_));
 AND2x2_ASAP7_75t_R _30872_ (.A(_16940_),
    .B(_10358_),
    .Y(_10407_));
 AO21x1_ASAP7_75t_R _30873_ (.A1(_10406_),
    .A2(_10363_),
    .B(_10407_),
    .Y(_03376_));
 NAND2x1_ASAP7_75t_R _30874_ (.A(_01203_),
    .B(_10365_),
    .Y(_10408_));
 OA21x2_ASAP7_75t_R _30875_ (.A1(_10248_),
    .A2(_10359_),
    .B(_10408_),
    .Y(_03377_));
 BUFx3_ASAP7_75t_R _30876_ (.A(_09471_),
    .Y(_10409_));
 AND2x2_ASAP7_75t_R _30877_ (.A(_17179_),
    .B(_10358_),
    .Y(_10410_));
 AO21x1_ASAP7_75t_R _30878_ (.A1(_10409_),
    .A2(_10363_),
    .B(_10410_),
    .Y(_03378_));
 NAND2x1_ASAP7_75t_R _30879_ (.A(_01187_),
    .B(_10295_),
    .Y(_10411_));
 OA21x2_ASAP7_75t_R _30880_ (.A1(_10248_),
    .A2(_10039_),
    .B(_10411_),
    .Y(_03379_));
 BUFx4f_ASAP7_75t_R _30881_ (.A(_09494_),
    .Y(_10412_));
 AND2x2_ASAP7_75t_R _30882_ (.A(_17310_),
    .B(_10358_),
    .Y(_10413_));
 AO21x1_ASAP7_75t_R _30883_ (.A1(_10412_),
    .A2(_10363_),
    .B(_10413_),
    .Y(_03380_));
 AND3x1_ASAP7_75t_R _30884_ (.A(_09508_),
    .B(_09511_),
    .C(_10363_),
    .Y(_10414_));
 AO21x1_ASAP7_75t_R _30885_ (.A1(_04337_),
    .A2(_10359_),
    .B(_10414_),
    .Y(_03381_));
 AND3x1_ASAP7_75t_R _30886_ (.A(_09539_),
    .B(_09542_),
    .C(_10363_),
    .Y(_10415_));
 AO21x1_ASAP7_75t_R _30887_ (.A1(_04467_),
    .A2(_10359_),
    .B(_10415_),
    .Y(_03382_));
 OR3x1_ASAP7_75t_R _30888_ (.A(_09578_),
    .B(_09572_),
    .C(_10365_),
    .Y(_10416_));
 OA21x2_ASAP7_75t_R _30889_ (.A1(_04577_),
    .A2(_10364_),
    .B(_10416_),
    .Y(_03383_));
 AND2x2_ASAP7_75t_R _30890_ (.A(_04691_),
    .B(_10358_),
    .Y(_10417_));
 AO21x1_ASAP7_75t_R _30891_ (.A1(net153),
    .A2(_10363_),
    .B(_10417_),
    .Y(_03384_));
 AND2x2_ASAP7_75t_R _30892_ (.A(_04756_),
    .B(_10358_),
    .Y(_10418_));
 AO21x1_ASAP7_75t_R _30893_ (.A1(net9),
    .A2(_10363_),
    .B(_10418_),
    .Y(_03385_));
 AND4x2_ASAP7_75t_R _30894_ (.A(_08329_),
    .B(_09773_),
    .C(_09834_),
    .D(_10271_),
    .Y(_10419_));
 BUFx16f_ASAP7_75t_R _30895_ (.A(_10419_),
    .Y(_10420_));
 INVx1_ASAP7_75t_R _30896_ (.A(_10420_),
    .Y(_10421_));
 OR4x2_ASAP7_75t_R _30897_ (.A(_08593_),
    .B(_08594_),
    .C(_09838_),
    .D(_10262_),
    .Y(_10422_));
 BUFx10_ASAP7_75t_R _30898_ (.A(_10422_),
    .Y(_10423_));
 NAND2x1_ASAP7_75t_R _30899_ (.A(_00433_),
    .B(_10423_),
    .Y(_10424_));
 OA21x2_ASAP7_75t_R _30900_ (.A1(_10162_),
    .A2(_10421_),
    .B(_10424_),
    .Y(_03386_));
 BUFx6f_ASAP7_75t_R _30901_ (.A(_10420_),
    .Y(_10425_));
 BUFx10_ASAP7_75t_R _30902_ (.A(_10419_),
    .Y(_10426_));
 NOR2x1_ASAP7_75t_R _30903_ (.A(_00386_),
    .B(_10426_),
    .Y(_10427_));
 AO21x1_ASAP7_75t_R _30904_ (.A1(_10361_),
    .A2(_10425_),
    .B(_10427_),
    .Y(_03387_));
 NAND2x1_ASAP7_75t_R _30905_ (.A(_00497_),
    .B(_10423_),
    .Y(_10428_));
 OA21x2_ASAP7_75t_R _30906_ (.A1(_10220_),
    .A2(_10423_),
    .B(_10428_),
    .Y(_03388_));
 NOR2x1_ASAP7_75t_R _30907_ (.A(_00528_),
    .B(_10426_),
    .Y(_10429_));
 AO21x1_ASAP7_75t_R _30908_ (.A1(_10368_),
    .A2(_10425_),
    .B(_10429_),
    .Y(_03389_));
 NAND2x1_ASAP7_75t_R _30909_ (.A(_01220_),
    .B(_10295_),
    .Y(_10430_));
 OA21x2_ASAP7_75t_R _30910_ (.A1(_09472_),
    .A2(_10039_),
    .B(_10430_),
    .Y(_03390_));
 AND2x2_ASAP7_75t_R _30911_ (.A(_14253_),
    .B(_10422_),
    .Y(_10431_));
 AO21x1_ASAP7_75t_R _30912_ (.A1(_10175_),
    .A2(_10425_),
    .B(_10431_),
    .Y(_03391_));
 NAND2x1_ASAP7_75t_R _30913_ (.A(_00590_),
    .B(_10423_),
    .Y(_10432_));
 OA21x2_ASAP7_75t_R _30914_ (.A1(_10177_),
    .A2(_10423_),
    .B(_10432_),
    .Y(_03392_));
 NOR2x1_ASAP7_75t_R _30915_ (.A(_00620_),
    .B(_10426_),
    .Y(_10433_));
 AO21x1_ASAP7_75t_R _30916_ (.A1(_10373_),
    .A2(_10425_),
    .B(_10433_),
    .Y(_03393_));
 NOR2x1_ASAP7_75t_R _30917_ (.A(_00650_),
    .B(_10426_),
    .Y(_10434_));
 AO21x1_ASAP7_75t_R _30918_ (.A1(_10375_),
    .A2(_10425_),
    .B(_10434_),
    .Y(_03394_));
 NAND2x1_ASAP7_75t_R _30919_ (.A(_14492_),
    .B(_10423_),
    .Y(_10435_));
 OAI21x1_ASAP7_75t_R _30920_ (.A1(_10279_),
    .A2(_10421_),
    .B(_10435_),
    .Y(_03395_));
 BUFx4f_ASAP7_75t_R _30921_ (.A(_08942_),
    .Y(_10436_));
 BUFx12f_ASAP7_75t_R _30922_ (.A(_10420_),
    .Y(_10437_));
 NOR2x1_ASAP7_75t_R _30923_ (.A(_00710_),
    .B(_10437_),
    .Y(_10438_));
 AO21x1_ASAP7_75t_R _30924_ (.A1(_10436_),
    .A2(_10425_),
    .B(_10438_),
    .Y(_03396_));
 NOR2x1_ASAP7_75t_R _30925_ (.A(_00740_),
    .B(_10437_),
    .Y(_10439_));
 AO21x1_ASAP7_75t_R _30926_ (.A1(_10379_),
    .A2(_10425_),
    .B(_10439_),
    .Y(_03397_));
 NOR2x1_ASAP7_75t_R _30927_ (.A(_00770_),
    .B(_10437_),
    .Y(_10440_));
 AO21x1_ASAP7_75t_R _30928_ (.A1(_10381_),
    .A2(_10425_),
    .B(_10440_),
    .Y(_03398_));
 NOR2x1_ASAP7_75t_R _30929_ (.A(_00466_),
    .B(_10437_),
    .Y(_10441_));
 AO21x1_ASAP7_75t_R _30930_ (.A1(_10384_),
    .A2(_10425_),
    .B(_10441_),
    .Y(_03399_));
 NOR2x1_ASAP7_75t_R _30931_ (.A(_00841_),
    .B(_10437_),
    .Y(_10442_));
 AO21x1_ASAP7_75t_R _30932_ (.A1(_10387_),
    .A2(_10425_),
    .B(_10442_),
    .Y(_03400_));
 NAND2x1_ASAP7_75t_R _30933_ (.A(_01253_),
    .B(_10295_),
    .Y(_10443_));
 OA21x2_ASAP7_75t_R _30934_ (.A1(_09495_),
    .A2(_10039_),
    .B(_10443_),
    .Y(_03401_));
 BUFx4f_ASAP7_75t_R _30935_ (.A(_10420_),
    .Y(_10444_));
 NOR2x1_ASAP7_75t_R _30936_ (.A(_00874_),
    .B(_10437_),
    .Y(_10445_));
 AO21x1_ASAP7_75t_R _30937_ (.A1(_10389_),
    .A2(_10444_),
    .B(_10445_),
    .Y(_03402_));
 NOR2x1_ASAP7_75t_R _30938_ (.A(_00907_),
    .B(_10437_),
    .Y(_10446_));
 AO21x1_ASAP7_75t_R _30939_ (.A1(_10391_),
    .A2(_10444_),
    .B(_10446_),
    .Y(_03403_));
 AND2x2_ASAP7_75t_R _30940_ (.A(_16085_),
    .B(_10422_),
    .Y(_10447_));
 AO21x1_ASAP7_75t_R _30941_ (.A1(_10238_),
    .A2(_10444_),
    .B(_10447_),
    .Y(_03404_));
 NOR2x1_ASAP7_75t_R _30942_ (.A(_00973_),
    .B(_10437_),
    .Y(_10448_));
 AO21x1_ASAP7_75t_R _30943_ (.A1(_10395_),
    .A2(_10444_),
    .B(_10448_),
    .Y(_03405_));
 NOR2x1_ASAP7_75t_R _30944_ (.A(_01006_),
    .B(_10437_),
    .Y(_10449_));
 AO21x1_ASAP7_75t_R _30945_ (.A1(_10397_),
    .A2(_10444_),
    .B(_10449_),
    .Y(_03406_));
 NOR2x1_ASAP7_75t_R _30946_ (.A(_01039_),
    .B(_10437_),
    .Y(_10450_));
 AO21x1_ASAP7_75t_R _30947_ (.A1(_10399_),
    .A2(_10444_),
    .B(_10450_),
    .Y(_03407_));
 NOR2x1_ASAP7_75t_R _30948_ (.A(_01072_),
    .B(_10420_),
    .Y(_10451_));
 AO21x1_ASAP7_75t_R _30949_ (.A1(_10401_),
    .A2(_10444_),
    .B(_10451_),
    .Y(_03408_));
 NOR2x1_ASAP7_75t_R _30950_ (.A(_01105_),
    .B(_10420_),
    .Y(_10452_));
 AO21x1_ASAP7_75t_R _30951_ (.A1(_10403_),
    .A2(_10444_),
    .B(_10452_),
    .Y(_03409_));
 BUFx4f_ASAP7_75t_R _30952_ (.A(_09389_),
    .Y(_10453_));
 NOR2x1_ASAP7_75t_R _30953_ (.A(_01138_),
    .B(_10420_),
    .Y(_10454_));
 AO21x1_ASAP7_75t_R _30954_ (.A1(_10453_),
    .A2(_10444_),
    .B(_10454_),
    .Y(_03410_));
 NOR2x1_ASAP7_75t_R _30955_ (.A(_01171_),
    .B(_10420_),
    .Y(_10455_));
 AO21x1_ASAP7_75t_R _30956_ (.A1(_10406_),
    .A2(_10444_),
    .B(_10455_),
    .Y(_03411_));
 NOR2x1_ASAP7_75t_R _30957_ (.A(_01286_),
    .B(_10098_),
    .Y(_10456_));
 AO21x1_ASAP7_75t_R _30958_ (.A1(_10305_),
    .A2(_10098_),
    .B(_10456_),
    .Y(_03412_));
 NAND2x1_ASAP7_75t_R _30959_ (.A(_01787_),
    .B(_09106_),
    .Y(_10457_));
 OA21x2_ASAP7_75t_R _30960_ (.A1(_08591_),
    .A2(_08762_),
    .B(_10457_),
    .Y(_03413_));
 NAND2x1_ASAP7_75t_R _30961_ (.A(_01204_),
    .B(_10423_),
    .Y(_10458_));
 OA21x2_ASAP7_75t_R _30962_ (.A1(_10248_),
    .A2(_10423_),
    .B(_10458_),
    .Y(_03414_));
 NOR2x1_ASAP7_75t_R _30963_ (.A(_01237_),
    .B(_10420_),
    .Y(_10459_));
 AO21x1_ASAP7_75t_R _30964_ (.A1(_10409_),
    .A2(_10426_),
    .B(_10459_),
    .Y(_03415_));
 NOR2x1_ASAP7_75t_R _30965_ (.A(_01270_),
    .B(_10420_),
    .Y(_10460_));
 AO21x1_ASAP7_75t_R _30966_ (.A1(_10412_),
    .A2(_10426_),
    .B(_10460_),
    .Y(_03416_));
 AND2x2_ASAP7_75t_R _30967_ (.A(_04334_),
    .B(_10422_),
    .Y(_10461_));
 AO21x1_ASAP7_75t_R _30968_ (.A1(_10305_),
    .A2(_10426_),
    .B(_10461_),
    .Y(_03417_));
 AND2x2_ASAP7_75t_R _30969_ (.A(_04464_),
    .B(_10422_),
    .Y(_10462_));
 AO21x1_ASAP7_75t_R _30970_ (.A1(_10253_),
    .A2(_10426_),
    .B(_10462_),
    .Y(_03418_));
 NAND2x1_ASAP7_75t_R _30971_ (.A(_01369_),
    .B(_10423_),
    .Y(_10463_));
 OA21x2_ASAP7_75t_R _30972_ (.A1(_10255_),
    .A2(_10423_),
    .B(_10463_),
    .Y(_03419_));
 AND2x2_ASAP7_75t_R _30973_ (.A(_04688_),
    .B(_10422_),
    .Y(_10464_));
 AO21x1_ASAP7_75t_R _30974_ (.A1(_10257_),
    .A2(_10426_),
    .B(_10464_),
    .Y(_03420_));
 AND2x2_ASAP7_75t_R _30975_ (.A(_04753_),
    .B(_10422_),
    .Y(_10465_));
 AO21x1_ASAP7_75t_R _30976_ (.A1(_10259_),
    .A2(_10426_),
    .B(_10465_),
    .Y(_03421_));
 OR3x2_ASAP7_75t_R _30977_ (.A(_14049_),
    .B(_14303_),
    .C(_14231_),
    .Y(_10466_));
 OR3x1_ASAP7_75t_R _30978_ (.A(_08677_),
    .B(_08588_),
    .C(_10466_),
    .Y(_10467_));
 BUFx6f_ASAP7_75t_R _30979_ (.A(_10467_),
    .Y(_10468_));
 BUFx6f_ASAP7_75t_R _30980_ (.A(_10468_),
    .Y(_10469_));
 BUFx10_ASAP7_75t_R _30981_ (.A(_10468_),
    .Y(_10470_));
 NAND2x1_ASAP7_75t_R _30982_ (.A(_00434_),
    .B(_10470_),
    .Y(_10471_));
 OA21x2_ASAP7_75t_R _30983_ (.A1(_10162_),
    .A2(_10469_),
    .B(_10471_),
    .Y(_03422_));
 NAND2x1_ASAP7_75t_R _30984_ (.A(_00387_),
    .B(_10470_),
    .Y(_10472_));
 OA21x2_ASAP7_75t_R _30985_ (.A1(_09676_),
    .A2(_10469_),
    .B(_10472_),
    .Y(_03423_));
 NOR2x1_ASAP7_75t_R _30986_ (.A(_01319_),
    .B(_10098_),
    .Y(_10473_));
 AO21x1_ASAP7_75t_R _30987_ (.A1(_10253_),
    .A2(_10098_),
    .B(_10473_),
    .Y(_03424_));
 NAND2x1_ASAP7_75t_R _30988_ (.A(_00498_),
    .B(_10470_),
    .Y(_10474_));
 OA21x2_ASAP7_75t_R _30989_ (.A1(_10220_),
    .A2(_10469_),
    .B(_10474_),
    .Y(_03425_));
 NAND2x1_ASAP7_75t_R _30990_ (.A(_00529_),
    .B(_10470_),
    .Y(_10475_));
 OA21x2_ASAP7_75t_R _30991_ (.A1(_09716_),
    .A2(_10469_),
    .B(_10475_),
    .Y(_03426_));
 AND3x4_ASAP7_75t_R _30992_ (.A(_14153_),
    .B(_14050_),
    .C(_14232_),
    .Y(_10476_));
 AND4x2_ASAP7_75t_R _30993_ (.A(_08593_),
    .B(_08594_),
    .C(_08595_),
    .D(_10476_),
    .Y(_10477_));
 BUFx6f_ASAP7_75t_R _30994_ (.A(_10477_),
    .Y(_10478_));
 NOR2x1_ASAP7_75t_R _30995_ (.A(_00559_),
    .B(_10478_),
    .Y(_10479_));
 AO21x1_ASAP7_75t_R _30996_ (.A1(_10175_),
    .A2(_10478_),
    .B(_10479_),
    .Y(_03427_));
 BUFx12_ASAP7_75t_R _30997_ (.A(_10468_),
    .Y(_10480_));
 NAND2x1_ASAP7_75t_R _30998_ (.A(_00591_),
    .B(_10480_),
    .Y(_10481_));
 OA21x2_ASAP7_75t_R _30999_ (.A1(_10177_),
    .A2(_10469_),
    .B(_10481_),
    .Y(_03428_));
 NAND2x1_ASAP7_75t_R _31000_ (.A(_00621_),
    .B(_10480_),
    .Y(_10482_));
 OA21x2_ASAP7_75t_R _31001_ (.A1(_08810_),
    .A2(_10469_),
    .B(_10482_),
    .Y(_03429_));
 NAND2x1_ASAP7_75t_R _31002_ (.A(_00651_),
    .B(_10480_),
    .Y(_10483_));
 OA21x2_ASAP7_75t_R _31003_ (.A1(_08851_),
    .A2(_10469_),
    .B(_10483_),
    .Y(_03430_));
 OR2x2_ASAP7_75t_R _31004_ (.A(_00681_),
    .B(_10477_),
    .Y(_10484_));
 OAI21x1_ASAP7_75t_R _31005_ (.A1(_10279_),
    .A2(_10469_),
    .B(_10484_),
    .Y(_03431_));
 NAND2x1_ASAP7_75t_R _31006_ (.A(_00711_),
    .B(_10480_),
    .Y(_10485_));
 OA21x2_ASAP7_75t_R _31007_ (.A1(_08943_),
    .A2(_10469_),
    .B(_10485_),
    .Y(_03432_));
 NAND2x1_ASAP7_75t_R _31008_ (.A(_00741_),
    .B(_10480_),
    .Y(_10486_));
 OA21x2_ASAP7_75t_R _31009_ (.A1(_08989_),
    .A2(_10469_),
    .B(_10486_),
    .Y(_03433_));
 BUFx6f_ASAP7_75t_R _31010_ (.A(_10468_),
    .Y(_10487_));
 NAND2x1_ASAP7_75t_R _31011_ (.A(_00771_),
    .B(_10480_),
    .Y(_10488_));
 OA21x2_ASAP7_75t_R _31012_ (.A1(_09728_),
    .A2(_10487_),
    .B(_10488_),
    .Y(_03434_));
 NAND2x1_ASAP7_75t_R _31013_ (.A(_01352_),
    .B(_10037_),
    .Y(_10489_));
 OA21x2_ASAP7_75t_R _31014_ (.A1(_10255_),
    .A2(_10039_),
    .B(_10489_),
    .Y(_03435_));
 NAND2x1_ASAP7_75t_R _31015_ (.A(_00467_),
    .B(_10480_),
    .Y(_10490_));
 OA21x2_ASAP7_75t_R _31016_ (.A1(_09074_),
    .A2(_10487_),
    .B(_10490_),
    .Y(_03436_));
 NAND2x1_ASAP7_75t_R _31017_ (.A(_00842_),
    .B(_10480_),
    .Y(_10491_));
 OA21x2_ASAP7_75t_R _31018_ (.A1(_09104_),
    .A2(_10487_),
    .B(_10491_),
    .Y(_03437_));
 NAND2x1_ASAP7_75t_R _31019_ (.A(_00875_),
    .B(_10480_),
    .Y(_10492_));
 OA21x2_ASAP7_75t_R _31020_ (.A1(_09144_),
    .A2(_10487_),
    .B(_10492_),
    .Y(_03438_));
 NAND2x1_ASAP7_75t_R _31021_ (.A(_00908_),
    .B(_10480_),
    .Y(_10493_));
 OA21x2_ASAP7_75t_R _31022_ (.A1(_09181_),
    .A2(_10487_),
    .B(_10493_),
    .Y(_03439_));
 NOR2x1_ASAP7_75t_R _31023_ (.A(_00941_),
    .B(_10478_),
    .Y(_10494_));
 AO21x1_ASAP7_75t_R _31024_ (.A1(_10238_),
    .A2(_10478_),
    .B(_10494_),
    .Y(_03440_));
 BUFx10_ASAP7_75t_R _31025_ (.A(_10468_),
    .Y(_10495_));
 NAND2x1_ASAP7_75t_R _31026_ (.A(_00974_),
    .B(_10495_),
    .Y(_10496_));
 OA21x2_ASAP7_75t_R _31027_ (.A1(_09245_),
    .A2(_10487_),
    .B(_10496_),
    .Y(_03441_));
 NAND2x1_ASAP7_75t_R _31028_ (.A(_01007_),
    .B(_10495_),
    .Y(_10497_));
 OA21x2_ASAP7_75t_R _31029_ (.A1(_09271_),
    .A2(_10487_),
    .B(_10497_),
    .Y(_03442_));
 NAND2x1_ASAP7_75t_R _31030_ (.A(_01040_),
    .B(_10495_),
    .Y(_10498_));
 OA21x2_ASAP7_75t_R _31031_ (.A1(_09299_),
    .A2(_10487_),
    .B(_10498_),
    .Y(_03443_));
 NAND2x1_ASAP7_75t_R _31032_ (.A(_01073_),
    .B(_10495_),
    .Y(_10499_));
 OA21x2_ASAP7_75t_R _31033_ (.A1(_09328_),
    .A2(_10487_),
    .B(_10499_),
    .Y(_03444_));
 NAND2x1_ASAP7_75t_R _31034_ (.A(_01106_),
    .B(_10495_),
    .Y(_10500_));
 OA21x2_ASAP7_75t_R _31035_ (.A1(_09357_),
    .A2(_10487_),
    .B(_10500_),
    .Y(_03445_));
 NOR2x1_ASAP7_75t_R _31036_ (.A(_01385_),
    .B(_10097_),
    .Y(_10501_));
 AO21x1_ASAP7_75t_R _31037_ (.A1(_10257_),
    .A2(_10098_),
    .B(_10501_),
    .Y(_03446_));
 NAND2x1_ASAP7_75t_R _31038_ (.A(_01139_),
    .B(_10495_),
    .Y(_10502_));
 OA21x2_ASAP7_75t_R _31039_ (.A1(_09390_),
    .A2(_10470_),
    .B(_10502_),
    .Y(_03447_));
 NAND2x1_ASAP7_75t_R _31040_ (.A(_01172_),
    .B(_10495_),
    .Y(_10503_));
 OA21x2_ASAP7_75t_R _31041_ (.A1(_09416_),
    .A2(_10470_),
    .B(_10503_),
    .Y(_03448_));
 NAND2x1_ASAP7_75t_R _31042_ (.A(_01205_),
    .B(_10495_),
    .Y(_10504_));
 OA21x2_ASAP7_75t_R _31043_ (.A1(_10248_),
    .A2(_10470_),
    .B(_10504_),
    .Y(_03449_));
 NAND2x1_ASAP7_75t_R _31044_ (.A(_01238_),
    .B(_10495_),
    .Y(_10505_));
 OA21x2_ASAP7_75t_R _31045_ (.A1(_09472_),
    .A2(_10470_),
    .B(_10505_),
    .Y(_03450_));
 NAND2x1_ASAP7_75t_R _31046_ (.A(_01271_),
    .B(_10495_),
    .Y(_10506_));
 OA21x2_ASAP7_75t_R _31047_ (.A1(_09495_),
    .A2(_10470_),
    .B(_10506_),
    .Y(_03451_));
 NOR2x1_ASAP7_75t_R _31048_ (.A(_01304_),
    .B(_10478_),
    .Y(_10507_));
 AO21x1_ASAP7_75t_R _31049_ (.A1(_10305_),
    .A2(_10478_),
    .B(_10507_),
    .Y(_03452_));
 NOR2x1_ASAP7_75t_R _31050_ (.A(_01337_),
    .B(_10478_),
    .Y(_10508_));
 AO21x1_ASAP7_75t_R _31051_ (.A1(_10253_),
    .A2(_10478_),
    .B(_10508_),
    .Y(_03453_));
 NAND2x1_ASAP7_75t_R _31052_ (.A(_01370_),
    .B(_10468_),
    .Y(_10509_));
 OA21x2_ASAP7_75t_R _31053_ (.A1(_10255_),
    .A2(_10470_),
    .B(_10509_),
    .Y(_03454_));
 NOR2x1_ASAP7_75t_R _31054_ (.A(_01403_),
    .B(_10477_),
    .Y(_10510_));
 AO21x1_ASAP7_75t_R _31055_ (.A1(_10257_),
    .A2(_10478_),
    .B(_10510_),
    .Y(_03455_));
 AND2x2_ASAP7_75t_R _31056_ (.A(_04853_),
    .B(_10468_),
    .Y(_10511_));
 AO21x1_ASAP7_75t_R _31057_ (.A1(_10259_),
    .A2(_10478_),
    .B(_10511_),
    .Y(_03456_));
 NOR2x1_ASAP7_75t_R _31058_ (.A(_01418_),
    .B(_10097_),
    .Y(_10512_));
 AO21x1_ASAP7_75t_R _31059_ (.A1(_10259_),
    .A2(_10098_),
    .B(_10512_),
    .Y(_03457_));
 NAND2x2_ASAP7_75t_R _31060_ (.A(_08341_),
    .B(_10476_),
    .Y(_10513_));
 OR3x1_ASAP7_75t_R _31061_ (.A(_09838_),
    .B(_08589_),
    .C(_10466_),
    .Y(_10514_));
 BUFx6f_ASAP7_75t_R _31062_ (.A(_10514_),
    .Y(_10515_));
 NAND2x1_ASAP7_75t_R _31063_ (.A(_00435_),
    .B(_10515_),
    .Y(_10516_));
 OA21x2_ASAP7_75t_R _31064_ (.A1(_10162_),
    .A2(_10513_),
    .B(_10516_),
    .Y(_03458_));
 AND4x1_ASAP7_75t_R _31065_ (.A(_14726_),
    .B(_08330_),
    .C(_08338_),
    .D(_10476_),
    .Y(_10517_));
 BUFx10_ASAP7_75t_R _31066_ (.A(_10517_),
    .Y(_10518_));
 BUFx6f_ASAP7_75t_R _31067_ (.A(_10518_),
    .Y(_10519_));
 BUFx10_ASAP7_75t_R _31068_ (.A(_10518_),
    .Y(_10520_));
 NOR2x1_ASAP7_75t_R _31069_ (.A(_00388_),
    .B(_10520_),
    .Y(_10521_));
 AO21x1_ASAP7_75t_R _31070_ (.A1(_10361_),
    .A2(_10519_),
    .B(_10521_),
    .Y(_03459_));
 NAND2x1_ASAP7_75t_R _31071_ (.A(_00499_),
    .B(_10515_),
    .Y(_10522_));
 OA21x2_ASAP7_75t_R _31072_ (.A1(_10220_),
    .A2(_10515_),
    .B(_10522_),
    .Y(_03460_));
 NOR2x1_ASAP7_75t_R _31073_ (.A(_00530_),
    .B(_10520_),
    .Y(_10523_));
 AO21x1_ASAP7_75t_R _31074_ (.A1(_10368_),
    .A2(_10519_),
    .B(_10523_),
    .Y(_03461_));
 NOR2x1_ASAP7_75t_R _31075_ (.A(_00560_),
    .B(_10520_),
    .Y(_10524_));
 AO21x1_ASAP7_75t_R _31076_ (.A1(_10175_),
    .A2(_10519_),
    .B(_10524_),
    .Y(_03462_));
 NAND2x1_ASAP7_75t_R _31077_ (.A(_00592_),
    .B(_10515_),
    .Y(_10525_));
 OA21x2_ASAP7_75t_R _31078_ (.A1(_10177_),
    .A2(_10515_),
    .B(_10525_),
    .Y(_03463_));
 NOR2x1_ASAP7_75t_R _31079_ (.A(_00622_),
    .B(_10520_),
    .Y(_10526_));
 AO21x1_ASAP7_75t_R _31080_ (.A1(_10373_),
    .A2(_10519_),
    .B(_10526_),
    .Y(_03464_));
 BUFx12f_ASAP7_75t_R _31081_ (.A(_10518_),
    .Y(_10527_));
 NOR2x1_ASAP7_75t_R _31082_ (.A(_00652_),
    .B(_10527_),
    .Y(_10528_));
 AO21x1_ASAP7_75t_R _31083_ (.A1(_10375_),
    .A2(_10519_),
    .B(_10528_),
    .Y(_03465_));
 OR2x2_ASAP7_75t_R _31084_ (.A(_00682_),
    .B(_10518_),
    .Y(_10529_));
 OAI21x1_ASAP7_75t_R _31085_ (.A1(_10279_),
    .A2(_10513_),
    .B(_10529_),
    .Y(_03466_));
 NOR2x1_ASAP7_75t_R _31086_ (.A(_00712_),
    .B(_10527_),
    .Y(_10530_));
 AO21x1_ASAP7_75t_R _31087_ (.A1(_10436_),
    .A2(_10519_),
    .B(_10530_),
    .Y(_03467_));
 AND4x1_ASAP7_75t_R _31088_ (.A(_14726_),
    .B(_09773_),
    .C(_14051_),
    .D(_08338_),
    .Y(_10531_));
 BUFx10_ASAP7_75t_R _31089_ (.A(_10531_),
    .Y(_10532_));
 INVx2_ASAP7_75t_R _31090_ (.A(_10532_),
    .Y(_10533_));
 OR4x1_ASAP7_75t_R _31091_ (.A(_08027_),
    .B(_08330_),
    .C(_08586_),
    .D(_08588_),
    .Y(_10534_));
 BUFx6f_ASAP7_75t_R _31092_ (.A(_10534_),
    .Y(_10535_));
 NAND2x1_ASAP7_75t_R _31093_ (.A(_00417_),
    .B(_10535_),
    .Y(_10536_));
 OA21x2_ASAP7_75t_R _31094_ (.A1(_10162_),
    .A2(_10533_),
    .B(_10536_),
    .Y(_03468_));
 NOR2x1_ASAP7_75t_R _31095_ (.A(_00742_),
    .B(_10527_),
    .Y(_10537_));
 AO21x1_ASAP7_75t_R _31096_ (.A1(_10379_),
    .A2(_10519_),
    .B(_10537_),
    .Y(_03469_));
 NOR2x1_ASAP7_75t_R _31097_ (.A(_00772_),
    .B(_10527_),
    .Y(_10538_));
 AO21x1_ASAP7_75t_R _31098_ (.A1(_10381_),
    .A2(_10519_),
    .B(_10538_),
    .Y(_03470_));
 NOR2x1_ASAP7_75t_R _31099_ (.A(_00468_),
    .B(_10527_),
    .Y(_10539_));
 AO21x1_ASAP7_75t_R _31100_ (.A1(_10384_),
    .A2(_10519_),
    .B(_10539_),
    .Y(_03471_));
 NOR2x1_ASAP7_75t_R _31101_ (.A(_00843_),
    .B(_10527_),
    .Y(_10540_));
 AO21x1_ASAP7_75t_R _31102_ (.A1(_10387_),
    .A2(_10519_),
    .B(_10540_),
    .Y(_03472_));
 BUFx4f_ASAP7_75t_R _31103_ (.A(_10518_),
    .Y(_10541_));
 NOR2x1_ASAP7_75t_R _31104_ (.A(_00876_),
    .B(_10527_),
    .Y(_10542_));
 AO21x1_ASAP7_75t_R _31105_ (.A1(_10389_),
    .A2(_10541_),
    .B(_10542_),
    .Y(_03473_));
 NOR2x1_ASAP7_75t_R _31106_ (.A(_00909_),
    .B(_10527_),
    .Y(_10543_));
 AO21x1_ASAP7_75t_R _31107_ (.A1(_10391_),
    .A2(_10541_),
    .B(_10543_),
    .Y(_03474_));
 NOR2x1_ASAP7_75t_R _31108_ (.A(_00942_),
    .B(_10527_),
    .Y(_10544_));
 AO21x1_ASAP7_75t_R _31109_ (.A1(_10238_),
    .A2(_10541_),
    .B(_10544_),
    .Y(_03475_));
 NOR2x1_ASAP7_75t_R _31110_ (.A(_00975_),
    .B(_10527_),
    .Y(_10545_));
 AO21x1_ASAP7_75t_R _31111_ (.A1(_10395_),
    .A2(_10541_),
    .B(_10545_),
    .Y(_03476_));
 BUFx10_ASAP7_75t_R _31112_ (.A(_10518_),
    .Y(_10546_));
 NOR2x1_ASAP7_75t_R _31113_ (.A(_01008_),
    .B(_10546_),
    .Y(_10547_));
 AO21x1_ASAP7_75t_R _31114_ (.A1(_10397_),
    .A2(_10541_),
    .B(_10547_),
    .Y(_03477_));
 NOR2x1_ASAP7_75t_R _31115_ (.A(_01041_),
    .B(_10546_),
    .Y(_10548_));
 AO21x1_ASAP7_75t_R _31116_ (.A1(_10399_),
    .A2(_10541_),
    .B(_10548_),
    .Y(_03478_));
 BUFx6f_ASAP7_75t_R _31117_ (.A(_10532_),
    .Y(_10549_));
 BUFx6f_ASAP7_75t_R _31118_ (.A(_10532_),
    .Y(_10550_));
 NOR2x1_ASAP7_75t_R _31119_ (.A(_00370_),
    .B(_10550_),
    .Y(_10551_));
 AO21x1_ASAP7_75t_R _31120_ (.A1(_10361_),
    .A2(_10549_),
    .B(_10551_),
    .Y(_03479_));
 NOR2x1_ASAP7_75t_R _31121_ (.A(_01074_),
    .B(_10546_),
    .Y(_10552_));
 AO21x1_ASAP7_75t_R _31122_ (.A1(_10401_),
    .A2(_10541_),
    .B(_10552_),
    .Y(_03480_));
 NOR2x1_ASAP7_75t_R _31123_ (.A(_01107_),
    .B(_10546_),
    .Y(_10553_));
 AO21x1_ASAP7_75t_R _31124_ (.A1(_10403_),
    .A2(_10541_),
    .B(_10553_),
    .Y(_03481_));
 NOR2x1_ASAP7_75t_R _31125_ (.A(_01140_),
    .B(_10546_),
    .Y(_10554_));
 AO21x1_ASAP7_75t_R _31126_ (.A1(_10453_),
    .A2(_10541_),
    .B(_10554_),
    .Y(_03482_));
 NOR2x1_ASAP7_75t_R _31127_ (.A(_01173_),
    .B(_10546_),
    .Y(_10555_));
 AO21x1_ASAP7_75t_R _31128_ (.A1(_10406_),
    .A2(_10541_),
    .B(_10555_),
    .Y(_03483_));
 NAND2x1_ASAP7_75t_R _31129_ (.A(_01206_),
    .B(_10515_),
    .Y(_10556_));
 OA21x2_ASAP7_75t_R _31130_ (.A1(_10248_),
    .A2(_10513_),
    .B(_10556_),
    .Y(_03484_));
 NOR2x1_ASAP7_75t_R _31131_ (.A(_01239_),
    .B(_10546_),
    .Y(_10557_));
 AO21x1_ASAP7_75t_R _31132_ (.A1(_10409_),
    .A2(_10520_),
    .B(_10557_),
    .Y(_03485_));
 NOR2x1_ASAP7_75t_R _31133_ (.A(_01272_),
    .B(_10546_),
    .Y(_10558_));
 AO21x1_ASAP7_75t_R _31134_ (.A1(_10412_),
    .A2(_10520_),
    .B(_10558_),
    .Y(_03486_));
 NOR2x1_ASAP7_75t_R _31135_ (.A(_01305_),
    .B(_10546_),
    .Y(_10559_));
 AO21x1_ASAP7_75t_R _31136_ (.A1(_10305_),
    .A2(_10520_),
    .B(_10559_),
    .Y(_03487_));
 NOR2x1_ASAP7_75t_R _31137_ (.A(_01338_),
    .B(_10546_),
    .Y(_10560_));
 AO21x1_ASAP7_75t_R _31138_ (.A1(_10253_),
    .A2(_10520_),
    .B(_10560_),
    .Y(_03488_));
 NAND2x1_ASAP7_75t_R _31139_ (.A(_01371_),
    .B(_10515_),
    .Y(_10561_));
 OA21x2_ASAP7_75t_R _31140_ (.A1(_10255_),
    .A2(_10515_),
    .B(_10561_),
    .Y(_03489_));
 NAND2x1_ASAP7_75t_R _31141_ (.A(_00481_),
    .B(_10535_),
    .Y(_10562_));
 OA21x2_ASAP7_75t_R _31142_ (.A1(_10220_),
    .A2(_10535_),
    .B(_10562_),
    .Y(_03490_));
 NOR2x1_ASAP7_75t_R _31143_ (.A(_01404_),
    .B(_10518_),
    .Y(_10563_));
 AO21x1_ASAP7_75t_R _31144_ (.A1(_10257_),
    .A2(_10520_),
    .B(_10563_),
    .Y(_03491_));
 AND2x2_ASAP7_75t_R _31145_ (.A(_04842_),
    .B(_10515_),
    .Y(_10564_));
 AO21x1_ASAP7_75t_R _31146_ (.A1(_10259_),
    .A2(_10520_),
    .B(_10564_),
    .Y(_03492_));
 OR3x1_ASAP7_75t_R _31147_ (.A(_09766_),
    .B(_09767_),
    .C(_10466_),
    .Y(_10565_));
 BUFx10_ASAP7_75t_R _31148_ (.A(_10565_),
    .Y(_10566_));
 BUFx6f_ASAP7_75t_R _31149_ (.A(_10566_),
    .Y(_10567_));
 NAND2x1_ASAP7_75t_R _31150_ (.A(_00436_),
    .B(_10567_),
    .Y(_10568_));
 OA21x2_ASAP7_75t_R _31151_ (.A1(_10162_),
    .A2(_10567_),
    .B(_10568_),
    .Y(_03493_));
 AND3x1_ASAP7_75t_R _31152_ (.A(_08339_),
    .B(_09774_),
    .C(_10476_),
    .Y(_10569_));
 BUFx10_ASAP7_75t_R _31153_ (.A(_10569_),
    .Y(_10570_));
 BUFx6f_ASAP7_75t_R _31154_ (.A(_10570_),
    .Y(_10571_));
 BUFx6f_ASAP7_75t_R _31155_ (.A(_10566_),
    .Y(_10572_));
 AND2x2_ASAP7_75t_R _31156_ (.A(_13522_),
    .B(_10572_),
    .Y(_10573_));
 AO21x1_ASAP7_75t_R _31157_ (.A1(_10361_),
    .A2(_10571_),
    .B(_10573_),
    .Y(_03494_));
 NAND2x1_ASAP7_75t_R _31158_ (.A(_00500_),
    .B(_10567_),
    .Y(_10574_));
 OA21x2_ASAP7_75t_R _31159_ (.A1(_10220_),
    .A2(_10567_),
    .B(_10574_),
    .Y(_03495_));
 AND2x2_ASAP7_75t_R _31160_ (.A(_14202_),
    .B(_10572_),
    .Y(_10575_));
 AO21x1_ASAP7_75t_R _31161_ (.A1(_10368_),
    .A2(_10571_),
    .B(_10575_),
    .Y(_03496_));
 AND2x2_ASAP7_75t_R _31162_ (.A(_14286_),
    .B(_10572_),
    .Y(_10576_));
 AO21x1_ASAP7_75t_R _31163_ (.A1(_10175_),
    .A2(_10571_),
    .B(_10576_),
    .Y(_03497_));
 NAND2x1_ASAP7_75t_R _31164_ (.A(_00593_),
    .B(_10567_),
    .Y(_10577_));
 OA21x2_ASAP7_75t_R _31165_ (.A1(_10177_),
    .A2(_10567_),
    .B(_10577_),
    .Y(_03498_));
 AND2x2_ASAP7_75t_R _31166_ (.A(_15158_),
    .B(_10572_),
    .Y(_10578_));
 AO21x1_ASAP7_75t_R _31167_ (.A1(_10373_),
    .A2(_10571_),
    .B(_10578_),
    .Y(_03499_));
 AND2x2_ASAP7_75t_R _31168_ (.A(_14444_),
    .B(_10572_),
    .Y(_10579_));
 AO21x1_ASAP7_75t_R _31169_ (.A1(_10375_),
    .A2(_10571_),
    .B(_10579_),
    .Y(_03500_));
 NOR2x1_ASAP7_75t_R _31170_ (.A(_00512_),
    .B(_10550_),
    .Y(_10580_));
 AO21x1_ASAP7_75t_R _31171_ (.A1(_10368_),
    .A2(_10549_),
    .B(_10580_),
    .Y(_03501_));
 OR3x1_ASAP7_75t_R _31172_ (.A(_09790_),
    .B(_09791_),
    .C(_10572_),
    .Y(_10581_));
 OAI21x1_ASAP7_75t_R _31173_ (.A1(_00683_),
    .A2(_10571_),
    .B(_10581_),
    .Y(_03502_));
 AND2x2_ASAP7_75t_R _31174_ (.A(_14597_),
    .B(_10572_),
    .Y(_10582_));
 AO21x1_ASAP7_75t_R _31175_ (.A1(_10436_),
    .A2(_10571_),
    .B(_10582_),
    .Y(_03503_));
 AND2x2_ASAP7_75t_R _31176_ (.A(_14624_),
    .B(_10572_),
    .Y(_10583_));
 AO21x1_ASAP7_75t_R _31177_ (.A1(_10379_),
    .A2(_10571_),
    .B(_10583_),
    .Y(_03504_));
 AND2x2_ASAP7_75t_R _31178_ (.A(_14675_),
    .B(_10572_),
    .Y(_10584_));
 AO21x1_ASAP7_75t_R _31179_ (.A1(_10381_),
    .A2(_10571_),
    .B(_10584_),
    .Y(_03505_));
 BUFx6f_ASAP7_75t_R _31180_ (.A(_10566_),
    .Y(_10585_));
 AND2x2_ASAP7_75t_R _31181_ (.A(_13974_),
    .B(_10585_),
    .Y(_10586_));
 AO21x1_ASAP7_75t_R _31182_ (.A1(_10384_),
    .A2(_10571_),
    .B(_10586_),
    .Y(_03506_));
 BUFx4f_ASAP7_75t_R _31183_ (.A(_10570_),
    .Y(_10587_));
 AND2x2_ASAP7_75t_R _31184_ (.A(_15636_),
    .B(_10585_),
    .Y(_10588_));
 AO21x1_ASAP7_75t_R _31185_ (.A1(_10387_),
    .A2(_10587_),
    .B(_10588_),
    .Y(_03507_));
 AND2x2_ASAP7_75t_R _31186_ (.A(_15786_),
    .B(_10585_),
    .Y(_10589_));
 AO21x1_ASAP7_75t_R _31187_ (.A1(_10389_),
    .A2(_10587_),
    .B(_10589_),
    .Y(_03508_));
 AND2x2_ASAP7_75t_R _31188_ (.A(_15916_),
    .B(_10585_),
    .Y(_10590_));
 AO21x1_ASAP7_75t_R _31189_ (.A1(_10391_),
    .A2(_10587_),
    .B(_10590_),
    .Y(_03509_));
 AND3x1_ASAP7_75t_R _31190_ (.A(_09204_),
    .B(_09212_),
    .C(_10570_),
    .Y(_10591_));
 AO21x1_ASAP7_75t_R _31191_ (.A1(_16064_),
    .A2(_10567_),
    .B(_10591_),
    .Y(_03510_));
 AND2x2_ASAP7_75t_R _31192_ (.A(_16181_),
    .B(_10585_),
    .Y(_10592_));
 AO21x1_ASAP7_75t_R _31193_ (.A1(_10395_),
    .A2(_10587_),
    .B(_10592_),
    .Y(_03511_));
 NOR2x1_ASAP7_75t_R _31194_ (.A(_00542_),
    .B(_10550_),
    .Y(_10593_));
 AO21x1_ASAP7_75t_R _31195_ (.A1(_10175_),
    .A2(_10549_),
    .B(_10593_),
    .Y(_03512_));
 AND2x2_ASAP7_75t_R _31196_ (.A(_16325_),
    .B(_10585_),
    .Y(_10594_));
 AO21x1_ASAP7_75t_R _31197_ (.A1(_10397_),
    .A2(_10587_),
    .B(_10594_),
    .Y(_03513_));
 AND2x2_ASAP7_75t_R _31198_ (.A(_16438_),
    .B(_10585_),
    .Y(_10595_));
 AO21x1_ASAP7_75t_R _31199_ (.A1(_10399_),
    .A2(_10587_),
    .B(_10595_),
    .Y(_03514_));
 AND2x2_ASAP7_75t_R _31200_ (.A(_16564_),
    .B(_10585_),
    .Y(_10596_));
 AO21x1_ASAP7_75t_R _31201_ (.A1(_10401_),
    .A2(_10587_),
    .B(_10596_),
    .Y(_03515_));
 AND2x2_ASAP7_75t_R _31202_ (.A(_16678_),
    .B(_10585_),
    .Y(_10597_));
 AO21x1_ASAP7_75t_R _31203_ (.A1(_10403_),
    .A2(_10587_),
    .B(_10597_),
    .Y(_03516_));
 AND2x2_ASAP7_75t_R _31204_ (.A(_16808_),
    .B(_10585_),
    .Y(_10598_));
 AO21x1_ASAP7_75t_R _31205_ (.A1(_10453_),
    .A2(_10587_),
    .B(_10598_),
    .Y(_03517_));
 AND2x2_ASAP7_75t_R _31206_ (.A(_16918_),
    .B(_10566_),
    .Y(_10599_));
 AO21x1_ASAP7_75t_R _31207_ (.A1(_10406_),
    .A2(_10587_),
    .B(_10599_),
    .Y(_03518_));
 NAND2x1_ASAP7_75t_R _31208_ (.A(_01207_),
    .B(_10567_),
    .Y(_10600_));
 OA21x2_ASAP7_75t_R _31209_ (.A1(_10248_),
    .A2(_10567_),
    .B(_10600_),
    .Y(_03519_));
 AND2x2_ASAP7_75t_R _31210_ (.A(_17157_),
    .B(_10566_),
    .Y(_10601_));
 AO21x1_ASAP7_75t_R _31211_ (.A1(_10409_),
    .A2(_10570_),
    .B(_10601_),
    .Y(_03520_));
 AND2x2_ASAP7_75t_R _31212_ (.A(_17288_),
    .B(_10566_),
    .Y(_10602_));
 AO21x1_ASAP7_75t_R _31213_ (.A1(_10412_),
    .A2(_10570_),
    .B(_10602_),
    .Y(_03521_));
 AND2x2_ASAP7_75t_R _31214_ (.A(_04315_),
    .B(_10566_),
    .Y(_10603_));
 AO21x1_ASAP7_75t_R _31215_ (.A1(_10305_),
    .A2(_10570_),
    .B(_10603_),
    .Y(_03522_));
 NAND2x1_ASAP7_75t_R _31216_ (.A(_00574_),
    .B(_10535_),
    .Y(_10604_));
 OA21x2_ASAP7_75t_R _31217_ (.A1(_10177_),
    .A2(_10535_),
    .B(_10604_),
    .Y(_03523_));
 NAND2x1_ASAP7_75t_R _31218_ (.A(_01786_),
    .B(_09106_),
    .Y(_10605_));
 OA21x2_ASAP7_75t_R _31219_ (.A1(_08591_),
    .A2(_08810_),
    .B(_10605_),
    .Y(_03524_));
 AND2x2_ASAP7_75t_R _31220_ (.A(_04445_),
    .B(_10566_),
    .Y(_10606_));
 AO21x1_ASAP7_75t_R _31221_ (.A1(_10253_),
    .A2(_10570_),
    .B(_10606_),
    .Y(_03525_));
 NAND2x1_ASAP7_75t_R _31222_ (.A(_01372_),
    .B(_10572_),
    .Y(_10607_));
 OA21x2_ASAP7_75t_R _31223_ (.A1(_10255_),
    .A2(_10567_),
    .B(_10607_),
    .Y(_03526_));
 AND2x2_ASAP7_75t_R _31224_ (.A(_04669_),
    .B(_10566_),
    .Y(_10608_));
 AO21x1_ASAP7_75t_R _31225_ (.A1(net153),
    .A2(_10570_),
    .B(_10608_),
    .Y(_03527_));
 AND2x2_ASAP7_75t_R _31226_ (.A(_04779_),
    .B(_10566_),
    .Y(_10609_));
 AO21x1_ASAP7_75t_R _31227_ (.A1(net9),
    .A2(_10570_),
    .B(_10609_),
    .Y(_03528_));
 AND4x2_ASAP7_75t_R _31228_ (.A(_08329_),
    .B(_09773_),
    .C(_09834_),
    .D(_10476_),
    .Y(_10610_));
 BUFx10_ASAP7_75t_R _31229_ (.A(_10610_),
    .Y(_10611_));
 INVx1_ASAP7_75t_R _31230_ (.A(_10611_),
    .Y(_10612_));
 OR4x2_ASAP7_75t_R _31231_ (.A(_08027_),
    .B(_08330_),
    .C(_09766_),
    .D(_10466_),
    .Y(_10613_));
 BUFx10_ASAP7_75t_R _31232_ (.A(_10613_),
    .Y(_10614_));
 NAND2x1_ASAP7_75t_R _31233_ (.A(_00437_),
    .B(_10614_),
    .Y(_10615_));
 OA21x2_ASAP7_75t_R _31234_ (.A1(_08585_),
    .A2(_10612_),
    .B(_10615_),
    .Y(_03529_));
 BUFx12f_ASAP7_75t_R _31235_ (.A(_10610_),
    .Y(_10616_));
 BUFx6f_ASAP7_75t_R _31236_ (.A(_10616_),
    .Y(_10617_));
 NOR2x1_ASAP7_75t_R _31237_ (.A(_00390_),
    .B(_10611_),
    .Y(_10618_));
 AO21x1_ASAP7_75t_R _31238_ (.A1(_10361_),
    .A2(_10617_),
    .B(_10618_),
    .Y(_03530_));
 NAND2x1_ASAP7_75t_R _31239_ (.A(_00501_),
    .B(_10614_),
    .Y(_10619_));
 OA21x2_ASAP7_75t_R _31240_ (.A1(_10220_),
    .A2(_10614_),
    .B(_10619_),
    .Y(_03531_));
 NOR2x1_ASAP7_75t_R _31241_ (.A(_00532_),
    .B(_10611_),
    .Y(_10620_));
 AO21x1_ASAP7_75t_R _31242_ (.A1(_10368_),
    .A2(_10617_),
    .B(_10620_),
    .Y(_03532_));
 AND2x2_ASAP7_75t_R _31243_ (.A(_14289_),
    .B(_10614_),
    .Y(_10621_));
 AO21x1_ASAP7_75t_R _31244_ (.A1(_08676_),
    .A2(_10617_),
    .B(_10621_),
    .Y(_03533_));
 NAND2x1_ASAP7_75t_R _31245_ (.A(_00594_),
    .B(_10614_),
    .Y(_10622_));
 OA21x2_ASAP7_75t_R _31246_ (.A1(_08763_),
    .A2(_10614_),
    .B(_10622_),
    .Y(_03534_));
 NOR2x1_ASAP7_75t_R _31247_ (.A(_00604_),
    .B(_10550_),
    .Y(_10623_));
 AO21x1_ASAP7_75t_R _31248_ (.A1(_10373_),
    .A2(_10549_),
    .B(_10623_),
    .Y(_03535_));
 BUFx12f_ASAP7_75t_R _31249_ (.A(_10610_),
    .Y(_10624_));
 NOR2x1_ASAP7_75t_R _31250_ (.A(_00624_),
    .B(_10624_),
    .Y(_10625_));
 AO21x1_ASAP7_75t_R _31251_ (.A1(_10373_),
    .A2(_10617_),
    .B(_10625_),
    .Y(_03536_));
 NOR2x1_ASAP7_75t_R _31252_ (.A(_00654_),
    .B(_10624_),
    .Y(_10626_));
 AO21x1_ASAP7_75t_R _31253_ (.A1(_10375_),
    .A2(_10617_),
    .B(_10626_),
    .Y(_03537_));
 OR3x1_ASAP7_75t_R _31254_ (.A(_09790_),
    .B(_09791_),
    .C(_10614_),
    .Y(_10627_));
 OAI21x1_ASAP7_75t_R _31255_ (.A1(_00684_),
    .A2(_10617_),
    .B(_10627_),
    .Y(_03538_));
 NOR2x1_ASAP7_75t_R _31256_ (.A(_00714_),
    .B(_10624_),
    .Y(_10628_));
 AO21x1_ASAP7_75t_R _31257_ (.A1(_10436_),
    .A2(_10617_),
    .B(_10628_),
    .Y(_03539_));
 NOR2x1_ASAP7_75t_R _31258_ (.A(_00744_),
    .B(_10624_),
    .Y(_10629_));
 AO21x1_ASAP7_75t_R _31259_ (.A1(_10379_),
    .A2(_10617_),
    .B(_10629_),
    .Y(_03540_));
 NOR2x1_ASAP7_75t_R _31260_ (.A(_00774_),
    .B(_10624_),
    .Y(_10630_));
 AO21x1_ASAP7_75t_R _31261_ (.A1(_10381_),
    .A2(_10617_),
    .B(_10630_),
    .Y(_03541_));
 NOR2x1_ASAP7_75t_R _31262_ (.A(_00470_),
    .B(_10624_),
    .Y(_10631_));
 AO21x1_ASAP7_75t_R _31263_ (.A1(_10384_),
    .A2(_10617_),
    .B(_10631_),
    .Y(_03542_));
 BUFx4f_ASAP7_75t_R _31264_ (.A(_10616_),
    .Y(_10632_));
 NOR2x1_ASAP7_75t_R _31265_ (.A(_00845_),
    .B(_10624_),
    .Y(_10633_));
 AO21x1_ASAP7_75t_R _31266_ (.A1(_10387_),
    .A2(_10632_),
    .B(_10633_),
    .Y(_03543_));
 NOR2x1_ASAP7_75t_R _31267_ (.A(_00878_),
    .B(_10624_),
    .Y(_10634_));
 AO21x1_ASAP7_75t_R _31268_ (.A1(_10389_),
    .A2(_10632_),
    .B(_10634_),
    .Y(_03544_));
 NOR2x1_ASAP7_75t_R _31269_ (.A(_00911_),
    .B(_10624_),
    .Y(_10635_));
 AO21x1_ASAP7_75t_R _31270_ (.A1(_10391_),
    .A2(_10632_),
    .B(_10635_),
    .Y(_03545_));
 BUFx10_ASAP7_75t_R _31271_ (.A(_10532_),
    .Y(_10636_));
 NOR2x1_ASAP7_75t_R _31272_ (.A(_00634_),
    .B(_10636_),
    .Y(_10637_));
 AO21x1_ASAP7_75t_R _31273_ (.A1(_10375_),
    .A2(_10549_),
    .B(_10637_),
    .Y(_03546_));
 AND2x2_ASAP7_75t_R _31274_ (.A(_16061_),
    .B(_10613_),
    .Y(_10638_));
 AO21x1_ASAP7_75t_R _31275_ (.A1(_10238_),
    .A2(_10632_),
    .B(_10638_),
    .Y(_03547_));
 NOR2x1_ASAP7_75t_R _31276_ (.A(_00977_),
    .B(_10624_),
    .Y(_10639_));
 AO21x1_ASAP7_75t_R _31277_ (.A1(_10395_),
    .A2(_10632_),
    .B(_10639_),
    .Y(_03548_));
 NOR2x1_ASAP7_75t_R _31278_ (.A(_01010_),
    .B(_10616_),
    .Y(_10640_));
 AO21x1_ASAP7_75t_R _31279_ (.A1(_10397_),
    .A2(_10632_),
    .B(_10640_),
    .Y(_03549_));
 NOR2x1_ASAP7_75t_R _31280_ (.A(_01043_),
    .B(_10616_),
    .Y(_10641_));
 AO21x1_ASAP7_75t_R _31281_ (.A1(_10399_),
    .A2(_10632_),
    .B(_10641_),
    .Y(_03550_));
 NOR2x1_ASAP7_75t_R _31282_ (.A(_01076_),
    .B(_10616_),
    .Y(_10642_));
 AO21x1_ASAP7_75t_R _31283_ (.A1(_10401_),
    .A2(_10632_),
    .B(_10642_),
    .Y(_03551_));
 NOR2x1_ASAP7_75t_R _31284_ (.A(_01109_),
    .B(_10616_),
    .Y(_10643_));
 AO21x1_ASAP7_75t_R _31285_ (.A1(_10403_),
    .A2(_10632_),
    .B(_10643_),
    .Y(_03552_));
 NOR2x1_ASAP7_75t_R _31286_ (.A(_01142_),
    .B(_10616_),
    .Y(_10644_));
 AO21x1_ASAP7_75t_R _31287_ (.A1(_10453_),
    .A2(_10632_),
    .B(_10644_),
    .Y(_03553_));
 NOR2x1_ASAP7_75t_R _31288_ (.A(_01175_),
    .B(_10616_),
    .Y(_10645_));
 AO21x1_ASAP7_75t_R _31289_ (.A1(_10406_),
    .A2(_10611_),
    .B(_10645_),
    .Y(_03554_));
 NAND2x1_ASAP7_75t_R _31290_ (.A(_01208_),
    .B(_10614_),
    .Y(_10646_));
 OA21x2_ASAP7_75t_R _31291_ (.A1(_10248_),
    .A2(_10612_),
    .B(_10646_),
    .Y(_03555_));
 NOR2x1_ASAP7_75t_R _31292_ (.A(_01241_),
    .B(_10616_),
    .Y(_10647_));
 AO21x1_ASAP7_75t_R _31293_ (.A1(_10409_),
    .A2(_10611_),
    .B(_10647_),
    .Y(_03556_));
 OR2x2_ASAP7_75t_R _31294_ (.A(_00664_),
    .B(_10532_),
    .Y(_10648_));
 OAI21x1_ASAP7_75t_R _31295_ (.A1(_10279_),
    .A2(_10533_),
    .B(_10648_),
    .Y(_03557_));
 NOR2x1_ASAP7_75t_R _31296_ (.A(_01274_),
    .B(_10616_),
    .Y(_10649_));
 AO21x1_ASAP7_75t_R _31297_ (.A1(_10412_),
    .A2(_10611_),
    .B(_10649_),
    .Y(_03558_));
 AND2x2_ASAP7_75t_R _31298_ (.A(_04312_),
    .B(_10613_),
    .Y(_10650_));
 AO21x1_ASAP7_75t_R _31299_ (.A1(_10305_),
    .A2(_10611_),
    .B(_10650_),
    .Y(_03559_));
 AND2x2_ASAP7_75t_R _31300_ (.A(_04442_),
    .B(_10613_),
    .Y(_10651_));
 AO21x1_ASAP7_75t_R _31301_ (.A1(_10253_),
    .A2(_10611_),
    .B(_10651_),
    .Y(_03560_));
 NAND2x1_ASAP7_75t_R _31302_ (.A(_01373_),
    .B(_10614_),
    .Y(_10652_));
 OA21x2_ASAP7_75t_R _31303_ (.A1(_10255_),
    .A2(_10614_),
    .B(_10652_),
    .Y(_03561_));
 AND2x2_ASAP7_75t_R _31304_ (.A(_04666_),
    .B(_10613_),
    .Y(_10653_));
 AO21x1_ASAP7_75t_R _31305_ (.A1(net153),
    .A2(_10611_),
    .B(_10653_),
    .Y(_03562_));
 AND2x2_ASAP7_75t_R _31306_ (.A(_04776_),
    .B(_10613_),
    .Y(_10654_));
 AO21x1_ASAP7_75t_R _31307_ (.A1(net9),
    .A2(_10611_),
    .B(_10654_),
    .Y(_03563_));
 OR3x2_ASAP7_75t_R _31308_ (.A(_14153_),
    .B(_14050_),
    .C(_14231_),
    .Y(_10655_));
 OR3x4_ASAP7_75t_R _31309_ (.A(_08677_),
    .B(_09766_),
    .C(_10655_),
    .Y(_10656_));
 BUFx6f_ASAP7_75t_R _31310_ (.A(_10656_),
    .Y(_10657_));
 BUFx10_ASAP7_75t_R _31311_ (.A(_10656_),
    .Y(_10658_));
 NAND2x1_ASAP7_75t_R _31312_ (.A(_00438_),
    .B(_10658_),
    .Y(_10659_));
 OA21x2_ASAP7_75t_R _31313_ (.A1(_08585_),
    .A2(_10657_),
    .B(_10659_),
    .Y(_03564_));
 AND3x2_ASAP7_75t_R _31314_ (.A(_14049_),
    .B(_14303_),
    .C(_14232_),
    .Y(_10660_));
 AND4x2_ASAP7_75t_R _31315_ (.A(_08593_),
    .B(_08594_),
    .C(_08595_),
    .D(_10660_),
    .Y(_10661_));
 BUFx6f_ASAP7_75t_R _31316_ (.A(_10661_),
    .Y(_10662_));
 BUFx10_ASAP7_75t_R _31317_ (.A(_10656_),
    .Y(_10663_));
 AND2x2_ASAP7_75t_R _31318_ (.A(_13534_),
    .B(_10663_),
    .Y(_10664_));
 AO21x1_ASAP7_75t_R _31319_ (.A1(_10361_),
    .A2(_10662_),
    .B(_10664_),
    .Y(_03565_));
 NAND2x1_ASAP7_75t_R _31320_ (.A(_00502_),
    .B(_10658_),
    .Y(_10665_));
 OA21x2_ASAP7_75t_R _31321_ (.A1(_09696_),
    .A2(_10657_),
    .B(_10665_),
    .Y(_03566_));
 NAND2x1_ASAP7_75t_R _31322_ (.A(_00533_),
    .B(_10658_),
    .Y(_10666_));
 OA21x2_ASAP7_75t_R _31323_ (.A1(_09716_),
    .A2(_10657_),
    .B(_10666_),
    .Y(_03567_));
 NOR2x1_ASAP7_75t_R _31324_ (.A(_00694_),
    .B(_10636_),
    .Y(_10667_));
 AO21x1_ASAP7_75t_R _31325_ (.A1(_10436_),
    .A2(_10549_),
    .B(_10667_),
    .Y(_03568_));
 NOR2x1_ASAP7_75t_R _31326_ (.A(_00563_),
    .B(_10661_),
    .Y(_10668_));
 AO21x1_ASAP7_75t_R _31327_ (.A1(_08676_),
    .A2(_10662_),
    .B(_10668_),
    .Y(_03569_));
 NAND2x1_ASAP7_75t_R _31328_ (.A(_00595_),
    .B(_10658_),
    .Y(_10669_));
 OA21x2_ASAP7_75t_R _31329_ (.A1(_08763_),
    .A2(_10657_),
    .B(_10669_),
    .Y(_03570_));
 NAND2x1_ASAP7_75t_R _31330_ (.A(_00625_),
    .B(_10658_),
    .Y(_10670_));
 OA21x2_ASAP7_75t_R _31331_ (.A1(_08810_),
    .A2(_10657_),
    .B(_10670_),
    .Y(_03571_));
 NAND2x1_ASAP7_75t_R _31332_ (.A(_00655_),
    .B(_10658_),
    .Y(_10671_));
 OA21x2_ASAP7_75t_R _31333_ (.A1(_08851_),
    .A2(_10657_),
    .B(_10671_),
    .Y(_03572_));
 NAND2x1_ASAP7_75t_R _31334_ (.A(_15320_),
    .B(_10658_),
    .Y(_10672_));
 OAI21x1_ASAP7_75t_R _31335_ (.A1(_10279_),
    .A2(_10657_),
    .B(_10672_),
    .Y(_03573_));
 NAND2x1_ASAP7_75t_R _31336_ (.A(_00715_),
    .B(_10658_),
    .Y(_10673_));
 OA21x2_ASAP7_75t_R _31337_ (.A1(_08943_),
    .A2(_10657_),
    .B(_10673_),
    .Y(_03574_));
 NAND2x1_ASAP7_75t_R _31338_ (.A(_00745_),
    .B(_10663_),
    .Y(_10674_));
 OA21x2_ASAP7_75t_R _31339_ (.A1(_08989_),
    .A2(_10657_),
    .B(_10674_),
    .Y(_03575_));
 NAND2x1_ASAP7_75t_R _31340_ (.A(_00775_),
    .B(_10663_),
    .Y(_10675_));
 OA21x2_ASAP7_75t_R _31341_ (.A1(_09728_),
    .A2(_10657_),
    .B(_10675_),
    .Y(_03576_));
 AND2x2_ASAP7_75t_R _31342_ (.A(_13997_),
    .B(_10663_),
    .Y(_10676_));
 AO21x1_ASAP7_75t_R _31343_ (.A1(_10384_),
    .A2(_10662_),
    .B(_10676_),
    .Y(_03577_));
 AND2x2_ASAP7_75t_R _31344_ (.A(_15650_),
    .B(_10663_),
    .Y(_10677_));
 AO21x1_ASAP7_75t_R _31345_ (.A1(_10387_),
    .A2(_10662_),
    .B(_10677_),
    .Y(_03578_));
 NOR2x1_ASAP7_75t_R _31346_ (.A(_00724_),
    .B(_10636_),
    .Y(_10678_));
 AO21x1_ASAP7_75t_R _31347_ (.A1(_10379_),
    .A2(_10549_),
    .B(_10678_),
    .Y(_03579_));
 AND2x2_ASAP7_75t_R _31348_ (.A(_15798_),
    .B(_10663_),
    .Y(_10679_));
 AO21x1_ASAP7_75t_R _31349_ (.A1(_10389_),
    .A2(_10662_),
    .B(_10679_),
    .Y(_03580_));
 AND2x2_ASAP7_75t_R _31350_ (.A(_15932_),
    .B(_10663_),
    .Y(_10680_));
 AO21x1_ASAP7_75t_R _31351_ (.A1(_10391_),
    .A2(_10662_),
    .B(_10680_),
    .Y(_03581_));
 AND2x2_ASAP7_75t_R _31352_ (.A(_16076_),
    .B(_10663_),
    .Y(_10681_));
 AO21x1_ASAP7_75t_R _31353_ (.A1(_10238_),
    .A2(_10662_),
    .B(_10681_),
    .Y(_03582_));
 BUFx4f_ASAP7_75t_R _31354_ (.A(_10656_),
    .Y(_10682_));
 AND2x2_ASAP7_75t_R _31355_ (.A(_16193_),
    .B(_10682_),
    .Y(_10683_));
 AO21x1_ASAP7_75t_R _31356_ (.A1(_10395_),
    .A2(_10662_),
    .B(_10683_),
    .Y(_03583_));
 AND2x2_ASAP7_75t_R _31357_ (.A(_16337_),
    .B(_10682_),
    .Y(_10684_));
 AO21x1_ASAP7_75t_R _31358_ (.A1(_10397_),
    .A2(_10662_),
    .B(_10684_),
    .Y(_03584_));
 AND2x2_ASAP7_75t_R _31359_ (.A(_16450_),
    .B(_10682_),
    .Y(_10685_));
 AO21x1_ASAP7_75t_R _31360_ (.A1(_10399_),
    .A2(_10662_),
    .B(_10685_),
    .Y(_03585_));
 BUFx4f_ASAP7_75t_R _31361_ (.A(_10661_),
    .Y(_10686_));
 AND2x2_ASAP7_75t_R _31362_ (.A(_16576_),
    .B(_10682_),
    .Y(_10687_));
 AO21x1_ASAP7_75t_R _31363_ (.A1(_10401_),
    .A2(_10686_),
    .B(_10687_),
    .Y(_03586_));
 AND2x2_ASAP7_75t_R _31364_ (.A(_16690_),
    .B(_10682_),
    .Y(_10688_));
 AO21x1_ASAP7_75t_R _31365_ (.A1(_10403_),
    .A2(_10686_),
    .B(_10688_),
    .Y(_03587_));
 AND2x2_ASAP7_75t_R _31366_ (.A(_16820_),
    .B(_10682_),
    .Y(_10689_));
 AO21x1_ASAP7_75t_R _31367_ (.A1(_10453_),
    .A2(_10686_),
    .B(_10689_),
    .Y(_03588_));
 AND2x2_ASAP7_75t_R _31368_ (.A(_16930_),
    .B(_10682_),
    .Y(_10690_));
 AO21x1_ASAP7_75t_R _31369_ (.A1(_10406_),
    .A2(_10686_),
    .B(_10690_),
    .Y(_03589_));
 NOR2x1_ASAP7_75t_R _31370_ (.A(_00754_),
    .B(_10636_),
    .Y(_10691_));
 AO21x1_ASAP7_75t_R _31371_ (.A1(_10381_),
    .A2(_10549_),
    .B(_10691_),
    .Y(_03590_));
 NAND2x1_ASAP7_75t_R _31372_ (.A(_01209_),
    .B(_10663_),
    .Y(_10692_));
 OA21x2_ASAP7_75t_R _31373_ (.A1(_09442_),
    .A2(_10658_),
    .B(_10692_),
    .Y(_03591_));
 AND2x2_ASAP7_75t_R _31374_ (.A(_17169_),
    .B(_10682_),
    .Y(_10693_));
 AO21x1_ASAP7_75t_R _31375_ (.A1(_10409_),
    .A2(_10686_),
    .B(_10693_),
    .Y(_03592_));
 AND2x2_ASAP7_75t_R _31376_ (.A(_17300_),
    .B(_10682_),
    .Y(_10694_));
 AO21x1_ASAP7_75t_R _31377_ (.A1(_10412_),
    .A2(_10686_),
    .B(_10694_),
    .Y(_03593_));
 AND2x2_ASAP7_75t_R _31378_ (.A(_04327_),
    .B(_10682_),
    .Y(_10695_));
 AO21x1_ASAP7_75t_R _31379_ (.A1(_10305_),
    .A2(_10686_),
    .B(_10695_),
    .Y(_03594_));
 AND2x2_ASAP7_75t_R _31380_ (.A(_04457_),
    .B(_10656_),
    .Y(_10696_));
 AO21x1_ASAP7_75t_R _31381_ (.A1(_10253_),
    .A2(_10686_),
    .B(_10696_),
    .Y(_03595_));
 NAND2x1_ASAP7_75t_R _31382_ (.A(_01374_),
    .B(_10663_),
    .Y(_10697_));
 OA21x2_ASAP7_75t_R _31383_ (.A1(_10255_),
    .A2(_10658_),
    .B(_10697_),
    .Y(_03596_));
 AND2x2_ASAP7_75t_R _31384_ (.A(_04681_),
    .B(_10656_),
    .Y(_10698_));
 AO21x1_ASAP7_75t_R _31385_ (.A1(net151),
    .A2(_10686_),
    .B(_10698_),
    .Y(_03597_));
 AND2x2_ASAP7_75t_R _31386_ (.A(_04830_),
    .B(_10656_),
    .Y(_10699_));
 AO21x1_ASAP7_75t_R _31387_ (.A1(net7),
    .A2(_10686_),
    .B(_10699_),
    .Y(_03598_));
 OR3x1_ASAP7_75t_R _31388_ (.A(_08588_),
    .B(_08589_),
    .C(_10655_),
    .Y(_10700_));
 BUFx6f_ASAP7_75t_R _31389_ (.A(_10700_),
    .Y(_10701_));
 BUFx6f_ASAP7_75t_R _31390_ (.A(_10701_),
    .Y(_10702_));
 AND3x1_ASAP7_75t_R _31391_ (.A(_08595_),
    .B(_09651_),
    .C(_10660_),
    .Y(_10703_));
 BUFx4f_ASAP7_75t_R _31392_ (.A(_10703_),
    .Y(_10704_));
 OA211x2_ASAP7_75t_R _31393_ (.A1(_08346_),
    .A2(_08556_),
    .B(_08583_),
    .C(_10704_),
    .Y(_10705_));
 AOI21x1_ASAP7_75t_R _31394_ (.A1(_00439_),
    .A2(_10702_),
    .B(_10705_),
    .Y(_03599_));
 BUFx10_ASAP7_75t_R _31395_ (.A(_10701_),
    .Y(_10706_));
 NAND2x1_ASAP7_75t_R _31396_ (.A(_00392_),
    .B(_10706_),
    .Y(_10707_));
 OA21x2_ASAP7_75t_R _31397_ (.A1(_09676_),
    .A2(_10702_),
    .B(_10707_),
    .Y(_03600_));
 NOR2x1_ASAP7_75t_R _31398_ (.A(_00450_),
    .B(_10636_),
    .Y(_10708_));
 AO21x1_ASAP7_75t_R _31399_ (.A1(_10384_),
    .A2(_10549_),
    .B(_10708_),
    .Y(_03601_));
 NAND2x1_ASAP7_75t_R _31400_ (.A(_00503_),
    .B(_10706_),
    .Y(_10709_));
 OA21x2_ASAP7_75t_R _31401_ (.A1(_09696_),
    .A2(_10702_),
    .B(_10709_),
    .Y(_03602_));
 NAND2x1_ASAP7_75t_R _31402_ (.A(_00534_),
    .B(_10706_),
    .Y(_10710_));
 OA21x2_ASAP7_75t_R _31403_ (.A1(_09716_),
    .A2(_10702_),
    .B(_10710_),
    .Y(_03603_));
 AND2x4_ASAP7_75t_R _31404_ (.A(_08341_),
    .B(_10660_),
    .Y(_10711_));
 NOR2x1_ASAP7_75t_R _31405_ (.A(_00564_),
    .B(_10704_),
    .Y(_10712_));
 AO21x1_ASAP7_75t_R _31406_ (.A1(_08676_),
    .A2(_10711_),
    .B(_10712_),
    .Y(_03604_));
 NAND2x1_ASAP7_75t_R _31407_ (.A(_00596_),
    .B(_10706_),
    .Y(_10713_));
 OA21x2_ASAP7_75t_R _31408_ (.A1(_08763_),
    .A2(_10702_),
    .B(_10713_),
    .Y(_03605_));
 BUFx12f_ASAP7_75t_R _31409_ (.A(_10701_),
    .Y(_10714_));
 NAND2x1_ASAP7_75t_R _31410_ (.A(_00626_),
    .B(_10714_),
    .Y(_10715_));
 OA21x2_ASAP7_75t_R _31411_ (.A1(_08810_),
    .A2(_10702_),
    .B(_10715_),
    .Y(_03606_));
 NAND2x1_ASAP7_75t_R _31412_ (.A(_00656_),
    .B(_10714_),
    .Y(_10716_));
 OA21x2_ASAP7_75t_R _31413_ (.A1(_08851_),
    .A2(_10702_),
    .B(_10716_),
    .Y(_03607_));
 OR3x1_ASAP7_75t_R _31414_ (.A(_09790_),
    .B(_09791_),
    .C(_10701_),
    .Y(_10717_));
 OAI21x1_ASAP7_75t_R _31415_ (.A1(_00686_),
    .A2(_10704_),
    .B(_10717_),
    .Y(_03608_));
 NAND2x1_ASAP7_75t_R _31416_ (.A(_00716_),
    .B(_10714_),
    .Y(_10718_));
 OA21x2_ASAP7_75t_R _31417_ (.A1(_08943_),
    .A2(_10702_),
    .B(_10718_),
    .Y(_03609_));
 NAND2x1_ASAP7_75t_R _31418_ (.A(_00746_),
    .B(_10714_),
    .Y(_10719_));
 OA21x2_ASAP7_75t_R _31419_ (.A1(_08989_),
    .A2(_10702_),
    .B(_10719_),
    .Y(_03610_));
 NAND2x1_ASAP7_75t_R _31420_ (.A(_00776_),
    .B(_10714_),
    .Y(_10720_));
 OA21x2_ASAP7_75t_R _31421_ (.A1(_09728_),
    .A2(_10702_),
    .B(_10720_),
    .Y(_03611_));
 NOR2x1_ASAP7_75t_R _31422_ (.A(_00825_),
    .B(_10636_),
    .Y(_10721_));
 AO21x1_ASAP7_75t_R _31423_ (.A1(_10387_),
    .A2(_10549_),
    .B(_10721_),
    .Y(_03612_));
 BUFx6f_ASAP7_75t_R _31424_ (.A(_10701_),
    .Y(_10722_));
 NAND2x1_ASAP7_75t_R _31425_ (.A(_00472_),
    .B(_10714_),
    .Y(_10723_));
 OA21x2_ASAP7_75t_R _31426_ (.A1(_09074_),
    .A2(_10722_),
    .B(_10723_),
    .Y(_03613_));
 NAND2x1_ASAP7_75t_R _31427_ (.A(_00847_),
    .B(_10714_),
    .Y(_10724_));
 OA21x2_ASAP7_75t_R _31428_ (.A1(_09104_),
    .A2(_10722_),
    .B(_10724_),
    .Y(_03614_));
 NAND2x1_ASAP7_75t_R _31429_ (.A(_00880_),
    .B(_10714_),
    .Y(_10725_));
 OA21x2_ASAP7_75t_R _31430_ (.A1(_09144_),
    .A2(_10722_),
    .B(_10725_),
    .Y(_03615_));
 NAND2x1_ASAP7_75t_R _31431_ (.A(_00913_),
    .B(_10714_),
    .Y(_10726_));
 OA21x2_ASAP7_75t_R _31432_ (.A1(_09181_),
    .A2(_10722_),
    .B(_10726_),
    .Y(_03616_));
 NAND2x1_ASAP7_75t_R _31433_ (.A(_00946_),
    .B(_10714_),
    .Y(_10727_));
 OA21x2_ASAP7_75t_R _31434_ (.A1(_09738_),
    .A2(_10722_),
    .B(_10727_),
    .Y(_03617_));
 BUFx10_ASAP7_75t_R _31435_ (.A(_10701_),
    .Y(_10728_));
 NAND2x1_ASAP7_75t_R _31436_ (.A(_00979_),
    .B(_10728_),
    .Y(_10729_));
 OA21x2_ASAP7_75t_R _31437_ (.A1(_09245_),
    .A2(_10722_),
    .B(_10729_),
    .Y(_03618_));
 NAND2x1_ASAP7_75t_R _31438_ (.A(_01012_),
    .B(_10728_),
    .Y(_10730_));
 OA21x2_ASAP7_75t_R _31439_ (.A1(_09271_),
    .A2(_10722_),
    .B(_10730_),
    .Y(_03619_));
 NAND2x1_ASAP7_75t_R _31440_ (.A(_01045_),
    .B(_10728_),
    .Y(_10731_));
 OA21x2_ASAP7_75t_R _31441_ (.A1(_09299_),
    .A2(_10722_),
    .B(_10731_),
    .Y(_03620_));
 NAND2x1_ASAP7_75t_R _31442_ (.A(_01078_),
    .B(_10728_),
    .Y(_10732_));
 OA21x2_ASAP7_75t_R _31443_ (.A1(_09328_),
    .A2(_10722_),
    .B(_10732_),
    .Y(_03621_));
 NAND2x1_ASAP7_75t_R _31444_ (.A(_01111_),
    .B(_10728_),
    .Y(_10733_));
 OA21x2_ASAP7_75t_R _31445_ (.A1(_09357_),
    .A2(_10722_),
    .B(_10733_),
    .Y(_03622_));
 BUFx4f_ASAP7_75t_R _31446_ (.A(_10532_),
    .Y(_10734_));
 NOR2x1_ASAP7_75t_R _31447_ (.A(_00858_),
    .B(_10636_),
    .Y(_10735_));
 AO21x1_ASAP7_75t_R _31448_ (.A1(_10389_),
    .A2(_10734_),
    .B(_10735_),
    .Y(_03623_));
 NAND2x1_ASAP7_75t_R _31449_ (.A(_01144_),
    .B(_10728_),
    .Y(_10736_));
 OA21x2_ASAP7_75t_R _31450_ (.A1(_09390_),
    .A2(_10706_),
    .B(_10736_),
    .Y(_03624_));
 NAND2x1_ASAP7_75t_R _31451_ (.A(_01177_),
    .B(_10728_),
    .Y(_10737_));
 OA21x2_ASAP7_75t_R _31452_ (.A1(_09416_),
    .A2(_10706_),
    .B(_10737_),
    .Y(_03625_));
 NAND2x1_ASAP7_75t_R _31453_ (.A(_01210_),
    .B(_10728_),
    .Y(_10738_));
 OA21x2_ASAP7_75t_R _31454_ (.A1(_09442_),
    .A2(_10706_),
    .B(_10738_),
    .Y(_03626_));
 NAND2x1_ASAP7_75t_R _31455_ (.A(_01243_),
    .B(_10728_),
    .Y(_10739_));
 OA21x2_ASAP7_75t_R _31456_ (.A1(_09472_),
    .A2(_10706_),
    .B(_10739_),
    .Y(_03627_));
 NAND2x1_ASAP7_75t_R _31457_ (.A(_01276_),
    .B(_10728_),
    .Y(_10740_));
 OA21x2_ASAP7_75t_R _31458_ (.A1(_09495_),
    .A2(_10706_),
    .B(_10740_),
    .Y(_03628_));
 NOR2x1_ASAP7_75t_R _31459_ (.A(_01309_),
    .B(_10704_),
    .Y(_10741_));
 AO21x1_ASAP7_75t_R _31460_ (.A1(_10305_),
    .A2(_10711_),
    .B(_10741_),
    .Y(_03629_));
 NOR2x1_ASAP7_75t_R _31461_ (.A(_01342_),
    .B(_10704_),
    .Y(_10742_));
 AO21x1_ASAP7_75t_R _31462_ (.A1(net95),
    .A2(_10711_),
    .B(_10742_),
    .Y(_03630_));
 NAND2x1_ASAP7_75t_R _31463_ (.A(_01375_),
    .B(_10701_),
    .Y(_10743_));
 OA21x2_ASAP7_75t_R _31464_ (.A1(net6),
    .A2(_10706_),
    .B(_10743_),
    .Y(_03631_));
 NOR2x1_ASAP7_75t_R _31465_ (.A(_01408_),
    .B(_10704_),
    .Y(_10744_));
 AO21x1_ASAP7_75t_R _31466_ (.A1(net151),
    .A2(_10711_),
    .B(_10744_),
    .Y(_03632_));
 AND2x2_ASAP7_75t_R _31467_ (.A(_04826_),
    .B(_10701_),
    .Y(_10745_));
 AO21x1_ASAP7_75t_R _31468_ (.A1(net7),
    .A2(_10711_),
    .B(_10745_),
    .Y(_03633_));
 NOR2x1_ASAP7_75t_R _31469_ (.A(_00891_),
    .B(_10636_),
    .Y(_10746_));
 AO21x1_ASAP7_75t_R _31470_ (.A1(_10391_),
    .A2(_10734_),
    .B(_10746_),
    .Y(_03634_));
 NAND2x1_ASAP7_75t_R _31471_ (.A(_01785_),
    .B(_09106_),
    .Y(_10747_));
 OA21x2_ASAP7_75t_R _31472_ (.A1(_08591_),
    .A2(_09788_),
    .B(_10747_),
    .Y(_03635_));
 OR3x1_ASAP7_75t_R _31473_ (.A(_09766_),
    .B(_09767_),
    .C(_10655_),
    .Y(_10748_));
 BUFx6f_ASAP7_75t_R _31474_ (.A(_10748_),
    .Y(_10749_));
 BUFx12_ASAP7_75t_R _31475_ (.A(_10749_),
    .Y(_10750_));
 BUFx6f_ASAP7_75t_R _31476_ (.A(_10749_),
    .Y(_10751_));
 NAND2x1_ASAP7_75t_R _31477_ (.A(_00440_),
    .B(_10751_),
    .Y(_10752_));
 OA21x2_ASAP7_75t_R _31478_ (.A1(_08585_),
    .A2(_10750_),
    .B(_10752_),
    .Y(_03636_));
 BUFx16f_ASAP7_75t_R _31479_ (.A(_10749_),
    .Y(_10753_));
 NAND2x1_ASAP7_75t_R _31480_ (.A(_00393_),
    .B(_10753_),
    .Y(_10754_));
 OA21x2_ASAP7_75t_R _31481_ (.A1(_09676_),
    .A2(_10750_),
    .B(_10754_),
    .Y(_03637_));
 NAND2x1_ASAP7_75t_R _31482_ (.A(_00504_),
    .B(_10753_),
    .Y(_10755_));
 OA21x2_ASAP7_75t_R _31483_ (.A1(_09696_),
    .A2(_10750_),
    .B(_10755_),
    .Y(_03638_));
 AND3x1_ASAP7_75t_R _31484_ (.A(_08339_),
    .B(_09774_),
    .C(_10660_),
    .Y(_10756_));
 BUFx6f_ASAP7_75t_R _31485_ (.A(_10756_),
    .Y(_10757_));
 BUFx6f_ASAP7_75t_R _31486_ (.A(_10757_),
    .Y(_10758_));
 BUFx10_ASAP7_75t_R _31487_ (.A(_10749_),
    .Y(_10759_));
 AND2x2_ASAP7_75t_R _31488_ (.A(_14972_),
    .B(_10759_),
    .Y(_10760_));
 AO21x1_ASAP7_75t_R _31489_ (.A1(_10368_),
    .A2(_10758_),
    .B(_10760_),
    .Y(_03639_));
 AND2x2_ASAP7_75t_R _31490_ (.A(_14279_),
    .B(_10759_),
    .Y(_10761_));
 AO21x1_ASAP7_75t_R _31491_ (.A1(_08676_),
    .A2(_10758_),
    .B(_10761_),
    .Y(_03640_));
 NAND2x1_ASAP7_75t_R _31492_ (.A(_00597_),
    .B(_10753_),
    .Y(_10762_));
 OA21x2_ASAP7_75t_R _31493_ (.A1(_08763_),
    .A2(_10750_),
    .B(_10762_),
    .Y(_03641_));
 AND2x2_ASAP7_75t_R _31494_ (.A(_14399_),
    .B(_10759_),
    .Y(_10763_));
 AO21x1_ASAP7_75t_R _31495_ (.A1(_10373_),
    .A2(_10758_),
    .B(_10763_),
    .Y(_03642_));
 AND2x2_ASAP7_75t_R _31496_ (.A(_15229_),
    .B(_10749_),
    .Y(_10764_));
 AO21x1_ASAP7_75t_R _31497_ (.A1(_10375_),
    .A2(_10758_),
    .B(_10764_),
    .Y(_03643_));
 OR2x2_ASAP7_75t_R _31498_ (.A(_00687_),
    .B(_10757_),
    .Y(_10765_));
 OAI21x1_ASAP7_75t_R _31499_ (.A1(_10279_),
    .A2(_10750_),
    .B(_10765_),
    .Y(_03644_));
 AND2x2_ASAP7_75t_R _31500_ (.A(_15385_),
    .B(_10749_),
    .Y(_10766_));
 AO21x1_ASAP7_75t_R _31501_ (.A1(_10436_),
    .A2(_10758_),
    .B(_10766_),
    .Y(_03645_));
 NOR2x1_ASAP7_75t_R _31502_ (.A(_00924_),
    .B(_10636_),
    .Y(_10767_));
 AO21x1_ASAP7_75t_R _31503_ (.A1(_10238_),
    .A2(_10734_),
    .B(_10767_),
    .Y(_03646_));
 AND2x2_ASAP7_75t_R _31504_ (.A(_14631_),
    .B(_10749_),
    .Y(_10768_));
 AO21x1_ASAP7_75t_R _31505_ (.A1(_10379_),
    .A2(_10758_),
    .B(_10768_),
    .Y(_03647_));
 AND2x2_ASAP7_75t_R _31506_ (.A(_14692_),
    .B(_10749_),
    .Y(_10769_));
 AO21x1_ASAP7_75t_R _31507_ (.A1(_10381_),
    .A2(_10758_),
    .B(_10769_),
    .Y(_03648_));
 NAND2x1_ASAP7_75t_R _31508_ (.A(_00473_),
    .B(_10753_),
    .Y(_10770_));
 OA21x2_ASAP7_75t_R _31509_ (.A1(_09074_),
    .A2(_10750_),
    .B(_10770_),
    .Y(_03649_));
 NAND2x1_ASAP7_75t_R _31510_ (.A(_00848_),
    .B(_10753_),
    .Y(_10771_));
 OA21x2_ASAP7_75t_R _31511_ (.A1(_09104_),
    .A2(_10750_),
    .B(_10771_),
    .Y(_03650_));
 NAND2x1_ASAP7_75t_R _31512_ (.A(_00881_),
    .B(_10753_),
    .Y(_10772_));
 OA21x2_ASAP7_75t_R _31513_ (.A1(_09144_),
    .A2(_10750_),
    .B(_10772_),
    .Y(_03651_));
 NAND2x1_ASAP7_75t_R _31514_ (.A(_00914_),
    .B(_10753_),
    .Y(_10773_));
 OA21x2_ASAP7_75t_R _31515_ (.A1(_09181_),
    .A2(_10750_),
    .B(_10773_),
    .Y(_03652_));
 NOR2x1_ASAP7_75t_R _31516_ (.A(_00947_),
    .B(_10757_),
    .Y(_10774_));
 AO21x1_ASAP7_75t_R _31517_ (.A1(_09213_),
    .A2(_10758_),
    .B(_10774_),
    .Y(_03653_));
 NAND2x1_ASAP7_75t_R _31518_ (.A(_00980_),
    .B(_10753_),
    .Y(_10775_));
 OA21x2_ASAP7_75t_R _31519_ (.A1(_09245_),
    .A2(_10750_),
    .B(_10775_),
    .Y(_03654_));
 NAND2x1_ASAP7_75t_R _31520_ (.A(_01013_),
    .B(_10753_),
    .Y(_10776_));
 OA21x2_ASAP7_75t_R _31521_ (.A1(_09271_),
    .A2(_10751_),
    .B(_10776_),
    .Y(_03655_));
 NAND2x1_ASAP7_75t_R _31522_ (.A(_01046_),
    .B(_10753_),
    .Y(_10777_));
 OA21x2_ASAP7_75t_R _31523_ (.A1(_09299_),
    .A2(_10751_),
    .B(_10777_),
    .Y(_03656_));
 NOR2x1_ASAP7_75t_R _31524_ (.A(_00957_),
    .B(_10636_),
    .Y(_10778_));
 AO21x1_ASAP7_75t_R _31525_ (.A1(_10395_),
    .A2(_10734_),
    .B(_10778_),
    .Y(_03657_));
 NAND2x1_ASAP7_75t_R _31526_ (.A(_01079_),
    .B(_10759_),
    .Y(_10779_));
 OA21x2_ASAP7_75t_R _31527_ (.A1(_09328_),
    .A2(_10751_),
    .B(_10779_),
    .Y(_03658_));
 NAND2x1_ASAP7_75t_R _31528_ (.A(_01112_),
    .B(_10759_),
    .Y(_10780_));
 OA21x2_ASAP7_75t_R _31529_ (.A1(_09357_),
    .A2(_10751_),
    .B(_10780_),
    .Y(_03659_));
 NOR2x1_ASAP7_75t_R _31530_ (.A(_01145_),
    .B(_10757_),
    .Y(_10781_));
 AO21x1_ASAP7_75t_R _31531_ (.A1(_10453_),
    .A2(_10758_),
    .B(_10781_),
    .Y(_03660_));
 NAND2x1_ASAP7_75t_R _31532_ (.A(_01178_),
    .B(_10759_),
    .Y(_10782_));
 OA21x2_ASAP7_75t_R _31533_ (.A1(_09416_),
    .A2(_10751_),
    .B(_10782_),
    .Y(_03661_));
 NAND2x1_ASAP7_75t_R _31534_ (.A(_01211_),
    .B(_10759_),
    .Y(_10783_));
 OA21x2_ASAP7_75t_R _31535_ (.A1(_09442_),
    .A2(_10751_),
    .B(_10783_),
    .Y(_03662_));
 NAND2x1_ASAP7_75t_R _31536_ (.A(_01244_),
    .B(_10759_),
    .Y(_10784_));
 OA21x2_ASAP7_75t_R _31537_ (.A1(_09472_),
    .A2(_10751_),
    .B(_10784_),
    .Y(_03663_));
 NAND2x1_ASAP7_75t_R _31538_ (.A(_01277_),
    .B(_10759_),
    .Y(_10785_));
 OA21x2_ASAP7_75t_R _31539_ (.A1(_09495_),
    .A2(_10751_),
    .B(_10785_),
    .Y(_03664_));
 NOR2x1_ASAP7_75t_R _31540_ (.A(_01310_),
    .B(_10757_),
    .Y(_10786_));
 AO21x1_ASAP7_75t_R _31541_ (.A1(_09512_),
    .A2(_10758_),
    .B(_10786_),
    .Y(_03665_));
 NOR2x1_ASAP7_75t_R _31542_ (.A(_01343_),
    .B(_10757_),
    .Y(_10787_));
 AO21x1_ASAP7_75t_R _31543_ (.A1(_09544_),
    .A2(_10757_),
    .B(_10787_),
    .Y(_03666_));
 NAND2x1_ASAP7_75t_R _31544_ (.A(_01376_),
    .B(_10759_),
    .Y(_10788_));
 OA21x2_ASAP7_75t_R _31545_ (.A1(net6),
    .A2(_10751_),
    .B(_10788_),
    .Y(_03667_));
 BUFx6f_ASAP7_75t_R _31546_ (.A(_10532_),
    .Y(_10789_));
 NOR2x1_ASAP7_75t_R _31547_ (.A(_00990_),
    .B(_10789_),
    .Y(_10790_));
 AO21x1_ASAP7_75t_R _31548_ (.A1(_10397_),
    .A2(_10734_),
    .B(_10790_),
    .Y(_03668_));
 NOR2x1_ASAP7_75t_R _31549_ (.A(_01409_),
    .B(_10757_),
    .Y(_10791_));
 AO21x1_ASAP7_75t_R _31550_ (.A1(_09622_),
    .A2(_10757_),
    .B(_10791_),
    .Y(_03669_));
 AND2x2_ASAP7_75t_R _31551_ (.A(_04771_),
    .B(_10749_),
    .Y(_10792_));
 AO21x1_ASAP7_75t_R _31552_ (.A1(_09648_),
    .A2(_10757_),
    .B(_10792_),
    .Y(_03670_));
 AND4x2_ASAP7_75t_R _31553_ (.A(_08329_),
    .B(_09773_),
    .C(_09834_),
    .D(_10660_),
    .Y(_10793_));
 BUFx6f_ASAP7_75t_R _31554_ (.A(_10793_),
    .Y(_10794_));
 INVx1_ASAP7_75t_R _31555_ (.A(_10794_),
    .Y(_10795_));
 OR4x2_ASAP7_75t_R _31556_ (.A(_08027_),
    .B(_08330_),
    .C(_08588_),
    .D(_10655_),
    .Y(_10796_));
 BUFx12_ASAP7_75t_R _31557_ (.A(_10796_),
    .Y(_10797_));
 NAND2x1_ASAP7_75t_R _31558_ (.A(_00441_),
    .B(_10797_),
    .Y(_10798_));
 OA21x2_ASAP7_75t_R _31559_ (.A1(_08585_),
    .A2(_10795_),
    .B(_10798_),
    .Y(_03671_));
 BUFx10_ASAP7_75t_R _31560_ (.A(_10793_),
    .Y(_10799_));
 BUFx6f_ASAP7_75t_R _31561_ (.A(_10799_),
    .Y(_10800_));
 NOR2x1_ASAP7_75t_R _31562_ (.A(_00394_),
    .B(_10794_),
    .Y(_10801_));
 AO21x1_ASAP7_75t_R _31563_ (.A1(_10361_),
    .A2(_10800_),
    .B(_10801_),
    .Y(_03672_));
 NAND2x1_ASAP7_75t_R _31564_ (.A(_00505_),
    .B(_10797_),
    .Y(_10802_));
 OA21x2_ASAP7_75t_R _31565_ (.A1(_09696_),
    .A2(_10797_),
    .B(_10802_),
    .Y(_03673_));
 NOR2x1_ASAP7_75t_R _31566_ (.A(_00536_),
    .B(_10794_),
    .Y(_10803_));
 AO21x1_ASAP7_75t_R _31567_ (.A1(_10368_),
    .A2(_10800_),
    .B(_10803_),
    .Y(_03674_));
 AND2x2_ASAP7_75t_R _31568_ (.A(_14282_),
    .B(_10796_),
    .Y(_10804_));
 AO21x1_ASAP7_75t_R _31569_ (.A1(_08676_),
    .A2(_10800_),
    .B(_10804_),
    .Y(_03675_));
 NAND2x1_ASAP7_75t_R _31570_ (.A(_00598_),
    .B(_10797_),
    .Y(_10805_));
 OA21x2_ASAP7_75t_R _31571_ (.A1(_08763_),
    .A2(_10797_),
    .B(_10805_),
    .Y(_03676_));
 BUFx12f_ASAP7_75t_R _31572_ (.A(_10793_),
    .Y(_10806_));
 NOR2x1_ASAP7_75t_R _31573_ (.A(_00628_),
    .B(_10806_),
    .Y(_10807_));
 AO21x1_ASAP7_75t_R _31574_ (.A1(_10373_),
    .A2(_10800_),
    .B(_10807_),
    .Y(_03677_));
 NOR2x1_ASAP7_75t_R _31575_ (.A(_00658_),
    .B(_10806_),
    .Y(_10808_));
 AO21x1_ASAP7_75t_R _31576_ (.A1(_10375_),
    .A2(_10800_),
    .B(_10808_),
    .Y(_03678_));
 NOR2x1_ASAP7_75t_R _31577_ (.A(_01023_),
    .B(_10789_),
    .Y(_10809_));
 AO21x1_ASAP7_75t_R _31578_ (.A1(_10399_),
    .A2(_10734_),
    .B(_10809_),
    .Y(_03679_));
 OR3x1_ASAP7_75t_R _31579_ (.A(_09790_),
    .B(_09791_),
    .C(_10797_),
    .Y(_10810_));
 OAI21x1_ASAP7_75t_R _31580_ (.A1(_00688_),
    .A2(_10800_),
    .B(_10810_),
    .Y(_03680_));
 NOR2x1_ASAP7_75t_R _31581_ (.A(_00718_),
    .B(_10806_),
    .Y(_10811_));
 AO21x1_ASAP7_75t_R _31582_ (.A1(_10436_),
    .A2(_10800_),
    .B(_10811_),
    .Y(_03681_));
 NOR2x1_ASAP7_75t_R _31583_ (.A(_00748_),
    .B(_10806_),
    .Y(_10812_));
 AO21x1_ASAP7_75t_R _31584_ (.A1(_10379_),
    .A2(_10800_),
    .B(_10812_),
    .Y(_03682_));
 NOR2x1_ASAP7_75t_R _31585_ (.A(_00778_),
    .B(_10806_),
    .Y(_10813_));
 AO21x1_ASAP7_75t_R _31586_ (.A1(_10381_),
    .A2(_10800_),
    .B(_10813_),
    .Y(_03683_));
 NOR2x1_ASAP7_75t_R _31587_ (.A(_00474_),
    .B(_10806_),
    .Y(_10814_));
 AO21x1_ASAP7_75t_R _31588_ (.A1(_10384_),
    .A2(_10800_),
    .B(_10814_),
    .Y(_03684_));
 BUFx4f_ASAP7_75t_R _31589_ (.A(_10799_),
    .Y(_10815_));
 NOR2x1_ASAP7_75t_R _31590_ (.A(_00849_),
    .B(_10806_),
    .Y(_10816_));
 AO21x1_ASAP7_75t_R _31591_ (.A1(_10387_),
    .A2(_10815_),
    .B(_10816_),
    .Y(_03685_));
 NOR2x1_ASAP7_75t_R _31592_ (.A(_00882_),
    .B(_10806_),
    .Y(_10817_));
 AO21x1_ASAP7_75t_R _31593_ (.A1(_10389_),
    .A2(_10815_),
    .B(_10817_),
    .Y(_03686_));
 NOR2x1_ASAP7_75t_R _31594_ (.A(_00915_),
    .B(_10806_),
    .Y(_10818_));
 AO21x1_ASAP7_75t_R _31595_ (.A1(_10391_),
    .A2(_10815_),
    .B(_10818_),
    .Y(_03687_));
 AND2x2_ASAP7_75t_R _31596_ (.A(_16080_),
    .B(_10796_),
    .Y(_10819_));
 AO21x1_ASAP7_75t_R _31597_ (.A1(_09213_),
    .A2(_10815_),
    .B(_10819_),
    .Y(_03688_));
 NOR2x1_ASAP7_75t_R _31598_ (.A(_00981_),
    .B(_10806_),
    .Y(_10820_));
 AO21x1_ASAP7_75t_R _31599_ (.A1(_10395_),
    .A2(_10815_),
    .B(_10820_),
    .Y(_03689_));
 NOR2x1_ASAP7_75t_R _31600_ (.A(_01056_),
    .B(_10789_),
    .Y(_10821_));
 AO21x1_ASAP7_75t_R _31601_ (.A1(_10401_),
    .A2(_10734_),
    .B(_10821_),
    .Y(_03690_));
 NOR2x1_ASAP7_75t_R _31602_ (.A(_01014_),
    .B(_10799_),
    .Y(_10822_));
 AO21x1_ASAP7_75t_R _31603_ (.A1(_10397_),
    .A2(_10815_),
    .B(_10822_),
    .Y(_03691_));
 NOR2x1_ASAP7_75t_R _31604_ (.A(_01047_),
    .B(_10799_),
    .Y(_10823_));
 AO21x1_ASAP7_75t_R _31605_ (.A1(_10399_),
    .A2(_10815_),
    .B(_10823_),
    .Y(_03692_));
 NOR2x1_ASAP7_75t_R _31606_ (.A(_01080_),
    .B(_10799_),
    .Y(_10824_));
 AO21x1_ASAP7_75t_R _31607_ (.A1(_10401_),
    .A2(_10815_),
    .B(_10824_),
    .Y(_03693_));
 NOR2x1_ASAP7_75t_R _31608_ (.A(_01113_),
    .B(_10799_),
    .Y(_10825_));
 AO21x1_ASAP7_75t_R _31609_ (.A1(_10403_),
    .A2(_10815_),
    .B(_10825_),
    .Y(_03694_));
 NOR2x1_ASAP7_75t_R _31610_ (.A(_01146_),
    .B(_10799_),
    .Y(_10826_));
 AO21x1_ASAP7_75t_R _31611_ (.A1(_10453_),
    .A2(_10815_),
    .B(_10826_),
    .Y(_03695_));
 NOR2x1_ASAP7_75t_R _31612_ (.A(_01179_),
    .B(_10799_),
    .Y(_10827_));
 AO21x1_ASAP7_75t_R _31613_ (.A1(_10406_),
    .A2(_10794_),
    .B(_10827_),
    .Y(_03696_));
 NAND2x1_ASAP7_75t_R _31614_ (.A(_01212_),
    .B(_10797_),
    .Y(_10828_));
 OA21x2_ASAP7_75t_R _31615_ (.A1(_09442_),
    .A2(_10797_),
    .B(_10828_),
    .Y(_03697_));
 NOR2x1_ASAP7_75t_R _31616_ (.A(_01245_),
    .B(_10799_),
    .Y(_10829_));
 AO21x1_ASAP7_75t_R _31617_ (.A1(_10409_),
    .A2(_10794_),
    .B(_10829_),
    .Y(_03698_));
 NOR2x1_ASAP7_75t_R _31618_ (.A(_01278_),
    .B(_10799_),
    .Y(_10830_));
 AO21x1_ASAP7_75t_R _31619_ (.A1(_10412_),
    .A2(_10794_),
    .B(_10830_),
    .Y(_03699_));
 AND2x2_ASAP7_75t_R _31620_ (.A(_04330_),
    .B(_10796_),
    .Y(_10831_));
 AO21x1_ASAP7_75t_R _31621_ (.A1(_09512_),
    .A2(_10794_),
    .B(_10831_),
    .Y(_03700_));
 NOR2x1_ASAP7_75t_R _31622_ (.A(_01089_),
    .B(_10789_),
    .Y(_10832_));
 AO21x1_ASAP7_75t_R _31623_ (.A1(_10403_),
    .A2(_10734_),
    .B(_10832_),
    .Y(_03701_));
 AND2x2_ASAP7_75t_R _31624_ (.A(_04460_),
    .B(_10796_),
    .Y(_10833_));
 AO21x1_ASAP7_75t_R _31625_ (.A1(_09544_),
    .A2(_10794_),
    .B(_10833_),
    .Y(_03702_));
 NAND2x1_ASAP7_75t_R _31626_ (.A(_01377_),
    .B(_10797_),
    .Y(_10834_));
 OA21x2_ASAP7_75t_R _31627_ (.A1(net6),
    .A2(_10797_),
    .B(_10834_),
    .Y(_03703_));
 AND2x2_ASAP7_75t_R _31628_ (.A(_04684_),
    .B(_10796_),
    .Y(_10835_));
 AO21x1_ASAP7_75t_R _31629_ (.A1(_09622_),
    .A2(_10794_),
    .B(_10835_),
    .Y(_03704_));
 AND2x2_ASAP7_75t_R _31630_ (.A(_04768_),
    .B(_10796_),
    .Y(_10836_));
 AO21x1_ASAP7_75t_R _31631_ (.A1(_09648_),
    .A2(_10794_),
    .B(_10836_),
    .Y(_03705_));
 OR3x2_ASAP7_75t_R _31632_ (.A(_14049_),
    .B(_14050_),
    .C(_14231_),
    .Y(_10837_));
 OR3x1_ASAP7_75t_R _31633_ (.A(_08677_),
    .B(_08588_),
    .C(_10837_),
    .Y(_10838_));
 BUFx10_ASAP7_75t_R _31634_ (.A(_10838_),
    .Y(_10839_));
 BUFx6f_ASAP7_75t_R _31635_ (.A(_10839_),
    .Y(_10840_));
 BUFx12f_ASAP7_75t_R _31636_ (.A(_10839_),
    .Y(_10841_));
 NAND2x1_ASAP7_75t_R _31637_ (.A(_00442_),
    .B(_10841_),
    .Y(_10842_));
 OA21x2_ASAP7_75t_R _31638_ (.A1(_08585_),
    .A2(_10840_),
    .B(_10842_),
    .Y(_03706_));
 NAND2x1_ASAP7_75t_R _31639_ (.A(_00395_),
    .B(_10841_),
    .Y(_10843_));
 OA21x2_ASAP7_75t_R _31640_ (.A1(_09676_),
    .A2(_10840_),
    .B(_10843_),
    .Y(_03707_));
 NAND2x1_ASAP7_75t_R _31641_ (.A(_00506_),
    .B(_10841_),
    .Y(_10844_));
 OA21x2_ASAP7_75t_R _31642_ (.A1(_09696_),
    .A2(_10840_),
    .B(_10844_),
    .Y(_03708_));
 BUFx12f_ASAP7_75t_R _31643_ (.A(_10839_),
    .Y(_10845_));
 NAND2x1_ASAP7_75t_R _31644_ (.A(_00537_),
    .B(_10845_),
    .Y(_10846_));
 OA21x2_ASAP7_75t_R _31645_ (.A1(_09716_),
    .A2(_10840_),
    .B(_10846_),
    .Y(_03709_));
 AND3x4_ASAP7_75t_R _31646_ (.A(_14153_),
    .B(_14303_),
    .C(_14232_),
    .Y(_10847_));
 AND4x2_ASAP7_75t_R _31647_ (.A(_08593_),
    .B(_08594_),
    .C(_08595_),
    .D(_10847_),
    .Y(_10848_));
 BUFx6f_ASAP7_75t_R _31648_ (.A(_10848_),
    .Y(_10849_));
 NOR2x1_ASAP7_75t_R _31649_ (.A(_00567_),
    .B(_10849_),
    .Y(_10850_));
 AO21x1_ASAP7_75t_R _31650_ (.A1(_08676_),
    .A2(_10849_),
    .B(_10850_),
    .Y(_03710_));
 NAND2x1_ASAP7_75t_R _31651_ (.A(_00599_),
    .B(_10845_),
    .Y(_10851_));
 OA21x2_ASAP7_75t_R _31652_ (.A1(_08763_),
    .A2(_10840_),
    .B(_10851_),
    .Y(_03711_));
 NOR2x1_ASAP7_75t_R _31653_ (.A(_01122_),
    .B(_10789_),
    .Y(_10852_));
 AO21x1_ASAP7_75t_R _31654_ (.A1(_10453_),
    .A2(_10734_),
    .B(_10852_),
    .Y(_03712_));
 NAND2x1_ASAP7_75t_R _31655_ (.A(_00629_),
    .B(_10845_),
    .Y(_10853_));
 OA21x2_ASAP7_75t_R _31656_ (.A1(_08810_),
    .A2(_10840_),
    .B(_10853_),
    .Y(_03713_));
 NAND2x1_ASAP7_75t_R _31657_ (.A(_00659_),
    .B(_10845_),
    .Y(_10854_));
 OA21x2_ASAP7_75t_R _31658_ (.A1(_08851_),
    .A2(_10840_),
    .B(_10854_),
    .Y(_03714_));
 NAND2x1_ASAP7_75t_R _31659_ (.A(_14501_),
    .B(_10841_),
    .Y(_10855_));
 OAI21x1_ASAP7_75t_R _31660_ (.A1(_10279_),
    .A2(_10840_),
    .B(_10855_),
    .Y(_03715_));
 AND2x2_ASAP7_75t_R _31661_ (.A(_14576_),
    .B(_10839_),
    .Y(_10856_));
 AO21x1_ASAP7_75t_R _31662_ (.A1(_10436_),
    .A2(_10849_),
    .B(_10856_),
    .Y(_03716_));
 NAND2x1_ASAP7_75t_R _31663_ (.A(_00749_),
    .B(_10845_),
    .Y(_10857_));
 OA21x2_ASAP7_75t_R _31664_ (.A1(_08989_),
    .A2(_10840_),
    .B(_10857_),
    .Y(_03717_));
 NAND2x1_ASAP7_75t_R _31665_ (.A(_00779_),
    .B(_10845_),
    .Y(_10858_));
 OA21x2_ASAP7_75t_R _31666_ (.A1(_09728_),
    .A2(_10840_),
    .B(_10858_),
    .Y(_03718_));
 BUFx6f_ASAP7_75t_R _31667_ (.A(_10839_),
    .Y(_10859_));
 NAND2x1_ASAP7_75t_R _31668_ (.A(_00475_),
    .B(_10845_),
    .Y(_10860_));
 OA21x2_ASAP7_75t_R _31669_ (.A1(_09074_),
    .A2(_10859_),
    .B(_10860_),
    .Y(_03719_));
 NAND2x1_ASAP7_75t_R _31670_ (.A(_00850_),
    .B(_10845_),
    .Y(_10861_));
 OA21x2_ASAP7_75t_R _31671_ (.A1(_09104_),
    .A2(_10859_),
    .B(_10861_),
    .Y(_03720_));
 NAND2x1_ASAP7_75t_R _31672_ (.A(_00883_),
    .B(_10845_),
    .Y(_10862_));
 OA21x2_ASAP7_75t_R _31673_ (.A1(_09144_),
    .A2(_10859_),
    .B(_10862_),
    .Y(_03721_));
 NAND2x1_ASAP7_75t_R _31674_ (.A(_00916_),
    .B(_10845_),
    .Y(_10863_));
 OA21x2_ASAP7_75t_R _31675_ (.A1(_09181_),
    .A2(_10859_),
    .B(_10863_),
    .Y(_03722_));
 NOR2x1_ASAP7_75t_R _31676_ (.A(_01155_),
    .B(_10789_),
    .Y(_10864_));
 AO21x1_ASAP7_75t_R _31677_ (.A1(_10406_),
    .A2(_10734_),
    .B(_10864_),
    .Y(_03723_));
 NOR2x1_ASAP7_75t_R _31678_ (.A(_00949_),
    .B(_10849_),
    .Y(_10865_));
 AO21x1_ASAP7_75t_R _31679_ (.A1(_09213_),
    .A2(_10849_),
    .B(_10865_),
    .Y(_03724_));
 BUFx12_ASAP7_75t_R _31680_ (.A(_10839_),
    .Y(_10866_));
 NAND2x1_ASAP7_75t_R _31681_ (.A(_00982_),
    .B(_10866_),
    .Y(_10867_));
 OA21x2_ASAP7_75t_R _31682_ (.A1(_09245_),
    .A2(_10859_),
    .B(_10867_),
    .Y(_03725_));
 NAND2x1_ASAP7_75t_R _31683_ (.A(_01015_),
    .B(_10866_),
    .Y(_10868_));
 OA21x2_ASAP7_75t_R _31684_ (.A1(_09271_),
    .A2(_10859_),
    .B(_10868_),
    .Y(_03726_));
 NAND2x1_ASAP7_75t_R _31685_ (.A(_01048_),
    .B(_10866_),
    .Y(_10869_));
 OA21x2_ASAP7_75t_R _31686_ (.A1(_09299_),
    .A2(_10859_),
    .B(_10869_),
    .Y(_03727_));
 NAND2x1_ASAP7_75t_R _31687_ (.A(_01081_),
    .B(_10866_),
    .Y(_10870_));
 OA21x2_ASAP7_75t_R _31688_ (.A1(_09328_),
    .A2(_10859_),
    .B(_10870_),
    .Y(_03728_));
 NAND2x1_ASAP7_75t_R _31689_ (.A(_01114_),
    .B(_10866_),
    .Y(_10871_));
 OA21x2_ASAP7_75t_R _31690_ (.A1(_09357_),
    .A2(_10859_),
    .B(_10871_),
    .Y(_03729_));
 NAND2x1_ASAP7_75t_R _31691_ (.A(_01147_),
    .B(_10866_),
    .Y(_10872_));
 OA21x2_ASAP7_75t_R _31692_ (.A1(_09390_),
    .A2(_10859_),
    .B(_10872_),
    .Y(_03730_));
 NAND2x1_ASAP7_75t_R _31693_ (.A(_01180_),
    .B(_10866_),
    .Y(_10873_));
 OA21x2_ASAP7_75t_R _31694_ (.A1(_09416_),
    .A2(_10841_),
    .B(_10873_),
    .Y(_03731_));
 NAND2x1_ASAP7_75t_R _31695_ (.A(_01213_),
    .B(_10866_),
    .Y(_10874_));
 OA21x2_ASAP7_75t_R _31696_ (.A1(_09442_),
    .A2(_10841_),
    .B(_10874_),
    .Y(_03732_));
 NAND2x1_ASAP7_75t_R _31697_ (.A(_01246_),
    .B(_10866_),
    .Y(_10875_));
 OA21x2_ASAP7_75t_R _31698_ (.A1(_09472_),
    .A2(_10841_),
    .B(_10875_),
    .Y(_03733_));
 NAND2x1_ASAP7_75t_R _31699_ (.A(_01188_),
    .B(_10535_),
    .Y(_10876_));
 OA21x2_ASAP7_75t_R _31700_ (.A1(_09442_),
    .A2(_10533_),
    .B(_10876_),
    .Y(_03734_));
 NAND2x1_ASAP7_75t_R _31701_ (.A(_01279_),
    .B(_10866_),
    .Y(_10877_));
 OA21x2_ASAP7_75t_R _31702_ (.A1(_09495_),
    .A2(_10841_),
    .B(_10877_),
    .Y(_03735_));
 INVx1_ASAP7_75t_R _31703_ (.A(_01312_),
    .Y(_10878_));
 AND3x1_ASAP7_75t_R _31704_ (.A(_09508_),
    .B(_09511_),
    .C(_10848_),
    .Y(_10879_));
 AO21x1_ASAP7_75t_R _31705_ (.A1(_10878_),
    .A2(_10841_),
    .B(_10879_),
    .Y(_03736_));
 NOR2x1_ASAP7_75t_R _31706_ (.A(_01345_),
    .B(_10849_),
    .Y(_10880_));
 AO21x1_ASAP7_75t_R _31707_ (.A1(_09544_),
    .A2(_10849_),
    .B(_10880_),
    .Y(_03737_));
 NAND2x1_ASAP7_75t_R _31708_ (.A(_01378_),
    .B(_10839_),
    .Y(_10881_));
 OA21x2_ASAP7_75t_R _31709_ (.A1(net6),
    .A2(_10841_),
    .B(_10881_),
    .Y(_03738_));
 NOR2x1_ASAP7_75t_R _31710_ (.A(_01411_),
    .B(_10849_),
    .Y(_10882_));
 AO21x1_ASAP7_75t_R _31711_ (.A1(_09622_),
    .A2(_10849_),
    .B(_10882_),
    .Y(_03739_));
 NOR2x1_ASAP7_75t_R _31712_ (.A(_01444_),
    .B(_10848_),
    .Y(_10883_));
 AO21x1_ASAP7_75t_R _31713_ (.A1(_09648_),
    .A2(_10849_),
    .B(_10883_),
    .Y(_03740_));
 NAND2x2_ASAP7_75t_R _31714_ (.A(_08341_),
    .B(_10847_),
    .Y(_10884_));
 OR3x2_ASAP7_75t_R _31715_ (.A(_09838_),
    .B(_08589_),
    .C(_10837_),
    .Y(_10885_));
 BUFx10_ASAP7_75t_R _31716_ (.A(_10885_),
    .Y(_10886_));
 NAND2x1_ASAP7_75t_R _31717_ (.A(_00443_),
    .B(_10886_),
    .Y(_10887_));
 OA21x2_ASAP7_75t_R _31718_ (.A1(_08585_),
    .A2(_10884_),
    .B(_10887_),
    .Y(_03741_));
 AND4x1_ASAP7_75t_R _31719_ (.A(_08329_),
    .B(_08330_),
    .C(_09834_),
    .D(_10847_),
    .Y(_10888_));
 BUFx10_ASAP7_75t_R _31720_ (.A(_10888_),
    .Y(_10889_));
 BUFx6f_ASAP7_75t_R _31721_ (.A(_10889_),
    .Y(_10890_));
 BUFx10_ASAP7_75t_R _31722_ (.A(_10889_),
    .Y(_10891_));
 NOR2x1_ASAP7_75t_R _31723_ (.A(_00396_),
    .B(_10891_),
    .Y(_10892_));
 AO21x1_ASAP7_75t_R _31724_ (.A1(_10361_),
    .A2(_10890_),
    .B(_10892_),
    .Y(_03742_));
 NAND2x1_ASAP7_75t_R _31725_ (.A(_00507_),
    .B(_10886_),
    .Y(_10893_));
 OA21x2_ASAP7_75t_R _31726_ (.A1(_09696_),
    .A2(_10886_),
    .B(_10893_),
    .Y(_03743_));
 NOR2x1_ASAP7_75t_R _31727_ (.A(_00538_),
    .B(_10891_),
    .Y(_10894_));
 AO21x1_ASAP7_75t_R _31728_ (.A1(_10368_),
    .A2(_10890_),
    .B(_10894_),
    .Y(_03744_));
 NOR2x1_ASAP7_75t_R _31729_ (.A(_01221_),
    .B(_10789_),
    .Y(_10895_));
 AO21x1_ASAP7_75t_R _31730_ (.A1(_10409_),
    .A2(_10550_),
    .B(_10895_),
    .Y(_03745_));
 OR2x2_ASAP7_75t_R _31731_ (.A(_01784_),
    .B(_09796_),
    .Y(_10896_));
 OAI21x1_ASAP7_75t_R _31732_ (.A1(_08342_),
    .A2(_08898_),
    .B(_10896_),
    .Y(_03746_));
 AND2x2_ASAP7_75t_R _31733_ (.A(_14244_),
    .B(_10885_),
    .Y(_10897_));
 AO21x1_ASAP7_75t_R _31734_ (.A1(_08676_),
    .A2(_10890_),
    .B(_10897_),
    .Y(_03747_));
 NAND2x1_ASAP7_75t_R _31735_ (.A(_00600_),
    .B(_10886_),
    .Y(_10898_));
 OA21x2_ASAP7_75t_R _31736_ (.A1(_08763_),
    .A2(_10886_),
    .B(_10898_),
    .Y(_03748_));
 NOR2x1_ASAP7_75t_R _31737_ (.A(_00630_),
    .B(_10891_),
    .Y(_10899_));
 AO21x1_ASAP7_75t_R _31738_ (.A1(_10373_),
    .A2(_10890_),
    .B(_10899_),
    .Y(_03749_));
 NOR2x1_ASAP7_75t_R _31739_ (.A(_00660_),
    .B(_10891_),
    .Y(_10900_));
 AO21x1_ASAP7_75t_R _31740_ (.A1(_10375_),
    .A2(_10890_),
    .B(_10900_),
    .Y(_03750_));
 NAND2x1_ASAP7_75t_R _31741_ (.A(_14530_),
    .B(_10886_),
    .Y(_10901_));
 OAI21x1_ASAP7_75t_R _31742_ (.A1(_10279_),
    .A2(_10884_),
    .B(_10901_),
    .Y(_03751_));
 BUFx12f_ASAP7_75t_R _31743_ (.A(_10889_),
    .Y(_10902_));
 NOR2x1_ASAP7_75t_R _31744_ (.A(_00720_),
    .B(_10902_),
    .Y(_10903_));
 AO21x1_ASAP7_75t_R _31745_ (.A1(_10436_),
    .A2(_10890_),
    .B(_10903_),
    .Y(_03752_));
 NOR2x1_ASAP7_75t_R _31746_ (.A(_00750_),
    .B(_10902_),
    .Y(_10904_));
 AO21x1_ASAP7_75t_R _31747_ (.A1(_10379_),
    .A2(_10890_),
    .B(_10904_),
    .Y(_03753_));
 NOR2x1_ASAP7_75t_R _31748_ (.A(_00780_),
    .B(_10902_),
    .Y(_10905_));
 AO21x1_ASAP7_75t_R _31749_ (.A1(_10381_),
    .A2(_10890_),
    .B(_10905_),
    .Y(_03754_));
 NOR2x1_ASAP7_75t_R _31750_ (.A(_00476_),
    .B(_10902_),
    .Y(_10906_));
 AO21x1_ASAP7_75t_R _31751_ (.A1(_10384_),
    .A2(_10890_),
    .B(_10906_),
    .Y(_03755_));
 NOR2x1_ASAP7_75t_R _31752_ (.A(_00851_),
    .B(_10902_),
    .Y(_10907_));
 AO21x1_ASAP7_75t_R _31753_ (.A1(_10387_),
    .A2(_10890_),
    .B(_10907_),
    .Y(_03756_));
 NOR2x1_ASAP7_75t_R _31754_ (.A(_01254_),
    .B(_10789_),
    .Y(_10908_));
 AO21x1_ASAP7_75t_R _31755_ (.A1(_10412_),
    .A2(_10550_),
    .B(_10908_),
    .Y(_03757_));
 BUFx4f_ASAP7_75t_R _31756_ (.A(_10889_),
    .Y(_10909_));
 NOR2x1_ASAP7_75t_R _31757_ (.A(_00884_),
    .B(_10902_),
    .Y(_10910_));
 AO21x1_ASAP7_75t_R _31758_ (.A1(_10389_),
    .A2(_10909_),
    .B(_10910_),
    .Y(_03758_));
 NOR2x1_ASAP7_75t_R _31759_ (.A(_00917_),
    .B(_10902_),
    .Y(_10911_));
 AO21x1_ASAP7_75t_R _31760_ (.A1(_10391_),
    .A2(_10909_),
    .B(_10911_),
    .Y(_03759_));
 NOR2x1_ASAP7_75t_R _31761_ (.A(_00950_),
    .B(_10902_),
    .Y(_10912_));
 AO21x1_ASAP7_75t_R _31762_ (.A1(_09213_),
    .A2(_10909_),
    .B(_10912_),
    .Y(_03760_));
 NOR2x1_ASAP7_75t_R _31763_ (.A(_00983_),
    .B(_10902_),
    .Y(_10913_));
 AO21x1_ASAP7_75t_R _31764_ (.A1(_10395_),
    .A2(_10909_),
    .B(_10913_),
    .Y(_03761_));
 NOR2x1_ASAP7_75t_R _31765_ (.A(_01016_),
    .B(_10902_),
    .Y(_10914_));
 AO21x1_ASAP7_75t_R _31766_ (.A1(_10397_),
    .A2(_10909_),
    .B(_10914_),
    .Y(_03762_));
 BUFx12_ASAP7_75t_R _31767_ (.A(_10889_),
    .Y(_10915_));
 NOR2x1_ASAP7_75t_R _31768_ (.A(_01049_),
    .B(_10915_),
    .Y(_10916_));
 AO21x1_ASAP7_75t_R _31769_ (.A1(_10399_),
    .A2(_10909_),
    .B(_10916_),
    .Y(_03763_));
 NOR2x1_ASAP7_75t_R _31770_ (.A(_01082_),
    .B(_10915_),
    .Y(_10917_));
 AO21x1_ASAP7_75t_R _31771_ (.A1(_10401_),
    .A2(_10909_),
    .B(_10917_),
    .Y(_03764_));
 NOR2x1_ASAP7_75t_R _31772_ (.A(_01115_),
    .B(_10915_),
    .Y(_10918_));
 AO21x1_ASAP7_75t_R _31773_ (.A1(_10403_),
    .A2(_10909_),
    .B(_10918_),
    .Y(_03765_));
 NOR2x1_ASAP7_75t_R _31774_ (.A(_01148_),
    .B(_10915_),
    .Y(_10919_));
 AO21x1_ASAP7_75t_R _31775_ (.A1(_10453_),
    .A2(_10909_),
    .B(_10919_),
    .Y(_03766_));
 NOR2x1_ASAP7_75t_R _31776_ (.A(_01181_),
    .B(_10915_),
    .Y(_10920_));
 AO21x1_ASAP7_75t_R _31777_ (.A1(_10406_),
    .A2(_10909_),
    .B(_10920_),
    .Y(_03767_));
 NOR2x1_ASAP7_75t_R _31778_ (.A(_01287_),
    .B(_10789_),
    .Y(_10921_));
 AO21x1_ASAP7_75t_R _31779_ (.A1(_09512_),
    .A2(_10550_),
    .B(_10921_),
    .Y(_03768_));
 NAND2x1_ASAP7_75t_R _31780_ (.A(_01214_),
    .B(_10886_),
    .Y(_10922_));
 OA21x2_ASAP7_75t_R _31781_ (.A1(_09442_),
    .A2(_10886_),
    .B(_10922_),
    .Y(_03769_));
 NOR2x1_ASAP7_75t_R _31782_ (.A(_01247_),
    .B(_10915_),
    .Y(_10923_));
 AO21x1_ASAP7_75t_R _31783_ (.A1(_10409_),
    .A2(_10891_),
    .B(_10923_),
    .Y(_03770_));
 NOR2x1_ASAP7_75t_R _31784_ (.A(_01280_),
    .B(_10915_),
    .Y(_10924_));
 AO21x1_ASAP7_75t_R _31785_ (.A1(_10412_),
    .A2(_10891_),
    .B(_10924_),
    .Y(_03771_));
 NOR2x1_ASAP7_75t_R _31786_ (.A(_01313_),
    .B(_10915_),
    .Y(_10925_));
 AO21x1_ASAP7_75t_R _31787_ (.A1(_09512_),
    .A2(_10891_),
    .B(_10925_),
    .Y(_03772_));
 NOR2x1_ASAP7_75t_R _31788_ (.A(_01346_),
    .B(_10915_),
    .Y(_10926_));
 AO21x1_ASAP7_75t_R _31789_ (.A1(net95),
    .A2(_10891_),
    .B(_10926_),
    .Y(_03773_));
 NAND2x1_ASAP7_75t_R _31790_ (.A(_01379_),
    .B(_10886_),
    .Y(_10927_));
 OA21x2_ASAP7_75t_R _31791_ (.A1(_09580_),
    .A2(_10886_),
    .B(_10927_),
    .Y(_03774_));
 NOR2x1_ASAP7_75t_R _31792_ (.A(_01412_),
    .B(_10915_),
    .Y(_10928_));
 AO21x1_ASAP7_75t_R _31793_ (.A1(net151),
    .A2(_10891_),
    .B(_10928_),
    .Y(_03775_));
 NOR2x1_ASAP7_75t_R _31794_ (.A(_01445_),
    .B(_10889_),
    .Y(_10929_));
 AO21x1_ASAP7_75t_R _31795_ (.A1(net7),
    .A2(_10891_),
    .B(_10929_),
    .Y(_03776_));
 OR3x1_ASAP7_75t_R _31796_ (.A(_09766_),
    .B(_09767_),
    .C(_10837_),
    .Y(_10930_));
 BUFx10_ASAP7_75t_R _31797_ (.A(_10930_),
    .Y(_10931_));
 BUFx12_ASAP7_75t_R _31798_ (.A(_10931_),
    .Y(_10932_));
 NAND2x1_ASAP7_75t_R _31799_ (.A(_00444_),
    .B(_10932_),
    .Y(_10933_));
 OA21x2_ASAP7_75t_R _31800_ (.A1(_08585_),
    .A2(_10932_),
    .B(_10933_),
    .Y(_03777_));
 AND3x1_ASAP7_75t_R _31801_ (.A(_08339_),
    .B(_09774_),
    .C(_10847_),
    .Y(_10934_));
 BUFx10_ASAP7_75t_R _31802_ (.A(_10934_),
    .Y(_10935_));
 BUFx6f_ASAP7_75t_R _31803_ (.A(_10935_),
    .Y(_10936_));
 BUFx6f_ASAP7_75t_R _31804_ (.A(_10931_),
    .Y(_10937_));
 AND2x2_ASAP7_75t_R _31805_ (.A(_13529_),
    .B(_10937_),
    .Y(_10938_));
 AO21x1_ASAP7_75t_R _31806_ (.A1(_10361_),
    .A2(_10936_),
    .B(_10938_),
    .Y(_03778_));
 NOR2x1_ASAP7_75t_R _31807_ (.A(_01320_),
    .B(_10789_),
    .Y(_10939_));
 AO21x1_ASAP7_75t_R _31808_ (.A1(_09544_),
    .A2(_10550_),
    .B(_10939_),
    .Y(_03779_));
 NAND2x1_ASAP7_75t_R _31809_ (.A(_00508_),
    .B(_10932_),
    .Y(_10940_));
 OA21x2_ASAP7_75t_R _31810_ (.A1(_09696_),
    .A2(_10932_),
    .B(_10940_),
    .Y(_03780_));
 AND2x2_ASAP7_75t_R _31811_ (.A(_14175_),
    .B(_10937_),
    .Y(_10941_));
 AO21x1_ASAP7_75t_R _31812_ (.A1(_10368_),
    .A2(_10936_),
    .B(_10941_),
    .Y(_03781_));
 AND2x2_ASAP7_75t_R _31813_ (.A(_14237_),
    .B(_10937_),
    .Y(_10942_));
 AO21x1_ASAP7_75t_R _31814_ (.A1(_08676_),
    .A2(_10936_),
    .B(_10942_),
    .Y(_03782_));
 NAND2x1_ASAP7_75t_R _31815_ (.A(_00601_),
    .B(_10932_),
    .Y(_10943_));
 OA21x2_ASAP7_75t_R _31816_ (.A1(_08763_),
    .A2(_10932_),
    .B(_10943_),
    .Y(_03783_));
 AND2x2_ASAP7_75t_R _31817_ (.A(_14396_),
    .B(_10937_),
    .Y(_10944_));
 AO21x1_ASAP7_75t_R _31818_ (.A1(_10373_),
    .A2(_10936_),
    .B(_10944_),
    .Y(_03784_));
 AND2x2_ASAP7_75t_R _31819_ (.A(_15216_),
    .B(_10937_),
    .Y(_10945_));
 AO21x1_ASAP7_75t_R _31820_ (.A1(_10375_),
    .A2(_10936_),
    .B(_10945_),
    .Y(_03785_));
 OR3x1_ASAP7_75t_R _31821_ (.A(_09790_),
    .B(_09791_),
    .C(_10932_),
    .Y(_10946_));
 OAI21x1_ASAP7_75t_R _31822_ (.A1(_00691_),
    .A2(_10936_),
    .B(_10946_),
    .Y(_03786_));
 AND2x2_ASAP7_75t_R _31823_ (.A(_14573_),
    .B(_10937_),
    .Y(_10947_));
 AO21x1_ASAP7_75t_R _31824_ (.A1(_10436_),
    .A2(_10936_),
    .B(_10947_),
    .Y(_03787_));
 AND2x2_ASAP7_75t_R _31825_ (.A(_14637_),
    .B(_10937_),
    .Y(_10948_));
 AO21x1_ASAP7_75t_R _31826_ (.A1(_10379_),
    .A2(_10936_),
    .B(_10948_),
    .Y(_03788_));
 AND2x2_ASAP7_75t_R _31827_ (.A(_14704_),
    .B(_10937_),
    .Y(_10949_));
 AO21x1_ASAP7_75t_R _31828_ (.A1(_10381_),
    .A2(_10936_),
    .B(_10949_),
    .Y(_03789_));
 NAND2x1_ASAP7_75t_R _31829_ (.A(_01353_),
    .B(_10535_),
    .Y(_10950_));
 OA21x2_ASAP7_75t_R _31830_ (.A1(net6),
    .A2(_10533_),
    .B(_10950_),
    .Y(_03790_));
 BUFx6f_ASAP7_75t_R _31831_ (.A(_10935_),
    .Y(_10951_));
 AND2x2_ASAP7_75t_R _31832_ (.A(_13992_),
    .B(_10937_),
    .Y(_10952_));
 AO21x1_ASAP7_75t_R _31833_ (.A1(_10384_),
    .A2(_10951_),
    .B(_10952_),
    .Y(_03791_));
 BUFx4f_ASAP7_75t_R _31834_ (.A(_10931_),
    .Y(_10953_));
 AND2x2_ASAP7_75t_R _31835_ (.A(_15643_),
    .B(_10953_),
    .Y(_10954_));
 AO21x1_ASAP7_75t_R _31836_ (.A1(_10387_),
    .A2(_10951_),
    .B(_10954_),
    .Y(_03792_));
 AND2x2_ASAP7_75t_R _31837_ (.A(_15793_),
    .B(_10953_),
    .Y(_10955_));
 AO21x1_ASAP7_75t_R _31838_ (.A1(_10389_),
    .A2(_10951_),
    .B(_10955_),
    .Y(_03793_));
 AND2x2_ASAP7_75t_R _31839_ (.A(_15924_),
    .B(_10953_),
    .Y(_10956_));
 AO21x1_ASAP7_75t_R _31840_ (.A1(_10391_),
    .A2(_10951_),
    .B(_10956_),
    .Y(_03794_));
 AND3x1_ASAP7_75t_R _31841_ (.A(_09204_),
    .B(_09212_),
    .C(_10935_),
    .Y(_10957_));
 AO21x1_ASAP7_75t_R _31842_ (.A1(_16071_),
    .A2(_10932_),
    .B(_10957_),
    .Y(_03795_));
 AND2x2_ASAP7_75t_R _31843_ (.A(_16188_),
    .B(_10953_),
    .Y(_10958_));
 AO21x1_ASAP7_75t_R _31844_ (.A1(_10395_),
    .A2(_10951_),
    .B(_10958_),
    .Y(_03796_));
 AND2x2_ASAP7_75t_R _31845_ (.A(_16332_),
    .B(_10953_),
    .Y(_10959_));
 AO21x1_ASAP7_75t_R _31846_ (.A1(_10397_),
    .A2(_10951_),
    .B(_10959_),
    .Y(_03797_));
 AND2x2_ASAP7_75t_R _31847_ (.A(_16445_),
    .B(_10953_),
    .Y(_10960_));
 AO21x1_ASAP7_75t_R _31848_ (.A1(_10399_),
    .A2(_10951_),
    .B(_10960_),
    .Y(_03798_));
 AND2x2_ASAP7_75t_R _31849_ (.A(_16571_),
    .B(_10953_),
    .Y(_10961_));
 AO21x1_ASAP7_75t_R _31850_ (.A1(_10401_),
    .A2(_10951_),
    .B(_10961_),
    .Y(_03799_));
 AND2x2_ASAP7_75t_R _31851_ (.A(_16685_),
    .B(_10953_),
    .Y(_10962_));
 AO21x1_ASAP7_75t_R _31852_ (.A1(_10403_),
    .A2(_10951_),
    .B(_10962_),
    .Y(_03800_));
 NOR2x1_ASAP7_75t_R _31853_ (.A(_01386_),
    .B(_10532_),
    .Y(_10963_));
 AO21x1_ASAP7_75t_R _31854_ (.A1(_09622_),
    .A2(_10550_),
    .B(_10963_),
    .Y(_03801_));
 AND2x2_ASAP7_75t_R _31855_ (.A(_16815_),
    .B(_10953_),
    .Y(_10964_));
 AO21x1_ASAP7_75t_R _31856_ (.A1(_10453_),
    .A2(_10951_),
    .B(_10964_),
    .Y(_03802_));
 AND2x2_ASAP7_75t_R _31857_ (.A(_16925_),
    .B(_10953_),
    .Y(_10965_));
 AO21x1_ASAP7_75t_R _31858_ (.A1(_10406_),
    .A2(_10935_),
    .B(_10965_),
    .Y(_03803_));
 NAND2x1_ASAP7_75t_R _31859_ (.A(_01215_),
    .B(_10932_),
    .Y(_10966_));
 OA21x2_ASAP7_75t_R _31860_ (.A1(_09442_),
    .A2(_10932_),
    .B(_10966_),
    .Y(_03804_));
 AND2x2_ASAP7_75t_R _31861_ (.A(_17164_),
    .B(_10931_),
    .Y(_10967_));
 AO21x1_ASAP7_75t_R _31862_ (.A1(_10409_),
    .A2(_10935_),
    .B(_10967_),
    .Y(_03805_));
 AND2x2_ASAP7_75t_R _31863_ (.A(_17295_),
    .B(_10931_),
    .Y(_10968_));
 AO21x1_ASAP7_75t_R _31864_ (.A1(_10412_),
    .A2(_10935_),
    .B(_10968_),
    .Y(_03806_));
 AND2x2_ASAP7_75t_R _31865_ (.A(_04322_),
    .B(_10931_),
    .Y(_10969_));
 AO21x1_ASAP7_75t_R _31866_ (.A1(_09512_),
    .A2(_10935_),
    .B(_10969_),
    .Y(_03807_));
 AND2x2_ASAP7_75t_R _31867_ (.A(_04452_),
    .B(_10931_),
    .Y(_10970_));
 AO21x1_ASAP7_75t_R _31868_ (.A1(net95),
    .A2(_10935_),
    .B(_10970_),
    .Y(_03808_));
 OR3x1_ASAP7_75t_R _31869_ (.A(_09578_),
    .B(_09572_),
    .C(_10937_),
    .Y(_10971_));
 OA21x2_ASAP7_75t_R _31870_ (.A1(_04562_),
    .A2(_10936_),
    .B(_10971_),
    .Y(_03809_));
 AND2x2_ASAP7_75t_R _31871_ (.A(_04676_),
    .B(_10931_),
    .Y(_10972_));
 AO21x1_ASAP7_75t_R _31872_ (.A1(net151),
    .A2(_10935_),
    .B(_10972_),
    .Y(_03810_));
 AND2x2_ASAP7_75t_R _31873_ (.A(_04794_),
    .B(_10931_),
    .Y(_10973_));
 AO21x1_ASAP7_75t_R _31874_ (.A1(net7),
    .A2(_10935_),
    .B(_10973_),
    .Y(_03811_));
 AND2x2_ASAP7_75t_R _31875_ (.A(_04835_),
    .B(_10535_),
    .Y(_10974_));
 AO21x1_ASAP7_75t_R _31876_ (.A1(_09648_),
    .A2(_10550_),
    .B(_10974_),
    .Y(_03812_));
 AND4x2_ASAP7_75t_R _31877_ (.A(_08329_),
    .B(_09773_),
    .C(_09834_),
    .D(_10847_),
    .Y(_10975_));
 BUFx10_ASAP7_75t_R _31878_ (.A(_10975_),
    .Y(_10976_));
 INVx1_ASAP7_75t_R _31879_ (.A(_10976_),
    .Y(_10977_));
 OR4x2_ASAP7_75t_R _31880_ (.A(_08593_),
    .B(_08594_),
    .C(_09838_),
    .D(_10837_),
    .Y(_10978_));
 BUFx12_ASAP7_75t_R _31881_ (.A(_10978_),
    .Y(_10979_));
 NAND2x1_ASAP7_75t_R _31882_ (.A(_00445_),
    .B(_10979_),
    .Y(_10980_));
 OA21x2_ASAP7_75t_R _31883_ (.A1(_08585_),
    .A2(_10977_),
    .B(_10980_),
    .Y(_03813_));
 BUFx4f_ASAP7_75t_R _31884_ (.A(_10976_),
    .Y(_10981_));
 BUFx6f_ASAP7_75t_R _31885_ (.A(_10975_),
    .Y(_10982_));
 NOR2x1_ASAP7_75t_R _31886_ (.A(_00398_),
    .B(_10982_),
    .Y(_10983_));
 AO21x1_ASAP7_75t_R _31887_ (.A1(_09675_),
    .A2(_10981_),
    .B(_10983_),
    .Y(_03814_));
 NAND2x1_ASAP7_75t_R _31888_ (.A(_00509_),
    .B(_10979_),
    .Y(_10984_));
 OA21x2_ASAP7_75t_R _31889_ (.A1(_09696_),
    .A2(_10979_),
    .B(_10984_),
    .Y(_03815_));
 NOR2x1_ASAP7_75t_R _31890_ (.A(_00540_),
    .B(_10982_),
    .Y(_10985_));
 AO21x1_ASAP7_75t_R _31891_ (.A1(_09715_),
    .A2(_10981_),
    .B(_10985_),
    .Y(_03816_));
 AND2x2_ASAP7_75t_R _31892_ (.A(_14241_),
    .B(_10978_),
    .Y(_10986_));
 AO21x1_ASAP7_75t_R _31893_ (.A1(_08676_),
    .A2(_10981_),
    .B(_10986_),
    .Y(_03817_));
 NAND2x1_ASAP7_75t_R _31894_ (.A(_00602_),
    .B(_10979_),
    .Y(_10987_));
 OA21x2_ASAP7_75t_R _31895_ (.A1(_08763_),
    .A2(_10979_),
    .B(_10987_),
    .Y(_03818_));
 NOR2x1_ASAP7_75t_R _31896_ (.A(_00632_),
    .B(_10982_),
    .Y(_10988_));
 AO21x1_ASAP7_75t_R _31897_ (.A1(_08809_),
    .A2(_10981_),
    .B(_10988_),
    .Y(_03819_));
 NOR2x1_ASAP7_75t_R _31898_ (.A(_00662_),
    .B(_10982_),
    .Y(_10989_));
 AO21x1_ASAP7_75t_R _31899_ (.A1(_08850_),
    .A2(_10981_),
    .B(_10989_),
    .Y(_03820_));
 NAND2x1_ASAP7_75t_R _31900_ (.A(_14516_),
    .B(_10979_),
    .Y(_10990_));
 OAI21x1_ASAP7_75t_R _31901_ (.A1(_08897_),
    .A2(_10977_),
    .B(_10990_),
    .Y(_03821_));
 BUFx12_ASAP7_75t_R _31902_ (.A(_10976_),
    .Y(_10991_));
 NOR2x1_ASAP7_75t_R _31903_ (.A(_00722_),
    .B(_10991_),
    .Y(_10992_));
 AO21x1_ASAP7_75t_R _31904_ (.A1(_08942_),
    .A2(_10981_),
    .B(_10992_),
    .Y(_03822_));
 NAND2x1_ASAP7_75t_R _31905_ (.A(_00418_),
    .B(_09358_),
    .Y(_10993_));
 OA21x2_ASAP7_75t_R _31906_ (.A1(_08585_),
    .A2(_08764_),
    .B(_10993_),
    .Y(_03823_));
 NOR2x1_ASAP7_75t_R _31907_ (.A(_00752_),
    .B(_10991_),
    .Y(_10994_));
 AO21x1_ASAP7_75t_R _31908_ (.A1(_08988_),
    .A2(_10981_),
    .B(_10994_),
    .Y(_03824_));
 NOR2x1_ASAP7_75t_R _31909_ (.A(_00782_),
    .B(_10991_),
    .Y(_10995_));
 AO21x1_ASAP7_75t_R _31910_ (.A1(_09036_),
    .A2(_10981_),
    .B(_10995_),
    .Y(_03825_));
 NOR2x1_ASAP7_75t_R _31911_ (.A(_00478_),
    .B(_10991_),
    .Y(_10996_));
 AO21x1_ASAP7_75t_R _31912_ (.A1(_09073_),
    .A2(_10981_),
    .B(_10996_),
    .Y(_03826_));
 NOR2x1_ASAP7_75t_R _31913_ (.A(_00853_),
    .B(_10991_),
    .Y(_10997_));
 AO21x1_ASAP7_75t_R _31914_ (.A1(_09103_),
    .A2(_10981_),
    .B(_10997_),
    .Y(_03827_));
 BUFx4f_ASAP7_75t_R _31915_ (.A(_10976_),
    .Y(_10998_));
 NOR2x1_ASAP7_75t_R _31916_ (.A(_00886_),
    .B(_10991_),
    .Y(_10999_));
 AO21x1_ASAP7_75t_R _31917_ (.A1(_09143_),
    .A2(_10998_),
    .B(_10999_),
    .Y(_03828_));
 NOR2x1_ASAP7_75t_R _31918_ (.A(_00919_),
    .B(_10991_),
    .Y(_11000_));
 AO21x1_ASAP7_75t_R _31919_ (.A1(_09180_),
    .A2(_10998_),
    .B(_11000_),
    .Y(_03829_));
 AND2x2_ASAP7_75t_R _31920_ (.A(_16068_),
    .B(_10978_),
    .Y(_11001_));
 AO21x1_ASAP7_75t_R _31921_ (.A1(_09213_),
    .A2(_10998_),
    .B(_11001_),
    .Y(_03830_));
 NOR2x1_ASAP7_75t_R _31922_ (.A(_00985_),
    .B(_10991_),
    .Y(_11002_));
 AO21x1_ASAP7_75t_R _31923_ (.A1(_09244_),
    .A2(_10998_),
    .B(_11002_),
    .Y(_03831_));
 NOR2x1_ASAP7_75t_R _31924_ (.A(_01018_),
    .B(_10991_),
    .Y(_11003_));
 AO21x1_ASAP7_75t_R _31925_ (.A1(_09270_),
    .A2(_10998_),
    .B(_11003_),
    .Y(_03832_));
 NOR2x1_ASAP7_75t_R _31926_ (.A(_01051_),
    .B(_10991_),
    .Y(_11004_));
 AO21x1_ASAP7_75t_R _31927_ (.A1(_09298_),
    .A2(_10998_),
    .B(_11004_),
    .Y(_03833_));
 NAND2x1_ASAP7_75t_R _31928_ (.A(_00371_),
    .B(_09358_),
    .Y(_11005_));
 OA21x2_ASAP7_75t_R _31929_ (.A1(_08764_),
    .A2(_09772_),
    .B(_11005_),
    .Y(_03834_));
 NOR2x1_ASAP7_75t_R _31930_ (.A(_01084_),
    .B(_10976_),
    .Y(_11006_));
 AO21x1_ASAP7_75t_R _31931_ (.A1(_09327_),
    .A2(_10998_),
    .B(_11006_),
    .Y(_03835_));
 NOR2x1_ASAP7_75t_R _31932_ (.A(_01117_),
    .B(_10976_),
    .Y(_11007_));
 AO21x1_ASAP7_75t_R _31933_ (.A1(_09356_),
    .A2(_10998_),
    .B(_11007_),
    .Y(_03836_));
 NOR2x1_ASAP7_75t_R _31934_ (.A(_01150_),
    .B(_10976_),
    .Y(_11008_));
 AO21x1_ASAP7_75t_R _31935_ (.A1(_09389_),
    .A2(_10998_),
    .B(_11008_),
    .Y(_03837_));
 NOR2x1_ASAP7_75t_R _31936_ (.A(_01183_),
    .B(_10976_),
    .Y(_11009_));
 AO21x1_ASAP7_75t_R _31937_ (.A1(_09415_),
    .A2(_10998_),
    .B(_11009_),
    .Y(_03838_));
 NAND2x1_ASAP7_75t_R _31938_ (.A(_01216_),
    .B(_10979_),
    .Y(_11010_));
 OA21x2_ASAP7_75t_R _31939_ (.A1(_09442_),
    .A2(_10979_),
    .B(_11010_),
    .Y(_03839_));
 NOR2x1_ASAP7_75t_R _31940_ (.A(_01249_),
    .B(_10976_),
    .Y(_11011_));
 AO21x1_ASAP7_75t_R _31941_ (.A1(_09471_),
    .A2(_10982_),
    .B(_11011_),
    .Y(_03840_));
 NOR2x1_ASAP7_75t_R _31942_ (.A(_01282_),
    .B(_10976_),
    .Y(_11012_));
 AO21x1_ASAP7_75t_R _31943_ (.A1(_09494_),
    .A2(_10982_),
    .B(_11012_),
    .Y(_03841_));
 AND2x2_ASAP7_75t_R _31944_ (.A(_04319_),
    .B(_10978_),
    .Y(_11013_));
 AO21x1_ASAP7_75t_R _31945_ (.A1(_09512_),
    .A2(_10982_),
    .B(_11013_),
    .Y(_03842_));
 AND2x2_ASAP7_75t_R _31946_ (.A(_04449_),
    .B(_10978_),
    .Y(_11014_));
 AO21x1_ASAP7_75t_R _31947_ (.A1(_09544_),
    .A2(_10982_),
    .B(_11014_),
    .Y(_03843_));
 NAND2x1_ASAP7_75t_R _31948_ (.A(_01381_),
    .B(_10979_),
    .Y(_11015_));
 OA21x2_ASAP7_75t_R _31949_ (.A1(_09580_),
    .A2(_10979_),
    .B(_11015_),
    .Y(_03844_));
 NAND2x1_ASAP7_75t_R _31950_ (.A(_00482_),
    .B(_09358_),
    .Y(_11016_));
 OA21x2_ASAP7_75t_R _31951_ (.A1(_08764_),
    .A2(_09695_),
    .B(_11016_),
    .Y(_03845_));
 AND2x2_ASAP7_75t_R _31952_ (.A(_04673_),
    .B(_10978_),
    .Y(_11017_));
 AO21x1_ASAP7_75t_R _31953_ (.A1(_09622_),
    .A2(_10982_),
    .B(_11017_),
    .Y(_03846_));
 AND2x2_ASAP7_75t_R _31954_ (.A(_04791_),
    .B(_10978_),
    .Y(_11018_));
 AO21x1_ASAP7_75t_R _31955_ (.A1(_09648_),
    .A2(_10982_),
    .B(_11018_),
    .Y(_03847_));
 NAND2x1_ASAP7_75t_R _31956_ (.A(_00513_),
    .B(_08680_),
    .Y(_11019_));
 OA21x2_ASAP7_75t_R _31957_ (.A1(_08764_),
    .A2(_09782_),
    .B(_11019_),
    .Y(_03848_));
 NAND2x1_ASAP7_75t_R _31958_ (.A(_01783_),
    .B(_09106_),
    .Y(_11020_));
 OA21x2_ASAP7_75t_R _31959_ (.A1(_08591_),
    .A2(_08943_),
    .B(_11020_),
    .Y(_03849_));
 AND5x1_ASAP7_75t_R _31960_ (.A(_05066_),
    .B(_05069_),
    .C(_05071_),
    .D(_05325_),
    .E(_05408_),
    .Y(_11021_));
 INVx1_ASAP7_75t_R _31961_ (.A(_11021_),
    .Y(_11022_));
 AO21x1_ASAP7_75t_R _31962_ (.A1(_13407_),
    .A2(_05379_),
    .B(net105),
    .Y(_11023_));
 AND2x4_ASAP7_75t_R _31963_ (.A(_04945_),
    .B(_11023_),
    .Y(_11024_));
 OAI21x1_ASAP7_75t_R _31964_ (.A1(_07221_),
    .A2(_07224_),
    .B(_11024_),
    .Y(_11025_));
 AND3x1_ASAP7_75t_R _31965_ (.A(_05077_),
    .B(_11022_),
    .C(_11025_),
    .Y(_11026_));
 NOR2x1_ASAP7_75t_R _31966_ (.A(_04935_),
    .B(_05421_),
    .Y(_11027_));
 INVx1_ASAP7_75t_R _31967_ (.A(_01455_),
    .Y(_11028_));
 OR4x2_ASAP7_75t_R _31968_ (.A(net105),
    .B(_11028_),
    .C(_05379_),
    .D(_05437_),
    .Y(_11029_));
 NAND2x1_ASAP7_75t_R _31969_ (.A(_04934_),
    .B(_11029_),
    .Y(_11030_));
 NOR2x1_ASAP7_75t_R _31970_ (.A(_05340_),
    .B(_11024_),
    .Y(_11031_));
 AND2x2_ASAP7_75t_R _31971_ (.A(_04935_),
    .B(_11031_),
    .Y(_11032_));
 AO221x1_ASAP7_75t_R _31972_ (.A1(_04934_),
    .A2(_05421_),
    .B1(_11027_),
    .B2(_11030_),
    .C(_11032_),
    .Y(_11033_));
 AO21x1_ASAP7_75t_R _31973_ (.A1(_04932_),
    .A2(_11033_),
    .B(_05381_),
    .Y(_11034_));
 BUFx10_ASAP7_75t_R _31974_ (.A(_04938_),
    .Y(_11035_));
 BUFx3_ASAP7_75t_R _31975_ (.A(_11035_),
    .Y(_11036_));
 INVx1_ASAP7_75t_R _31976_ (.A(_06834_),
    .Y(_11037_));
 OA21x2_ASAP7_75t_R _31977_ (.A1(_14039_),
    .A2(_05071_),
    .B(_05069_),
    .Y(_11038_));
 AND4x2_ASAP7_75t_R _31978_ (.A(_13479_),
    .B(net12),
    .C(_13484_),
    .D(_02308_),
    .Y(_11039_));
 NAND2x1_ASAP7_75t_R _31979_ (.A(_02310_),
    .B(_14038_),
    .Y(_11040_));
 NOR3x1_ASAP7_75t_R _31980_ (.A(_02308_),
    .B(_14062_),
    .C(_11040_),
    .Y(_11041_));
 AO21x1_ASAP7_75t_R _31981_ (.A1(_05080_),
    .A2(_11039_),
    .B(_11041_),
    .Y(_11042_));
 AND4x1_ASAP7_75t_R _31982_ (.A(_14037_),
    .B(_14070_),
    .C(_04940_),
    .D(_11042_),
    .Y(_11043_));
 OR4x1_ASAP7_75t_R _31983_ (.A(_11037_),
    .B(_05067_),
    .C(_11038_),
    .D(_11043_),
    .Y(_11044_));
 AOI21x1_ASAP7_75t_R _31984_ (.A1(_05089_),
    .A2(_05090_),
    .B(_11044_),
    .Y(_11045_));
 NAND2x1_ASAP7_75t_R _31985_ (.A(_06859_),
    .B(_11024_),
    .Y(_11046_));
 AND3x1_ASAP7_75t_R _31986_ (.A(_11036_),
    .B(_11045_),
    .C(_11046_),
    .Y(_11047_));
 AND2x2_ASAP7_75t_R _31987_ (.A(_04932_),
    .B(_04936_),
    .Y(_11048_));
 OA21x2_ASAP7_75t_R _31988_ (.A1(_04934_),
    .A2(_05421_),
    .B(_11048_),
    .Y(_11049_));
 INVx1_ASAP7_75t_R _31989_ (.A(_11049_),
    .Y(_11050_));
 AND2x2_ASAP7_75t_R _31990_ (.A(_06859_),
    .B(_11050_),
    .Y(_11051_));
 AND2x2_ASAP7_75t_R _31991_ (.A(_05376_),
    .B(_05437_),
    .Y(_11052_));
 AND3x1_ASAP7_75t_R _31992_ (.A(_04935_),
    .B(_05374_),
    .C(_11031_),
    .Y(_11053_));
 INVx1_ASAP7_75t_R _31993_ (.A(_11053_),
    .Y(_11054_));
 OA33x2_ASAP7_75t_R _31994_ (.A1(_11026_),
    .A2(_11034_),
    .A3(_11047_),
    .B1(_11051_),
    .B2(_11052_),
    .B3(_11054_),
    .Y(_03850_));
 AND2x2_ASAP7_75t_R _31995_ (.A(_05077_),
    .B(_11025_),
    .Y(_11055_));
 AO21x1_ASAP7_75t_R _31996_ (.A1(_06859_),
    .A2(_11052_),
    .B(_04936_),
    .Y(_11056_));
 INVx1_ASAP7_75t_R _31997_ (.A(_11045_),
    .Y(_11057_));
 AO21x1_ASAP7_75t_R _31998_ (.A1(_11046_),
    .A2(_11056_),
    .B(_11057_),
    .Y(_11058_));
 INVx1_ASAP7_75t_R _31999_ (.A(_11029_),
    .Y(_11059_));
 OA211x2_ASAP7_75t_R _32000_ (.A1(_05421_),
    .A2(_11059_),
    .B(_11048_),
    .C(_04934_),
    .Y(_11060_));
 AO21x1_ASAP7_75t_R _32001_ (.A1(_11052_),
    .A2(_11053_),
    .B(_11060_),
    .Y(_11061_));
 AO221x1_ASAP7_75t_R _32002_ (.A1(_11021_),
    .A2(_11055_),
    .B1(_11058_),
    .B2(_11036_),
    .C(_11061_),
    .Y(_03851_));
 OA21x2_ASAP7_75t_R _32003_ (.A1(_11057_),
    .A2(_11046_),
    .B(_11036_),
    .Y(_11062_));
 AO21x1_ASAP7_75t_R _32004_ (.A1(_05075_),
    .A2(_11032_),
    .B(_11027_),
    .Y(_11063_));
 AND2x2_ASAP7_75t_R _32005_ (.A(_04933_),
    .B(_04935_),
    .Y(_11064_));
 AO21x1_ASAP7_75t_R _32006_ (.A1(_04932_),
    .A2(_05340_),
    .B(_11064_),
    .Y(_11065_));
 AO222x2_ASAP7_75t_R _32007_ (.A1(_04932_),
    .A2(_11063_),
    .B1(_11065_),
    .B2(_04934_),
    .C1(_05335_),
    .C2(_11026_),
    .Y(_11066_));
 OR3x1_ASAP7_75t_R _32008_ (.A(_05075_),
    .B(_05421_),
    .C(_11029_),
    .Y(_11067_));
 AO21x1_ASAP7_75t_R _32009_ (.A1(_04932_),
    .A2(_11067_),
    .B(_05380_),
    .Y(_11068_));
 OA21x2_ASAP7_75t_R _32010_ (.A1(_11062_),
    .A2(_11066_),
    .B(_11068_),
    .Y(_03852_));
 AOI21x1_ASAP7_75t_R _32011_ (.A1(_05335_),
    .A2(_11025_),
    .B(_05340_),
    .Y(_11069_));
 AO21x1_ASAP7_75t_R _32012_ (.A1(_06831_),
    .A2(_11045_),
    .B(_05421_),
    .Y(_11070_));
 OR3x2_ASAP7_75t_R _32013_ (.A(_06787_),
    .B(_06827_),
    .C(_06829_),
    .Y(_11071_));
 BUFx6f_ASAP7_75t_R _32014_ (.A(_11071_),
    .Y(_11072_));
 INVx1_ASAP7_75t_R _32015_ (.A(_11052_),
    .Y(_11073_));
 OA211x2_ASAP7_75t_R _32016_ (.A1(_11072_),
    .A2(_11073_),
    .B(_04933_),
    .C(_05340_),
    .Y(_11074_));
 AO221x1_ASAP7_75t_R _32017_ (.A1(_11024_),
    .A2(_11070_),
    .B1(_11074_),
    .B2(_11045_),
    .C(_04936_),
    .Y(_11075_));
 OA211x2_ASAP7_75t_R _32018_ (.A1(_04935_),
    .A2(_11069_),
    .B(_11075_),
    .C(_05374_),
    .Y(_03853_));
 OR3x1_ASAP7_75t_R _32019_ (.A(net105),
    .B(_05379_),
    .C(_05340_),
    .Y(_11076_));
 AND2x2_ASAP7_75t_R _32020_ (.A(_05381_),
    .B(_11076_),
    .Y(_11077_));
 OA21x2_ASAP7_75t_R _32021_ (.A1(_11028_),
    .A2(_11077_),
    .B(_05418_),
    .Y(_03854_));
 AO22x1_ASAP7_75t_R _32022_ (.A1(net194),
    .A2(_05377_),
    .B1(_07230_),
    .B2(_07761_),
    .Y(_03855_));
 OA21x2_ASAP7_75t_R _32023_ (.A1(_08347_),
    .A2(_08350_),
    .B(_13570_),
    .Y(_11078_));
 OR3x1_ASAP7_75t_R _32024_ (.A(_14026_),
    .B(_05321_),
    .C(_11078_),
    .Y(_11079_));
 AO21x1_ASAP7_75t_R _32025_ (.A1(_04928_),
    .A2(_11079_),
    .B(_06785_),
    .Y(_11080_));
 INVx1_ASAP7_75t_R _32026_ (.A(_06783_),
    .Y(_11081_));
 AOI21x1_ASAP7_75t_R _32027_ (.A1(_04940_),
    .A2(_11081_),
    .B(_01776_),
    .Y(_11082_));
 AO21x1_ASAP7_75t_R _32028_ (.A1(_05753_),
    .A2(_11080_),
    .B(_11082_),
    .Y(_03856_));
 NAND2x2_ASAP7_75t_R _32029_ (.A(_05105_),
    .B(_05132_),
    .Y(_11083_));
 BUFx6f_ASAP7_75t_R _32030_ (.A(_11083_),
    .Y(_11084_));
 AND2x4_ASAP7_75t_R _32031_ (.A(_04875_),
    .B(_04876_),
    .Y(_11085_));
 NAND2x2_ASAP7_75t_R _32032_ (.A(_11085_),
    .B(_05295_),
    .Y(_11086_));
 BUFx4f_ASAP7_75t_R _32033_ (.A(_11086_),
    .Y(_11087_));
 BUFx4f_ASAP7_75t_R _32034_ (.A(_11087_),
    .Y(_11088_));
 BUFx4f_ASAP7_75t_R _32035_ (.A(_05296_),
    .Y(_11089_));
 OR2x2_ASAP7_75t_R _32036_ (.A(_05672_),
    .B(_11089_),
    .Y(_11090_));
 OA211x2_ASAP7_75t_R _32037_ (.A1(net52),
    .A2(_11088_),
    .B(_11090_),
    .C(_05108_),
    .Y(_11091_));
 AOI21x1_ASAP7_75t_R _32038_ (.A1(_01775_),
    .A2(_11084_),
    .B(_11091_),
    .Y(_03857_));
 BUFx6f_ASAP7_75t_R _32039_ (.A(_11083_),
    .Y(_11092_));
 BUFx4f_ASAP7_75t_R _32040_ (.A(_11086_),
    .Y(_11093_));
 OR2x2_ASAP7_75t_R _32041_ (.A(_14666_),
    .B(_05297_),
    .Y(_11094_));
 BUFx3_ASAP7_75t_R _32042_ (.A(_05107_),
    .Y(_11095_));
 OA211x2_ASAP7_75t_R _32043_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_11093_),
    .B(_11094_),
    .C(_11095_),
    .Y(_11096_));
 AO21x1_ASAP7_75t_R _32044_ (.A1(_05584_),
    .A2(_11092_),
    .B(_11096_),
    .Y(_03858_));
 BUFx4f_ASAP7_75t_R _32045_ (.A(_05296_),
    .Y(_11097_));
 NAND2x1_ASAP7_75t_R _32046_ (.A(\alu_adder_result_ex[11] ),
    .B(_11097_),
    .Y(_11098_));
 OA211x2_ASAP7_75t_R _32047_ (.A1(_05589_),
    .A2(_11097_),
    .B(_11098_),
    .C(_05108_),
    .Y(_11099_));
 AOI21x1_ASAP7_75t_R _32048_ (.A1(_01773_),
    .A2(_11084_),
    .B(_11099_),
    .Y(_03859_));
 OR2x2_ASAP7_75t_R _32049_ (.A(_05261_),
    .B(_05297_),
    .Y(_11100_));
 BUFx3_ASAP7_75t_R _32050_ (.A(_05107_),
    .Y(_11101_));
 OA211x2_ASAP7_75t_R _32051_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_11093_),
    .B(_11100_),
    .C(_11101_),
    .Y(_11102_));
 AO21x1_ASAP7_75t_R _32052_ (.A1(_05702_),
    .A2(_11092_),
    .B(_11102_),
    .Y(_03860_));
 AO21x1_ASAP7_75t_R _32053_ (.A1(_15632_),
    .A2(_15670_),
    .B(_11097_),
    .Y(_11103_));
 OA211x2_ASAP7_75t_R _32054_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_11093_),
    .B(_11103_),
    .C(_11101_),
    .Y(_11104_));
 AO21x1_ASAP7_75t_R _32055_ (.A1(_05599_),
    .A2(_11092_),
    .B(_11104_),
    .Y(_03861_));
 NAND2x1_ASAP7_75t_R _32056_ (.A(_15816_),
    .B(_11087_),
    .Y(_11105_));
 OA211x2_ASAP7_75t_R _32057_ (.A1(_16028_),
    .A2(_11088_),
    .B(_11105_),
    .C(_05108_),
    .Y(_11106_));
 AOI21x1_ASAP7_75t_R _32058_ (.A1(_01770_),
    .A2(_11084_),
    .B(_11106_),
    .Y(_03862_));
 BUFx4f_ASAP7_75t_R _32059_ (.A(_11083_),
    .Y(_11107_));
 NAND2x1_ASAP7_75t_R _32060_ (.A(_04875_),
    .B(_04876_),
    .Y(_11108_));
 INVx1_ASAP7_75t_R _32061_ (.A(_05295_),
    .Y(_11109_));
 OR3x1_ASAP7_75t_R _32062_ (.A(\alu_adder_result_ex[15] ),
    .B(_11108_),
    .C(_11109_),
    .Y(_11110_));
 OA211x2_ASAP7_75t_R _32063_ (.A1(_15950_),
    .A2(_11097_),
    .B(_11110_),
    .C(_11101_),
    .Y(_11111_));
 AO21x1_ASAP7_75t_R _32064_ (.A1(_05610_),
    .A2(_11107_),
    .B(_11111_),
    .Y(_03863_));
 AO21x1_ASAP7_75t_R _32065_ (.A1(_16060_),
    .A2(_16093_),
    .B(_11089_),
    .Y(_11112_));
 OA211x2_ASAP7_75t_R _32066_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_11093_),
    .B(_11112_),
    .C(_11101_),
    .Y(_11113_));
 AO21x1_ASAP7_75t_R _32067_ (.A1(_05615_),
    .A2(_11107_),
    .B(_11113_),
    .Y(_03864_));
 INVx1_ASAP7_75t_R _32068_ (.A(_16209_),
    .Y(_11114_));
 NAND2x1_ASAP7_75t_R _32069_ (.A(\alu_adder_result_ex[17] ),
    .B(_11097_),
    .Y(_11115_));
 OA211x2_ASAP7_75t_R _32070_ (.A1(_11114_),
    .A2(_11097_),
    .B(_11115_),
    .C(_05108_),
    .Y(_11116_));
 AOI21x1_ASAP7_75t_R _32071_ (.A1(_01767_),
    .A2(_11084_),
    .B(_11116_),
    .Y(_03865_));
 AO21x1_ASAP7_75t_R _32072_ (.A1(_16320_),
    .A2(_16353_),
    .B(_11089_),
    .Y(_11117_));
 OA211x2_ASAP7_75t_R _32073_ (.A1(\alu_adder_result_ex[18] ),
    .A2(_11093_),
    .B(_11117_),
    .C(_11101_),
    .Y(_11118_));
 AO21x1_ASAP7_75t_R _32074_ (.A1(_05717_),
    .A2(_11107_),
    .B(_11118_),
    .Y(_03866_));
 AO21x1_ASAP7_75t_R _32075_ (.A1(_16434_),
    .A2(_16465_),
    .B(_11089_),
    .Y(_11119_));
 OA211x2_ASAP7_75t_R _32076_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_11093_),
    .B(_11119_),
    .C(_11101_),
    .Y(_11120_));
 AO21x1_ASAP7_75t_R _32077_ (.A1(_05624_),
    .A2(_11107_),
    .B(_11120_),
    .Y(_03867_));
 OR2x2_ASAP7_75t_R _32078_ (.A(_05528_),
    .B(_11089_),
    .Y(_11121_));
 OA211x2_ASAP7_75t_R _32079_ (.A1(_18764_),
    .A2(_11088_),
    .B(_11121_),
    .C(_05108_),
    .Y(_11122_));
 AOI21x1_ASAP7_75t_R _32080_ (.A1(_01764_),
    .A2(_11084_),
    .B(_11122_),
    .Y(_03868_));
 OR2x2_ASAP7_75t_R _32081_ (.A(_16592_),
    .B(_11089_),
    .Y(_11123_));
 OA211x2_ASAP7_75t_R _32082_ (.A1(_16777_),
    .A2(_11088_),
    .B(_11123_),
    .C(_05108_),
    .Y(_11124_));
 AOI21x1_ASAP7_75t_R _32083_ (.A1(_01763_),
    .A2(_11084_),
    .B(_11124_),
    .Y(_03869_));
 NAND2x1_ASAP7_75t_R _32084_ (.A(\alu_adder_result_ex[21] ),
    .B(_11097_),
    .Y(_11125_));
 OA211x2_ASAP7_75t_R _32085_ (.A1(_16706_),
    .A2(_11097_),
    .B(_11125_),
    .C(_05108_),
    .Y(_11126_));
 AOI21x1_ASAP7_75t_R _32086_ (.A1(_01762_),
    .A2(_11084_),
    .B(_11126_),
    .Y(_03870_));
 OR2x2_ASAP7_75t_R _32087_ (.A(_16836_),
    .B(_11089_),
    .Y(_11127_));
 OA211x2_ASAP7_75t_R _32088_ (.A1(_17017_),
    .A2(_11088_),
    .B(_11127_),
    .C(_05108_),
    .Y(_11128_));
 AOI21x1_ASAP7_75t_R _32089_ (.A1(_01761_),
    .A2(_11084_),
    .B(_11128_),
    .Y(_03871_));
 AO21x1_ASAP7_75t_R _32090_ (.A1(_16914_),
    .A2(_16945_),
    .B(_11089_),
    .Y(_11129_));
 OA211x2_ASAP7_75t_R _32091_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_11093_),
    .B(_11129_),
    .C(_11101_),
    .Y(_11130_));
 AO21x1_ASAP7_75t_R _32092_ (.A1(_05726_),
    .A2(_11107_),
    .B(_11130_),
    .Y(_03872_));
 OR2x2_ASAP7_75t_R _32093_ (.A(_17076_),
    .B(_11089_),
    .Y(_11131_));
 OA211x2_ASAP7_75t_R _32094_ (.A1(_17257_),
    .A2(_11088_),
    .B(_11131_),
    .C(_05108_),
    .Y(_11132_));
 AOI21x1_ASAP7_75t_R _32095_ (.A1(_01759_),
    .A2(_11084_),
    .B(_11132_),
    .Y(_03873_));
 INVx1_ASAP7_75t_R _32096_ (.A(_01758_),
    .Y(_11133_));
 NAND2x1_ASAP7_75t_R _32097_ (.A(_17185_),
    .B(_11087_),
    .Y(_11134_));
 OA211x2_ASAP7_75t_R _32098_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_11087_),
    .B(_11134_),
    .C(_11101_),
    .Y(_11135_));
 AO21x1_ASAP7_75t_R _32099_ (.A1(_11133_),
    .A2(_11107_),
    .B(_11135_),
    .Y(_03874_));
 OR2x2_ASAP7_75t_R _32100_ (.A(_17316_),
    .B(_11089_),
    .Y(_11136_));
 OA211x2_ASAP7_75t_R _32101_ (.A1(_04414_),
    .A2(_11088_),
    .B(_11136_),
    .C(_11095_),
    .Y(_11137_));
 AOI21x1_ASAP7_75t_R _32102_ (.A1(_01757_),
    .A2(_11084_),
    .B(_11137_),
    .Y(_03875_));
 NAND2x1_ASAP7_75t_R _32103_ (.A(\alu_adder_result_ex[27] ),
    .B(_11097_),
    .Y(_11138_));
 OA211x2_ASAP7_75t_R _32104_ (.A1(_04343_),
    .A2(_11097_),
    .B(_11138_),
    .C(_11095_),
    .Y(_11139_));
 AOI21x1_ASAP7_75t_R _32105_ (.A1(_01756_),
    .A2(_11092_),
    .B(_11139_),
    .Y(_03876_));
 OR2x2_ASAP7_75t_R _32106_ (.A(_04473_),
    .B(_05297_),
    .Y(_11140_));
 OA211x2_ASAP7_75t_R _32107_ (.A1(_05135_),
    .A2(_11088_),
    .B(_11140_),
    .C(_11095_),
    .Y(_11141_));
 AOI21x1_ASAP7_75t_R _32108_ (.A1(_01755_),
    .A2(_11092_),
    .B(_11141_),
    .Y(_03877_));
 INVx1_ASAP7_75t_R _32109_ (.A(\alu_adder_result_ex[29] ),
    .Y(_11142_));
 OR2x2_ASAP7_75t_R _32110_ (.A(_04583_),
    .B(_05297_),
    .Y(_11143_));
 OA211x2_ASAP7_75t_R _32111_ (.A1(_11142_),
    .A2(_11088_),
    .B(_11143_),
    .C(_11095_),
    .Y(_11144_));
 AOI21x1_ASAP7_75t_R _32112_ (.A1(_01754_),
    .A2(_11092_),
    .B(_11144_),
    .Y(_03878_));
 OR2x2_ASAP7_75t_R _32113_ (.A(_14148_),
    .B(_05297_),
    .Y(_11145_));
 OA211x2_ASAP7_75t_R _32114_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_11087_),
    .B(_11145_),
    .C(_11101_),
    .Y(_11146_));
 AO21x1_ASAP7_75t_R _32115_ (.A1(_05678_),
    .A2(_11107_),
    .B(_11146_),
    .Y(_03879_));
 OR2x2_ASAP7_75t_R _32116_ (.A(_04697_),
    .B(_05297_),
    .Y(_11147_));
 OA211x2_ASAP7_75t_R _32117_ (.A1(_04917_),
    .A2(_11088_),
    .B(_11147_),
    .C(_11095_),
    .Y(_11148_));
 AOI21x1_ASAP7_75t_R _32118_ (.A1(_01752_),
    .A2(_11092_),
    .B(_11148_),
    .Y(_03880_));
 INVx1_ASAP7_75t_R _32119_ (.A(_01751_),
    .Y(_11149_));
 OA211x2_ASAP7_75t_R _32120_ (.A1(\alu_adder_result_ex[31] ),
    .A2(_11109_),
    .B(_11095_),
    .C(_11085_),
    .Y(_11150_));
 AO21x1_ASAP7_75t_R _32121_ (.A1(_11149_),
    .A2(_11107_),
    .B(_11150_),
    .Y(_03881_));
 AND3x2_ASAP7_75t_R _32122_ (.A(_05523_),
    .B(_02212_),
    .C(_05525_),
    .Y(_11151_));
 BUFx4f_ASAP7_75t_R _32123_ (.A(_11151_),
    .Y(_11152_));
 AND3x4_ASAP7_75t_R _32124_ (.A(_13566_),
    .B(_05304_),
    .C(_08135_),
    .Y(_11153_));
 BUFx6f_ASAP7_75t_R _32125_ (.A(_11153_),
    .Y(_11154_));
 BUFx4f_ASAP7_75t_R _32126_ (.A(_11154_),
    .Y(_11155_));
 NAND2x1_ASAP7_75t_R _32127_ (.A(_00447_),
    .B(_08298_),
    .Y(_11156_));
 OA21x2_ASAP7_75t_R _32128_ (.A1(\alu_adder_result_ex[0] ),
    .A2(_08272_),
    .B(_11156_),
    .Y(_11157_));
 AND2x2_ASAP7_75t_R _32129_ (.A(_05100_),
    .B(_05101_),
    .Y(_11158_));
 NAND2x1_ASAP7_75t_R _32130_ (.A(_00071_),
    .B(_11154_),
    .Y(_11159_));
 AO21x1_ASAP7_75t_R _32131_ (.A1(_11158_),
    .A2(_08285_),
    .B(_11159_),
    .Y(_11160_));
 INVx2_ASAP7_75t_R _32132_ (.A(_02217_),
    .Y(_11161_));
 OA211x2_ASAP7_75t_R _32133_ (.A1(_11155_),
    .A2(_11157_),
    .B(_11160_),
    .C(_11161_),
    .Y(_11162_));
 AO22x1_ASAP7_75t_R _32134_ (.A1(_05138_),
    .A2(\alu_adder_result_ex[0] ),
    .B1(_08240_),
    .B2(_05105_),
    .Y(_11163_));
 XOR2x1_ASAP7_75t_R _32135_ (.A(_05101_),
    .Y(_11164_),
    .B(_02317_));
 BUFx3_ASAP7_75t_R _32136_ (.A(_08143_),
    .Y(_11165_));
 NAND2x1_ASAP7_75t_R _32137_ (.A(_08143_),
    .B(_00120_),
    .Y(_11166_));
 OA211x2_ASAP7_75t_R _32138_ (.A1(_11165_),
    .A2(_08178_),
    .B(_11166_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11167_));
 BUFx4f_ASAP7_75t_R _32139_ (.A(_02316_),
    .Y(_11168_));
 NAND2x1_ASAP7_75t_R _32140_ (.A(_08143_),
    .B(_00119_),
    .Y(_11169_));
 OA211x2_ASAP7_75t_R _32141_ (.A1(_11168_),
    .A2(_08181_),
    .B(_11169_),
    .C(_05162_),
    .Y(_11170_));
 OR3x1_ASAP7_75t_R _32142_ (.A(_08150_),
    .B(_11167_),
    .C(_11170_),
    .Y(_11171_));
 XNOR2x2_ASAP7_75t_R _32143_ (.A(_05094_),
    .B(_08149_),
    .Y(_11172_));
 NAND2x1_ASAP7_75t_R _32144_ (.A(_08143_),
    .B(_00112_),
    .Y(_11173_));
 OA211x2_ASAP7_75t_R _32145_ (.A1(_11165_),
    .A2(_08244_),
    .B(_11173_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11174_));
 NAND2x1_ASAP7_75t_R _32146_ (.A(_08143_),
    .B(_00111_),
    .Y(_11175_));
 OA211x2_ASAP7_75t_R _32147_ (.A1(_11168_),
    .A2(_08247_),
    .B(_11175_),
    .C(_05162_),
    .Y(_11176_));
 OR3x1_ASAP7_75t_R _32148_ (.A(_11172_),
    .B(_11174_),
    .C(_11176_),
    .Y(_11177_));
 AND3x1_ASAP7_75t_R _32149_ (.A(_11164_),
    .B(_11171_),
    .C(_11177_),
    .Y(_11178_));
 NAND2x1_ASAP7_75t_R _32150_ (.A(_08144_),
    .B(_00114_),
    .Y(_11179_));
 OA211x2_ASAP7_75t_R _32151_ (.A1(_08144_),
    .A2(_08170_),
    .B(_11179_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11180_));
 NAND2x1_ASAP7_75t_R _32152_ (.A(_11168_),
    .B(_00115_),
    .Y(_11181_));
 OA211x2_ASAP7_75t_R _32153_ (.A1(_11165_),
    .A2(_08256_),
    .B(_11181_),
    .C(_05162_),
    .Y(_11182_));
 OR3x1_ASAP7_75t_R _32154_ (.A(_08150_),
    .B(_11180_),
    .C(_11182_),
    .Y(_11183_));
 NAND2x1_ASAP7_75t_R _32155_ (.A(_00106_),
    .B(_08144_),
    .Y(_11184_));
 OA211x2_ASAP7_75t_R _32156_ (.A1(_08235_),
    .A2(_08144_),
    .B(_11184_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11185_));
 NAND2x1_ASAP7_75t_R _32157_ (.A(_00107_),
    .B(_11168_),
    .Y(_11186_));
 OA211x2_ASAP7_75t_R _32158_ (.A1(_08202_),
    .A2(_11165_),
    .B(_11186_),
    .C(_05162_),
    .Y(_11187_));
 OR3x1_ASAP7_75t_R _32159_ (.A(_11172_),
    .B(_11185_),
    .C(_11187_),
    .Y(_11188_));
 AND3x1_ASAP7_75t_R _32160_ (.A(_08146_),
    .B(_11183_),
    .C(_11188_),
    .Y(_11189_));
 NOR2x1_ASAP7_75t_R _32161_ (.A(_11178_),
    .B(_11189_),
    .Y(_11190_));
 XNOR2x1_ASAP7_75t_R _32162_ (.B(_08157_),
    .Y(_11191_),
    .A(_08155_));
 NAND2x1_ASAP7_75t_R _32163_ (.A(_11190_),
    .B(_11191_),
    .Y(_11192_));
 NOR2x1_ASAP7_75t_R _32164_ (.A(_11165_),
    .B(_00125_),
    .Y(_11193_));
 AO21x1_ASAP7_75t_R _32165_ (.A1(_11165_),
    .A2(_08216_),
    .B(_11193_),
    .Y(_11194_));
 NAND2x1_ASAP7_75t_R _32166_ (.A(_11168_),
    .B(_00128_),
    .Y(_11195_));
 OA211x2_ASAP7_75t_R _32167_ (.A1(_11165_),
    .A2(_08205_),
    .B(_11195_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11196_));
 AO21x1_ASAP7_75t_R _32168_ (.A1(_05162_),
    .A2(_11194_),
    .B(_11196_),
    .Y(_11197_));
 NAND2x1_ASAP7_75t_R _32169_ (.A(_08143_),
    .B(_00136_),
    .Y(_11198_));
 OA211x2_ASAP7_75t_R _32170_ (.A1(_11168_),
    .A2(_08229_),
    .B(_11198_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11199_));
 NAND2x1_ASAP7_75t_R _32171_ (.A(_08143_),
    .B(_00135_),
    .Y(_11200_));
 OA211x2_ASAP7_75t_R _32172_ (.A1(_11168_),
    .A2(_08232_),
    .B(_11200_),
    .C(_05162_),
    .Y(_11201_));
 OR3x1_ASAP7_75t_R _32173_ (.A(_08150_),
    .B(_11199_),
    .C(_11201_),
    .Y(_11202_));
 OA211x2_ASAP7_75t_R _32174_ (.A1(_11172_),
    .A2(_11197_),
    .B(_11202_),
    .C(_11164_),
    .Y(_11203_));
 NOR2x1_ASAP7_75t_R _32175_ (.A(_11165_),
    .B(_00121_),
    .Y(_11204_));
 AO21x1_ASAP7_75t_R _32176_ (.A1(_11165_),
    .A2(_08199_),
    .B(_11204_),
    .Y(_11205_));
 NAND2x1_ASAP7_75t_R _32177_ (.A(_11168_),
    .B(_00124_),
    .Y(_11206_));
 OA211x2_ASAP7_75t_R _32178_ (.A1(_11165_),
    .A2(_08191_),
    .B(_11206_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11207_));
 AO21x1_ASAP7_75t_R _32179_ (.A1(_05162_),
    .A2(_11205_),
    .B(_11207_),
    .Y(_11208_));
 INVx1_ASAP7_75t_R _32180_ (.A(_00130_),
    .Y(_11209_));
 NAND2x1_ASAP7_75t_R _32181_ (.A(_08143_),
    .B(_00132_),
    .Y(_11210_));
 OA211x2_ASAP7_75t_R _32182_ (.A1(_11168_),
    .A2(_11209_),
    .B(_11210_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_11211_));
 NAND2x1_ASAP7_75t_R _32183_ (.A(_08143_),
    .B(_00131_),
    .Y(_11212_));
 OA211x2_ASAP7_75t_R _32184_ (.A1(_11168_),
    .A2(_08221_),
    .B(_11212_),
    .C(_05162_),
    .Y(_11213_));
 OR3x1_ASAP7_75t_R _32185_ (.A(_08150_),
    .B(_11211_),
    .C(_11213_),
    .Y(_11214_));
 OA211x2_ASAP7_75t_R _32186_ (.A1(_11172_),
    .A2(_11208_),
    .B(_11214_),
    .C(_08146_),
    .Y(_11215_));
 OR3x1_ASAP7_75t_R _32187_ (.A(_11191_),
    .B(_11203_),
    .C(_11215_),
    .Y(_11216_));
 AND3x1_ASAP7_75t_R _32188_ (.A(_05091_),
    .B(_11192_),
    .C(_11216_),
    .Y(_11217_));
 OR4x1_ASAP7_75t_R _32189_ (.A(_11152_),
    .B(_11162_),
    .C(_11163_),
    .D(_11217_),
    .Y(_11218_));
 OR3x4_ASAP7_75t_R _32190_ (.A(_04871_),
    .B(_05105_),
    .C(_04870_),
    .Y(_11219_));
 AND3x1_ASAP7_75t_R _32191_ (.A(_05296_),
    .B(_08161_),
    .C(_11153_),
    .Y(_11220_));
 AO21x1_ASAP7_75t_R _32192_ (.A1(_11086_),
    .A2(_08166_),
    .B(_11220_),
    .Y(_11221_));
 AO221x1_ASAP7_75t_R _32193_ (.A1(_08166_),
    .A2(_08136_),
    .B1(_11221_),
    .B2(_01817_),
    .C(_00408_),
    .Y(_11222_));
 OA21x2_ASAP7_75t_R _32194_ (.A1(_05133_),
    .A2(_11219_),
    .B(_11222_),
    .Y(_11223_));
 OA211x2_ASAP7_75t_R _32195_ (.A1(net2004),
    .A2(_11223_),
    .B(_05097_),
    .C(_05514_),
    .Y(_11224_));
 BUFx6f_ASAP7_75t_R _32196_ (.A(_11224_),
    .Y(_11225_));
 AND2x2_ASAP7_75t_R _32197_ (.A(_05096_),
    .B(_11225_),
    .Y(_11226_));
 BUFx4f_ASAP7_75t_R _32198_ (.A(_11226_),
    .Y(_11227_));
 OR2x2_ASAP7_75t_R _32199_ (.A(_11219_),
    .B(_11153_),
    .Y(_11228_));
 BUFx4f_ASAP7_75t_R _32200_ (.A(_11228_),
    .Y(_11229_));
 BUFx4f_ASAP7_75t_R _32201_ (.A(_11229_),
    .Y(_11230_));
 AO21x1_ASAP7_75t_R _32202_ (.A1(_13901_),
    .A2(_13941_),
    .B(_11230_),
    .Y(_11231_));
 NAND2x2_ASAP7_75t_R _32203_ (.A(_11225_),
    .B(_08551_),
    .Y(_11232_));
 NAND2x1_ASAP7_75t_R _32204_ (.A(_00447_),
    .B(_11232_),
    .Y(_11233_));
 BUFx6f_ASAP7_75t_R _32205_ (.A(_05096_),
    .Y(_11234_));
 BUFx4f_ASAP7_75t_R _32206_ (.A(_11234_),
    .Y(_11235_));
 BUFx4f_ASAP7_75t_R _32207_ (.A(_08551_),
    .Y(_11236_));
 AND2x4_ASAP7_75t_R _32208_ (.A(_11225_),
    .B(_11236_),
    .Y(_11237_));
 OAI21x1_ASAP7_75t_R _32209_ (.A1(_00104_),
    .A2(_11235_),
    .B(_11237_),
    .Y(_11238_));
 AO32x1_ASAP7_75t_R _32210_ (.A1(_11218_),
    .A2(_11227_),
    .A3(_11231_),
    .B1(_11233_),
    .B2(_11238_),
    .Y(_03882_));
 BUFx4f_ASAP7_75t_R _32211_ (.A(_08136_),
    .Y(_11239_));
 BUFx4f_ASAP7_75t_R _32212_ (.A(_08298_),
    .Y(_11240_));
 BUFx4f_ASAP7_75t_R _32213_ (.A(_08271_),
    .Y(_11241_));
 NAND2x1_ASAP7_75t_R _32214_ (.A(_00414_),
    .B(_11241_),
    .Y(_11242_));
 OA21x2_ASAP7_75t_R _32215_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_11240_),
    .B(_11242_),
    .Y(_11243_));
 AOI21x1_ASAP7_75t_R _32216_ (.A1(_00072_),
    .A2(_08299_),
    .B(_08137_),
    .Y(_11244_));
 AO21x1_ASAP7_75t_R _32217_ (.A1(_11239_),
    .A2(_11243_),
    .B(_11244_),
    .Y(_11245_));
 BUFx3_ASAP7_75t_R _32218_ (.A(_11161_),
    .Y(_11246_));
 AO21x1_ASAP7_75t_R _32219_ (.A1(_05139_),
    .A2(\alu_adder_result_ex[1] ),
    .B(_11152_),
    .Y(_11247_));
 AO221x1_ASAP7_75t_R _32220_ (.A1(_05092_),
    .A2(_11157_),
    .B1(_11245_),
    .B2(_11246_),
    .C(_11247_),
    .Y(_11248_));
 OA21x2_ASAP7_75t_R _32221_ (.A1(_05531_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11249_));
 OR3x1_ASAP7_75t_R _32222_ (.A(_00137_),
    .B(_11234_),
    .C(_11232_),
    .Y(_11250_));
 OAI21x1_ASAP7_75t_R _32223_ (.A1(_00414_),
    .A2(_11237_),
    .B(_11250_),
    .Y(_11251_));
 AO21x1_ASAP7_75t_R _32224_ (.A1(_11248_),
    .A2(_11249_),
    .B(_11251_),
    .Y(_03883_));
 BUFx4f_ASAP7_75t_R _32225_ (.A(_11232_),
    .Y(_11252_));
 NAND2x1_ASAP7_75t_R _32226_ (.A(_00073_),
    .B(_11155_),
    .Y(_11253_));
 AO21x1_ASAP7_75t_R _32227_ (.A1(_11158_),
    .A2(_08293_),
    .B(_11253_),
    .Y(_11254_));
 BUFx3_ASAP7_75t_R _32228_ (.A(_08262_),
    .Y(_11255_));
 BUFx3_ASAP7_75t_R _32229_ (.A(_08263_),
    .Y(_11256_));
 AO21x1_ASAP7_75t_R _32230_ (.A1(_11255_),
    .A2(_11256_),
    .B(_05677_),
    .Y(_11257_));
 OA21x2_ASAP7_75t_R _32231_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_11241_),
    .B(_11257_),
    .Y(_11258_));
 OA21x2_ASAP7_75t_R _32232_ (.A1(_11155_),
    .A2(_11258_),
    .B(_11246_),
    .Y(_11259_));
 AO21x1_ASAP7_75t_R _32233_ (.A1(_05555_),
    .A2(\alu_adder_result_ex[2] ),
    .B(_11152_),
    .Y(_11260_));
 AO221x1_ASAP7_75t_R _32234_ (.A1(_05092_),
    .A2(_11243_),
    .B1(_11254_),
    .B2(_11259_),
    .C(_11260_),
    .Y(_11261_));
 OA21x2_ASAP7_75t_R _32235_ (.A1(_05196_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11262_));
 INVx1_ASAP7_75t_R _32236_ (.A(_00140_),
    .Y(_11263_));
 BUFx4f_ASAP7_75t_R _32237_ (.A(_09361_),
    .Y(_11264_));
 AND3x1_ASAP7_75t_R _32238_ (.A(_11263_),
    .B(_11264_),
    .C(_11237_),
    .Y(_11265_));
 AO221x1_ASAP7_75t_R _32239_ (.A1(_05677_),
    .A2(_11252_),
    .B1(_11261_),
    .B2(_11262_),
    .C(_11265_),
    .Y(_03884_));
 NAND2x1_ASAP7_75t_R _32240_ (.A(_00075_),
    .B(_11155_),
    .Y(_11266_));
 AO21x1_ASAP7_75t_R _32241_ (.A1(_11158_),
    .A2(_08296_),
    .B(_11266_),
    .Y(_11267_));
 BUFx4f_ASAP7_75t_R _32242_ (.A(_11154_),
    .Y(_11268_));
 AO21x1_ASAP7_75t_R _32243_ (.A1(_11255_),
    .A2(_11256_),
    .B(_05545_),
    .Y(_11269_));
 OA21x2_ASAP7_75t_R _32244_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_11240_),
    .B(_11269_),
    .Y(_11270_));
 OA21x2_ASAP7_75t_R _32245_ (.A1(_11268_),
    .A2(_11270_),
    .B(_11246_),
    .Y(_11271_));
 BUFx4f_ASAP7_75t_R _32246_ (.A(_04871_),
    .Y(_11272_));
 AO221x1_ASAP7_75t_R _32247_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[3] ),
    .B1(_11258_),
    .B2(_05092_),
    .C(_11152_),
    .Y(_11273_));
 AO21x1_ASAP7_75t_R _32248_ (.A1(_11267_),
    .A2(_11271_),
    .B(_11273_),
    .Y(_11274_));
 OA21x2_ASAP7_75t_R _32249_ (.A1(_05204_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11275_));
 AND3x1_ASAP7_75t_R _32250_ (.A(_09708_),
    .B(_11264_),
    .C(_11237_),
    .Y(_11276_));
 AO221x1_ASAP7_75t_R _32251_ (.A1(_05545_),
    .A2(_11252_),
    .B1(_11274_),
    .B2(_11275_),
    .C(_11276_),
    .Y(_03885_));
 NAND2x1_ASAP7_75t_R _32252_ (.A(_00076_),
    .B(_11155_),
    .Y(_11277_));
 AO21x1_ASAP7_75t_R _32253_ (.A1(_08285_),
    .A2(_08319_),
    .B(_11277_),
    .Y(_11278_));
 AO21x1_ASAP7_75t_R _32254_ (.A1(_11255_),
    .A2(_11256_),
    .B(_05683_),
    .Y(_11279_));
 OA21x2_ASAP7_75t_R _32255_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_11240_),
    .B(_11279_),
    .Y(_11280_));
 OA21x2_ASAP7_75t_R _32256_ (.A1(_11268_),
    .A2(_11280_),
    .B(_11246_),
    .Y(_11281_));
 AO221x1_ASAP7_75t_R _32257_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[4] ),
    .B1(_11270_),
    .B2(_05092_),
    .C(_11152_),
    .Y(_11282_));
 AO21x1_ASAP7_75t_R _32258_ (.A1(_11278_),
    .A2(_11281_),
    .B(_11282_),
    .Y(_11283_));
 OA21x2_ASAP7_75t_R _32259_ (.A1(_05210_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11284_));
 AND3x1_ASAP7_75t_R _32260_ (.A(_08610_),
    .B(_11264_),
    .C(_11237_),
    .Y(_11285_));
 AO221x1_ASAP7_75t_R _32261_ (.A1(_05683_),
    .A2(_11252_),
    .B1(_11283_),
    .B2(_11284_),
    .C(_11285_),
    .Y(_03886_));
 NAND2x1_ASAP7_75t_R _32262_ (.A(_00077_),
    .B(_11155_),
    .Y(_11286_));
 AO21x1_ASAP7_75t_R _32263_ (.A1(_08319_),
    .A2(_08290_),
    .B(_11286_),
    .Y(_11287_));
 INVx1_ASAP7_75t_R _32264_ (.A(\alu_adder_result_ex[5] ),
    .Y(_11288_));
 BUFx4f_ASAP7_75t_R _32265_ (.A(_08262_),
    .Y(_11289_));
 BUFx4f_ASAP7_75t_R _32266_ (.A(_08263_),
    .Y(_11290_));
 AND3x1_ASAP7_75t_R _32267_ (.A(_11288_),
    .B(_11289_),
    .C(_11290_),
    .Y(_11291_));
 AO21x1_ASAP7_75t_R _32268_ (.A1(_00801_),
    .A2(_08272_),
    .B(_11291_),
    .Y(_11292_));
 AOI21x1_ASAP7_75t_R _32269_ (.A1(_08138_),
    .A2(_11292_),
    .B(_05157_),
    .Y(_11293_));
 AO221x1_ASAP7_75t_R _32270_ (.A1(_05139_),
    .A2(\alu_adder_result_ex[5] ),
    .B1(_11280_),
    .B2(_05092_),
    .C(_11152_),
    .Y(_11294_));
 AO21x1_ASAP7_75t_R _32271_ (.A1(_11287_),
    .A2(_11293_),
    .B(_11294_),
    .Y(_11295_));
 OA21x2_ASAP7_75t_R _32272_ (.A1(_05553_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11296_));
 OR3x1_ASAP7_75t_R _32273_ (.A(_00158_),
    .B(_11234_),
    .C(_11232_),
    .Y(_11297_));
 OAI21x1_ASAP7_75t_R _32274_ (.A1(_00801_),
    .A2(_11237_),
    .B(_11297_),
    .Y(_11298_));
 AO21x1_ASAP7_75t_R _32275_ (.A1(_11295_),
    .A2(_11296_),
    .B(_11298_),
    .Y(_03887_));
 OR2x2_ASAP7_75t_R _32276_ (.A(_14225_),
    .B(_05297_),
    .Y(_11299_));
 OA211x2_ASAP7_75t_R _32277_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_11087_),
    .B(_11299_),
    .C(_11101_),
    .Y(_11300_));
 AO21x1_ASAP7_75t_R _32278_ (.A1(_05546_),
    .A2(_11107_),
    .B(_11300_),
    .Y(_03888_));
 BUFx4f_ASAP7_75t_R _32279_ (.A(_11225_),
    .Y(_11301_));
 AO21x1_ASAP7_75t_R _32280_ (.A1(_08319_),
    .A2(_08293_),
    .B(_08323_),
    .Y(_11302_));
 AND3x1_ASAP7_75t_R _32281_ (.A(_15272_),
    .B(_08262_),
    .C(_08263_),
    .Y(_11303_));
 AO21x1_ASAP7_75t_R _32282_ (.A1(_00804_),
    .A2(_08298_),
    .B(_11303_),
    .Y(_11304_));
 NAND2x1_ASAP7_75t_R _32283_ (.A(_08136_),
    .B(_11304_),
    .Y(_11305_));
 OA211x2_ASAP7_75t_R _32284_ (.A1(_08137_),
    .A2(_11302_),
    .B(_11305_),
    .C(_11246_),
    .Y(_11306_));
 BUFx4f_ASAP7_75t_R _32285_ (.A(_11219_),
    .Y(_11307_));
 BUFx4f_ASAP7_75t_R _32286_ (.A(_11153_),
    .Y(_11308_));
 NOR2x2_ASAP7_75t_R _32287_ (.A(_11307_),
    .B(_11308_),
    .Y(_11309_));
 OA21x2_ASAP7_75t_R _32288_ (.A1(_05523_),
    .A2(_15272_),
    .B(_11219_),
    .Y(_11310_));
 OA21x2_ASAP7_75t_R _32289_ (.A1(_05159_),
    .A2(_11292_),
    .B(_11310_),
    .Y(_11311_));
 AOI21x1_ASAP7_75t_R _32290_ (.A1(_05559_),
    .A2(_11309_),
    .B(_11311_),
    .Y(_11312_));
 OR3x1_ASAP7_75t_R _32291_ (.A(_11264_),
    .B(_11306_),
    .C(_11312_),
    .Y(_11313_));
 BUFx4f_ASAP7_75t_R _32292_ (.A(_11234_),
    .Y(_11314_));
 AO21x1_ASAP7_75t_R _32293_ (.A1(_11236_),
    .A2(_08773_),
    .B(_11314_),
    .Y(_11315_));
 AO32x1_ASAP7_75t_R _32294_ (.A1(_11301_),
    .A2(_11313_),
    .A3(_11315_),
    .B1(_11252_),
    .B2(_05688_),
    .Y(_03889_));
 NAND2x1_ASAP7_75t_R _32295_ (.A(_00079_),
    .B(_11155_),
    .Y(_11316_));
 AO21x1_ASAP7_75t_R _32296_ (.A1(_08319_),
    .A2(_08296_),
    .B(_11316_),
    .Y(_11317_));
 AND3x1_ASAP7_75t_R _32297_ (.A(_15247_),
    .B(_11289_),
    .C(_11290_),
    .Y(_11318_));
 AO21x1_ASAP7_75t_R _32298_ (.A1(_00807_),
    .A2(_08272_),
    .B(_11318_),
    .Y(_11319_));
 AOI21x1_ASAP7_75t_R _32299_ (.A1(_08138_),
    .A2(_11319_),
    .B(_05157_),
    .Y(_11320_));
 OA21x2_ASAP7_75t_R _32300_ (.A1(_05523_),
    .A2(_15247_),
    .B(_11307_),
    .Y(_11321_));
 OA21x2_ASAP7_75t_R _32301_ (.A1(_05160_),
    .A2(_11304_),
    .B(_11321_),
    .Y(_11322_));
 NOR2x1_ASAP7_75t_R _32302_ (.A(_05568_),
    .B(_11229_),
    .Y(_11323_));
 OAI21x1_ASAP7_75t_R _32303_ (.A1(_11322_),
    .A2(_11323_),
    .B(_11234_),
    .Y(_11324_));
 AO21x1_ASAP7_75t_R _32304_ (.A1(_11317_),
    .A2(_11320_),
    .B(_11324_),
    .Y(_11325_));
 AO21x1_ASAP7_75t_R _32305_ (.A1(_11236_),
    .A2(_08826_),
    .B(_11314_),
    .Y(_11326_));
 AO32x1_ASAP7_75t_R _32306_ (.A1(_11301_),
    .A2(_11325_),
    .A3(_11326_),
    .B1(_11252_),
    .B2(_05566_),
    .Y(_03890_));
 AND3x1_ASAP7_75t_R _32307_ (.A(\alu_adder_result_ex[8] ),
    .B(_11289_),
    .C(_11290_),
    .Y(_11327_));
 AO21x1_ASAP7_75t_R _32308_ (.A1(_05571_),
    .A2(_11241_),
    .B(_11327_),
    .Y(_11328_));
 INVx1_ASAP7_75t_R _32309_ (.A(_00080_),
    .Y(_11329_));
 AND4x1_ASAP7_75t_R _32310_ (.A(_05095_),
    .B(_08284_),
    .C(_11158_),
    .D(_08264_),
    .Y(_11330_));
 OR3x1_ASAP7_75t_R _32311_ (.A(_11329_),
    .B(_08136_),
    .C(_11330_),
    .Y(_11331_));
 OA211x2_ASAP7_75t_R _32312_ (.A1(_11155_),
    .A2(_11328_),
    .B(_11331_),
    .C(_11246_),
    .Y(_11332_));
 OA21x2_ASAP7_75t_R _32313_ (.A1(_05523_),
    .A2(_15417_),
    .B(_11219_),
    .Y(_11333_));
 OA21x2_ASAP7_75t_R _32314_ (.A1(_05159_),
    .A2(_11319_),
    .B(_11333_),
    .Y(_11334_));
 AOI21x1_ASAP7_75t_R _32315_ (.A1(_05692_),
    .A2(_11309_),
    .B(_11334_),
    .Y(_11335_));
 OR3x1_ASAP7_75t_R _32316_ (.A(_11264_),
    .B(_11332_),
    .C(_11335_),
    .Y(_11336_));
 AO21x1_ASAP7_75t_R _32317_ (.A1(_11236_),
    .A2(_08866_),
    .B(_11314_),
    .Y(_11337_));
 AO32x1_ASAP7_75t_R _32318_ (.A1(_11301_),
    .A2(_11336_),
    .A3(_11337_),
    .B1(_11252_),
    .B2(_05571_),
    .Y(_03891_));
 AO21x1_ASAP7_75t_R _32319_ (.A1(_11255_),
    .A2(_11256_),
    .B(_05579_),
    .Y(_11338_));
 OA21x2_ASAP7_75t_R _32320_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_08273_),
    .B(_11338_),
    .Y(_11339_));
 AOI21x1_ASAP7_75t_R _32321_ (.A1(_00081_),
    .A2(_08327_),
    .B(_11239_),
    .Y(_11340_));
 AO21x1_ASAP7_75t_R _32322_ (.A1(_08138_),
    .A2(_11339_),
    .B(_11340_),
    .Y(_11341_));
 AO221x1_ASAP7_75t_R _32323_ (.A1(_05139_),
    .A2(\alu_adder_result_ex[9] ),
    .B1(_11328_),
    .B2(_05092_),
    .C(_11152_),
    .Y(_11342_));
 AO21x1_ASAP7_75t_R _32324_ (.A1(_11246_),
    .A2(_11341_),
    .B(_11342_),
    .Y(_11343_));
 AND2x2_ASAP7_75t_R _32325_ (.A(_15365_),
    .B(_15390_),
    .Y(_11344_));
 OA21x2_ASAP7_75t_R _32326_ (.A1(_11344_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11345_));
 OR3x1_ASAP7_75t_R _32327_ (.A(_11234_),
    .B(_08935_),
    .C(_11232_),
    .Y(_11346_));
 OAI21x1_ASAP7_75t_R _32328_ (.A1(_00812_),
    .A2(_11237_),
    .B(_11346_),
    .Y(_11347_));
 AO21x1_ASAP7_75t_R _32329_ (.A1(_11343_),
    .A2(_11345_),
    .B(_11347_),
    .Y(_03892_));
 BUFx4f_ASAP7_75t_R _32330_ (.A(_09361_),
    .Y(_11348_));
 OAI21x1_ASAP7_75t_R _32331_ (.A1(_09186_),
    .A2(_08985_),
    .B(_11348_),
    .Y(_11349_));
 AND5x2_ASAP7_75t_R _32332_ (.A(_15483_),
    .B(_15488_),
    .C(_15489_),
    .D(_11289_),
    .E(_11290_),
    .Y(_11350_));
 AOI21x1_ASAP7_75t_R _32333_ (.A1(_00815_),
    .A2(_11240_),
    .B(_11350_),
    .Y(_11351_));
 OR4x1_ASAP7_75t_R _32334_ (.A(_08148_),
    .B(_08270_),
    .C(_05102_),
    .D(_08298_),
    .Y(_11352_));
 AOI21x1_ASAP7_75t_R _32335_ (.A1(_00082_),
    .A2(_11352_),
    .B(_08137_),
    .Y(_11353_));
 AO21x1_ASAP7_75t_R _32336_ (.A1(_11239_),
    .A2(_11351_),
    .B(_11353_),
    .Y(_11354_));
 BUFx3_ASAP7_75t_R _32337_ (.A(_11151_),
    .Y(_11355_));
 AO21x1_ASAP7_75t_R _32338_ (.A1(_15440_),
    .A2(_15463_),
    .B(_11154_),
    .Y(_11356_));
 AO221x1_ASAP7_75t_R _32339_ (.A1(_05138_),
    .A2(\alu_adder_result_ex[10] ),
    .B1(_11355_),
    .B2(_11356_),
    .C(_09361_),
    .Y(_11357_));
 AO221x1_ASAP7_75t_R _32340_ (.A1(_05092_),
    .A2(_11339_),
    .B1(_11354_),
    .B2(_11246_),
    .C(_11357_),
    .Y(_11358_));
 AO32x1_ASAP7_75t_R _32341_ (.A1(_11301_),
    .A2(_11349_),
    .A3(_11358_),
    .B1(_11252_),
    .B2(_05583_),
    .Y(_03893_));
 OR3x1_ASAP7_75t_R _32342_ (.A(_11314_),
    .B(_09186_),
    .C(_09028_),
    .Y(_11359_));
 AO221x1_ASAP7_75t_R _32343_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[11] ),
    .B1(_11351_),
    .B2(_05091_),
    .C(_11355_),
    .Y(_11360_));
 BUFx6f_ASAP7_75t_R _32344_ (.A(_11229_),
    .Y(_11361_));
 AO21x1_ASAP7_75t_R _32345_ (.A1(_14775_),
    .A2(_14803_),
    .B(_11361_),
    .Y(_11362_));
 AO21x1_ASAP7_75t_R _32346_ (.A1(_11360_),
    .A2(_11362_),
    .B(_11264_),
    .Y(_11363_));
 AND3x2_ASAP7_75t_R _32347_ (.A(_13567_),
    .B(_11161_),
    .C(_05516_),
    .Y(_11364_));
 NOR2x1_ASAP7_75t_R _32348_ (.A(\alu_adder_result_ex[11] ),
    .B(_11240_),
    .Y(_11365_));
 AO21x1_ASAP7_75t_R _32349_ (.A1(_05506_),
    .A2(_08273_),
    .B(_11365_),
    .Y(_11366_));
 OR4x1_ASAP7_75t_R _32350_ (.A(_08148_),
    .B(_08275_),
    .C(_05103_),
    .D(_11240_),
    .Y(_11367_));
 AO21x1_ASAP7_75t_R _32351_ (.A1(_00083_),
    .A2(_11367_),
    .B(_11239_),
    .Y(_11368_));
 OAI21x1_ASAP7_75t_R _32352_ (.A1(_11268_),
    .A2(_11366_),
    .B(_11368_),
    .Y(_11369_));
 AOI22x1_ASAP7_75t_R _32353_ (.A1(_11359_),
    .A2(_11363_),
    .B1(_11364_),
    .B2(_11369_),
    .Y(_11370_));
 BUFx6f_ASAP7_75t_R _32354_ (.A(_11225_),
    .Y(_11371_));
 AOI22x1_ASAP7_75t_R _32355_ (.A1(_05506_),
    .A2(_11252_),
    .B1(_11370_),
    .B2(_11371_),
    .Y(_03894_));
 AND4x1_ASAP7_75t_R _32356_ (.A(_15737_),
    .B(_15744_),
    .C(_08262_),
    .D(_08263_),
    .Y(_11372_));
 AO21x1_ASAP7_75t_R _32357_ (.A1(_00821_),
    .A2(_11241_),
    .B(_11372_),
    .Y(_11373_));
 OA211x2_ASAP7_75t_R _32358_ (.A1(_08259_),
    .A2(_08278_),
    .B(_11308_),
    .C(_00084_),
    .Y(_11374_));
 AO21x1_ASAP7_75t_R _32359_ (.A1(_11239_),
    .A2(_11373_),
    .B(_11374_),
    .Y(_11375_));
 AOI211x1_ASAP7_75t_R _32360_ (.A1(_05506_),
    .A2(_08273_),
    .B(_11365_),
    .C(_05160_),
    .Y(_11376_));
 AO21x1_ASAP7_75t_R _32361_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[12] ),
    .B(_11355_),
    .Y(_11377_));
 OAI22x1_ASAP7_75t_R _32362_ (.A1(_05700_),
    .A2(_11361_),
    .B1(_11376_),
    .B2(_11377_),
    .Y(_11378_));
 OA211x2_ASAP7_75t_R _32363_ (.A1(_05157_),
    .A2(_11375_),
    .B(_11378_),
    .C(_11226_),
    .Y(_11379_));
 AND3x1_ASAP7_75t_R _32364_ (.A(_11348_),
    .B(_09068_),
    .C(_11237_),
    .Y(_11380_));
 AOI211x1_ASAP7_75t_R _32365_ (.A1(_00821_),
    .A2(_11252_),
    .B(_11379_),
    .C(_11380_),
    .Y(_03895_));
 AND3x1_ASAP7_75t_R _32366_ (.A(_15733_),
    .B(_11289_),
    .C(_11290_),
    .Y(_11381_));
 AO21x1_ASAP7_75t_R _32367_ (.A1(_00854_),
    .A2(_08272_),
    .B(_11381_),
    .Y(_11382_));
 OA211x2_ASAP7_75t_R _32368_ (.A1(_05093_),
    .A2(_08278_),
    .B(_11308_),
    .C(_00085_),
    .Y(_11383_));
 AOI211x1_ASAP7_75t_R _32369_ (.A1(_11239_),
    .A2(_11382_),
    .B(_11383_),
    .C(_05156_),
    .Y(_11384_));
 OA21x2_ASAP7_75t_R _32370_ (.A1(_05523_),
    .A2(_15733_),
    .B(_11219_),
    .Y(_11385_));
 OAI21x1_ASAP7_75t_R _32371_ (.A1(_05160_),
    .A2(_11373_),
    .B(_11385_),
    .Y(_11386_));
 OA21x2_ASAP7_75t_R _32372_ (.A1(_05597_),
    .A2(_11229_),
    .B(_11386_),
    .Y(_11387_));
 OR3x1_ASAP7_75t_R _32373_ (.A(_09361_),
    .B(_11384_),
    .C(_11387_),
    .Y(_11388_));
 AO21x1_ASAP7_75t_R _32374_ (.A1(_11236_),
    .A2(_09084_),
    .B(_11314_),
    .Y(_11389_));
 AO32x1_ASAP7_75t_R _32375_ (.A1(_11301_),
    .A2(_11388_),
    .A3(_11389_),
    .B1(_11252_),
    .B2(_05598_),
    .Y(_03896_));
 OAI21x1_ASAP7_75t_R _32376_ (.A1(_08270_),
    .A2(_08278_),
    .B(_00086_),
    .Y(_11390_));
 AND3x1_ASAP7_75t_R _32377_ (.A(\alu_adder_result_ex[14] ),
    .B(_08262_),
    .C(_08263_),
    .Y(_11391_));
 AO21x1_ASAP7_75t_R _32378_ (.A1(_05604_),
    .A2(_08271_),
    .B(_11391_),
    .Y(_11392_));
 OR2x2_ASAP7_75t_R _32379_ (.A(_11154_),
    .B(_11392_),
    .Y(_11393_));
 OA211x2_ASAP7_75t_R _32380_ (.A1(_08137_),
    .A2(_11390_),
    .B(_11393_),
    .C(_11161_),
    .Y(_11394_));
 OA21x2_ASAP7_75t_R _32381_ (.A1(_05523_),
    .A2(_16028_),
    .B(_11219_),
    .Y(_11395_));
 OAI21x1_ASAP7_75t_R _32382_ (.A1(_05159_),
    .A2(_11382_),
    .B(_11395_),
    .Y(_11396_));
 OA21x2_ASAP7_75t_R _32383_ (.A1(_05603_),
    .A2(_11229_),
    .B(_11396_),
    .Y(_11397_));
 OR3x1_ASAP7_75t_R _32384_ (.A(_09361_),
    .B(_11394_),
    .C(_11397_),
    .Y(_11398_));
 OAI21x1_ASAP7_75t_R _32385_ (.A1(_09186_),
    .A2(_09128_),
    .B(_11348_),
    .Y(_11399_));
 AO32x1_ASAP7_75t_R _32386_ (.A1(_11301_),
    .A2(_11398_),
    .A3(_11399_),
    .B1(_11232_),
    .B2(_05604_),
    .Y(_03897_));
 AO21x1_ASAP7_75t_R _32387_ (.A1(_11236_),
    .A2(_09157_),
    .B(_11314_),
    .Y(_11400_));
 NOR2x1_ASAP7_75t_R _32388_ (.A(\alu_adder_result_ex[15] ),
    .B(_11241_),
    .Y(_11401_));
 AO21x1_ASAP7_75t_R _32389_ (.A1(_00920_),
    .A2(_11240_),
    .B(_11401_),
    .Y(_11402_));
 OA211x2_ASAP7_75t_R _32390_ (.A1(_08275_),
    .A2(_08278_),
    .B(_11154_),
    .C(_00087_),
    .Y(_11403_));
 AOI21x1_ASAP7_75t_R _32391_ (.A1(_11239_),
    .A2(_11402_),
    .B(_11403_),
    .Y(_11404_));
 AO21x1_ASAP7_75t_R _32392_ (.A1(_15978_),
    .A2(_16002_),
    .B(_11154_),
    .Y(_11405_));
 AO221x1_ASAP7_75t_R _32393_ (.A1(_05138_),
    .A2(\alu_adder_result_ex[15] ),
    .B1(_11355_),
    .B2(_11405_),
    .C(_09361_),
    .Y(_11406_));
 AO221x1_ASAP7_75t_R _32394_ (.A1(_05092_),
    .A2(_11392_),
    .B1(_11404_),
    .B2(_11246_),
    .C(_11406_),
    .Y(_11407_));
 AO32x1_ASAP7_75t_R _32395_ (.A1(_11301_),
    .A2(_11400_),
    .A3(_11407_),
    .B1(_11232_),
    .B2(_05609_),
    .Y(_03898_));
 OR2x2_ASAP7_75t_R _32396_ (.A(_14295_),
    .B(_05296_),
    .Y(_11408_));
 OA211x2_ASAP7_75t_R _32397_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_11087_),
    .B(_11408_),
    .C(_05107_),
    .Y(_11409_));
 AO21x1_ASAP7_75t_R _32398_ (.A1(_05684_),
    .A2(_11107_),
    .B(_11409_),
    .Y(_03899_));
 NOR2x1_ASAP7_75t_R _32399_ (.A(_13595_),
    .B(_11223_),
    .Y(_11410_));
 OR3x1_ASAP7_75t_R _32400_ (.A(_05141_),
    .B(_05143_),
    .C(_11410_),
    .Y(_11411_));
 BUFx3_ASAP7_75t_R _32401_ (.A(_11411_),
    .Y(_11412_));
 BUFx4f_ASAP7_75t_R _32402_ (.A(_11412_),
    .Y(_11413_));
 INVx1_ASAP7_75t_R _32403_ (.A(\alu_adder_result_ex[16] ),
    .Y(_11414_));
 AND3x1_ASAP7_75t_R _32404_ (.A(_11414_),
    .B(_11289_),
    .C(_11290_),
    .Y(_11415_));
 AO21x1_ASAP7_75t_R _32405_ (.A1(_05180_),
    .A2(_11241_),
    .B(_11415_),
    .Y(_11416_));
 NAND2x1_ASAP7_75t_R _32406_ (.A(_08285_),
    .B(_08286_),
    .Y(_11417_));
 AND2x2_ASAP7_75t_R _32407_ (.A(_00088_),
    .B(_11155_),
    .Y(_11418_));
 AO221x1_ASAP7_75t_R _32408_ (.A1(_11239_),
    .A2(_11416_),
    .B1(_11417_),
    .B2(_11418_),
    .C(_05156_),
    .Y(_11419_));
 OA21x2_ASAP7_75t_R _32409_ (.A1(_05622_),
    .A2(_11414_),
    .B(_11307_),
    .Y(_11420_));
 OA21x2_ASAP7_75t_R _32410_ (.A1(_05160_),
    .A2(_11402_),
    .B(_11420_),
    .Y(_11421_));
 OAI21x1_ASAP7_75t_R _32411_ (.A1(_05169_),
    .A2(_11230_),
    .B(_11235_),
    .Y(_11422_));
 AO21x1_ASAP7_75t_R _32412_ (.A1(_11419_),
    .A2(_11421_),
    .B(_11422_),
    .Y(_11423_));
 AOI21x1_ASAP7_75t_R _32413_ (.A1(_11348_),
    .A2(_09193_),
    .B(_11413_),
    .Y(_11424_));
 AOI22x1_ASAP7_75t_R _32414_ (.A1(_05180_),
    .A2(_11413_),
    .B1(_11423_),
    .B2(_11424_),
    .Y(_03900_));
 INVx1_ASAP7_75t_R _32415_ (.A(_09238_),
    .Y(_11425_));
 AOI21x1_ASAP7_75t_R _32416_ (.A1(_05138_),
    .A2(\alu_adder_result_ex[17] ),
    .B(_11151_),
    .Y(_11426_));
 OAI21x1_ASAP7_75t_R _32417_ (.A1(_05160_),
    .A2(_11416_),
    .B(_11426_),
    .Y(_11427_));
 OA211x2_ASAP7_75t_R _32418_ (.A1(_05189_),
    .A2(_11361_),
    .B(_11427_),
    .C(_11234_),
    .Y(_11428_));
 AO21x1_ASAP7_75t_R _32419_ (.A1(_11348_),
    .A2(_11425_),
    .B(_11428_),
    .Y(_11429_));
 NAND2x1_ASAP7_75t_R _32420_ (.A(_00089_),
    .B(_11268_),
    .Y(_11430_));
 AO21x1_ASAP7_75t_R _32421_ (.A1(_08286_),
    .A2(_08290_),
    .B(_11430_),
    .Y(_11431_));
 AO21x1_ASAP7_75t_R _32422_ (.A1(_11289_),
    .A2(_11290_),
    .B(_05710_),
    .Y(_11432_));
 OA21x2_ASAP7_75t_R _32423_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_11241_),
    .B(_11432_),
    .Y(_11433_));
 OA21x2_ASAP7_75t_R _32424_ (.A1(_11268_),
    .A2(_11433_),
    .B(_11364_),
    .Y(_11434_));
 AO21x1_ASAP7_75t_R _32425_ (.A1(_11431_),
    .A2(_11434_),
    .B(_11412_),
    .Y(_11435_));
 OA22x2_ASAP7_75t_R _32426_ (.A1(_05710_),
    .A2(_11371_),
    .B1(_11429_),
    .B2(_11435_),
    .Y(_03901_));
 AOI211x1_ASAP7_75t_R _32427_ (.A1(_08286_),
    .A2(_08293_),
    .B(_08294_),
    .C(_08138_),
    .Y(_11436_));
 AND3x1_ASAP7_75t_R _32428_ (.A(_16531_),
    .B(_11289_),
    .C(_11290_),
    .Y(_11437_));
 AO21x1_ASAP7_75t_R _32429_ (.A1(_01019_),
    .A2(_08272_),
    .B(_11437_),
    .Y(_11438_));
 AO21x1_ASAP7_75t_R _32430_ (.A1(_08138_),
    .A2(_11438_),
    .B(_05157_),
    .Y(_11439_));
 AND2x2_ASAP7_75t_R _32431_ (.A(_05091_),
    .B(_11433_),
    .Y(_11440_));
 AO21x1_ASAP7_75t_R _32432_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[18] ),
    .B(_11355_),
    .Y(_11441_));
 OAI22x1_ASAP7_75t_R _32433_ (.A1(_05715_),
    .A2(_11361_),
    .B1(_11440_),
    .B2(_11441_),
    .Y(_11442_));
 OA211x2_ASAP7_75t_R _32434_ (.A1(_11436_),
    .A2(_11439_),
    .B(_11442_),
    .C(_11235_),
    .Y(_11443_));
 AO21x1_ASAP7_75t_R _32435_ (.A1(_11348_),
    .A2(_09266_),
    .B(_11413_),
    .Y(_11444_));
 OAI22x1_ASAP7_75t_R _32436_ (.A1(_01019_),
    .A2(_11371_),
    .B1(_11443_),
    .B2(_11444_),
    .Y(_03902_));
 AO21x1_ASAP7_75t_R _32437_ (.A1(_11255_),
    .A2(_11256_),
    .B(_05623_),
    .Y(_11445_));
 OA21x2_ASAP7_75t_R _32438_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_11240_),
    .B(_11445_),
    .Y(_11446_));
 NAND2x1_ASAP7_75t_R _32439_ (.A(_00091_),
    .B(_11154_),
    .Y(_11447_));
 AO21x1_ASAP7_75t_R _32440_ (.A1(_08286_),
    .A2(_08296_),
    .B(_11447_),
    .Y(_11448_));
 OA211x2_ASAP7_75t_R _32441_ (.A1(_11155_),
    .A2(_11446_),
    .B(_11448_),
    .C(_11246_),
    .Y(_11449_));
 NAND2x1_ASAP7_75t_R _32442_ (.A(_04871_),
    .B(\alu_adder_result_ex[19] ),
    .Y(_11450_));
 OA211x2_ASAP7_75t_R _32443_ (.A1(_05159_),
    .A2(_11438_),
    .B(_11450_),
    .C(_11307_),
    .Y(_11451_));
 NOR2x1_ASAP7_75t_R _32444_ (.A(_05621_),
    .B(_11229_),
    .Y(_11452_));
 OAI21x1_ASAP7_75t_R _32445_ (.A1(_11451_),
    .A2(_11452_),
    .B(_11234_),
    .Y(_11453_));
 NAND2x1_ASAP7_75t_R _32446_ (.A(_09361_),
    .B(_09280_),
    .Y(_11454_));
 OA211x2_ASAP7_75t_R _32447_ (.A1(_11449_),
    .A2(_11453_),
    .B(_11454_),
    .C(_11225_),
    .Y(_11455_));
 AO21x1_ASAP7_75t_R _32448_ (.A1(_05623_),
    .A2(_11413_),
    .B(_11455_),
    .Y(_03903_));
 INVx1_ASAP7_75t_R _32449_ (.A(_05315_),
    .Y(_11456_));
 NOR2x2_ASAP7_75t_R _32450_ (.A(_05100_),
    .B(_05101_),
    .Y(_11457_));
 NAND2x1_ASAP7_75t_R _32451_ (.A(_00092_),
    .B(_11154_),
    .Y(_11458_));
 AO21x1_ASAP7_75t_R _32452_ (.A1(_08285_),
    .A2(_11457_),
    .B(_11458_),
    .Y(_11459_));
 AND3x1_ASAP7_75t_R _32453_ (.A(_16777_),
    .B(_11289_),
    .C(_11290_),
    .Y(_11460_));
 AO21x1_ASAP7_75t_R _32454_ (.A1(_05315_),
    .A2(_08272_),
    .B(_11460_),
    .Y(_11461_));
 AOI21x1_ASAP7_75t_R _32455_ (.A1(_08137_),
    .A2(_11461_),
    .B(_05156_),
    .Y(_11462_));
 AO21x1_ASAP7_75t_R _32456_ (.A1(_05138_),
    .A2(\alu_adder_result_ex[20] ),
    .B(_11355_),
    .Y(_11463_));
 AO221x1_ASAP7_75t_R _32457_ (.A1(_05091_),
    .A2(_11446_),
    .B1(_11459_),
    .B2(_11462_),
    .C(_11463_),
    .Y(_11464_));
 OA21x2_ASAP7_75t_R _32458_ (.A1(_05631_),
    .A2(_11361_),
    .B(_11234_),
    .Y(_11465_));
 AO221x1_ASAP7_75t_R _32459_ (.A1(_11264_),
    .A2(_09315_),
    .B1(_11464_),
    .B2(_11465_),
    .C(_11412_),
    .Y(_11466_));
 OA21x2_ASAP7_75t_R _32460_ (.A1(_11456_),
    .A2(_11371_),
    .B(_11466_),
    .Y(_03904_));
 NOR2x1_ASAP7_75t_R _32461_ (.A(_05160_),
    .B(_11461_),
    .Y(_11467_));
 AO21x1_ASAP7_75t_R _32462_ (.A1(_05138_),
    .A2(\alu_adder_result_ex[21] ),
    .B(_11355_),
    .Y(_11468_));
 OA22x2_ASAP7_75t_R _32463_ (.A1(_05217_),
    .A2(_11361_),
    .B1(_11467_),
    .B2(_11468_),
    .Y(_11469_));
 NOR2x1_ASAP7_75t_R _32464_ (.A(_11314_),
    .B(_09343_),
    .Y(_11470_));
 AO21x1_ASAP7_75t_R _32465_ (.A1(_11235_),
    .A2(_11469_),
    .B(_11470_),
    .Y(_11471_));
 NAND2x1_ASAP7_75t_R _32466_ (.A(_00093_),
    .B(_11268_),
    .Y(_11472_));
 AO21x1_ASAP7_75t_R _32467_ (.A1(_08290_),
    .A2(_11457_),
    .B(_11472_),
    .Y(_11473_));
 AO21x1_ASAP7_75t_R _32468_ (.A1(_11255_),
    .A2(_11256_),
    .B(_05722_),
    .Y(_11474_));
 OA21x2_ASAP7_75t_R _32469_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_11241_),
    .B(_11474_),
    .Y(_11475_));
 OA21x2_ASAP7_75t_R _32470_ (.A1(_11268_),
    .A2(_11475_),
    .B(_11364_),
    .Y(_11476_));
 AO21x1_ASAP7_75t_R _32471_ (.A1(_11473_),
    .A2(_11476_),
    .B(_11412_),
    .Y(_11477_));
 OA22x2_ASAP7_75t_R _32472_ (.A1(_05722_),
    .A2(_11371_),
    .B1(_11471_),
    .B2(_11477_),
    .Y(_03905_));
 AND3x1_ASAP7_75t_R _32473_ (.A(_17017_),
    .B(_11255_),
    .C(_11256_),
    .Y(_11478_));
 AO21x1_ASAP7_75t_R _32474_ (.A1(_05316_),
    .A2(_11240_),
    .B(_11478_),
    .Y(_11479_));
 NAND2x1_ASAP7_75t_R _32475_ (.A(_08293_),
    .B(_11457_),
    .Y(_11480_));
 AND2x2_ASAP7_75t_R _32476_ (.A(_00094_),
    .B(_11308_),
    .Y(_11481_));
 AO221x1_ASAP7_75t_R _32477_ (.A1(_11239_),
    .A2(_11479_),
    .B1(_11480_),
    .B2(_11481_),
    .C(_05156_),
    .Y(_11482_));
 AO221x1_ASAP7_75t_R _32478_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[22] ),
    .B1(_11475_),
    .B2(_05091_),
    .C(_11355_),
    .Y(_11483_));
 OAI21x1_ASAP7_75t_R _32479_ (.A1(_05225_),
    .A2(_11361_),
    .B(_11483_),
    .Y(_11484_));
 AND3x1_ASAP7_75t_R _32480_ (.A(_11235_),
    .B(_11482_),
    .C(_11484_),
    .Y(_11485_));
 AO21x1_ASAP7_75t_R _32481_ (.A1(_11348_),
    .A2(_09369_),
    .B(_11412_),
    .Y(_11486_));
 OAI22x1_ASAP7_75t_R _32482_ (.A1(_05316_),
    .A2(_11371_),
    .B1(_11485_),
    .B2(_11486_),
    .Y(_03906_));
 AND3x1_ASAP7_75t_R _32483_ (.A(_17002_),
    .B(_11255_),
    .C(_11256_),
    .Y(_11487_));
 AND2x2_ASAP7_75t_R _32484_ (.A(_01184_),
    .B(_08298_),
    .Y(_11488_));
 OA21x2_ASAP7_75t_R _32485_ (.A1(_11487_),
    .A2(_11488_),
    .B(_08137_),
    .Y(_11489_));
 INVx1_ASAP7_75t_R _32486_ (.A(_00095_),
    .Y(_11490_));
 AOI211x1_ASAP7_75t_R _32487_ (.A1(_08296_),
    .A2(_11457_),
    .B(_11490_),
    .C(_08137_),
    .Y(_11491_));
 OR3x1_ASAP7_75t_R _32488_ (.A(_05156_),
    .B(_11489_),
    .C(_11491_),
    .Y(_11492_));
 OA21x2_ASAP7_75t_R _32489_ (.A1(_05544_),
    .A2(_17002_),
    .B(_11307_),
    .Y(_11493_));
 OA211x2_ASAP7_75t_R _32490_ (.A1(_05160_),
    .A2(_11479_),
    .B(_11492_),
    .C(_11493_),
    .Y(_11494_));
 OAI21x1_ASAP7_75t_R _32491_ (.A1(_05234_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11495_));
 OA21x2_ASAP7_75t_R _32492_ (.A1(_11314_),
    .A2(_09397_),
    .B(_11225_),
    .Y(_11496_));
 AO21x1_ASAP7_75t_R _32493_ (.A1(_01184_),
    .A2(_11413_),
    .B(_11496_),
    .Y(_11497_));
 OAI21x1_ASAP7_75t_R _32494_ (.A1(_11494_),
    .A2(_11495_),
    .B(_11497_),
    .Y(_03907_));
 AND3x1_ASAP7_75t_R _32495_ (.A(_17257_),
    .B(_11255_),
    .C(_11256_),
    .Y(_11498_));
 AO21x1_ASAP7_75t_R _32496_ (.A1(_05317_),
    .A2(_11240_),
    .B(_11498_),
    .Y(_11499_));
 OA211x2_ASAP7_75t_R _32497_ (.A1(_08259_),
    .A2(_08307_),
    .B(_11308_),
    .C(_00096_),
    .Y(_11500_));
 AO21x1_ASAP7_75t_R _32498_ (.A1(_08138_),
    .A2(_11499_),
    .B(_11500_),
    .Y(_11501_));
 OR3x1_ASAP7_75t_R _32499_ (.A(_05159_),
    .B(_11487_),
    .C(_11488_),
    .Y(_11502_));
 NAND2x1_ASAP7_75t_R _32500_ (.A(_11272_),
    .B(\alu_adder_result_ex[24] ),
    .Y(_11503_));
 INVx1_ASAP7_75t_R _32501_ (.A(_05241_),
    .Y(_11504_));
 AO32x1_ASAP7_75t_R _32502_ (.A1(_11307_),
    .A2(_11502_),
    .A3(_11503_),
    .B1(_11309_),
    .B2(_11504_),
    .Y(_11505_));
 OA211x2_ASAP7_75t_R _32503_ (.A1(_05157_),
    .A2(_11501_),
    .B(_11505_),
    .C(_11235_),
    .Y(_11506_));
 OAI21x1_ASAP7_75t_R _32504_ (.A1(_11235_),
    .A2(_09424_),
    .B(_11301_),
    .Y(_11507_));
 OAI22x1_ASAP7_75t_R _32505_ (.A1(_05317_),
    .A2(_11371_),
    .B1(_11506_),
    .B2(_11507_),
    .Y(_03908_));
 AO21x1_ASAP7_75t_R _32506_ (.A1(_08932_),
    .A2(_09466_),
    .B(_09468_),
    .Y(_11508_));
 NOR2x1_ASAP7_75t_R _32507_ (.A(_05645_),
    .B(_11301_),
    .Y(_11509_));
 NOR2x1_ASAP7_75t_R _32508_ (.A(\alu_adder_result_ex[25] ),
    .B(_08272_),
    .Y(_11510_));
 AND2x2_ASAP7_75t_R _32509_ (.A(_01250_),
    .B(_08298_),
    .Y(_11511_));
 OA21x2_ASAP7_75t_R _32510_ (.A1(_11510_),
    .A2(_11511_),
    .B(_08137_),
    .Y(_11512_));
 OA211x2_ASAP7_75t_R _32511_ (.A1(_05093_),
    .A2(_08307_),
    .B(_11308_),
    .C(_00097_),
    .Y(_11513_));
 OR3x1_ASAP7_75t_R _32512_ (.A(_05156_),
    .B(_11512_),
    .C(_11513_),
    .Y(_11514_));
 NOR2x1_ASAP7_75t_R _32513_ (.A(_05160_),
    .B(_11499_),
    .Y(_11515_));
 AO21x1_ASAP7_75t_R _32514_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[25] ),
    .B(_11152_),
    .Y(_11516_));
 OAI22x1_ASAP7_75t_R _32515_ (.A1(_05249_),
    .A2(_11361_),
    .B1(_11515_),
    .B2(_11516_),
    .Y(_11517_));
 AND3x1_ASAP7_75t_R _32516_ (.A(_11227_),
    .B(_11514_),
    .C(_11517_),
    .Y(_11518_));
 AOI211x1_ASAP7_75t_R _32517_ (.A1(_11301_),
    .A2(_11508_),
    .B(_11509_),
    .C(_11518_),
    .Y(_03909_));
 OR2x2_ASAP7_75t_R _32518_ (.A(_14371_),
    .B(_05297_),
    .Y(_11519_));
 OA211x2_ASAP7_75t_R _32519_ (.A1(_11288_),
    .A2(_11093_),
    .B(_11519_),
    .C(_11095_),
    .Y(_11520_));
 AOI21x1_ASAP7_75t_R _32520_ (.A1(_01748_),
    .A2(_11092_),
    .B(_11520_),
    .Y(_03910_));
 NAND2x1_ASAP7_75t_R _32521_ (.A(_05318_),
    .B(_08298_),
    .Y(_11521_));
 OAI21x1_ASAP7_75t_R _32522_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_08273_),
    .B(_11521_),
    .Y(_11522_));
 OA211x2_ASAP7_75t_R _32523_ (.A1(_08270_),
    .A2(_08307_),
    .B(_11308_),
    .C(_00098_),
    .Y(_11523_));
 AO21x1_ASAP7_75t_R _32524_ (.A1(_08138_),
    .A2(_11522_),
    .B(_11523_),
    .Y(_11524_));
 OR3x1_ASAP7_75t_R _32525_ (.A(_05159_),
    .B(_11510_),
    .C(_11511_),
    .Y(_11525_));
 NAND2x1_ASAP7_75t_R _32526_ (.A(_11272_),
    .B(\alu_adder_result_ex[26] ),
    .Y(_11526_));
 AO32x1_ASAP7_75t_R _32527_ (.A1(_11307_),
    .A2(_11525_),
    .A3(_11526_),
    .B1(_11309_),
    .B2(_05649_),
    .Y(_11527_));
 OA211x2_ASAP7_75t_R _32528_ (.A1(_05157_),
    .A2(_11524_),
    .B(_11527_),
    .C(_11235_),
    .Y(_11528_));
 AO21x1_ASAP7_75t_R _32529_ (.A1(_11348_),
    .A2(_09487_),
    .B(_11412_),
    .Y(_11529_));
 OAI22x1_ASAP7_75t_R _32530_ (.A1(_05318_),
    .A2(_11371_),
    .B1(_11528_),
    .B2(_11529_),
    .Y(_03911_));
 AO21x1_ASAP7_75t_R _32531_ (.A1(_11255_),
    .A2(_11256_),
    .B(_05738_),
    .Y(_11530_));
 OAI21x1_ASAP7_75t_R _32532_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_08273_),
    .B(_11530_),
    .Y(_11531_));
 OA211x2_ASAP7_75t_R _32533_ (.A1(_08275_),
    .A2(_08307_),
    .B(_11308_),
    .C(_00099_),
    .Y(_11532_));
 AOI211x1_ASAP7_75t_R _32534_ (.A1(_11239_),
    .A2(_11531_),
    .B(_11532_),
    .C(_05156_),
    .Y(_11533_));
 OA211x2_ASAP7_75t_R _32535_ (.A1(\alu_adder_result_ex[26] ),
    .A2(_11241_),
    .B(_11521_),
    .C(_05091_),
    .Y(_11534_));
 AO21x1_ASAP7_75t_R _32536_ (.A1(_05138_),
    .A2(\alu_adder_result_ex[27] ),
    .B(_11355_),
    .Y(_11535_));
 OA22x2_ASAP7_75t_R _32537_ (.A1(_05265_),
    .A2(_11229_),
    .B1(_11534_),
    .B2(_11535_),
    .Y(_11536_));
 OR3x1_ASAP7_75t_R _32538_ (.A(_11264_),
    .B(_11533_),
    .C(_11536_),
    .Y(_11537_));
 AND2x2_ASAP7_75t_R _32539_ (.A(_09500_),
    .B(_09501_),
    .Y(_11538_));
 OA21x2_ASAP7_75t_R _32540_ (.A1(_11314_),
    .A2(_11538_),
    .B(_11225_),
    .Y(_11539_));
 AO22x1_ASAP7_75t_R _32541_ (.A1(_05738_),
    .A2(_11413_),
    .B1(_11537_),
    .B2(_11539_),
    .Y(_03912_));
 OA211x2_ASAP7_75t_R _32542_ (.A1(_08259_),
    .A2(_08312_),
    .B(_11268_),
    .C(_00100_),
    .Y(_11540_));
 NAND2x1_ASAP7_75t_R _32543_ (.A(_05319_),
    .B(_11241_),
    .Y(_11541_));
 OAI21x1_ASAP7_75t_R _32544_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_08273_),
    .B(_11541_),
    .Y(_11542_));
 AO21x1_ASAP7_75t_R _32545_ (.A1(_08138_),
    .A2(_11542_),
    .B(_05157_),
    .Y(_11543_));
 OA21x2_ASAP7_75t_R _32546_ (.A1(_05622_),
    .A2(_05135_),
    .B(_11307_),
    .Y(_11544_));
 OA21x2_ASAP7_75t_R _32547_ (.A1(_05160_),
    .A2(_11531_),
    .B(_11544_),
    .Y(_11545_));
 OAI21x1_ASAP7_75t_R _32548_ (.A1(_11540_),
    .A2(_11543_),
    .B(_11545_),
    .Y(_11546_));
 OA21x2_ASAP7_75t_R _32549_ (.A1(_05273_),
    .A2(_11230_),
    .B(_11227_),
    .Y(_11547_));
 NOR2x1_ASAP7_75t_R _32550_ (.A(_05319_),
    .B(_11225_),
    .Y(_11548_));
 AO221x1_ASAP7_75t_R _32551_ (.A1(_05145_),
    .A2(_09520_),
    .B1(_11546_),
    .B2(_11547_),
    .C(_11548_),
    .Y(_03913_));
 AND3x1_ASAP7_75t_R _32552_ (.A(_11142_),
    .B(_11289_),
    .C(_11290_),
    .Y(_11549_));
 AO21x1_ASAP7_75t_R _32553_ (.A1(_01382_),
    .A2(_08272_),
    .B(_11549_),
    .Y(_11550_));
 OA211x2_ASAP7_75t_R _32554_ (.A1(_05093_),
    .A2(_08312_),
    .B(_11308_),
    .C(_00101_),
    .Y(_11551_));
 AO21x1_ASAP7_75t_R _32555_ (.A1(_08138_),
    .A2(_11550_),
    .B(_11551_),
    .Y(_11552_));
 OA211x2_ASAP7_75t_R _32556_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_08273_),
    .B(_11541_),
    .C(_05091_),
    .Y(_11553_));
 AO21x1_ASAP7_75t_R _32557_ (.A1(_11272_),
    .A2(\alu_adder_result_ex[29] ),
    .B(_11355_),
    .Y(_11554_));
 OAI22x1_ASAP7_75t_R _32558_ (.A1(_05281_),
    .A2(_11361_),
    .B1(_11553_),
    .B2(_11554_),
    .Y(_11555_));
 OA211x2_ASAP7_75t_R _32559_ (.A1(_05157_),
    .A2(_11552_),
    .B(_11555_),
    .C(_11314_),
    .Y(_11556_));
 AO21x1_ASAP7_75t_R _32560_ (.A1(_11348_),
    .A2(_09564_),
    .B(_11412_),
    .Y(_11557_));
 OAI22x1_ASAP7_75t_R _32561_ (.A1(_01382_),
    .A2(_11371_),
    .B1(_11556_),
    .B2(_11557_),
    .Y(_03914_));
 OA211x2_ASAP7_75t_R _32562_ (.A1(_08270_),
    .A2(_08312_),
    .B(_11308_),
    .C(_00102_),
    .Y(_11558_));
 AND3x1_ASAP7_75t_R _32563_ (.A(_04917_),
    .B(_08262_),
    .C(_08263_),
    .Y(_11559_));
 AO21x1_ASAP7_75t_R _32564_ (.A1(_05320_),
    .A2(_08298_),
    .B(_11559_),
    .Y(_11560_));
 AO21x1_ASAP7_75t_R _32565_ (.A1(_08137_),
    .A2(_11560_),
    .B(_05156_),
    .Y(_11561_));
 OA21x2_ASAP7_75t_R _32566_ (.A1(_05523_),
    .A2(_04917_),
    .B(_11307_),
    .Y(_11562_));
 OA21x2_ASAP7_75t_R _32567_ (.A1(_05159_),
    .A2(_11550_),
    .B(_11562_),
    .Y(_11563_));
 NOR2x1_ASAP7_75t_R _32568_ (.A(_05289_),
    .B(_11229_),
    .Y(_11564_));
 OA221x2_ASAP7_75t_R _32569_ (.A1(_11558_),
    .A2(_11561_),
    .B1(_11563_),
    .B2(_11564_),
    .C(_11234_),
    .Y(_11565_));
 AND2x2_ASAP7_75t_R _32570_ (.A(_08551_),
    .B(_09586_),
    .Y(_11566_));
 OA21x2_ASAP7_75t_R _32571_ (.A1(_09587_),
    .A2(_11566_),
    .B(_09361_),
    .Y(_11567_));
 OR3x1_ASAP7_75t_R _32572_ (.A(_11412_),
    .B(_11565_),
    .C(_11567_),
    .Y(_11568_));
 OAI21x1_ASAP7_75t_R _32573_ (.A1(_05320_),
    .A2(_11371_),
    .B(_11568_),
    .Y(_03915_));
 AO21x1_ASAP7_75t_R _32574_ (.A1(_04898_),
    .A2(_04908_),
    .B(_04868_),
    .Y(_11569_));
 OR4x1_ASAP7_75t_R _32575_ (.A(_08148_),
    .B(_00067_),
    .C(_08271_),
    .D(_08301_),
    .Y(_11570_));
 AND2x2_ASAP7_75t_R _32576_ (.A(_00103_),
    .B(_11154_),
    .Y(_11571_));
 AO221x1_ASAP7_75t_R _32577_ (.A1(_08136_),
    .A2(_11569_),
    .B1(_11570_),
    .B2(_11571_),
    .C(_05156_),
    .Y(_11572_));
 OR2x2_ASAP7_75t_R _32578_ (.A(_05159_),
    .B(_11560_),
    .Y(_11573_));
 AO21x1_ASAP7_75t_R _32579_ (.A1(_04898_),
    .A2(_04908_),
    .B(_05622_),
    .Y(_11574_));
 AND4x1_ASAP7_75t_R _32580_ (.A(_11307_),
    .B(_11572_),
    .C(_11573_),
    .D(_11574_),
    .Y(_11575_));
 NOR2x1_ASAP7_75t_R _32581_ (.A(_04861_),
    .B(_11361_),
    .Y(_11576_));
 OR3x1_ASAP7_75t_R _32582_ (.A(_11348_),
    .B(_11575_),
    .C(_11576_),
    .Y(_11577_));
 XNOR2x1_ASAP7_75t_R _32583_ (.B(_09630_),
    .Y(_11578_),
    .A(_00274_));
 NOR2x1_ASAP7_75t_R _32584_ (.A(_11236_),
    .B(_09157_),
    .Y(_11579_));
 AO21x1_ASAP7_75t_R _32585_ (.A1(_11236_),
    .A2(_11578_),
    .B(_11579_),
    .Y(_11580_));
 OA21x2_ASAP7_75t_R _32586_ (.A1(_11235_),
    .A2(_11580_),
    .B(_11225_),
    .Y(_11581_));
 AOI22x1_ASAP7_75t_R _32587_ (.A1(_04868_),
    .A2(_11413_),
    .B1(_11577_),
    .B2(_11581_),
    .Y(_03916_));
 INVx1_ASAP7_75t_R _32588_ (.A(_00275_),
    .Y(_11582_));
 AOI21x1_ASAP7_75t_R _32589_ (.A1(_09583_),
    .A2(_09585_),
    .B(_11582_),
    .Y(_11583_));
 OA21x2_ASAP7_75t_R _32590_ (.A1(_00274_),
    .A2(_11583_),
    .B(_00281_),
    .Y(_11584_));
 XOR2x1_ASAP7_75t_R _32591_ (.A(_00280_),
    .Y(_11585_),
    .B(_11584_));
 AND3x1_ASAP7_75t_R _32592_ (.A(_11264_),
    .B(_11236_),
    .C(_11585_),
    .Y(_11586_));
 AO32x1_ASAP7_75t_R _32593_ (.A1(_04869_),
    .A2(_05092_),
    .A3(\alu_adder_result_ex[31] ),
    .B1(_11152_),
    .B2(_11268_),
    .Y(_11587_));
 AO21x1_ASAP7_75t_R _32594_ (.A1(_11235_),
    .A2(_11587_),
    .B(_11412_),
    .Y(_11588_));
 NAND2x1_ASAP7_75t_R _32595_ (.A(_01747_),
    .B(_11413_),
    .Y(_11589_));
 OA21x2_ASAP7_75t_R _32596_ (.A1(_11586_),
    .A2(_11588_),
    .B(_11589_),
    .Y(_03917_));
 OA21x2_ASAP7_75t_R _32597_ (.A1(_00274_),
    .A2(_09630_),
    .B(_00281_),
    .Y(_11590_));
 OA21x2_ASAP7_75t_R _32598_ (.A1(_00280_),
    .A2(_11590_),
    .B(_00287_),
    .Y(_11591_));
 XOR2x1_ASAP7_75t_R _32599_ (.A(_18260_),
    .Y(_11592_),
    .B(_02233_));
 XNOR2x1_ASAP7_75t_R _32600_ (.B(_11592_),
    .Y(_11593_),
    .A(_02250_));
 XOR2x1_ASAP7_75t_R _32601_ (.A(net1),
    .Y(_11594_),
    .B(_00286_));
 XNOR2x1_ASAP7_75t_R _32602_ (.B(_00229_),
    .Y(_11595_),
    .A(_00283_));
 XNOR2x1_ASAP7_75t_R _32603_ (.B(_11595_),
    .Y(_11596_),
    .A(_11594_));
 XNOR2x1_ASAP7_75t_R _32604_ (.B(_00282_),
    .Y(_11597_),
    .A(_18227_));
 XNOR2x1_ASAP7_75t_R _32605_ (.B(_11597_),
    .Y(_11598_),
    .A(_11596_));
 XOR2x1_ASAP7_75t_R _32606_ (.A(_00285_),
    .Y(_11599_),
    .B(_00276_));
 XNOR2x1_ASAP7_75t_R _32607_ (.B(_00284_),
    .Y(_11600_),
    .A(_18302_));
 XNOR2x1_ASAP7_75t_R _32608_ (.B(_11600_),
    .Y(_11601_),
    .A(_11599_));
 XNOR2x1_ASAP7_75t_R _32609_ (.B(_02230_),
    .Y(_11602_),
    .A(_02234_));
 XNOR2x1_ASAP7_75t_R _32610_ (.B(_02231_),
    .Y(_11603_),
    .A(_18286_));
 XNOR2x1_ASAP7_75t_R _32611_ (.B(_11603_),
    .Y(_11604_),
    .A(_11602_));
 XNOR2x1_ASAP7_75t_R _32612_ (.B(_11604_),
    .Y(_11605_),
    .A(_11601_));
 XNOR2x1_ASAP7_75t_R _32613_ (.B(_11605_),
    .Y(_11606_),
    .A(_11598_));
 XNOR2x1_ASAP7_75t_R _32614_ (.B(_11606_),
    .Y(_11607_),
    .A(_11593_));
 OA21x2_ASAP7_75t_R _32615_ (.A1(_00232_),
    .A2(_05152_),
    .B(_05312_),
    .Y(_11608_));
 XNOR2x1_ASAP7_75t_R _32616_ (.B(_11608_),
    .Y(_11609_),
    .A(_11607_));
 XNOR2x1_ASAP7_75t_R _32617_ (.B(_11609_),
    .Y(_11610_),
    .A(_11591_));
 AO32x1_ASAP7_75t_R _32618_ (.A1(_11264_),
    .A2(_11236_),
    .A3(_11610_),
    .B1(_11152_),
    .B2(_11268_),
    .Y(_11611_));
 NAND2x1_ASAP7_75t_R _32619_ (.A(_00232_),
    .B(_11413_),
    .Y(_11612_));
 OA21x2_ASAP7_75t_R _32620_ (.A1(_11413_),
    .A2(_11611_),
    .B(_11612_),
    .Y(_03918_));
 OR2x2_ASAP7_75t_R _32621_ (.A(_05558_),
    .B(_05297_),
    .Y(_11613_));
 OA211x2_ASAP7_75t_R _32622_ (.A1(_15272_),
    .A2(_11093_),
    .B(_11613_),
    .C(_11095_),
    .Y(_11614_));
 AOI21x1_ASAP7_75t_R _32623_ (.A1(_01746_),
    .A2(_11092_),
    .B(_11614_),
    .Y(_03919_));
 OR2x2_ASAP7_75t_R _32624_ (.A(_14486_),
    .B(_05296_),
    .Y(_11615_));
 OA211x2_ASAP7_75t_R _32625_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_11087_),
    .B(_11615_),
    .C(_05107_),
    .Y(_11616_));
 AO21x1_ASAP7_75t_R _32626_ (.A1(_05567_),
    .A2(_11083_),
    .B(_11616_),
    .Y(_03920_));
 NAND2x1_ASAP7_75t_R _32627_ (.A(_05230_),
    .B(_11087_),
    .Y(_11617_));
 OA211x2_ASAP7_75t_R _32628_ (.A1(_15417_),
    .A2(_11093_),
    .B(_11617_),
    .C(_11095_),
    .Y(_11618_));
 AOI21x1_ASAP7_75t_R _32629_ (.A1(_01744_),
    .A2(_11092_),
    .B(_11618_),
    .Y(_03921_));
 INVx1_ASAP7_75t_R _32630_ (.A(_02222_),
    .Y(_11619_));
 OR2x2_ASAP7_75t_R _32631_ (.A(_14603_),
    .B(_05296_),
    .Y(_11620_));
 OA211x2_ASAP7_75t_R _32632_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_11087_),
    .B(_11620_),
    .C(_05107_),
    .Y(_11621_));
 AO21x1_ASAP7_75t_R _32633_ (.A1(_11619_),
    .A2(_11083_),
    .B(_11621_),
    .Y(_03922_));
 NAND2x2_ASAP7_75t_R _32634_ (.A(_05467_),
    .B(_05513_),
    .Y(_11622_));
 BUFx6f_ASAP7_75t_R _32635_ (.A(_11622_),
    .Y(_11623_));
 BUFx4f_ASAP7_75t_R _32636_ (.A(_11623_),
    .Y(_11624_));
 AO31x2_ASAP7_75t_R _32637_ (.A1(_15483_),
    .A2(_15488_),
    .A3(_15489_),
    .B(_05422_),
    .Y(_11625_));
 OR2x2_ASAP7_75t_R _32638_ (.A(_11028_),
    .B(_05325_),
    .Y(_11626_));
 AO21x1_ASAP7_75t_R _32639_ (.A1(_04931_),
    .A2(_11626_),
    .B(_05436_),
    .Y(_11627_));
 BUFx4f_ASAP7_75t_R _32640_ (.A(_11627_),
    .Y(_11628_));
 OA222x2_ASAP7_75t_R _32641_ (.A1(_01977_),
    .A2(_05411_),
    .B1(_05415_),
    .B2(_02074_),
    .C1(_11628_),
    .C2(_01467_),
    .Y(_11629_));
 NAND2x1_ASAP7_75t_R _32642_ (.A(net23),
    .B(_05432_),
    .Y(_11630_));
 AND3x4_ASAP7_75t_R _32643_ (.A(_05385_),
    .B(_11629_),
    .C(_11630_),
    .Y(_11631_));
 AND2x2_ASAP7_75t_R _32644_ (.A(_01742_),
    .B(_05465_),
    .Y(_11632_));
 AO21x1_ASAP7_75t_R _32645_ (.A1(_11625_),
    .A2(_11631_),
    .B(_11632_),
    .Y(_11633_));
 OR3x1_ASAP7_75t_R _32646_ (.A(_01950_),
    .B(_05408_),
    .C(_05409_),
    .Y(_11634_));
 OA211x2_ASAP7_75t_R _32647_ (.A1(_01464_),
    .A2(_05416_),
    .B(_07531_),
    .C(_11634_),
    .Y(_11635_));
 OA31x2_ASAP7_75t_R _32648_ (.A1(_15270_),
    .A2(_15271_),
    .A3(_05422_),
    .B1(_11635_),
    .Y(_11636_));
 OA22x2_ASAP7_75t_R _32649_ (.A1(_01716_),
    .A2(_05386_),
    .B1(_05433_),
    .B2(_11636_),
    .Y(_11637_));
 OA22x2_ASAP7_75t_R _32650_ (.A1(_01952_),
    .A2(_05412_),
    .B1(_05416_),
    .B2(_01462_),
    .Y(_11638_));
 OA211x2_ASAP7_75t_R _32651_ (.A1(_05423_),
    .A2(_05128_),
    .B(_07515_),
    .C(_11638_),
    .Y(_11639_));
 OR2x4_ASAP7_75t_R _32652_ (.A(_05433_),
    .B(_11639_),
    .Y(_11640_));
 OA21x2_ASAP7_75t_R _32653_ (.A1(_01718_),
    .A2(_05387_),
    .B(_11640_),
    .Y(_11641_));
 OAI22x1_ASAP7_75t_R _32654_ (.A1(_01951_),
    .A2(_05411_),
    .B1(_05416_),
    .B2(_01463_),
    .Y(_11642_));
 AOI211x1_ASAP7_75t_R _32655_ (.A1(_11035_),
    .A2(\alu_adder_result_ex[5] ),
    .B(_07525_),
    .C(_11642_),
    .Y(_11643_));
 OR2x2_ASAP7_75t_R _32656_ (.A(_05433_),
    .B(_11643_),
    .Y(_11644_));
 BUFx3_ASAP7_75t_R _32657_ (.A(_11644_),
    .Y(_11645_));
 OA21x2_ASAP7_75t_R _32658_ (.A1(_01717_),
    .A2(_05387_),
    .B(_11645_),
    .Y(_11646_));
 OR4x1_ASAP7_75t_R _32659_ (.A(_02292_),
    .B(_11637_),
    .C(_11641_),
    .D(_11646_),
    .Y(_11647_));
 BUFx4f_ASAP7_75t_R _32660_ (.A(_11647_),
    .Y(_11648_));
 OA222x2_ASAP7_75t_R _32661_ (.A1(_01948_),
    .A2(_05410_),
    .B1(_05415_),
    .B2(_02050_),
    .C1(_11628_),
    .C2(_01465_),
    .Y(_11649_));
 INVx1_ASAP7_75t_R _32662_ (.A(_11649_),
    .Y(_11650_));
 AND2x2_ASAP7_75t_R _32663_ (.A(net45),
    .B(_05432_),
    .Y(_11651_));
 OR3x4_ASAP7_75t_R _32664_ (.A(_05425_),
    .B(_11650_),
    .C(_11651_),
    .Y(_11652_));
 AO31x2_ASAP7_75t_R _32665_ (.A1(_15414_),
    .A2(_15416_),
    .A3(_11035_),
    .B(_11652_),
    .Y(_11653_));
 NAND2x2_ASAP7_75t_R _32666_ (.A(_01713_),
    .B(_05425_),
    .Y(_11654_));
 OA22x2_ASAP7_75t_R _32667_ (.A1(_02049_),
    .A2(_05066_),
    .B1(_05408_),
    .B2(_01947_),
    .Y(_11655_));
 OAI22x1_ASAP7_75t_R _32668_ (.A1(_01466_),
    .A2(_11628_),
    .B1(_11655_),
    .B2(_05409_),
    .Y(_11656_));
 AO221x1_ASAP7_75t_R _32669_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_04938_),
    .B1(_05432_),
    .B2(net46),
    .C(_11656_),
    .Y(_11657_));
 OR2x4_ASAP7_75t_R _32670_ (.A(_05425_),
    .B(_11657_),
    .Y(_11658_));
 NAND2x2_ASAP7_75t_R _32671_ (.A(_01714_),
    .B(_05425_),
    .Y(_11659_));
 NAND2x2_ASAP7_75t_R _32672_ (.A(_01715_),
    .B(_05425_),
    .Y(_11660_));
 OAI22x1_ASAP7_75t_R _32673_ (.A1(_01949_),
    .A2(_05410_),
    .B1(_05415_),
    .B2(_02051_),
    .Y(_11661_));
 AND2x2_ASAP7_75t_R _32674_ (.A(\alu_adder_result_ex[7] ),
    .B(_04938_),
    .Y(_11662_));
 OR4x2_ASAP7_75t_R _32675_ (.A(_05425_),
    .B(_05432_),
    .C(_11661_),
    .D(_11662_),
    .Y(_11663_));
 AND5x1_ASAP7_75t_R _32676_ (.A(_11654_),
    .B(_11658_),
    .C(_11659_),
    .D(_11660_),
    .E(_11663_),
    .Y(_11664_));
 NAND2x1_ASAP7_75t_R _32677_ (.A(_11653_),
    .B(_11664_),
    .Y(_11665_));
 NOR2x1_ASAP7_75t_R _32678_ (.A(_11648_),
    .B(_11665_),
    .Y(_11666_));
 XNOR2x1_ASAP7_75t_R _32679_ (.B(_11666_),
    .Y(_11667_),
    .A(_11633_));
 BUFx6f_ASAP7_75t_R _32680_ (.A(_11622_),
    .Y(_11668_));
 NOR2x1_ASAP7_75t_R _32681_ (.A(_01742_),
    .B(_11668_),
    .Y(_11669_));
 AO21x1_ASAP7_75t_R _32682_ (.A1(_11624_),
    .A2(_11667_),
    .B(_11669_),
    .Y(_03923_));
 NAND2x1_ASAP7_75t_R _32683_ (.A(\alu_adder_result_ex[11] ),
    .B(_11035_),
    .Y(_11670_));
 NAND2x1_ASAP7_75t_R _32684_ (.A(net24),
    .B(_05432_),
    .Y(_11671_));
 AO21x1_ASAP7_75t_R _32685_ (.A1(_04931_),
    .A2(_05325_),
    .B(_05436_),
    .Y(_11672_));
 AND2x4_ASAP7_75t_R _32686_ (.A(_05430_),
    .B(_11672_),
    .Y(_11673_));
 OA21x2_ASAP7_75t_R _32687_ (.A1(_04945_),
    .A2(_07786_),
    .B(_05430_),
    .Y(_11674_));
 AND2x2_ASAP7_75t_R _32688_ (.A(_00785_),
    .B(_11674_),
    .Y(_11675_));
 OA222x2_ASAP7_75t_R _32689_ (.A1(_01976_),
    .A2(_05411_),
    .B1(_11673_),
    .B2(_11675_),
    .C1(_05415_),
    .C2(_02073_),
    .Y(_11676_));
 AND4x2_ASAP7_75t_R _32690_ (.A(_05386_),
    .B(_11670_),
    .C(_11671_),
    .D(_11676_),
    .Y(_11677_));
 AOI21x1_ASAP7_75t_R _32691_ (.A1(_01741_),
    .A2(_05466_),
    .B(_11677_),
    .Y(_11678_));
 BUFx6f_ASAP7_75t_R _32692_ (.A(_05432_),
    .Y(_11679_));
 BUFx4f_ASAP7_75t_R _32693_ (.A(_11679_),
    .Y(_11680_));
 OA31x2_ASAP7_75t_R _32694_ (.A1(_11680_),
    .A2(_11639_),
    .A3(_11645_),
    .B1(_05387_),
    .Y(_11681_));
 AND2x2_ASAP7_75t_R _32695_ (.A(_01717_),
    .B(_11645_),
    .Y(_11682_));
 OA21x2_ASAP7_75t_R _32696_ (.A1(_05433_),
    .A2(_11639_),
    .B(_01718_),
    .Y(_11683_));
 OR3x1_ASAP7_75t_R _32697_ (.A(_02290_),
    .B(_05464_),
    .C(_11637_),
    .Y(_11684_));
 OR4x2_ASAP7_75t_R _32698_ (.A(_11681_),
    .B(_11682_),
    .C(_11683_),
    .D(_11684_),
    .Y(_11685_));
 OR3x1_ASAP7_75t_R _32699_ (.A(_11633_),
    .B(_11665_),
    .C(_11685_),
    .Y(_11686_));
 XNOR2x1_ASAP7_75t_R _32700_ (.B(_11686_),
    .Y(_11687_),
    .A(_11678_));
 NOR2x1_ASAP7_75t_R _32701_ (.A(_01741_),
    .B(_11668_),
    .Y(_11688_));
 AO21x1_ASAP7_75t_R _32702_ (.A1(_11624_),
    .A2(_11687_),
    .B(_11688_),
    .Y(_03924_));
 AO21x2_ASAP7_75t_R _32703_ (.A1(_15737_),
    .A2(_15744_),
    .B(_05422_),
    .Y(_11689_));
 OA222x2_ASAP7_75t_R _32704_ (.A1(_01975_),
    .A2(_05411_),
    .B1(_05415_),
    .B2(_02072_),
    .C1(_11628_),
    .C2(_00784_),
    .Y(_11690_));
 INVx1_ASAP7_75t_R _32705_ (.A(_11690_),
    .Y(_11691_));
 AND2x2_ASAP7_75t_R _32706_ (.A(net25),
    .B(_05432_),
    .Y(_11692_));
 OR3x1_ASAP7_75t_R _32707_ (.A(_05425_),
    .B(_11691_),
    .C(_11692_),
    .Y(_11693_));
 INVx2_ASAP7_75t_R _32708_ (.A(_11693_),
    .Y(_11694_));
 AND2x2_ASAP7_75t_R _32709_ (.A(_01740_),
    .B(_05425_),
    .Y(_11695_));
 AO21x1_ASAP7_75t_R _32710_ (.A1(_11689_),
    .A2(_11694_),
    .B(_11695_),
    .Y(_11696_));
 INVx1_ASAP7_75t_R _32711_ (.A(_11648_),
    .Y(_11697_));
 AOI21x1_ASAP7_75t_R _32712_ (.A1(_11625_),
    .A2(_11631_),
    .B(_11632_),
    .Y(_11698_));
 AND4x1_ASAP7_75t_R _32713_ (.A(_11698_),
    .B(_11653_),
    .C(_11664_),
    .D(_11678_),
    .Y(_11699_));
 AND2x2_ASAP7_75t_R _32714_ (.A(_11697_),
    .B(_11699_),
    .Y(_11700_));
 XNOR2x1_ASAP7_75t_R _32715_ (.B(_11700_),
    .Y(_11701_),
    .A(_11696_));
 NOR2x1_ASAP7_75t_R _32716_ (.A(_01740_),
    .B(_11668_),
    .Y(_11702_));
 AO21x1_ASAP7_75t_R _32717_ (.A1(_11624_),
    .A2(_11701_),
    .B(_11702_),
    .Y(_03925_));
 BUFx4f_ASAP7_75t_R _32718_ (.A(_05467_),
    .Y(_11703_));
 BUFx6f_ASAP7_75t_R _32719_ (.A(_11703_),
    .Y(_11704_));
 AO21x1_ASAP7_75t_R _32720_ (.A1(_01741_),
    .A2(_05465_),
    .B(_11677_),
    .Y(_11705_));
 OR4x2_ASAP7_75t_R _32721_ (.A(_11633_),
    .B(_11665_),
    .C(_11705_),
    .D(_11696_),
    .Y(_11706_));
 OR3x1_ASAP7_75t_R _32722_ (.A(_05513_),
    .B(_11685_),
    .C(_11706_),
    .Y(_11707_));
 XOR2x1_ASAP7_75t_R _32723_ (.A(_01739_),
    .Y(_11708_),
    .B(_11707_));
 BUFx6f_ASAP7_75t_R _32724_ (.A(_05390_),
    .Y(_11709_));
 OR2x2_ASAP7_75t_R _32725_ (.A(_11685_),
    .B(_11706_),
    .Y(_11710_));
 OA222x2_ASAP7_75t_R _32726_ (.A1(_01974_),
    .A2(_05411_),
    .B1(_05415_),
    .B2(_02071_),
    .C1(_11628_),
    .C2(_01468_),
    .Y(_11711_));
 INVx1_ASAP7_75t_R _32727_ (.A(_11711_),
    .Y(_11712_));
 AO221x2_ASAP7_75t_R _32728_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_11035_),
    .B1(_11679_),
    .B2(net26),
    .C(_11712_),
    .Y(_11713_));
 XNOR2x1_ASAP7_75t_R _32729_ (.B(_11713_),
    .Y(_11714_),
    .A(_11710_));
 AND2x2_ASAP7_75t_R _32730_ (.A(_11709_),
    .B(_11714_),
    .Y(_11715_));
 AO21x1_ASAP7_75t_R _32731_ (.A1(_11704_),
    .A2(_11708_),
    .B(_11715_),
    .Y(_03926_));
 OA222x2_ASAP7_75t_R _32732_ (.A1(_01973_),
    .A2(_05411_),
    .B1(_05416_),
    .B2(_02070_),
    .C1(_11628_),
    .C2(_01469_),
    .Y(_11716_));
 NAND2x1_ASAP7_75t_R _32733_ (.A(net27),
    .B(_11679_),
    .Y(_11717_));
 AND3x1_ASAP7_75t_R _32734_ (.A(_05386_),
    .B(_11716_),
    .C(_11717_),
    .Y(_11718_));
 OA21x2_ASAP7_75t_R _32735_ (.A1(_16028_),
    .A2(_05423_),
    .B(_11718_),
    .Y(_11719_));
 AND2x2_ASAP7_75t_R _32736_ (.A(_01738_),
    .B(_05465_),
    .Y(_11720_));
 NOR2x2_ASAP7_75t_R _32737_ (.A(_11719_),
    .B(_11720_),
    .Y(_11721_));
 NAND2x1_ASAP7_75t_R _32738_ (.A(_01739_),
    .B(_05465_),
    .Y(_11722_));
 OAI21x1_ASAP7_75t_R _32739_ (.A1(_05466_),
    .A2(_11713_),
    .B(_11722_),
    .Y(_11723_));
 OR3x1_ASAP7_75t_R _32740_ (.A(_11648_),
    .B(_11706_),
    .C(_11723_),
    .Y(_11724_));
 XNOR2x1_ASAP7_75t_R _32741_ (.B(_11724_),
    .Y(_11725_),
    .A(_11721_));
 NOR2x1_ASAP7_75t_R _32742_ (.A(_01738_),
    .B(_11668_),
    .Y(_11726_));
 AO21x1_ASAP7_75t_R _32743_ (.A1(_11624_),
    .A2(_11725_),
    .B(_11726_),
    .Y(_03927_));
 OR3x2_ASAP7_75t_R _32744_ (.A(_11719_),
    .B(_11720_),
    .C(_11723_),
    .Y(_11727_));
 NOR2x2_ASAP7_75t_R _32745_ (.A(_11710_),
    .B(_11727_),
    .Y(_11728_));
 AND2x2_ASAP7_75t_R _32746_ (.A(_18773_),
    .B(_11728_),
    .Y(_11729_));
 XNOR2x1_ASAP7_75t_R _32747_ (.B(_11729_),
    .Y(_11730_),
    .A(_01737_));
 BUFx4f_ASAP7_75t_R _32748_ (.A(_05389_),
    .Y(_11731_));
 OA222x2_ASAP7_75t_R _32749_ (.A1(_01972_),
    .A2(_05411_),
    .B1(_05415_),
    .B2(_02069_),
    .C1(_11628_),
    .C2(_01470_),
    .Y(_11732_));
 INVx1_ASAP7_75t_R _32750_ (.A(_11732_),
    .Y(_11733_));
 AO221x2_ASAP7_75t_R _32751_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_11035_),
    .B1(_11679_),
    .B2(net28),
    .C(_11733_),
    .Y(_11734_));
 XOR2x1_ASAP7_75t_R _32752_ (.A(_11728_),
    .Y(_11735_),
    .B(_11734_));
 AND2x2_ASAP7_75t_R _32753_ (.A(_11731_),
    .B(_11735_),
    .Y(_11736_));
 AO21x1_ASAP7_75t_R _32754_ (.A1(_11704_),
    .A2(_11730_),
    .B(_11736_),
    .Y(_03928_));
 AND2x2_ASAP7_75t_R _32755_ (.A(net29),
    .B(_05432_),
    .Y(_11737_));
 AND2x2_ASAP7_75t_R _32756_ (.A(_01471_),
    .B(_11674_),
    .Y(_11738_));
 OA222x2_ASAP7_75t_R _32757_ (.A1(_01971_),
    .A2(_05411_),
    .B1(_11673_),
    .B2(_11738_),
    .C1(_05415_),
    .C2(_02068_),
    .Y(_11739_));
 INVx1_ASAP7_75t_R _32758_ (.A(_11739_),
    .Y(_11740_));
 OR3x2_ASAP7_75t_R _32759_ (.A(_05465_),
    .B(_11737_),
    .C(_11740_),
    .Y(_11741_));
 OA31x2_ASAP7_75t_R _32760_ (.A1(_16279_),
    .A2(_16284_),
    .A3(_16289_),
    .B1(_11035_),
    .Y(_11742_));
 NAND2x1_ASAP7_75t_R _32761_ (.A(_01736_),
    .B(_05465_),
    .Y(_11743_));
 OA21x2_ASAP7_75t_R _32762_ (.A1(_11741_),
    .A2(_11742_),
    .B(_11743_),
    .Y(_11744_));
 AOI21x1_ASAP7_75t_R _32763_ (.A1(_11689_),
    .A2(_11694_),
    .B(_11695_),
    .Y(_11745_));
 OA21x2_ASAP7_75t_R _32764_ (.A1(_05466_),
    .A2(_11713_),
    .B(_11722_),
    .Y(_11746_));
 AND4x1_ASAP7_75t_R _32765_ (.A(_11745_),
    .B(_11699_),
    .C(_11721_),
    .D(_11746_),
    .Y(_11747_));
 NAND2x1_ASAP7_75t_R _32766_ (.A(_01737_),
    .B(_05465_),
    .Y(_11748_));
 OA21x2_ASAP7_75t_R _32767_ (.A1(_05465_),
    .A2(_11734_),
    .B(_11748_),
    .Y(_11749_));
 AND3x1_ASAP7_75t_R _32768_ (.A(_11697_),
    .B(_11747_),
    .C(_11749_),
    .Y(_11750_));
 XOR2x1_ASAP7_75t_R _32769_ (.A(_11744_),
    .Y(_11751_),
    .B(_11750_));
 NOR2x1_ASAP7_75t_R _32770_ (.A(_01736_),
    .B(_11668_),
    .Y(_11752_));
 AO21x1_ASAP7_75t_R _32771_ (.A1(_11624_),
    .A2(_11751_),
    .B(_11752_),
    .Y(_03929_));
 BUFx4f_ASAP7_75t_R _32772_ (.A(_11628_),
    .Y(_11753_));
 OA222x2_ASAP7_75t_R _32773_ (.A1(_01970_),
    .A2(_05412_),
    .B1(_05416_),
    .B2(_02067_),
    .C1(_11753_),
    .C2(_01472_),
    .Y(_11754_));
 AOI22x1_ASAP7_75t_R _32774_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_11035_),
    .B1(_11679_),
    .B2(net30),
    .Y(_11755_));
 AOI21x1_ASAP7_75t_R _32775_ (.A1(_11754_),
    .A2(_11755_),
    .B(_05465_),
    .Y(_11756_));
 INVx1_ASAP7_75t_R _32776_ (.A(_11756_),
    .Y(_11757_));
 OA21x2_ASAP7_75t_R _32777_ (.A1(_01735_),
    .A2(_05386_),
    .B(_11757_),
    .Y(_11758_));
 AND3x1_ASAP7_75t_R _32778_ (.A(_11728_),
    .B(_11744_),
    .C(_11749_),
    .Y(_11759_));
 XNOR2x1_ASAP7_75t_R _32779_ (.B(_11759_),
    .Y(_11760_),
    .A(_11758_));
 NOR2x1_ASAP7_75t_R _32780_ (.A(_01735_),
    .B(_11668_),
    .Y(_11761_));
 AO21x1_ASAP7_75t_R _32781_ (.A1(_11624_),
    .A2(_11760_),
    .B(_11761_),
    .Y(_03930_));
 OA222x2_ASAP7_75t_R _32782_ (.A1(_01969_),
    .A2(_05411_),
    .B1(_05416_),
    .B2(_02066_),
    .C1(_11628_),
    .C2(_01473_),
    .Y(_11762_));
 NAND2x1_ASAP7_75t_R _32783_ (.A(net31),
    .B(_11679_),
    .Y(_11763_));
 AND3x1_ASAP7_75t_R _32784_ (.A(_05386_),
    .B(_11762_),
    .C(_11763_),
    .Y(_11764_));
 OA21x2_ASAP7_75t_R _32785_ (.A1(_16531_),
    .A2(_05423_),
    .B(_11764_),
    .Y(_11765_));
 AO21x2_ASAP7_75t_R _32786_ (.A1(_01734_),
    .A2(_05466_),
    .B(_11765_),
    .Y(_11766_));
 NAND2x1_ASAP7_75t_R _32787_ (.A(_11744_),
    .B(_11749_),
    .Y(_11767_));
 NOR2x1_ASAP7_75t_R _32788_ (.A(_11758_),
    .B(_11767_),
    .Y(_11768_));
 AND3x1_ASAP7_75t_R _32789_ (.A(_11697_),
    .B(_11747_),
    .C(_11768_),
    .Y(_11769_));
 XNOR2x1_ASAP7_75t_R _32790_ (.B(_11769_),
    .Y(_11770_),
    .A(_11766_));
 NOR2x1_ASAP7_75t_R _32791_ (.A(_01734_),
    .B(_11668_),
    .Y(_11771_));
 AO21x1_ASAP7_75t_R _32792_ (.A1(_11624_),
    .A2(_11770_),
    .B(_11771_),
    .Y(_03931_));
 INVx1_ASAP7_75t_R _32793_ (.A(_01733_),
    .Y(_11772_));
 BUFx4f_ASAP7_75t_R _32794_ (.A(_05513_),
    .Y(_11773_));
 AND2x2_ASAP7_75t_R _32795_ (.A(_05467_),
    .B(_11773_),
    .Y(_11774_));
 OA222x2_ASAP7_75t_R _32796_ (.A1(_01968_),
    .A2(_05412_),
    .B1(_05417_),
    .B2(_02065_),
    .C1(_11753_),
    .C2(_01474_),
    .Y(_11775_));
 INVx1_ASAP7_75t_R _32797_ (.A(_11775_),
    .Y(_11776_));
 AO221x1_ASAP7_75t_R _32798_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_11036_),
    .B1(_11680_),
    .B2(net32),
    .C(_11776_),
    .Y(_11777_));
 NAND2x2_ASAP7_75t_R _32799_ (.A(_05387_),
    .B(_11777_),
    .Y(_11778_));
 OA21x2_ASAP7_75t_R _32800_ (.A1(_01733_),
    .A2(_05388_),
    .B(_11778_),
    .Y(_11779_));
 OR5x2_ASAP7_75t_R _32801_ (.A(_11706_),
    .B(_11727_),
    .C(_11758_),
    .D(_11767_),
    .E(_11766_),
    .Y(_11780_));
 OR3x4_ASAP7_75t_R _32802_ (.A(_11685_),
    .B(_11779_),
    .C(_11780_),
    .Y(_11781_));
 OAI21x1_ASAP7_75t_R _32803_ (.A1(_11685_),
    .A2(_11780_),
    .B(_11779_),
    .Y(_11782_));
 AND3x1_ASAP7_75t_R _32804_ (.A(_11623_),
    .B(_11781_),
    .C(_11782_),
    .Y(_11783_));
 AO21x1_ASAP7_75t_R _32805_ (.A1(_11772_),
    .A2(_11774_),
    .B(_11783_),
    .Y(_03932_));
 BUFx4f_ASAP7_75t_R _32806_ (.A(_11623_),
    .Y(_11784_));
 OR3x4_ASAP7_75t_R _32807_ (.A(_11648_),
    .B(_11779_),
    .C(_11780_),
    .Y(_11785_));
 INVx1_ASAP7_75t_R _32808_ (.A(_01732_),
    .Y(_11786_));
 NAND2x1_ASAP7_75t_R _32809_ (.A(net33),
    .B(_11679_),
    .Y(_11787_));
 AND2x2_ASAP7_75t_R _32810_ (.A(_01475_),
    .B(_11674_),
    .Y(_11788_));
 OA222x2_ASAP7_75t_R _32811_ (.A1(_01966_),
    .A2(_05412_),
    .B1(_11673_),
    .B2(_11788_),
    .C1(_05416_),
    .C2(_02064_),
    .Y(_11789_));
 AND3x2_ASAP7_75t_R _32812_ (.A(_05386_),
    .B(_11787_),
    .C(_11789_),
    .Y(_11790_));
 OAI21x1_ASAP7_75t_R _32813_ (.A1(_16777_),
    .A2(_05423_),
    .B(_11790_),
    .Y(_11791_));
 OA21x2_ASAP7_75t_R _32814_ (.A1(_11786_),
    .A2(_05389_),
    .B(_11791_),
    .Y(_11792_));
 XNOR2x1_ASAP7_75t_R _32815_ (.B(_11792_),
    .Y(_11793_),
    .A(_11785_));
 BUFx6f_ASAP7_75t_R _32816_ (.A(_05467_),
    .Y(_11794_));
 AND3x1_ASAP7_75t_R _32817_ (.A(_11786_),
    .B(_11794_),
    .C(_11773_),
    .Y(_11795_));
 AO21x1_ASAP7_75t_R _32818_ (.A1(_11784_),
    .A2(_11793_),
    .B(_11795_),
    .Y(_03933_));
 AND2x2_ASAP7_75t_R _32819_ (.A(_01731_),
    .B(_05467_),
    .Y(_11796_));
 INVx1_ASAP7_75t_R _32820_ (.A(_11792_),
    .Y(_11797_));
 OR3x1_ASAP7_75t_R _32821_ (.A(_11773_),
    .B(_11781_),
    .C(_11797_),
    .Y(_11798_));
 NOR2x1_ASAP7_75t_R _32822_ (.A(_11781_),
    .B(_11797_),
    .Y(_11799_));
 NAND2x2_ASAP7_75t_R _32823_ (.A(\alu_adder_result_ex[21] ),
    .B(_11035_),
    .Y(_11800_));
 OA222x2_ASAP7_75t_R _32824_ (.A1(_01965_),
    .A2(_05412_),
    .B1(_05416_),
    .B2(_02063_),
    .C1(_11753_),
    .C2(_01476_),
    .Y(_11801_));
 NAND2x1_ASAP7_75t_R _32825_ (.A(net34),
    .B(_11679_),
    .Y(_11802_));
 AND4x2_ASAP7_75t_R _32826_ (.A(_05386_),
    .B(_11800_),
    .C(_11801_),
    .D(_11802_),
    .Y(_11803_));
 OAI21x1_ASAP7_75t_R _32827_ (.A1(_11796_),
    .A2(_11803_),
    .B(_11799_),
    .Y(_11804_));
 OA211x2_ASAP7_75t_R _32828_ (.A1(_11799_),
    .A2(_11803_),
    .B(_11804_),
    .C(_11623_),
    .Y(_11805_));
 AOI21x1_ASAP7_75t_R _32829_ (.A1(_11796_),
    .A2(_11798_),
    .B(_11805_),
    .Y(_03934_));
 INVx1_ASAP7_75t_R _32830_ (.A(_01730_),
    .Y(_11806_));
 OA222x2_ASAP7_75t_R _32831_ (.A1(_01964_),
    .A2(_05413_),
    .B1(_05417_),
    .B2(_02062_),
    .C1(_11753_),
    .C2(_01477_),
    .Y(_11807_));
 NAND2x1_ASAP7_75t_R _32832_ (.A(net35),
    .B(_11679_),
    .Y(_11808_));
 AND3x1_ASAP7_75t_R _32833_ (.A(_05386_),
    .B(_11807_),
    .C(_11808_),
    .Y(_11809_));
 OAI21x1_ASAP7_75t_R _32834_ (.A1(_17017_),
    .A2(_05423_),
    .B(_11809_),
    .Y(_11810_));
 OA21x2_ASAP7_75t_R _32835_ (.A1(_11806_),
    .A2(_05388_),
    .B(_11810_),
    .Y(_11811_));
 NOR3x2_ASAP7_75t_R _32836_ (.B(_11779_),
    .C(_11780_),
    .Y(_11812_),
    .A(_11648_));
 AOI21x1_ASAP7_75t_R _32837_ (.A1(_01731_),
    .A2(_05466_),
    .B(_11803_),
    .Y(_11813_));
 OA211x2_ASAP7_75t_R _32838_ (.A1(_11786_),
    .A2(_05387_),
    .B(_11791_),
    .C(_11813_),
    .Y(_11814_));
 AND2x2_ASAP7_75t_R _32839_ (.A(_11812_),
    .B(_11814_),
    .Y(_11815_));
 XOR2x1_ASAP7_75t_R _32840_ (.A(_11811_),
    .Y(_11816_),
    .B(_11815_));
 AND3x1_ASAP7_75t_R _32841_ (.A(_11806_),
    .B(_11794_),
    .C(_11773_),
    .Y(_11817_));
 AO21x1_ASAP7_75t_R _32842_ (.A1(_11784_),
    .A2(_11816_),
    .B(_11817_),
    .Y(_03935_));
 OA222x2_ASAP7_75t_R _32843_ (.A1(_01963_),
    .A2(_05412_),
    .B1(_05417_),
    .B2(_02061_),
    .C1(_11753_),
    .C2(_01478_),
    .Y(_11818_));
 INVx1_ASAP7_75t_R _32844_ (.A(_11818_),
    .Y(_11819_));
 AO221x2_ASAP7_75t_R _32845_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_11035_),
    .B1(_11679_),
    .B2(net36),
    .C(_11819_),
    .Y(_11820_));
 NAND2x2_ASAP7_75t_R _32846_ (.A(_05387_),
    .B(_11820_),
    .Y(_11821_));
 OAI21x1_ASAP7_75t_R _32847_ (.A1(_01729_),
    .A2(_05388_),
    .B(_11821_),
    .Y(_11822_));
 INVx1_ASAP7_75t_R _32848_ (.A(_11781_),
    .Y(_11823_));
 AND3x1_ASAP7_75t_R _32849_ (.A(_11823_),
    .B(_11811_),
    .C(_11814_),
    .Y(_11824_));
 XOR2x1_ASAP7_75t_R _32850_ (.A(_11822_),
    .Y(_11825_),
    .B(_11824_));
 NOR2x1_ASAP7_75t_R _32851_ (.A(_01729_),
    .B(_11668_),
    .Y(_11826_));
 AO21x1_ASAP7_75t_R _32852_ (.A1(_11784_),
    .A2(_11825_),
    .B(_11826_),
    .Y(_03936_));
 NAND2x1_ASAP7_75t_R _32853_ (.A(_01728_),
    .B(_05466_),
    .Y(_11827_));
 OA222x2_ASAP7_75t_R _32854_ (.A1(_01962_),
    .A2(_05413_),
    .B1(_05417_),
    .B2(_02060_),
    .C1(_11753_),
    .C2(_01479_),
    .Y(_11828_));
 NAND2x1_ASAP7_75t_R _32855_ (.A(net37),
    .B(_11680_),
    .Y(_11829_));
 AND3x1_ASAP7_75t_R _32856_ (.A(_05387_),
    .B(_11828_),
    .C(_11829_),
    .Y(_11830_));
 OAI21x1_ASAP7_75t_R _32857_ (.A1(_17257_),
    .A2(_05423_),
    .B(_11830_),
    .Y(_11831_));
 AND3x2_ASAP7_75t_R _32858_ (.A(_11811_),
    .B(_11814_),
    .C(_11822_),
    .Y(_11832_));
 NAND2x2_ASAP7_75t_R _32859_ (.A(_11812_),
    .B(_11832_),
    .Y(_11833_));
 AO21x1_ASAP7_75t_R _32860_ (.A1(_11827_),
    .A2(_11831_),
    .B(_11833_),
    .Y(_11834_));
 AOI21x1_ASAP7_75t_R _32861_ (.A1(_11833_),
    .A2(_11831_),
    .B(_11774_),
    .Y(_11835_));
 OA211x2_ASAP7_75t_R _32862_ (.A1(_11773_),
    .A2(_11833_),
    .B(_01728_),
    .C(_11703_),
    .Y(_11836_));
 AOI21x1_ASAP7_75t_R _32863_ (.A1(_11834_),
    .A2(_11835_),
    .B(_11836_),
    .Y(_03937_));
 INVx1_ASAP7_75t_R _32864_ (.A(_01727_),
    .Y(_11837_));
 AND2x2_ASAP7_75t_R _32865_ (.A(_01480_),
    .B(_11674_),
    .Y(_11838_));
 OA222x2_ASAP7_75t_R _32866_ (.A1(_01961_),
    .A2(_05412_),
    .B1(_11673_),
    .B2(_11838_),
    .C1(_05417_),
    .C2(_02059_),
    .Y(_11839_));
 INVx1_ASAP7_75t_R _32867_ (.A(_11839_),
    .Y(_11840_));
 AO221x1_ASAP7_75t_R _32868_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_11036_),
    .B1(_11680_),
    .B2(net38),
    .C(_11840_),
    .Y(_11841_));
 AND2x2_ASAP7_75t_R _32869_ (.A(_05388_),
    .B(_11841_),
    .Y(_11842_));
 AOI21x1_ASAP7_75t_R _32870_ (.A1(_11837_),
    .A2(_05466_),
    .B(_11842_),
    .Y(_11843_));
 AND2x2_ASAP7_75t_R _32871_ (.A(_11827_),
    .B(_11831_),
    .Y(_11844_));
 AND2x2_ASAP7_75t_R _32872_ (.A(_11832_),
    .B(_11844_),
    .Y(_11845_));
 AND2x2_ASAP7_75t_R _32873_ (.A(_11823_),
    .B(_11845_),
    .Y(_11846_));
 XNOR2x1_ASAP7_75t_R _32874_ (.B(_11846_),
    .Y(_11847_),
    .A(_11843_));
 AND3x1_ASAP7_75t_R _32875_ (.A(_11837_),
    .B(_11703_),
    .C(_11773_),
    .Y(_11848_));
 AO21x1_ASAP7_75t_R _32876_ (.A1(_11784_),
    .A2(_11847_),
    .B(_11848_),
    .Y(_03938_));
 OA222x2_ASAP7_75t_R _32877_ (.A1(_01960_),
    .A2(_05413_),
    .B1(_05417_),
    .B2(_02058_),
    .C1(_11753_),
    .C2(_01481_),
    .Y(_11849_));
 NAND2x1_ASAP7_75t_R _32878_ (.A(net39),
    .B(_11680_),
    .Y(_11850_));
 OA211x2_ASAP7_75t_R _32879_ (.A1(_04414_),
    .A2(_05423_),
    .B(_11849_),
    .C(_11850_),
    .Y(_11851_));
 OR2x2_ASAP7_75t_R _32880_ (.A(_01726_),
    .B(_05387_),
    .Y(_11852_));
 OA21x2_ASAP7_75t_R _32881_ (.A1(_05466_),
    .A2(_11851_),
    .B(_11852_),
    .Y(_11853_));
 AO21x1_ASAP7_75t_R _32882_ (.A1(_11837_),
    .A2(_05466_),
    .B(_11842_),
    .Y(_11854_));
 AND3x1_ASAP7_75t_R _32883_ (.A(_11812_),
    .B(_11854_),
    .C(_11845_),
    .Y(_11855_));
 XNOR2x1_ASAP7_75t_R _32884_ (.B(_11855_),
    .Y(_11856_),
    .A(_11853_));
 NOR2x1_ASAP7_75t_R _32885_ (.A(_01726_),
    .B(_11668_),
    .Y(_11857_));
 AO21x1_ASAP7_75t_R _32886_ (.A1(_11784_),
    .A2(_11856_),
    .B(_11857_),
    .Y(_03939_));
 NAND3x1_ASAP7_75t_R _32887_ (.A(_11811_),
    .B(_11814_),
    .C(_11822_),
    .Y(_11858_));
 NAND2x1_ASAP7_75t_R _32888_ (.A(_11827_),
    .B(_11831_),
    .Y(_11859_));
 OR4x1_ASAP7_75t_R _32889_ (.A(_11858_),
    .B(_11843_),
    .C(_11859_),
    .D(_11853_),
    .Y(_11860_));
 AND2x2_ASAP7_75t_R _32890_ (.A(_00007_),
    .B(_11674_),
    .Y(_11861_));
 OA222x2_ASAP7_75t_R _32891_ (.A1(_01959_),
    .A2(_05412_),
    .B1(_11673_),
    .B2(_11861_),
    .C1(_05417_),
    .C2(_02057_),
    .Y(_11862_));
 INVx1_ASAP7_75t_R _32892_ (.A(_11862_),
    .Y(_11863_));
 AO221x2_ASAP7_75t_R _32893_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_11036_),
    .B1(_11680_),
    .B2(net40),
    .C(_11863_),
    .Y(_11864_));
 NAND2x2_ASAP7_75t_R _32894_ (.A(_05387_),
    .B(_11864_),
    .Y(_11865_));
 OA21x2_ASAP7_75t_R _32895_ (.A1(_11781_),
    .A2(_11860_),
    .B(_11865_),
    .Y(_11866_));
 OA21x2_ASAP7_75t_R _32896_ (.A1(_01725_),
    .A2(_05388_),
    .B(_11865_),
    .Y(_11867_));
 OR5x2_ASAP7_75t_R _32897_ (.A(_11858_),
    .B(_11843_),
    .C(_11859_),
    .D(_11853_),
    .E(_11867_),
    .Y(_11868_));
 NOR2x1_ASAP7_75t_R _32898_ (.A(_11781_),
    .B(_11868_),
    .Y(_11869_));
 AO21x1_ASAP7_75t_R _32899_ (.A1(_11709_),
    .A2(_11866_),
    .B(_11869_),
    .Y(_11870_));
 OA21x2_ASAP7_75t_R _32900_ (.A1(_11774_),
    .A2(_11866_),
    .B(_01725_),
    .Y(_11871_));
 AOI21x1_ASAP7_75t_R _32901_ (.A1(_11624_),
    .A2(_11870_),
    .B(_11871_),
    .Y(_03940_));
 AND2x2_ASAP7_75t_R _32902_ (.A(_00008_),
    .B(_11674_),
    .Y(_11872_));
 OA222x2_ASAP7_75t_R _32903_ (.A1(_01958_),
    .A2(_05413_),
    .B1(_11673_),
    .B2(_11872_),
    .C1(_05417_),
    .C2(_02056_),
    .Y(_11873_));
 INVx1_ASAP7_75t_R _32904_ (.A(_11873_),
    .Y(_11874_));
 AO221x2_ASAP7_75t_R _32905_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_11036_),
    .B1(_11680_),
    .B2(net41),
    .C(_11874_),
    .Y(_11875_));
 NOR2x1_ASAP7_75t_R _32906_ (.A(_01724_),
    .B(_05388_),
    .Y(_11876_));
 AOI21x1_ASAP7_75t_R _32907_ (.A1(_05388_),
    .A2(_11875_),
    .B(_11876_),
    .Y(_11877_));
 OR2x2_ASAP7_75t_R _32908_ (.A(_11785_),
    .B(_11868_),
    .Y(_11878_));
 XOR2x1_ASAP7_75t_R _32909_ (.A(_11877_),
    .Y(_11879_),
    .B(_11878_));
 NOR2x1_ASAP7_75t_R _32910_ (.A(_01724_),
    .B(_11623_),
    .Y(_11880_));
 AO21x1_ASAP7_75t_R _32911_ (.A1(_11784_),
    .A2(_11879_),
    .B(_11880_),
    .Y(_03941_));
 OA222x2_ASAP7_75t_R _32912_ (.A1(_01957_),
    .A2(_05413_),
    .B1(_05417_),
    .B2(_02055_),
    .C1(_11753_),
    .C2(_00009_),
    .Y(_11881_));
 INVx1_ASAP7_75t_R _32913_ (.A(_11881_),
    .Y(_11882_));
 AO221x2_ASAP7_75t_R _32914_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_11036_),
    .B1(_11680_),
    .B2(net42),
    .C(_11882_),
    .Y(_11883_));
 NAND2x2_ASAP7_75t_R _32915_ (.A(_05388_),
    .B(_11883_),
    .Y(_11884_));
 OA21x2_ASAP7_75t_R _32916_ (.A1(_01723_),
    .A2(_05389_),
    .B(_11884_),
    .Y(_11885_));
 OR3x2_ASAP7_75t_R _32917_ (.A(_11781_),
    .B(_11868_),
    .C(_11877_),
    .Y(_11886_));
 XOR2x1_ASAP7_75t_R _32918_ (.A(_11885_),
    .Y(_11887_),
    .B(_11886_));
 NOR2x1_ASAP7_75t_R _32919_ (.A(_01723_),
    .B(_11623_),
    .Y(_11888_));
 AO21x1_ASAP7_75t_R _32920_ (.A1(_11784_),
    .A2(_11887_),
    .B(_11888_),
    .Y(_03942_));
 BUFx6f_ASAP7_75t_R _32921_ (.A(_05467_),
    .Y(_11889_));
 AND3x1_ASAP7_75t_R _32922_ (.A(_01722_),
    .B(_11889_),
    .C(_11773_),
    .Y(_11890_));
 AOI21x1_ASAP7_75t_R _32923_ (.A1(_02291_),
    .A2(_11624_),
    .B(_11890_),
    .Y(_03943_));
 INVx1_ASAP7_75t_R _32924_ (.A(_01721_),
    .Y(_11891_));
 OA222x2_ASAP7_75t_R _32925_ (.A1(_01955_),
    .A2(_05413_),
    .B1(_05418_),
    .B2(_02053_),
    .C1(_11753_),
    .C2(_00010_),
    .Y(_11892_));
 INVx1_ASAP7_75t_R _32926_ (.A(_11892_),
    .Y(_11893_));
 AO221x1_ASAP7_75t_R _32927_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_11036_),
    .B1(_11680_),
    .B2(net43),
    .C(_11893_),
    .Y(_11894_));
 AND2x2_ASAP7_75t_R _32928_ (.A(_05389_),
    .B(_11894_),
    .Y(_11895_));
 AOI21x1_ASAP7_75t_R _32929_ (.A1(_11891_),
    .A2(_05467_),
    .B(_11895_),
    .Y(_11896_));
 OR4x1_ASAP7_75t_R _32930_ (.A(_11785_),
    .B(_11868_),
    .C(_11877_),
    .D(_11885_),
    .Y(_11897_));
 XOR2x1_ASAP7_75t_R _32931_ (.A(_11896_),
    .Y(_11898_),
    .B(_11897_));
 AND3x1_ASAP7_75t_R _32932_ (.A(_11891_),
    .B(_11703_),
    .C(_11773_),
    .Y(_11899_));
 AO21x1_ASAP7_75t_R _32933_ (.A1(_11784_),
    .A2(_11898_),
    .B(_11899_),
    .Y(_03944_));
 OA222x2_ASAP7_75t_R _32934_ (.A1(_01954_),
    .A2(_05413_),
    .B1(_05418_),
    .B2(_02052_),
    .C1(_11753_),
    .C2(_00011_),
    .Y(_11900_));
 INVx1_ASAP7_75t_R _32935_ (.A(_11900_),
    .Y(_11901_));
 AO221x2_ASAP7_75t_R _32936_ (.A1(_11036_),
    .A2(\alu_adder_result_ex[31] ),
    .B1(_11680_),
    .B2(net44),
    .C(_11901_),
    .Y(_11902_));
 NAND2x2_ASAP7_75t_R _32937_ (.A(_11902_),
    .B(_05389_),
    .Y(_11903_));
 OA21x2_ASAP7_75t_R _32938_ (.A1(_01720_),
    .A2(_05389_),
    .B(_11903_),
    .Y(_11904_));
 OR3x1_ASAP7_75t_R _32939_ (.A(_11885_),
    .B(_11886_),
    .C(_11896_),
    .Y(_11905_));
 XOR2x1_ASAP7_75t_R _32940_ (.A(_11904_),
    .Y(_11906_),
    .B(_11905_));
 NAND2x1_ASAP7_75t_R _32941_ (.A(_01720_),
    .B(_11774_),
    .Y(_11907_));
 OA21x2_ASAP7_75t_R _32942_ (.A1(_11774_),
    .A2(_11906_),
    .B(_11907_),
    .Y(_03945_));
 AND3x1_ASAP7_75t_R _32943_ (.A(_01719_),
    .B(_11889_),
    .C(_11773_),
    .Y(_11908_));
 AOI21x1_ASAP7_75t_R _32944_ (.A1(_02293_),
    .A2(_11624_),
    .B(_11908_),
    .Y(_03946_));
 INVx1_ASAP7_75t_R _32945_ (.A(_11640_),
    .Y(_11909_));
 NOR2x1_ASAP7_75t_R _32946_ (.A(_01718_),
    .B(_05389_),
    .Y(_11910_));
 OR3x1_ASAP7_75t_R _32947_ (.A(_05507_),
    .B(_02292_),
    .C(_05512_),
    .Y(_11911_));
 INVx1_ASAP7_75t_R _32948_ (.A(_02292_),
    .Y(_11912_));
 AO21x1_ASAP7_75t_R _32949_ (.A1(_01718_),
    .A2(_18773_),
    .B(_05390_),
    .Y(_11913_));
 AND3x1_ASAP7_75t_R _32950_ (.A(_11912_),
    .B(_11640_),
    .C(_11913_),
    .Y(_11914_));
 AO221x1_ASAP7_75t_R _32951_ (.A1(_02292_),
    .A2(_11909_),
    .B1(_11910_),
    .B2(_11911_),
    .C(_11914_),
    .Y(_03947_));
 INVx1_ASAP7_75t_R _32952_ (.A(_01717_),
    .Y(_11915_));
 OA211x2_ASAP7_75t_R _32953_ (.A1(_11909_),
    .A2(_11910_),
    .B(_18775_),
    .C(_18776_),
    .Y(_11916_));
 AND3x1_ASAP7_75t_R _32954_ (.A(_11915_),
    .B(_18773_),
    .C(_11916_),
    .Y(_11917_));
 AO21x1_ASAP7_75t_R _32955_ (.A1(_01717_),
    .A2(_11773_),
    .B(_11917_),
    .Y(_11918_));
 XOR2x1_ASAP7_75t_R _32956_ (.A(_11645_),
    .Y(_11919_),
    .B(_11916_));
 OA21x2_ASAP7_75t_R _32957_ (.A1(_01717_),
    .A2(_11709_),
    .B(_11919_),
    .Y(_11920_));
 AOI21x1_ASAP7_75t_R _32958_ (.A1(_11704_),
    .A2(_11918_),
    .B(_11920_),
    .Y(_03948_));
 OR3x1_ASAP7_75t_R _32959_ (.A(_02292_),
    .B(_11641_),
    .C(_11646_),
    .Y(_11921_));
 XOR2x1_ASAP7_75t_R _32960_ (.A(_11637_),
    .Y(_11922_),
    .B(_11921_));
 NOR2x1_ASAP7_75t_R _32961_ (.A(_01716_),
    .B(_11623_),
    .Y(_11923_));
 AO21x1_ASAP7_75t_R _32962_ (.A1(_11784_),
    .A2(_11922_),
    .B(_11923_),
    .Y(_03949_));
 NAND2x2_ASAP7_75t_R _32963_ (.A(_11660_),
    .B(_11663_),
    .Y(_11924_));
 XOR2x1_ASAP7_75t_R _32964_ (.A(_11924_),
    .Y(_11925_),
    .B(_11685_));
 NOR2x1_ASAP7_75t_R _32965_ (.A(_01715_),
    .B(_11623_),
    .Y(_11926_));
 AO21x1_ASAP7_75t_R _32966_ (.A1(_11784_),
    .A2(_11925_),
    .B(_11926_),
    .Y(_03950_));
 NOR2x2_ASAP7_75t_R _32967_ (.A(_11648_),
    .B(_11924_),
    .Y(_11927_));
 AOI21x1_ASAP7_75t_R _32968_ (.A1(_18773_),
    .A2(_11927_),
    .B(_11659_),
    .Y(_11928_));
 XNOR2x1_ASAP7_75t_R _32969_ (.B(_11927_),
    .Y(_11929_),
    .A(_11653_));
 AND3x1_ASAP7_75t_R _32970_ (.A(_11623_),
    .B(_11659_),
    .C(_11929_),
    .Y(_11930_));
 NOR2x1_ASAP7_75t_R _32971_ (.A(_11928_),
    .B(_11930_),
    .Y(_03951_));
 NAND2x2_ASAP7_75t_R _32972_ (.A(_11654_),
    .B(_11658_),
    .Y(_11931_));
 NAND2x1_ASAP7_75t_R _32973_ (.A(_11653_),
    .B(_11659_),
    .Y(_11932_));
 OR3x1_ASAP7_75t_R _32974_ (.A(_11932_),
    .B(_11924_),
    .C(_11685_),
    .Y(_11933_));
 XOR2x1_ASAP7_75t_R _32975_ (.A(_11931_),
    .Y(_11934_),
    .B(_11933_));
 NOR2x1_ASAP7_75t_R _32976_ (.A(_01713_),
    .B(_11623_),
    .Y(_11935_));
 AO21x1_ASAP7_75t_R _32977_ (.A1(_11668_),
    .A2(_11934_),
    .B(_11935_),
    .Y(_03952_));
 OR3x1_ASAP7_75t_R _32978_ (.A(_11024_),
    .B(_11044_),
    .C(_11052_),
    .Y(_11936_));
 INVx1_ASAP7_75t_R _32979_ (.A(_11936_),
    .Y(_11937_));
 AND2x2_ASAP7_75t_R _32980_ (.A(_05087_),
    .B(_11937_),
    .Y(_11938_));
 NAND2x1_ASAP7_75t_R _32981_ (.A(_04928_),
    .B(_11938_),
    .Y(_11939_));
 AND3x1_ASAP7_75t_R _32982_ (.A(_08332_),
    .B(_04925_),
    .C(_04926_),
    .Y(_11940_));
 OAI21x1_ASAP7_75t_R _32983_ (.A1(_05061_),
    .A2(_11940_),
    .B(_11938_),
    .Y(_11941_));
 OAI21x1_ASAP7_75t_R _32984_ (.A1(_05058_),
    .A2(_11939_),
    .B(_11941_),
    .Y(_11942_));
 AO21x2_ASAP7_75t_R _32985_ (.A1(_11031_),
    .A2(_11073_),
    .B(_04937_),
    .Y(_11943_));
 AO21x1_ASAP7_75t_R _32986_ (.A1(_05477_),
    .A2(_05481_),
    .B(_07310_),
    .Y(_11944_));
 OR2x2_ASAP7_75t_R _32987_ (.A(_05508_),
    .B(_11944_),
    .Y(_11945_));
 INVx2_ASAP7_75t_R _32988_ (.A(_02227_),
    .Y(_11946_));
 AND3x4_ASAP7_75t_R _32989_ (.A(net177),
    .B(_02223_),
    .C(_11946_),
    .Y(_11947_));
 NAND2x1_ASAP7_75t_R _32990_ (.A(_11944_),
    .B(_11947_),
    .Y(_11948_));
 INVx4_ASAP7_75t_R _32991_ (.A(_05508_),
    .Y(_11949_));
 NOR2x1_ASAP7_75t_R _32992_ (.A(_11949_),
    .B(_11947_),
    .Y(_11950_));
 INVx1_ASAP7_75t_R _32993_ (.A(_11944_),
    .Y(_11951_));
 AO32x2_ASAP7_75t_R _32994_ (.A1(_05486_),
    .A2(_11945_),
    .A3(_11948_),
    .B1(_11950_),
    .B2(_11951_),
    .Y(_11952_));
 NOR2x1_ASAP7_75t_R _32995_ (.A(_11049_),
    .B(_11952_),
    .Y(_11953_));
 OA21x2_ASAP7_75t_R _32996_ (.A1(_11942_),
    .A2(_11943_),
    .B(_11953_),
    .Y(_11954_));
 BUFx4f_ASAP7_75t_R _32997_ (.A(_11954_),
    .Y(_11955_));
 NAND2x1_ASAP7_75t_R _32998_ (.A(_06830_),
    .B(_11955_),
    .Y(_11956_));
 BUFx4f_ASAP7_75t_R _32999_ (.A(_11956_),
    .Y(_11957_));
 BUFx4f_ASAP7_75t_R _33000_ (.A(_05486_),
    .Y(_11958_));
 BUFx4f_ASAP7_75t_R _33001_ (.A(_11958_),
    .Y(_11959_));
 INVx1_ASAP7_75t_R _33002_ (.A(_05488_),
    .Y(_11960_));
 OA211x2_ASAP7_75t_R _33003_ (.A1(_05480_),
    .A2(_05491_),
    .B(_11960_),
    .C(_07312_),
    .Y(_11961_));
 BUFx3_ASAP7_75t_R _33004_ (.A(_11961_),
    .Y(_11962_));
 AND2x2_ASAP7_75t_R _33005_ (.A(net177),
    .B(_11946_),
    .Y(_11963_));
 NAND2x1_ASAP7_75t_R _33006_ (.A(_02223_),
    .B(_11963_),
    .Y(_11964_));
 OR3x1_ASAP7_75t_R _33007_ (.A(_11959_),
    .B(_11962_),
    .C(_11964_),
    .Y(_11965_));
 OAI21x1_ASAP7_75t_R _33008_ (.A1(_11942_),
    .A2(_11943_),
    .B(_11953_),
    .Y(_11966_));
 AND2x2_ASAP7_75t_R _33009_ (.A(_11959_),
    .B(_11947_),
    .Y(_11967_));
 OAI21x1_ASAP7_75t_R _33010_ (.A1(_11072_),
    .A2(_11966_),
    .B(_11967_),
    .Y(_11968_));
 OA21x2_ASAP7_75t_R _33011_ (.A1(_11957_),
    .A2(_11965_),
    .B(_11968_),
    .Y(_11969_));
 BUFx3_ASAP7_75t_R _33012_ (.A(_11969_),
    .Y(_11970_));
 OR2x2_ASAP7_75t_R _33013_ (.A(_05508_),
    .B(_11962_),
    .Y(_11971_));
 OR3x4_ASAP7_75t_R _33014_ (.A(_11072_),
    .B(_11966_),
    .C(_11971_),
    .Y(_11972_));
 BUFx3_ASAP7_75t_R _33015_ (.A(_11972_),
    .Y(_11973_));
 AND2x6_ASAP7_75t_R _33016_ (.A(_11962_),
    .B(_11967_),
    .Y(_11974_));
 BUFx6f_ASAP7_75t_R _33017_ (.A(_11974_),
    .Y(_11975_));
 NOR2x1_ASAP7_75t_R _33018_ (.A(_01712_),
    .B(_11975_),
    .Y(_11976_));
 BUFx4f_ASAP7_75t_R _33019_ (.A(_11949_),
    .Y(_11977_));
 BUFx6f_ASAP7_75t_R _33020_ (.A(_11977_),
    .Y(_11978_));
 BUFx6f_ASAP7_75t_R _33021_ (.A(_11978_),
    .Y(_11979_));
 BUFx4f_ASAP7_75t_R _33022_ (.A(_11979_),
    .Y(_11980_));
 BUFx4f_ASAP7_75t_R _33023_ (.A(_11979_),
    .Y(_11981_));
 NAND2x1_ASAP7_75t_R _33024_ (.A(_11981_),
    .B(_01711_),
    .Y(_11982_));
 OA21x2_ASAP7_75t_R _33025_ (.A1(net139),
    .A2(_11980_),
    .B(_11982_),
    .Y(_11983_));
 AND3x1_ASAP7_75t_R _33026_ (.A(_05493_),
    .B(_06830_),
    .C(_11955_),
    .Y(_11984_));
 NAND2x1_ASAP7_75t_R _33027_ (.A(_05508_),
    .B(_11965_),
    .Y(_11985_));
 OA31x2_ASAP7_75t_R _33028_ (.A1(_11962_),
    .A2(_11072_),
    .A3(_11966_),
    .B1(_11967_),
    .Y(_11986_));
 AO21x2_ASAP7_75t_R _33029_ (.A1(_11984_),
    .A2(_11985_),
    .B(_11986_),
    .Y(_11987_));
 BUFx2_ASAP7_75t_R _33030_ (.A(_11987_),
    .Y(_11988_));
 AO32x1_ASAP7_75t_R _33031_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_11976_),
    .B1(_11983_),
    .B2(_11988_),
    .Y(_03953_));
 OA211x2_ASAP7_75t_R _33032_ (.A1(_11942_),
    .A2(_11943_),
    .B(_05493_),
    .C(_11050_),
    .Y(_11989_));
 NAND2x1_ASAP7_75t_R _33033_ (.A(_06831_),
    .B(_11989_),
    .Y(_11990_));
 OR3x1_ASAP7_75t_R _33034_ (.A(_11959_),
    .B(_11979_),
    .C(_11964_),
    .Y(_11991_));
 BUFx6f_ASAP7_75t_R _33035_ (.A(_02226_),
    .Y(_11992_));
 NOR2x1_ASAP7_75t_R _33036_ (.A(_11992_),
    .B(_11952_),
    .Y(_11993_));
 AND2x6_ASAP7_75t_R _33037_ (.A(_11978_),
    .B(_11947_),
    .Y(_11994_));
 NOR2x1_ASAP7_75t_R _33038_ (.A(_11993_),
    .B(_11994_),
    .Y(_11995_));
 AND3x1_ASAP7_75t_R _33039_ (.A(_06831_),
    .B(_11989_),
    .C(_11995_),
    .Y(_11996_));
 AO21x1_ASAP7_75t_R _33040_ (.A1(_11990_),
    .A2(_11991_),
    .B(_11996_),
    .Y(_11997_));
 BUFx4f_ASAP7_75t_R _33041_ (.A(_11997_),
    .Y(_11998_));
 BUFx6f_ASAP7_75t_R _33042_ (.A(_11998_),
    .Y(_11999_));
 INVx4_ASAP7_75t_R _33043_ (.A(_11992_),
    .Y(_12000_));
 BUFx6f_ASAP7_75t_R _33044_ (.A(_12000_),
    .Y(_12001_));
 BUFx3_ASAP7_75t_R _33045_ (.A(_11992_),
    .Y(_12002_));
 AND2x2_ASAP7_75t_R _33046_ (.A(_05479_),
    .B(_12002_),
    .Y(_12003_));
 AO21x1_ASAP7_75t_R _33047_ (.A1(_01710_),
    .A2(_12001_),
    .B(_12003_),
    .Y(_12004_));
 AND3x1_ASAP7_75t_R _33048_ (.A(_05490_),
    .B(_05508_),
    .C(_11947_),
    .Y(_12005_));
 AND3x1_ASAP7_75t_R _33049_ (.A(_06831_),
    .B(_11989_),
    .C(_11993_),
    .Y(_12006_));
 AO21x1_ASAP7_75t_R _33050_ (.A1(_11990_),
    .A2(_12005_),
    .B(_12006_),
    .Y(_12007_));
 BUFx4f_ASAP7_75t_R _33051_ (.A(_12007_),
    .Y(_12008_));
 BUFx6f_ASAP7_75t_R _33052_ (.A(_12008_),
    .Y(_12009_));
 AND2x4_ASAP7_75t_R _33053_ (.A(_06831_),
    .B(_11989_),
    .Y(_12010_));
 AO21x1_ASAP7_75t_R _33054_ (.A1(_12010_),
    .A2(_11994_),
    .B(_01711_),
    .Y(_12011_));
 OAI22x1_ASAP7_75t_R _33055_ (.A1(_11999_),
    .A2(_12004_),
    .B1(_12009_),
    .B2(_12011_),
    .Y(_03954_));
 NAND2x2_ASAP7_75t_R _33056_ (.A(_11992_),
    .B(_11994_),
    .Y(_12012_));
 BUFx6f_ASAP7_75t_R _33057_ (.A(_12012_),
    .Y(_12013_));
 BUFx4f_ASAP7_75t_R _33058_ (.A(_12013_),
    .Y(_12014_));
 BUFx6f_ASAP7_75t_R _33059_ (.A(_12012_),
    .Y(_12015_));
 NAND2x1_ASAP7_75t_R _33060_ (.A(_01710_),
    .B(_12015_),
    .Y(_12016_));
 OA21x2_ASAP7_75t_R _33061_ (.A1(net139),
    .A2(_12014_),
    .B(_12016_),
    .Y(_03955_));
 BUFx6f_ASAP7_75t_R _33062_ (.A(_11956_),
    .Y(_12017_));
 BUFx6f_ASAP7_75t_R _33063_ (.A(_12017_),
    .Y(_12018_));
 AND3x1_ASAP7_75t_R _33064_ (.A(_05482_),
    .B(_06859_),
    .C(_11955_),
    .Y(_12019_));
 OAI22x1_ASAP7_75t_R _33065_ (.A1(_05493_),
    .A2(_12018_),
    .B1(_12019_),
    .B2(_07313_),
    .Y(_12020_));
 OA222x2_ASAP7_75t_R _33066_ (.A1(_18764_),
    .A2(_05423_),
    .B1(_07230_),
    .B2(_01967_),
    .C1(_00789_),
    .C2(_05418_),
    .Y(_12021_));
 NAND2x1_ASAP7_75t_R _33067_ (.A(_11709_),
    .B(_12021_),
    .Y(_12022_));
 OA21x2_ASAP7_75t_R _33068_ (.A1(_11709_),
    .A2(_12020_),
    .B(_12022_),
    .Y(_03956_));
 BUFx6f_ASAP7_75t_R _33069_ (.A(_11957_),
    .Y(_12023_));
 INVx1_ASAP7_75t_R _33070_ (.A(_01689_),
    .Y(_12024_));
 NAND2x2_ASAP7_75t_R _33071_ (.A(_00295_),
    .B(_12024_),
    .Y(_12025_));
 OR3x1_ASAP7_75t_R _33072_ (.A(_07383_),
    .B(_07378_),
    .C(_12025_),
    .Y(_12026_));
 OR2x4_ASAP7_75t_R _33073_ (.A(_01685_),
    .B(_12026_),
    .Y(_12027_));
 NOR2x1_ASAP7_75t_R _33074_ (.A(_12023_),
    .B(_12027_),
    .Y(_12028_));
 NAND2x1_ASAP7_75t_R _33075_ (.A(_01709_),
    .B(_11889_),
    .Y(_12029_));
 OR3x2_ASAP7_75t_R _33076_ (.A(_01682_),
    .B(_07397_),
    .C(_07392_),
    .Y(_12030_));
 OA211x2_ASAP7_75t_R _33077_ (.A1(_07255_),
    .A2(_12030_),
    .B(_05467_),
    .C(_01709_),
    .Y(_12031_));
 NOR2x1_ASAP7_75t_R _33078_ (.A(_11677_),
    .B(_12031_),
    .Y(_12032_));
 OR3x2_ASAP7_75t_R _33079_ (.A(_07255_),
    .B(_01709_),
    .C(_12030_),
    .Y(_12033_));
 OR4x1_ASAP7_75t_R _33080_ (.A(_11731_),
    .B(_12017_),
    .C(_12027_),
    .D(_12033_),
    .Y(_12034_));
 OA211x2_ASAP7_75t_R _33081_ (.A1(_12028_),
    .A2(_12029_),
    .B(_12032_),
    .C(_12034_),
    .Y(_03957_));
 OR2x2_ASAP7_75t_R _33082_ (.A(_00292_),
    .B(_18319_),
    .Y(_12035_));
 AO21x2_ASAP7_75t_R _33083_ (.A1(_00294_),
    .A2(_12035_),
    .B(_01689_),
    .Y(_12036_));
 OR4x1_ASAP7_75t_R _33084_ (.A(_01685_),
    .B(_07383_),
    .C(_07378_),
    .D(_12036_),
    .Y(_12037_));
 OR3x1_ASAP7_75t_R _33085_ (.A(_11072_),
    .B(_11966_),
    .C(_12037_),
    .Y(_12038_));
 BUFx6f_ASAP7_75t_R _33086_ (.A(_12038_),
    .Y(_12039_));
 AND2x2_ASAP7_75t_R _33087_ (.A(_01708_),
    .B(_11703_),
    .Y(_12040_));
 AO32x1_ASAP7_75t_R _33088_ (.A1(_01708_),
    .A2(_11703_),
    .A3(_12033_),
    .B1(_11694_),
    .B2(_11689_),
    .Y(_12041_));
 OR3x1_ASAP7_75t_R _33089_ (.A(_01708_),
    .B(_11731_),
    .C(_12033_),
    .Y(_12042_));
 NOR2x1_ASAP7_75t_R _33090_ (.A(_12039_),
    .B(_12042_),
    .Y(_12043_));
 AOI211x1_ASAP7_75t_R _33091_ (.A1(_12039_),
    .A2(_12040_),
    .B(_12041_),
    .C(_12043_),
    .Y(_03958_));
 BUFx4f_ASAP7_75t_R _33092_ (.A(_05468_),
    .Y(_12044_));
 BUFx4f_ASAP7_75t_R _33093_ (.A(_11957_),
    .Y(_12045_));
 OR3x1_ASAP7_75t_R _33094_ (.A(_01708_),
    .B(_12027_),
    .C(_12033_),
    .Y(_12046_));
 AND2x2_ASAP7_75t_R _33095_ (.A(_01707_),
    .B(_05468_),
    .Y(_12047_));
 OAI21x1_ASAP7_75t_R _33096_ (.A1(_12045_),
    .A2(_12046_),
    .B(_12047_),
    .Y(_12048_));
 OR4x1_ASAP7_75t_R _33097_ (.A(_01707_),
    .B(_05390_),
    .C(_11957_),
    .D(_12046_),
    .Y(_12049_));
 OA211x2_ASAP7_75t_R _33098_ (.A1(_12044_),
    .A2(_11713_),
    .B(_12048_),
    .C(_12049_),
    .Y(_03959_));
 OR3x2_ASAP7_75t_R _33099_ (.A(_01707_),
    .B(_01708_),
    .C(_12033_),
    .Y(_12050_));
 OR4x1_ASAP7_75t_R _33100_ (.A(_07276_),
    .B(_11731_),
    .C(_12039_),
    .D(_12050_),
    .Y(_12051_));
 NAND3x1_ASAP7_75t_R _33101_ (.A(_07276_),
    .B(_11794_),
    .C(_12039_),
    .Y(_12052_));
 AND3x1_ASAP7_75t_R _33102_ (.A(_07276_),
    .B(_05468_),
    .C(_12050_),
    .Y(_12053_));
 NOR2x1_ASAP7_75t_R _33103_ (.A(_11719_),
    .B(_12053_),
    .Y(_12054_));
 AND3x1_ASAP7_75t_R _33104_ (.A(_12051_),
    .B(_12052_),
    .C(_12054_),
    .Y(_03960_));
 OR3x1_ASAP7_75t_R _33105_ (.A(_07276_),
    .B(_12027_),
    .C(_12050_),
    .Y(_12055_));
 AND2x2_ASAP7_75t_R _33106_ (.A(_01705_),
    .B(_05468_),
    .Y(_12056_));
 OAI21x1_ASAP7_75t_R _33107_ (.A1(_12045_),
    .A2(_12055_),
    .B(_12056_),
    .Y(_12057_));
 OR4x1_ASAP7_75t_R _33108_ (.A(_01705_),
    .B(_05390_),
    .C(_11957_),
    .D(_12055_),
    .Y(_12058_));
 OA211x2_ASAP7_75t_R _33109_ (.A1(_12044_),
    .A2(_11734_),
    .B(_12057_),
    .C(_12058_),
    .Y(_03961_));
 OR3x2_ASAP7_75t_R _33110_ (.A(_01705_),
    .B(_07276_),
    .C(_12050_),
    .Y(_12059_));
 OR4x1_ASAP7_75t_R _33111_ (.A(_07286_),
    .B(_11731_),
    .C(_12039_),
    .D(_12059_),
    .Y(_12060_));
 NAND3x1_ASAP7_75t_R _33112_ (.A(_07286_),
    .B(_11794_),
    .C(_12039_),
    .Y(_12061_));
 NAND2x1_ASAP7_75t_R _33113_ (.A(_07286_),
    .B(_12059_),
    .Y(_12062_));
 OA22x2_ASAP7_75t_R _33114_ (.A1(_11741_),
    .A2(_11742_),
    .B1(_12062_),
    .B2(_11731_),
    .Y(_12063_));
 AND3x1_ASAP7_75t_R _33115_ (.A(_12060_),
    .B(_12061_),
    .C(_12063_),
    .Y(_03962_));
 INVx1_ASAP7_75t_R _33116_ (.A(_07293_),
    .Y(_12064_));
 AO21x2_ASAP7_75t_R _33117_ (.A1(_06859_),
    .A2(_11955_),
    .B(_05390_),
    .Y(_12065_));
 OR3x1_ASAP7_75t_R _33118_ (.A(_07286_),
    .B(_12027_),
    .C(_12059_),
    .Y(_12066_));
 OR4x1_ASAP7_75t_R _33119_ (.A(_07293_),
    .B(_11756_),
    .C(_11957_),
    .D(_12066_),
    .Y(_12067_));
 NAND2x1_ASAP7_75t_R _33120_ (.A(_07293_),
    .B(_12066_),
    .Y(_12068_));
 AO21x1_ASAP7_75t_R _33121_ (.A1(_11703_),
    .A2(_12068_),
    .B(_11756_),
    .Y(_12069_));
 OA211x2_ASAP7_75t_R _33122_ (.A1(_12064_),
    .A2(_12065_),
    .B(_12067_),
    .C(_12069_),
    .Y(_03963_));
 OR3x1_ASAP7_75t_R _33123_ (.A(_07286_),
    .B(_12037_),
    .C(_12059_),
    .Y(_12070_));
 NOR2x1_ASAP7_75t_R _33124_ (.A(_07293_),
    .B(_12070_),
    .Y(_12071_));
 AND3x1_ASAP7_75t_R _33125_ (.A(_06831_),
    .B(_11955_),
    .C(_12071_),
    .Y(_12072_));
 XOR2x1_ASAP7_75t_R _33126_ (.A(_01702_),
    .Y(_12073_),
    .B(_12072_));
 AOI21x1_ASAP7_75t_R _33127_ (.A1(_11704_),
    .A2(_12073_),
    .B(_11765_),
    .Y(_03964_));
 AND2x2_ASAP7_75t_R _33128_ (.A(_06830_),
    .B(_11955_),
    .Y(_12074_));
 BUFx6f_ASAP7_75t_R _33129_ (.A(_12074_),
    .Y(_12075_));
 OR3x4_ASAP7_75t_R _33130_ (.A(_01702_),
    .B(_07293_),
    .C(_12066_),
    .Y(_12076_));
 NOR2x1_ASAP7_75t_R _33131_ (.A(_07302_),
    .B(_12076_),
    .Y(_12077_));
 AO21x1_ASAP7_75t_R _33132_ (.A1(_12075_),
    .A2(_12077_),
    .B(_11709_),
    .Y(_12078_));
 AO22x1_ASAP7_75t_R _33133_ (.A1(_11889_),
    .A2(_12045_),
    .B1(_12076_),
    .B2(_11778_),
    .Y(_12079_));
 AOI22x1_ASAP7_75t_R _33134_ (.A1(_11778_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_07302_),
    .Y(_03965_));
 BUFx4f_ASAP7_75t_R _33135_ (.A(_12074_),
    .Y(_12080_));
 OR3x2_ASAP7_75t_R _33136_ (.A(_01702_),
    .B(_07293_),
    .C(_12070_),
    .Y(_12081_));
 NOR2x1_ASAP7_75t_R _33137_ (.A(_07302_),
    .B(_12081_),
    .Y(_12082_));
 NAND2x1_ASAP7_75t_R _33138_ (.A(_01700_),
    .B(_05468_),
    .Y(_12083_));
 AO21x1_ASAP7_75t_R _33139_ (.A1(_12080_),
    .A2(_12082_),
    .B(_12083_),
    .Y(_12084_));
 OR5x1_ASAP7_75t_R _33140_ (.A(_01700_),
    .B(_07302_),
    .C(_05390_),
    .D(_11957_),
    .E(_12081_),
    .Y(_12085_));
 AND3x1_ASAP7_75t_R _33141_ (.A(_11791_),
    .B(_12084_),
    .C(_12085_),
    .Y(_03966_));
 INVx1_ASAP7_75t_R _33142_ (.A(_00293_),
    .Y(_12086_));
 OR3x1_ASAP7_75t_R _33143_ (.A(_12086_),
    .B(_11072_),
    .C(_11966_),
    .Y(_12087_));
 AO21x1_ASAP7_75t_R _33144_ (.A1(_06859_),
    .A2(_11955_),
    .B(_18317_),
    .Y(_12088_));
 AO21x1_ASAP7_75t_R _33145_ (.A1(_12087_),
    .A2(_12088_),
    .B(_11709_),
    .Y(_12089_));
 NAND2x1_ASAP7_75t_R _33146_ (.A(_05434_),
    .B(_12089_),
    .Y(_03967_));
 OR2x2_ASAP7_75t_R _33147_ (.A(_01700_),
    .B(_07302_),
    .Y(_12090_));
 OR4x1_ASAP7_75t_R _33148_ (.A(_11072_),
    .B(_11966_),
    .C(_12076_),
    .D(_12090_),
    .Y(_12091_));
 XNOR2x1_ASAP7_75t_R _33149_ (.B(_12091_),
    .Y(_12092_),
    .A(_01699_));
 AOI21x1_ASAP7_75t_R _33150_ (.A1(_11704_),
    .A2(_12092_),
    .B(_11803_),
    .Y(_03968_));
 OR4x1_ASAP7_75t_R _33151_ (.A(_01698_),
    .B(_01699_),
    .C(_01700_),
    .D(_05389_),
    .Y(_12093_));
 OR4x1_ASAP7_75t_R _33152_ (.A(_07302_),
    .B(_12017_),
    .C(_12081_),
    .D(_12093_),
    .Y(_12094_));
 NAND2x1_ASAP7_75t_R _33153_ (.A(_01698_),
    .B(_05468_),
    .Y(_12095_));
 AO21x1_ASAP7_75t_R _33154_ (.A1(_12080_),
    .A2(_12082_),
    .B(_12095_),
    .Y(_12096_));
 OA21x2_ASAP7_75t_R _33155_ (.A1(_01699_),
    .A2(_01700_),
    .B(_01698_),
    .Y(_12097_));
 NAND2x1_ASAP7_75t_R _33156_ (.A(_11794_),
    .B(_12097_),
    .Y(_12098_));
 AND4x1_ASAP7_75t_R _33157_ (.A(_11810_),
    .B(_12094_),
    .C(_12096_),
    .D(_12098_),
    .Y(_03969_));
 OR3x2_ASAP7_75t_R _33158_ (.A(_01698_),
    .B(_01699_),
    .C(_12090_),
    .Y(_12099_));
 OR2x2_ASAP7_75t_R _33159_ (.A(_12076_),
    .B(_12099_),
    .Y(_12100_));
 OAI21x1_ASAP7_75t_R _33160_ (.A1(_12018_),
    .A2(_12100_),
    .B(_07333_),
    .Y(_12101_));
 OR4x1_ASAP7_75t_R _33161_ (.A(_07333_),
    .B(_12017_),
    .C(_12076_),
    .D(_12099_),
    .Y(_12102_));
 INVx1_ASAP7_75t_R _33162_ (.A(_11821_),
    .Y(_12103_));
 AO31x2_ASAP7_75t_R _33163_ (.A1(_11704_),
    .A2(_12101_),
    .A3(_12102_),
    .B(_12103_),
    .Y(_03970_));
 OR2x2_ASAP7_75t_R _33164_ (.A(_12081_),
    .B(_12099_),
    .Y(_12104_));
 OR5x1_ASAP7_75t_R _33165_ (.A(_01696_),
    .B(_07333_),
    .C(_05390_),
    .D(_11957_),
    .E(_12104_),
    .Y(_12105_));
 AND2x2_ASAP7_75t_R _33166_ (.A(_01696_),
    .B(_05468_),
    .Y(_12106_));
 OAI21x1_ASAP7_75t_R _33167_ (.A1(_07333_),
    .A2(_12045_),
    .B(_12106_),
    .Y(_12107_));
 AND3x1_ASAP7_75t_R _33168_ (.A(_01696_),
    .B(_05468_),
    .C(_12104_),
    .Y(_12108_));
 INVx1_ASAP7_75t_R _33169_ (.A(_12108_),
    .Y(_12109_));
 AND4x1_ASAP7_75t_R _33170_ (.A(_11831_),
    .B(_12105_),
    .C(_12107_),
    .D(_12109_),
    .Y(_03971_));
 OR4x2_ASAP7_75t_R _33171_ (.A(_01696_),
    .B(_07333_),
    .C(_12076_),
    .D(_12099_),
    .Y(_12110_));
 OR3x2_ASAP7_75t_R _33172_ (.A(_11072_),
    .B(_11966_),
    .C(_12110_),
    .Y(_12111_));
 OA21x2_ASAP7_75t_R _33173_ (.A1(_01695_),
    .A2(_12111_),
    .B(_11794_),
    .Y(_12112_));
 INVx1_ASAP7_75t_R _33174_ (.A(_12110_),
    .Y(_12113_));
 OA21x2_ASAP7_75t_R _33175_ (.A1(_11842_),
    .A2(_12113_),
    .B(_12065_),
    .Y(_12114_));
 INVx1_ASAP7_75t_R _33176_ (.A(_01695_),
    .Y(_12115_));
 OA22x2_ASAP7_75t_R _33177_ (.A1(_11842_),
    .A2(_12112_),
    .B1(_12114_),
    .B2(_12115_),
    .Y(_03972_));
 OR2x2_ASAP7_75t_R _33178_ (.A(_05467_),
    .B(_11851_),
    .Y(_12116_));
 BUFx6f_ASAP7_75t_R _33179_ (.A(_12017_),
    .Y(_12117_));
 OR3x4_ASAP7_75t_R _33180_ (.A(_01696_),
    .B(_07333_),
    .C(_12104_),
    .Y(_12118_));
 OR3x1_ASAP7_75t_R _33181_ (.A(_01694_),
    .B(_01695_),
    .C(_12118_),
    .Y(_12119_));
 OAI21x1_ASAP7_75t_R _33182_ (.A1(_12117_),
    .A2(_12119_),
    .B(_12044_),
    .Y(_12120_));
 OA21x2_ASAP7_75t_R _33183_ (.A1(_01695_),
    .A2(_12118_),
    .B(_12116_),
    .Y(_12121_));
 AO21x1_ASAP7_75t_R _33184_ (.A1(_12044_),
    .A2(_12045_),
    .B(_12121_),
    .Y(_12122_));
 AOI22x1_ASAP7_75t_R _33185_ (.A1(_12116_),
    .A2(_12120_),
    .B1(_12122_),
    .B2(_01694_),
    .Y(_03973_));
 OR3x1_ASAP7_75t_R _33186_ (.A(_01694_),
    .B(_01695_),
    .C(_12110_),
    .Y(_12123_));
 AO22x1_ASAP7_75t_R _33187_ (.A1(_11889_),
    .A2(_12023_),
    .B1(_12123_),
    .B2(_11865_),
    .Y(_12124_));
 OR3x4_ASAP7_75t_R _33188_ (.A(_01693_),
    .B(_01694_),
    .C(_01695_),
    .Y(_12125_));
 OAI21x1_ASAP7_75t_R _33189_ (.A1(_12111_),
    .A2(_12125_),
    .B(_11704_),
    .Y(_12126_));
 AOI22x1_ASAP7_75t_R _33190_ (.A1(_01693_),
    .A2(_12124_),
    .B1(_12126_),
    .B2(_11865_),
    .Y(_03974_));
 INVx1_ASAP7_75t_R _33191_ (.A(_01692_),
    .Y(_12127_));
 AND2x2_ASAP7_75t_R _33192_ (.A(_05389_),
    .B(_11875_),
    .Y(_12128_));
 OR2x2_ASAP7_75t_R _33193_ (.A(_01692_),
    .B(_12125_),
    .Y(_12129_));
 OR4x1_ASAP7_75t_R _33194_ (.A(_12128_),
    .B(_12017_),
    .C(_12118_),
    .D(_12129_),
    .Y(_12130_));
 OAI21x1_ASAP7_75t_R _33195_ (.A1(_12118_),
    .A2(_12125_),
    .B(_01692_),
    .Y(_12131_));
 AO21x1_ASAP7_75t_R _33196_ (.A1(_11703_),
    .A2(_12131_),
    .B(_12128_),
    .Y(_12132_));
 OA211x2_ASAP7_75t_R _33197_ (.A1(_12127_),
    .A2(_12065_),
    .B(_12130_),
    .C(_12132_),
    .Y(_03975_));
 OA21x2_ASAP7_75t_R _33198_ (.A1(_12110_),
    .A2(_12129_),
    .B(_11884_),
    .Y(_12133_));
 AO21x1_ASAP7_75t_R _33199_ (.A1(_12044_),
    .A2(_12045_),
    .B(_12133_),
    .Y(_12134_));
 OR3x1_ASAP7_75t_R _33200_ (.A(_01691_),
    .B(_01692_),
    .C(_12125_),
    .Y(_12135_));
 OAI21x1_ASAP7_75t_R _33201_ (.A1(_12111_),
    .A2(_12135_),
    .B(_11704_),
    .Y(_12136_));
 AOI22x1_ASAP7_75t_R _33202_ (.A1(_01691_),
    .A2(_12134_),
    .B1(_12136_),
    .B2(_11884_),
    .Y(_03976_));
 INVx1_ASAP7_75t_R _33203_ (.A(_01690_),
    .Y(_12137_));
 OR3x1_ASAP7_75t_R _33204_ (.A(_01690_),
    .B(_01691_),
    .C(_12129_),
    .Y(_12138_));
 OR4x1_ASAP7_75t_R _33205_ (.A(_11895_),
    .B(_12017_),
    .C(_12118_),
    .D(_12138_),
    .Y(_12139_));
 OR3x1_ASAP7_75t_R _33206_ (.A(_01691_),
    .B(_12118_),
    .C(_12129_),
    .Y(_12140_));
 NAND2x1_ASAP7_75t_R _33207_ (.A(_01690_),
    .B(_12140_),
    .Y(_12141_));
 AO21x1_ASAP7_75t_R _33208_ (.A1(_11703_),
    .A2(_12141_),
    .B(_11895_),
    .Y(_12142_));
 OA211x2_ASAP7_75t_R _33209_ (.A1(_12137_),
    .A2(_12065_),
    .B(_12139_),
    .C(_12142_),
    .Y(_03977_));
 INVx1_ASAP7_75t_R _33210_ (.A(_00295_),
    .Y(_12143_));
 OR2x2_ASAP7_75t_R _33211_ (.A(_05433_),
    .B(_05463_),
    .Y(_12144_));
 AO22x1_ASAP7_75t_R _33212_ (.A1(_12143_),
    .A2(_12144_),
    .B1(_12045_),
    .B2(_11794_),
    .Y(_12145_));
 OAI21x1_ASAP7_75t_R _33213_ (.A1(_12117_),
    .A2(_12025_),
    .B(_11704_),
    .Y(_12146_));
 AOI22x1_ASAP7_75t_R _33214_ (.A1(_01689_),
    .A2(_12145_),
    .B1(_12146_),
    .B2(_12144_),
    .Y(_03978_));
 OR3x1_ASAP7_75t_R _33215_ (.A(_01688_),
    .B(_12110_),
    .C(_12138_),
    .Y(_12147_));
 OAI21x1_ASAP7_75t_R _33216_ (.A1(_12117_),
    .A2(_12147_),
    .B(_12044_),
    .Y(_12148_));
 OA21x2_ASAP7_75t_R _33217_ (.A1(_12110_),
    .A2(_12138_),
    .B(_11903_),
    .Y(_12149_));
 AO21x1_ASAP7_75t_R _33218_ (.A1(_12044_),
    .A2(_12045_),
    .B(_12149_),
    .Y(_12150_));
 AOI22x1_ASAP7_75t_R _33219_ (.A1(_11903_),
    .A2(_12148_),
    .B1(_12150_),
    .B2(_01688_),
    .Y(_03979_));
 NOR2x1_ASAP7_75t_R _33220_ (.A(_07378_),
    .B(_12036_),
    .Y(_12151_));
 AO21x1_ASAP7_75t_R _33221_ (.A1(_12075_),
    .A2(_12151_),
    .B(_11709_),
    .Y(_12152_));
 AO22x1_ASAP7_75t_R _33222_ (.A1(_11889_),
    .A2(_12045_),
    .B1(_12036_),
    .B2(_11640_),
    .Y(_12153_));
 AOI22x1_ASAP7_75t_R _33223_ (.A1(_11640_),
    .A2(_12152_),
    .B1(_12153_),
    .B2(_07378_),
    .Y(_03980_));
 BUFx6f_ASAP7_75t_R _33224_ (.A(_12017_),
    .Y(_12154_));
 OAI21x1_ASAP7_75t_R _33225_ (.A1(_12154_),
    .A2(_12026_),
    .B(_12044_),
    .Y(_12155_));
 OA21x2_ASAP7_75t_R _33226_ (.A1(_07378_),
    .A2(_12025_),
    .B(_11645_),
    .Y(_12156_));
 AO21x1_ASAP7_75t_R _33227_ (.A1(_12044_),
    .A2(_12045_),
    .B(_12156_),
    .Y(_12157_));
 AOI22x1_ASAP7_75t_R _33228_ (.A1(_11645_),
    .A2(_12155_),
    .B1(_12157_),
    .B2(_07383_),
    .Y(_03981_));
 OR3x1_ASAP7_75t_R _33229_ (.A(_07383_),
    .B(_07378_),
    .C(_12036_),
    .Y(_12158_));
 OR2x2_ASAP7_75t_R _33230_ (.A(_05433_),
    .B(_11636_),
    .Y(_12159_));
 AO22x1_ASAP7_75t_R _33231_ (.A1(_11794_),
    .A2(_12023_),
    .B1(_12158_),
    .B2(_12159_),
    .Y(_12160_));
 NAND2x1_ASAP7_75t_R _33232_ (.A(_12044_),
    .B(_12039_),
    .Y(_12161_));
 AOI22x1_ASAP7_75t_R _33233_ (.A1(_01685_),
    .A2(_12160_),
    .B1(_12161_),
    .B2(_12159_),
    .Y(_03982_));
 NAND2x1_ASAP7_75t_R _33234_ (.A(_07392_),
    .B(_11889_),
    .Y(_12162_));
 OR4x1_ASAP7_75t_R _33235_ (.A(_07392_),
    .B(_05390_),
    .C(_11957_),
    .D(_12027_),
    .Y(_12163_));
 OA211x2_ASAP7_75t_R _33236_ (.A1(_12028_),
    .A2(_12162_),
    .B(_12163_),
    .C(_11663_),
    .Y(_03983_));
 NAND3x1_ASAP7_75t_R _33237_ (.A(_07397_),
    .B(_11794_),
    .C(_12039_),
    .Y(_12164_));
 OR4x1_ASAP7_75t_R _33238_ (.A(_07397_),
    .B(_07392_),
    .C(_05390_),
    .D(_12038_),
    .Y(_12165_));
 NAND3x1_ASAP7_75t_R _33239_ (.A(_07397_),
    .B(_07392_),
    .C(_11703_),
    .Y(_12166_));
 AND4x1_ASAP7_75t_R _33240_ (.A(_11653_),
    .B(_12164_),
    .C(_12165_),
    .D(_12166_),
    .Y(_03984_));
 NAND2x1_ASAP7_75t_R _33241_ (.A(_01682_),
    .B(_11889_),
    .Y(_12167_));
 OAI21x1_ASAP7_75t_R _33242_ (.A1(_07397_),
    .A2(_07392_),
    .B(_01682_),
    .Y(_12168_));
 OA21x2_ASAP7_75t_R _33243_ (.A1(_11731_),
    .A2(_12168_),
    .B(_11658_),
    .Y(_12169_));
 OR4x1_ASAP7_75t_R _33244_ (.A(_11731_),
    .B(_12017_),
    .C(_12027_),
    .D(_12030_),
    .Y(_12170_));
 OA211x2_ASAP7_75t_R _33245_ (.A1(_12028_),
    .A2(_12167_),
    .B(_12169_),
    .C(_12170_),
    .Y(_03985_));
 NAND3x1_ASAP7_75t_R _33246_ (.A(_07255_),
    .B(_11794_),
    .C(_12039_),
    .Y(_12171_));
 OR4x1_ASAP7_75t_R _33247_ (.A(_07255_),
    .B(_11731_),
    .C(_12030_),
    .D(_12039_),
    .Y(_12172_));
 AND2x2_ASAP7_75t_R _33248_ (.A(_07255_),
    .B(_12030_),
    .Y(_12173_));
 AOI22x1_ASAP7_75t_R _33249_ (.A1(_11625_),
    .A2(_11631_),
    .B1(_12173_),
    .B2(_11889_),
    .Y(_12174_));
 AND3x1_ASAP7_75t_R _33250_ (.A(_12171_),
    .B(_12172_),
    .C(_12174_),
    .Y(_03986_));
 NOR2x1_ASAP7_75t_R _33251_ (.A(_01680_),
    .B(_11975_),
    .Y(_12175_));
 NAND2x1_ASAP7_75t_R _33252_ (.A(_11977_),
    .B(_01655_),
    .Y(_12176_));
 OA21x2_ASAP7_75t_R _33253_ (.A1(net141),
    .A2(_11977_),
    .B(_12176_),
    .Y(_12177_));
 AO32x1_ASAP7_75t_R _33254_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12175_),
    .B1(_12177_),
    .B2(_11988_),
    .Y(_03987_));
 NOR2x1_ASAP7_75t_R _33255_ (.A(_01679_),
    .B(_11975_),
    .Y(_12178_));
 NAND2x1_ASAP7_75t_R _33256_ (.A(_11949_),
    .B(_01644_),
    .Y(_12179_));
 OA21x2_ASAP7_75t_R _33257_ (.A1(net142),
    .A2(_11977_),
    .B(_12179_),
    .Y(_12180_));
 AO32x1_ASAP7_75t_R _33258_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12178_),
    .B1(_12180_),
    .B2(_11988_),
    .Y(_03988_));
 NOR2x1_ASAP7_75t_R _33259_ (.A(_01678_),
    .B(_11975_),
    .Y(_12181_));
 BUFx4f_ASAP7_75t_R _33260_ (.A(_11949_),
    .Y(_12182_));
 NAND2x1_ASAP7_75t_R _33261_ (.A(_11977_),
    .B(_01643_),
    .Y(_12183_));
 OA21x2_ASAP7_75t_R _33262_ (.A1(net143),
    .A2(_12182_),
    .B(_12183_),
    .Y(_12184_));
 AO32x1_ASAP7_75t_R _33263_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12181_),
    .B1(_12184_),
    .B2(_11988_),
    .Y(_03989_));
 NOR2x1_ASAP7_75t_R _33264_ (.A(_01677_),
    .B(_11975_),
    .Y(_12185_));
 NAND2x1_ASAP7_75t_R _33265_ (.A(_12182_),
    .B(_01642_),
    .Y(_12186_));
 OA21x2_ASAP7_75t_R _33266_ (.A1(net144),
    .A2(_11978_),
    .B(_12186_),
    .Y(_12187_));
 AO32x1_ASAP7_75t_R _33267_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12185_),
    .B1(_12187_),
    .B2(_11988_),
    .Y(_03990_));
 NOR2x1_ASAP7_75t_R _33268_ (.A(_01676_),
    .B(_11975_),
    .Y(_12188_));
 NAND2x1_ASAP7_75t_R _33269_ (.A(_12182_),
    .B(_01641_),
    .Y(_12189_));
 OA21x2_ASAP7_75t_R _33270_ (.A1(net146),
    .A2(_11978_),
    .B(_12189_),
    .Y(_12190_));
 AO32x1_ASAP7_75t_R _33271_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12188_),
    .B1(_12190_),
    .B2(_11988_),
    .Y(_03991_));
 NOR2x1_ASAP7_75t_R _33272_ (.A(_01675_),
    .B(_11975_),
    .Y(_12191_));
 NAND2x1_ASAP7_75t_R _33273_ (.A(_11949_),
    .B(_01640_),
    .Y(_12192_));
 OA21x2_ASAP7_75t_R _33274_ (.A1(net147),
    .A2(_11977_),
    .B(_12192_),
    .Y(_12193_));
 AO32x1_ASAP7_75t_R _33275_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12191_),
    .B1(_12193_),
    .B2(_11988_),
    .Y(_03992_));
 NOR2x1_ASAP7_75t_R _33276_ (.A(_01674_),
    .B(_11975_),
    .Y(_12194_));
 NAND2x1_ASAP7_75t_R _33277_ (.A(_11978_),
    .B(_01639_),
    .Y(_12195_));
 OA21x2_ASAP7_75t_R _33278_ (.A1(net148),
    .A2(_11978_),
    .B(_12195_),
    .Y(_12196_));
 AO32x1_ASAP7_75t_R _33279_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12194_),
    .B1(_12196_),
    .B2(_11988_),
    .Y(_03993_));
 NOR2x1_ASAP7_75t_R _33280_ (.A(_01673_),
    .B(_11975_),
    .Y(_12197_));
 NAND2x1_ASAP7_75t_R _33281_ (.A(_11981_),
    .B(_01638_),
    .Y(_12198_));
 OA21x2_ASAP7_75t_R _33282_ (.A1(net149),
    .A2(_11980_),
    .B(_12198_),
    .Y(_12199_));
 AO32x1_ASAP7_75t_R _33283_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12197_),
    .B1(_12199_),
    .B2(_11988_),
    .Y(_03994_));
 NOR2x1_ASAP7_75t_R _33284_ (.A(_01672_),
    .B(_11975_),
    .Y(_12200_));
 BUFx6f_ASAP7_75t_R _33285_ (.A(_11979_),
    .Y(_12201_));
 NAND2x1_ASAP7_75t_R _33286_ (.A(_12201_),
    .B(_01637_),
    .Y(_12202_));
 OA21x2_ASAP7_75t_R _33287_ (.A1(net150),
    .A2(_11980_),
    .B(_12202_),
    .Y(_12203_));
 AO32x1_ASAP7_75t_R _33288_ (.A1(_11970_),
    .A2(_11973_),
    .A3(_12200_),
    .B1(_12203_),
    .B2(_11988_),
    .Y(_03995_));
 BUFx3_ASAP7_75t_R _33289_ (.A(_11969_),
    .Y(_12204_));
 BUFx3_ASAP7_75t_R _33290_ (.A(_11972_),
    .Y(_12205_));
 BUFx6f_ASAP7_75t_R _33291_ (.A(_11974_),
    .Y(_12206_));
 NOR2x1_ASAP7_75t_R _33292_ (.A(_01671_),
    .B(_12206_),
    .Y(_12207_));
 NAND2x1_ASAP7_75t_R _33293_ (.A(_12201_),
    .B(_01635_),
    .Y(_12208_));
 OA21x2_ASAP7_75t_R _33294_ (.A1(net154),
    .A2(_11980_),
    .B(_12208_),
    .Y(_12209_));
 BUFx3_ASAP7_75t_R _33295_ (.A(_11987_),
    .Y(_12210_));
 AO32x1_ASAP7_75t_R _33296_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12207_),
    .B1(_12209_),
    .B2(_12210_),
    .Y(_03996_));
 NOR2x1_ASAP7_75t_R _33297_ (.A(_01670_),
    .B(_12206_),
    .Y(_12211_));
 NAND2x1_ASAP7_75t_R _33298_ (.A(_12201_),
    .B(_01634_),
    .Y(_12212_));
 OA21x2_ASAP7_75t_R _33299_ (.A1(net155),
    .A2(_11980_),
    .B(_12212_),
    .Y(_12213_));
 AO32x1_ASAP7_75t_R _33300_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12211_),
    .B1(_12213_),
    .B2(_12210_),
    .Y(_03997_));
 NOR2x1_ASAP7_75t_R _33301_ (.A(_01669_),
    .B(_12206_),
    .Y(_12214_));
 NAND2x1_ASAP7_75t_R _33302_ (.A(_12182_),
    .B(_01654_),
    .Y(_12215_));
 OA21x2_ASAP7_75t_R _33303_ (.A1(net156),
    .A2(_12182_),
    .B(_12215_),
    .Y(_12216_));
 AO32x1_ASAP7_75t_R _33304_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12214_),
    .B1(_12216_),
    .B2(_12210_),
    .Y(_03998_));
 NOR2x1_ASAP7_75t_R _33305_ (.A(_01668_),
    .B(_12206_),
    .Y(_12217_));
 NAND2x1_ASAP7_75t_R _33306_ (.A(_12201_),
    .B(_01633_),
    .Y(_12218_));
 OA21x2_ASAP7_75t_R _33307_ (.A1(net157),
    .A2(_11980_),
    .B(_12218_),
    .Y(_12219_));
 AO32x1_ASAP7_75t_R _33308_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12217_),
    .B1(_12219_),
    .B2(_12210_),
    .Y(_03999_));
 NOR2x1_ASAP7_75t_R _33309_ (.A(_01667_),
    .B(_12206_),
    .Y(_12220_));
 NAND2x1_ASAP7_75t_R _33310_ (.A(_12201_),
    .B(_01632_),
    .Y(_12221_));
 OA21x2_ASAP7_75t_R _33311_ (.A1(net158),
    .A2(_11980_),
    .B(_12221_),
    .Y(_12222_));
 AO32x1_ASAP7_75t_R _33312_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12220_),
    .B1(_12222_),
    .B2(_12210_),
    .Y(_04000_));
 NOR2x1_ASAP7_75t_R _33313_ (.A(_01666_),
    .B(_12206_),
    .Y(_12223_));
 NAND2x1_ASAP7_75t_R _33314_ (.A(_12201_),
    .B(_01631_),
    .Y(_12224_));
 OA21x2_ASAP7_75t_R _33315_ (.A1(net159),
    .A2(_11980_),
    .B(_12224_),
    .Y(_12225_));
 AO32x1_ASAP7_75t_R _33316_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12223_),
    .B1(_12225_),
    .B2(_12210_),
    .Y(_04001_));
 NOR2x1_ASAP7_75t_R _33317_ (.A(_01665_),
    .B(_12206_),
    .Y(_12226_));
 NAND2x1_ASAP7_75t_R _33318_ (.A(_12201_),
    .B(_01630_),
    .Y(_12227_));
 OA21x2_ASAP7_75t_R _33319_ (.A1(net160),
    .A2(_11980_),
    .B(_12227_),
    .Y(_12228_));
 AO32x1_ASAP7_75t_R _33320_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12226_),
    .B1(_12228_),
    .B2(_12210_),
    .Y(_04002_));
 NOR2x1_ASAP7_75t_R _33321_ (.A(_01664_),
    .B(_12206_),
    .Y(_12229_));
 NAND2x1_ASAP7_75t_R _33322_ (.A(_12201_),
    .B(_01629_),
    .Y(_12230_));
 OA21x2_ASAP7_75t_R _33323_ (.A1(net161),
    .A2(_11981_),
    .B(_12230_),
    .Y(_12231_));
 AO32x1_ASAP7_75t_R _33324_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12229_),
    .B1(_12231_),
    .B2(_12210_),
    .Y(_04003_));
 NOR2x1_ASAP7_75t_R _33325_ (.A(_01663_),
    .B(_12206_),
    .Y(_12232_));
 NAND2x1_ASAP7_75t_R _33326_ (.A(_12201_),
    .B(_01628_),
    .Y(_12233_));
 OA21x2_ASAP7_75t_R _33327_ (.A1(net162),
    .A2(_11981_),
    .B(_12233_),
    .Y(_12234_));
 AO32x1_ASAP7_75t_R _33328_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12232_),
    .B1(_12234_),
    .B2(_12210_),
    .Y(_04004_));
 NOR2x1_ASAP7_75t_R _33329_ (.A(_01662_),
    .B(_12206_),
    .Y(_12235_));
 NAND2x1_ASAP7_75t_R _33330_ (.A(_12201_),
    .B(_01627_),
    .Y(_12236_));
 OA21x2_ASAP7_75t_R _33331_ (.A1(net163),
    .A2(_11981_),
    .B(_12236_),
    .Y(_12237_));
 AO32x1_ASAP7_75t_R _33332_ (.A1(_12204_),
    .A2(_12205_),
    .A3(_12235_),
    .B1(_12237_),
    .B2(_12210_),
    .Y(_04005_));
 BUFx3_ASAP7_75t_R _33333_ (.A(_11969_),
    .Y(_12238_));
 BUFx3_ASAP7_75t_R _33334_ (.A(_11972_),
    .Y(_12239_));
 BUFx6f_ASAP7_75t_R _33335_ (.A(_11974_),
    .Y(_12240_));
 NOR2x1_ASAP7_75t_R _33336_ (.A(_01661_),
    .B(_12240_),
    .Y(_12241_));
 NAND2x1_ASAP7_75t_R _33337_ (.A(_11979_),
    .B(_01626_),
    .Y(_12242_));
 OA21x2_ASAP7_75t_R _33338_ (.A1(net164),
    .A2(_11981_),
    .B(_12242_),
    .Y(_12243_));
 BUFx2_ASAP7_75t_R _33339_ (.A(_11987_),
    .Y(_12244_));
 AO32x1_ASAP7_75t_R _33340_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12241_),
    .B1(_12243_),
    .B2(_12244_),
    .Y(_04006_));
 NOR2x1_ASAP7_75t_R _33341_ (.A(_01660_),
    .B(_12240_),
    .Y(_12245_));
 NAND2x1_ASAP7_75t_R _33342_ (.A(_11979_),
    .B(_01624_),
    .Y(_12246_));
 OA21x2_ASAP7_75t_R _33343_ (.A1(net165),
    .A2(_11981_),
    .B(_12246_),
    .Y(_12247_));
 AO32x1_ASAP7_75t_R _33344_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12245_),
    .B1(_12247_),
    .B2(_12244_),
    .Y(_04007_));
 NOR2x1_ASAP7_75t_R _33345_ (.A(_01659_),
    .B(_12240_),
    .Y(_12248_));
 NAND2x1_ASAP7_75t_R _33346_ (.A(_11979_),
    .B(_01623_),
    .Y(_12249_));
 OA21x2_ASAP7_75t_R _33347_ (.A1(net166),
    .A2(_11981_),
    .B(_12249_),
    .Y(_12250_));
 AO32x1_ASAP7_75t_R _33348_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12248_),
    .B1(_12250_),
    .B2(_12244_),
    .Y(_04008_));
 NOR2x1_ASAP7_75t_R _33349_ (.A(_01658_),
    .B(_12240_),
    .Y(_12251_));
 INVx1_ASAP7_75t_R _33350_ (.A(net167),
    .Y(_12252_));
 AND2x2_ASAP7_75t_R _33351_ (.A(_12252_),
    .B(_05508_),
    .Y(_12253_));
 AO21x1_ASAP7_75t_R _33352_ (.A1(_11977_),
    .A2(_01653_),
    .B(_12253_),
    .Y(_12254_));
 INVx1_ASAP7_75t_R _33353_ (.A(_12254_),
    .Y(_12255_));
 AO32x1_ASAP7_75t_R _33354_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12251_),
    .B1(_12255_),
    .B2(_12244_),
    .Y(_04009_));
 NOR2x1_ASAP7_75t_R _33355_ (.A(_01657_),
    .B(_12240_),
    .Y(_12256_));
 NAND2x1_ASAP7_75t_R _33356_ (.A(_11979_),
    .B(_01622_),
    .Y(_12257_));
 OA21x2_ASAP7_75t_R _33357_ (.A1(net168),
    .A2(_11981_),
    .B(_12257_),
    .Y(_12258_));
 AO32x1_ASAP7_75t_R _33358_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12256_),
    .B1(_12258_),
    .B2(_12244_),
    .Y(_04010_));
 NOR2x1_ASAP7_75t_R _33359_ (.A(_01656_),
    .B(_12240_),
    .Y(_12259_));
 NAND2x1_ASAP7_75t_R _33360_ (.A(_11979_),
    .B(_01621_),
    .Y(_12260_));
 OA21x2_ASAP7_75t_R _33361_ (.A1(net169),
    .A2(_11981_),
    .B(_12260_),
    .Y(_12261_));
 AO32x1_ASAP7_75t_R _33362_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12259_),
    .B1(_12261_),
    .B2(_12244_),
    .Y(_04011_));
 BUFx6f_ASAP7_75t_R _33363_ (.A(_12000_),
    .Y(_12262_));
 BUFx6f_ASAP7_75t_R _33364_ (.A(_12000_),
    .Y(_12263_));
 NAND2x1_ASAP7_75t_R _33365_ (.A(_01620_),
    .B(_12263_),
    .Y(_12264_));
 OAI21x1_ASAP7_75t_R _33366_ (.A1(net141),
    .A2(_12262_),
    .B(_12264_),
    .Y(_12265_));
 BUFx4f_ASAP7_75t_R _33367_ (.A(_12010_),
    .Y(_12266_));
 BUFx4f_ASAP7_75t_R _33368_ (.A(_11994_),
    .Y(_12267_));
 AO21x1_ASAP7_75t_R _33369_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01655_),
    .Y(_12268_));
 OAI22x1_ASAP7_75t_R _33370_ (.A1(_11999_),
    .A2(_12265_),
    .B1(_12268_),
    .B2(_12009_),
    .Y(_04012_));
 NAND2x1_ASAP7_75t_R _33371_ (.A(_01619_),
    .B(_12263_),
    .Y(_12269_));
 OAI21x1_ASAP7_75t_R _33372_ (.A1(net156),
    .A2(_12262_),
    .B(_12269_),
    .Y(_12270_));
 AO21x1_ASAP7_75t_R _33373_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01654_),
    .Y(_12271_));
 OAI22x1_ASAP7_75t_R _33374_ (.A1(_11999_),
    .A2(_12270_),
    .B1(_12271_),
    .B2(_12009_),
    .Y(_04013_));
 AND2x2_ASAP7_75t_R _33375_ (.A(_12252_),
    .B(_12002_),
    .Y(_12272_));
 AO21x1_ASAP7_75t_R _33376_ (.A1(_01618_),
    .A2(_12001_),
    .B(_12272_),
    .Y(_12273_));
 AO21x1_ASAP7_75t_R _33377_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01653_),
    .Y(_12274_));
 OAI22x1_ASAP7_75t_R _33378_ (.A1(_11999_),
    .A2(_12273_),
    .B1(_12274_),
    .B2(_12009_),
    .Y(_04014_));
 NAND2x1_ASAP7_75t_R _33379_ (.A(_01617_),
    .B(_12263_),
    .Y(_12275_));
 OAI21x1_ASAP7_75t_R _33380_ (.A1(net170),
    .A2(_12262_),
    .B(_12275_),
    .Y(_12276_));
 AO21x1_ASAP7_75t_R _33381_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01652_),
    .Y(_12277_));
 OAI22x1_ASAP7_75t_R _33382_ (.A1(_11999_),
    .A2(_12276_),
    .B1(_12277_),
    .B2(_12009_),
    .Y(_04015_));
 NAND2x1_ASAP7_75t_R _33383_ (.A(_01616_),
    .B(_12263_),
    .Y(_12278_));
 OAI21x1_ASAP7_75t_R _33384_ (.A1(net171),
    .A2(_12262_),
    .B(_12278_),
    .Y(_12279_));
 AO21x1_ASAP7_75t_R _33385_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01651_),
    .Y(_12280_));
 OAI22x1_ASAP7_75t_R _33386_ (.A1(_11999_),
    .A2(_12279_),
    .B1(_12280_),
    .B2(_12009_),
    .Y(_04016_));
 NAND2x1_ASAP7_75t_R _33387_ (.A(_01615_),
    .B(_12263_),
    .Y(_12281_));
 OAI21x1_ASAP7_75t_R _33388_ (.A1(net172),
    .A2(_12262_),
    .B(_12281_),
    .Y(_12282_));
 AO21x1_ASAP7_75t_R _33389_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01650_),
    .Y(_12283_));
 OAI22x1_ASAP7_75t_R _33390_ (.A1(_11999_),
    .A2(_12282_),
    .B1(_12283_),
    .B2(_12009_),
    .Y(_04017_));
 NAND2x1_ASAP7_75t_R _33391_ (.A(_01613_),
    .B(_12263_),
    .Y(_12284_));
 OAI21x1_ASAP7_75t_R _33392_ (.A1(net173),
    .A2(_12262_),
    .B(_12284_),
    .Y(_12285_));
 AO21x1_ASAP7_75t_R _33393_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01649_),
    .Y(_12286_));
 OAI22x1_ASAP7_75t_R _33394_ (.A1(_11999_),
    .A2(_12285_),
    .B1(_12286_),
    .B2(_12009_),
    .Y(_04018_));
 BUFx6f_ASAP7_75t_R _33395_ (.A(_12000_),
    .Y(_12287_));
 NAND2x1_ASAP7_75t_R _33396_ (.A(_01612_),
    .B(_12287_),
    .Y(_12288_));
 OAI21x1_ASAP7_75t_R _33397_ (.A1(net174),
    .A2(_12262_),
    .B(_12288_),
    .Y(_12289_));
 AO21x1_ASAP7_75t_R _33398_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01648_),
    .Y(_12290_));
 OAI22x1_ASAP7_75t_R _33399_ (.A1(_11999_),
    .A2(_12289_),
    .B1(_12290_),
    .B2(_12009_),
    .Y(_04019_));
 NOR2x1_ASAP7_75t_R _33400_ (.A(_01647_),
    .B(_12240_),
    .Y(_12291_));
 NAND2x1_ASAP7_75t_R _33401_ (.A(_11977_),
    .B(_01652_),
    .Y(_12292_));
 OA21x2_ASAP7_75t_R _33402_ (.A1(net170),
    .A2(_12182_),
    .B(_12292_),
    .Y(_12293_));
 AO32x1_ASAP7_75t_R _33403_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12291_),
    .B1(_12293_),
    .B2(_12244_),
    .Y(_04020_));
 NAND2x1_ASAP7_75t_R _33404_ (.A(_01611_),
    .B(_12287_),
    .Y(_12294_));
 OAI21x1_ASAP7_75t_R _33405_ (.A1(net175),
    .A2(_12262_),
    .B(_12294_),
    .Y(_12295_));
 AO21x1_ASAP7_75t_R _33406_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01646_),
    .Y(_12296_));
 OAI22x1_ASAP7_75t_R _33407_ (.A1(_11999_),
    .A2(_12295_),
    .B1(_12296_),
    .B2(_12009_),
    .Y(_04021_));
 BUFx6f_ASAP7_75t_R _33408_ (.A(_11998_),
    .Y(_12297_));
 NAND2x1_ASAP7_75t_R _33409_ (.A(_01610_),
    .B(_12287_),
    .Y(_12298_));
 OAI21x1_ASAP7_75t_R _33410_ (.A1(net176),
    .A2(_12262_),
    .B(_12298_),
    .Y(_12299_));
 AO21x1_ASAP7_75t_R _33411_ (.A1(_12266_),
    .A2(_12267_),
    .B(_01645_),
    .Y(_12300_));
 BUFx6f_ASAP7_75t_R _33412_ (.A(_12008_),
    .Y(_12301_));
 OAI22x1_ASAP7_75t_R _33413_ (.A1(_12297_),
    .A2(_12299_),
    .B1(_12300_),
    .B2(_12301_),
    .Y(_04022_));
 NAND2x1_ASAP7_75t_R _33414_ (.A(_01609_),
    .B(_12287_),
    .Y(_12302_));
 OAI21x1_ASAP7_75t_R _33415_ (.A1(net142),
    .A2(_12262_),
    .B(_12302_),
    .Y(_12303_));
 BUFx4f_ASAP7_75t_R _33416_ (.A(_12010_),
    .Y(_12304_));
 BUFx4f_ASAP7_75t_R _33417_ (.A(_11994_),
    .Y(_12305_));
 AO21x1_ASAP7_75t_R _33418_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01644_),
    .Y(_12306_));
 OAI22x1_ASAP7_75t_R _33419_ (.A1(_12297_),
    .A2(_12303_),
    .B1(_12306_),
    .B2(_12301_),
    .Y(_04023_));
 NAND2x1_ASAP7_75t_R _33420_ (.A(_01608_),
    .B(_12287_),
    .Y(_12307_));
 OAI21x1_ASAP7_75t_R _33421_ (.A1(net143),
    .A2(_12001_),
    .B(_12307_),
    .Y(_12308_));
 AO21x1_ASAP7_75t_R _33422_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01643_),
    .Y(_12309_));
 OAI22x1_ASAP7_75t_R _33423_ (.A1(_12297_),
    .A2(_12308_),
    .B1(_12309_),
    .B2(_12301_),
    .Y(_04024_));
 NAND2x1_ASAP7_75t_R _33424_ (.A(_01607_),
    .B(_12287_),
    .Y(_12310_));
 OAI21x1_ASAP7_75t_R _33425_ (.A1(net144),
    .A2(_12001_),
    .B(_12310_),
    .Y(_12311_));
 AO21x1_ASAP7_75t_R _33426_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01642_),
    .Y(_12312_));
 OAI22x1_ASAP7_75t_R _33427_ (.A1(_12297_),
    .A2(_12311_),
    .B1(_12312_),
    .B2(_12301_),
    .Y(_04025_));
 NAND2x1_ASAP7_75t_R _33428_ (.A(_01606_),
    .B(_12287_),
    .Y(_12313_));
 OAI21x1_ASAP7_75t_R _33429_ (.A1(net146),
    .A2(_12001_),
    .B(_12313_),
    .Y(_12314_));
 AO21x1_ASAP7_75t_R _33430_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01641_),
    .Y(_12315_));
 OAI22x1_ASAP7_75t_R _33431_ (.A1(_12297_),
    .A2(_12314_),
    .B1(_12315_),
    .B2(_12301_),
    .Y(_04026_));
 NAND2x1_ASAP7_75t_R _33432_ (.A(_01605_),
    .B(_12287_),
    .Y(_12316_));
 OAI21x1_ASAP7_75t_R _33433_ (.A1(net147),
    .A2(_12001_),
    .B(_12316_),
    .Y(_12317_));
 AO21x1_ASAP7_75t_R _33434_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01640_),
    .Y(_12318_));
 OAI22x1_ASAP7_75t_R _33435_ (.A1(_12297_),
    .A2(_12317_),
    .B1(_12318_),
    .B2(_12301_),
    .Y(_04027_));
 NAND2x1_ASAP7_75t_R _33436_ (.A(_01604_),
    .B(_12287_),
    .Y(_12319_));
 OAI21x1_ASAP7_75t_R _33437_ (.A1(net148),
    .A2(_12001_),
    .B(_12319_),
    .Y(_12320_));
 AO21x1_ASAP7_75t_R _33438_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01639_),
    .Y(_12321_));
 OAI22x1_ASAP7_75t_R _33439_ (.A1(_12297_),
    .A2(_12320_),
    .B1(_12321_),
    .B2(_12301_),
    .Y(_04028_));
 NAND2x1_ASAP7_75t_R _33440_ (.A(_01602_),
    .B(_12287_),
    .Y(_12322_));
 OAI21x1_ASAP7_75t_R _33441_ (.A1(net149),
    .A2(_12001_),
    .B(_12322_),
    .Y(_12323_));
 AO21x1_ASAP7_75t_R _33442_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01638_),
    .Y(_12324_));
 OAI22x1_ASAP7_75t_R _33443_ (.A1(_12297_),
    .A2(_12323_),
    .B1(_12324_),
    .B2(_12301_),
    .Y(_04029_));
 NAND2x1_ASAP7_75t_R _33444_ (.A(_01601_),
    .B(_12000_),
    .Y(_12325_));
 OAI21x1_ASAP7_75t_R _33445_ (.A1(net150),
    .A2(_12001_),
    .B(_12325_),
    .Y(_12326_));
 AO21x1_ASAP7_75t_R _33446_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01637_),
    .Y(_12327_));
 OAI22x1_ASAP7_75t_R _33447_ (.A1(_12297_),
    .A2(_12326_),
    .B1(_12327_),
    .B2(_12301_),
    .Y(_04030_));
 NOR2x1_ASAP7_75t_R _33448_ (.A(_01636_),
    .B(_12240_),
    .Y(_12328_));
 NAND2x1_ASAP7_75t_R _33449_ (.A(_11977_),
    .B(_01651_),
    .Y(_12329_));
 OA21x2_ASAP7_75t_R _33450_ (.A1(net171),
    .A2(_12182_),
    .B(_12329_),
    .Y(_12330_));
 AO32x1_ASAP7_75t_R _33451_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12328_),
    .B1(_12330_),
    .B2(_12244_),
    .Y(_04031_));
 INVx1_ASAP7_75t_R _33452_ (.A(net154),
    .Y(_12331_));
 AND2x2_ASAP7_75t_R _33453_ (.A(_12331_),
    .B(_12002_),
    .Y(_12332_));
 AO21x1_ASAP7_75t_R _33454_ (.A1(_01600_),
    .A2(_12001_),
    .B(_12332_),
    .Y(_12333_));
 AO21x1_ASAP7_75t_R _33455_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01635_),
    .Y(_12334_));
 OAI22x1_ASAP7_75t_R _33456_ (.A1(_12297_),
    .A2(_12333_),
    .B1(_12334_),
    .B2(_12301_),
    .Y(_04032_));
 BUFx6f_ASAP7_75t_R _33457_ (.A(_11998_),
    .Y(_12335_));
 BUFx4f_ASAP7_75t_R _33458_ (.A(_12000_),
    .Y(_12336_));
 INVx1_ASAP7_75t_R _33459_ (.A(net155),
    .Y(_12337_));
 AND2x2_ASAP7_75t_R _33460_ (.A(_12337_),
    .B(_12002_),
    .Y(_12338_));
 AO21x1_ASAP7_75t_R _33461_ (.A1(_01599_),
    .A2(_12336_),
    .B(_12338_),
    .Y(_12339_));
 AO21x1_ASAP7_75t_R _33462_ (.A1(_12304_),
    .A2(_12305_),
    .B(_01634_),
    .Y(_12340_));
 BUFx6f_ASAP7_75t_R _33463_ (.A(_12008_),
    .Y(_12341_));
 OAI22x1_ASAP7_75t_R _33464_ (.A1(_12335_),
    .A2(_12339_),
    .B1(_12340_),
    .B2(_12341_),
    .Y(_04033_));
 INVx1_ASAP7_75t_R _33465_ (.A(net157),
    .Y(_12342_));
 AND2x2_ASAP7_75t_R _33466_ (.A(_12342_),
    .B(_12002_),
    .Y(_12343_));
 AO21x1_ASAP7_75t_R _33467_ (.A1(_01598_),
    .A2(_12336_),
    .B(_12343_),
    .Y(_12344_));
 BUFx3_ASAP7_75t_R _33468_ (.A(_12010_),
    .Y(_12345_));
 BUFx3_ASAP7_75t_R _33469_ (.A(_11994_),
    .Y(_12346_));
 AO21x1_ASAP7_75t_R _33470_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01633_),
    .Y(_12347_));
 OAI22x1_ASAP7_75t_R _33471_ (.A1(_12335_),
    .A2(_12344_),
    .B1(_12347_),
    .B2(_12341_),
    .Y(_04034_));
 INVx1_ASAP7_75t_R _33472_ (.A(net158),
    .Y(_12348_));
 AND2x2_ASAP7_75t_R _33473_ (.A(_12348_),
    .B(_12002_),
    .Y(_12349_));
 AO21x1_ASAP7_75t_R _33474_ (.A1(_01597_),
    .A2(_12336_),
    .B(_12349_),
    .Y(_12350_));
 AO21x1_ASAP7_75t_R _33475_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01632_),
    .Y(_12351_));
 OAI22x1_ASAP7_75t_R _33476_ (.A1(_12335_),
    .A2(_12350_),
    .B1(_12351_),
    .B2(_12341_),
    .Y(_04035_));
 INVx1_ASAP7_75t_R _33477_ (.A(net159),
    .Y(_12352_));
 AND2x2_ASAP7_75t_R _33478_ (.A(_12352_),
    .B(_12002_),
    .Y(_12353_));
 AO21x1_ASAP7_75t_R _33479_ (.A1(_01596_),
    .A2(_12336_),
    .B(_12353_),
    .Y(_12354_));
 AO21x1_ASAP7_75t_R _33480_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01631_),
    .Y(_12355_));
 OAI22x1_ASAP7_75t_R _33481_ (.A1(_12335_),
    .A2(_12354_),
    .B1(_12355_),
    .B2(_12341_),
    .Y(_04036_));
 INVx1_ASAP7_75t_R _33482_ (.A(net160),
    .Y(_12356_));
 AND2x2_ASAP7_75t_R _33483_ (.A(_12356_),
    .B(_12002_),
    .Y(_12357_));
 AO21x1_ASAP7_75t_R _33484_ (.A1(_01595_),
    .A2(_12336_),
    .B(_12357_),
    .Y(_12358_));
 AO21x1_ASAP7_75t_R _33485_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01630_),
    .Y(_12359_));
 OAI22x1_ASAP7_75t_R _33486_ (.A1(_12335_),
    .A2(_12358_),
    .B1(_12359_),
    .B2(_12341_),
    .Y(_04037_));
 INVx1_ASAP7_75t_R _33487_ (.A(net161),
    .Y(_12360_));
 AND2x2_ASAP7_75t_R _33488_ (.A(_12360_),
    .B(_12002_),
    .Y(_12361_));
 AO21x1_ASAP7_75t_R _33489_ (.A1(_01594_),
    .A2(_12336_),
    .B(_12361_),
    .Y(_12362_));
 AO21x1_ASAP7_75t_R _33490_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01629_),
    .Y(_12363_));
 OAI22x1_ASAP7_75t_R _33491_ (.A1(_12335_),
    .A2(_12362_),
    .B1(_12363_),
    .B2(_12341_),
    .Y(_04038_));
 INVx1_ASAP7_75t_R _33492_ (.A(net162),
    .Y(_12364_));
 AND2x2_ASAP7_75t_R _33493_ (.A(_12364_),
    .B(_12002_),
    .Y(_12365_));
 AO21x1_ASAP7_75t_R _33494_ (.A1(_01593_),
    .A2(_12336_),
    .B(_12365_),
    .Y(_12366_));
 AO21x1_ASAP7_75t_R _33495_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01628_),
    .Y(_12367_));
 OAI22x1_ASAP7_75t_R _33496_ (.A1(_12335_),
    .A2(_12366_),
    .B1(_12367_),
    .B2(_12341_),
    .Y(_04039_));
 INVx1_ASAP7_75t_R _33497_ (.A(net163),
    .Y(_12368_));
 AND2x2_ASAP7_75t_R _33498_ (.A(_12368_),
    .B(_11992_),
    .Y(_12369_));
 AO21x1_ASAP7_75t_R _33499_ (.A1(_01591_),
    .A2(_12336_),
    .B(_12369_),
    .Y(_12370_));
 AO21x1_ASAP7_75t_R _33500_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01627_),
    .Y(_12371_));
 OAI22x1_ASAP7_75t_R _33501_ (.A1(_12335_),
    .A2(_12370_),
    .B1(_12371_),
    .B2(_12341_),
    .Y(_04040_));
 INVx1_ASAP7_75t_R _33502_ (.A(net164),
    .Y(_12372_));
 AND2x2_ASAP7_75t_R _33503_ (.A(_12372_),
    .B(_11992_),
    .Y(_12373_));
 AO21x1_ASAP7_75t_R _33504_ (.A1(_01590_),
    .A2(_12336_),
    .B(_12373_),
    .Y(_12374_));
 AO21x1_ASAP7_75t_R _33505_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01626_),
    .Y(_12375_));
 OAI22x1_ASAP7_75t_R _33506_ (.A1(_12335_),
    .A2(_12374_),
    .B1(_12375_),
    .B2(_12341_),
    .Y(_04041_));
 NOR2x1_ASAP7_75t_R _33507_ (.A(_01625_),
    .B(_12240_),
    .Y(_12376_));
 NAND2x1_ASAP7_75t_R _33508_ (.A(_11978_),
    .B(_01650_),
    .Y(_12377_));
 OA21x2_ASAP7_75t_R _33509_ (.A1(net172),
    .A2(_11978_),
    .B(_12377_),
    .Y(_12378_));
 AO32x1_ASAP7_75t_R _33510_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12376_),
    .B1(_12378_),
    .B2(_12244_),
    .Y(_04042_));
 INVx1_ASAP7_75t_R _33511_ (.A(net165),
    .Y(_12379_));
 AND2x2_ASAP7_75t_R _33512_ (.A(_12379_),
    .B(_11992_),
    .Y(_12380_));
 AO21x1_ASAP7_75t_R _33513_ (.A1(_01589_),
    .A2(_12336_),
    .B(_12380_),
    .Y(_12381_));
 AO21x1_ASAP7_75t_R _33514_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01624_),
    .Y(_12382_));
 OAI22x1_ASAP7_75t_R _33515_ (.A1(_12335_),
    .A2(_12381_),
    .B1(_12382_),
    .B2(_12341_),
    .Y(_04043_));
 INVx1_ASAP7_75t_R _33516_ (.A(net166),
    .Y(_12383_));
 AND2x2_ASAP7_75t_R _33517_ (.A(_12383_),
    .B(_11992_),
    .Y(_12384_));
 AO21x1_ASAP7_75t_R _33518_ (.A1(_01588_),
    .A2(_12263_),
    .B(_12384_),
    .Y(_12385_));
 AO21x1_ASAP7_75t_R _33519_ (.A1(_12345_),
    .A2(_12346_),
    .B(_01623_),
    .Y(_12386_));
 OAI22x1_ASAP7_75t_R _33520_ (.A1(_11998_),
    .A2(_12385_),
    .B1(_12386_),
    .B2(_12008_),
    .Y(_04044_));
 INVx1_ASAP7_75t_R _33521_ (.A(net168),
    .Y(_12387_));
 AND2x2_ASAP7_75t_R _33522_ (.A(_12387_),
    .B(_11992_),
    .Y(_12388_));
 AO21x1_ASAP7_75t_R _33523_ (.A1(_01587_),
    .A2(_12263_),
    .B(_12388_),
    .Y(_12389_));
 AO21x1_ASAP7_75t_R _33524_ (.A1(_12010_),
    .A2(_11994_),
    .B(_01622_),
    .Y(_12390_));
 OAI22x1_ASAP7_75t_R _33525_ (.A1(_11998_),
    .A2(_12389_),
    .B1(_12390_),
    .B2(_12008_),
    .Y(_04045_));
 INVx1_ASAP7_75t_R _33526_ (.A(net169),
    .Y(_12391_));
 AND2x2_ASAP7_75t_R _33527_ (.A(_12391_),
    .B(_11992_),
    .Y(_12392_));
 AO21x1_ASAP7_75t_R _33528_ (.A1(_01586_),
    .A2(_12263_),
    .B(_12392_),
    .Y(_12393_));
 AO21x1_ASAP7_75t_R _33529_ (.A1(_12010_),
    .A2(_11994_),
    .B(_01621_),
    .Y(_12394_));
 OAI22x1_ASAP7_75t_R _33530_ (.A1(_11998_),
    .A2(_12393_),
    .B1(_12394_),
    .B2(_12008_),
    .Y(_04046_));
 NAND2x1_ASAP7_75t_R _33531_ (.A(_01620_),
    .B(_12015_),
    .Y(_12395_));
 OA21x2_ASAP7_75t_R _33532_ (.A1(net141),
    .A2(_12014_),
    .B(_12395_),
    .Y(_04047_));
 NAND2x1_ASAP7_75t_R _33533_ (.A(_01619_),
    .B(_12015_),
    .Y(_12396_));
 OA21x2_ASAP7_75t_R _33534_ (.A1(net156),
    .A2(_12014_),
    .B(_12396_),
    .Y(_04048_));
 NAND2x1_ASAP7_75t_R _33535_ (.A(_01618_),
    .B(_12015_),
    .Y(_12397_));
 OA21x2_ASAP7_75t_R _33536_ (.A1(net167),
    .A2(_12014_),
    .B(_12397_),
    .Y(_04049_));
 NAND2x1_ASAP7_75t_R _33537_ (.A(_01617_),
    .B(_12015_),
    .Y(_12398_));
 OA21x2_ASAP7_75t_R _33538_ (.A1(net170),
    .A2(_12014_),
    .B(_12398_),
    .Y(_04050_));
 NAND2x1_ASAP7_75t_R _33539_ (.A(_01616_),
    .B(_12015_),
    .Y(_12399_));
 OA21x2_ASAP7_75t_R _33540_ (.A1(net171),
    .A2(_12014_),
    .B(_12399_),
    .Y(_04051_));
 NAND2x1_ASAP7_75t_R _33541_ (.A(_01615_),
    .B(_12015_),
    .Y(_12400_));
 OA21x2_ASAP7_75t_R _33542_ (.A1(net172),
    .A2(_12014_),
    .B(_12400_),
    .Y(_04052_));
 NOR2x1_ASAP7_75t_R _33543_ (.A(_01614_),
    .B(_12240_),
    .Y(_12401_));
 NAND2x1_ASAP7_75t_R _33544_ (.A(_11978_),
    .B(_01649_),
    .Y(_12402_));
 OA21x2_ASAP7_75t_R _33545_ (.A1(net173),
    .A2(_11978_),
    .B(_12402_),
    .Y(_12403_));
 AO32x1_ASAP7_75t_R _33546_ (.A1(_12238_),
    .A2(_12239_),
    .A3(_12401_),
    .B1(_12403_),
    .B2(_12244_),
    .Y(_04053_));
 BUFx6f_ASAP7_75t_R _33547_ (.A(_12013_),
    .Y(_12404_));
 NAND2x1_ASAP7_75t_R _33548_ (.A(_01613_),
    .B(_12404_),
    .Y(_12405_));
 OA21x2_ASAP7_75t_R _33549_ (.A1(net173),
    .A2(_12014_),
    .B(_12405_),
    .Y(_04054_));
 NAND2x1_ASAP7_75t_R _33550_ (.A(_01612_),
    .B(_12404_),
    .Y(_12406_));
 OA21x2_ASAP7_75t_R _33551_ (.A1(net174),
    .A2(_12014_),
    .B(_12406_),
    .Y(_04055_));
 NAND2x1_ASAP7_75t_R _33552_ (.A(_01611_),
    .B(_12404_),
    .Y(_12407_));
 OA21x2_ASAP7_75t_R _33553_ (.A1(net175),
    .A2(_12014_),
    .B(_12407_),
    .Y(_04056_));
 BUFx4f_ASAP7_75t_R _33554_ (.A(_12013_),
    .Y(_12408_));
 NAND2x1_ASAP7_75t_R _33555_ (.A(_01610_),
    .B(_12404_),
    .Y(_12409_));
 OA21x2_ASAP7_75t_R _33556_ (.A1(net176),
    .A2(_12408_),
    .B(_12409_),
    .Y(_04057_));
 NAND2x1_ASAP7_75t_R _33557_ (.A(_01609_),
    .B(_12404_),
    .Y(_12410_));
 OA21x2_ASAP7_75t_R _33558_ (.A1(net142),
    .A2(_12408_),
    .B(_12410_),
    .Y(_04058_));
 NAND2x1_ASAP7_75t_R _33559_ (.A(_01608_),
    .B(_12404_),
    .Y(_12411_));
 OA21x2_ASAP7_75t_R _33560_ (.A1(net143),
    .A2(_12408_),
    .B(_12411_),
    .Y(_04059_));
 NAND2x1_ASAP7_75t_R _33561_ (.A(_01607_),
    .B(_12404_),
    .Y(_12412_));
 OA21x2_ASAP7_75t_R _33562_ (.A1(net144),
    .A2(_12408_),
    .B(_12412_),
    .Y(_04060_));
 NAND2x1_ASAP7_75t_R _33563_ (.A(_01606_),
    .B(_12404_),
    .Y(_12413_));
 OA21x2_ASAP7_75t_R _33564_ (.A1(net146),
    .A2(_12408_),
    .B(_12413_),
    .Y(_04061_));
 NAND2x1_ASAP7_75t_R _33565_ (.A(_01605_),
    .B(_12404_),
    .Y(_12414_));
 OA21x2_ASAP7_75t_R _33566_ (.A1(net147),
    .A2(_12408_),
    .B(_12414_),
    .Y(_04062_));
 NAND2x1_ASAP7_75t_R _33567_ (.A(_01604_),
    .B(_12404_),
    .Y(_12415_));
 OA21x2_ASAP7_75t_R _33568_ (.A1(net148),
    .A2(_12408_),
    .B(_12415_),
    .Y(_04063_));
 NOR2x1_ASAP7_75t_R _33569_ (.A(_01603_),
    .B(_11974_),
    .Y(_12416_));
 NAND2x1_ASAP7_75t_R _33570_ (.A(_11977_),
    .B(_01648_),
    .Y(_12417_));
 OA21x2_ASAP7_75t_R _33571_ (.A1(net174),
    .A2(_12182_),
    .B(_12417_),
    .Y(_12418_));
 AO32x1_ASAP7_75t_R _33572_ (.A1(_11969_),
    .A2(_11972_),
    .A3(_12416_),
    .B1(_12418_),
    .B2(_11987_),
    .Y(_04064_));
 BUFx6f_ASAP7_75t_R _33573_ (.A(_12012_),
    .Y(_12419_));
 NAND2x1_ASAP7_75t_R _33574_ (.A(_01602_),
    .B(_12419_),
    .Y(_12420_));
 OA21x2_ASAP7_75t_R _33575_ (.A1(net149),
    .A2(_12408_),
    .B(_12420_),
    .Y(_04065_));
 NAND2x1_ASAP7_75t_R _33576_ (.A(_01601_),
    .B(_12419_),
    .Y(_12421_));
 OA21x2_ASAP7_75t_R _33577_ (.A1(net150),
    .A2(_12408_),
    .B(_12421_),
    .Y(_04066_));
 NAND2x1_ASAP7_75t_R _33578_ (.A(_01600_),
    .B(_12419_),
    .Y(_12422_));
 OA21x2_ASAP7_75t_R _33579_ (.A1(net154),
    .A2(_12408_),
    .B(_12422_),
    .Y(_04067_));
 BUFx3_ASAP7_75t_R _33580_ (.A(_12013_),
    .Y(_12423_));
 NAND2x1_ASAP7_75t_R _33581_ (.A(_01599_),
    .B(_12419_),
    .Y(_12424_));
 OA21x2_ASAP7_75t_R _33582_ (.A1(net155),
    .A2(_12423_),
    .B(_12424_),
    .Y(_04068_));
 NAND2x1_ASAP7_75t_R _33583_ (.A(_01598_),
    .B(_12419_),
    .Y(_12425_));
 OA21x2_ASAP7_75t_R _33584_ (.A1(net157),
    .A2(_12423_),
    .B(_12425_),
    .Y(_04069_));
 NAND2x1_ASAP7_75t_R _33585_ (.A(_01597_),
    .B(_12419_),
    .Y(_12426_));
 OA21x2_ASAP7_75t_R _33586_ (.A1(net158),
    .A2(_12423_),
    .B(_12426_),
    .Y(_04070_));
 NAND2x1_ASAP7_75t_R _33587_ (.A(_01596_),
    .B(_12419_),
    .Y(_12427_));
 OA21x2_ASAP7_75t_R _33588_ (.A1(net159),
    .A2(_12423_),
    .B(_12427_),
    .Y(_04071_));
 NAND2x1_ASAP7_75t_R _33589_ (.A(_01595_),
    .B(_12419_),
    .Y(_12428_));
 OA21x2_ASAP7_75t_R _33590_ (.A1(net160),
    .A2(_12423_),
    .B(_12428_),
    .Y(_04072_));
 NAND2x1_ASAP7_75t_R _33591_ (.A(_01594_),
    .B(_12419_),
    .Y(_12429_));
 OA21x2_ASAP7_75t_R _33592_ (.A1(net161),
    .A2(_12423_),
    .B(_12429_),
    .Y(_04073_));
 NAND2x1_ASAP7_75t_R _33593_ (.A(_01593_),
    .B(_12419_),
    .Y(_12430_));
 OA21x2_ASAP7_75t_R _33594_ (.A1(net162),
    .A2(_12423_),
    .B(_12430_),
    .Y(_04074_));
 NOR2x1_ASAP7_75t_R _33595_ (.A(_01592_),
    .B(_11974_),
    .Y(_12431_));
 NAND2x1_ASAP7_75t_R _33596_ (.A(_11949_),
    .B(_01646_),
    .Y(_12432_));
 OA21x2_ASAP7_75t_R _33597_ (.A1(net175),
    .A2(_11949_),
    .B(_12432_),
    .Y(_12433_));
 AO32x1_ASAP7_75t_R _33598_ (.A1(_11969_),
    .A2(_11972_),
    .A3(_12431_),
    .B1(_12433_),
    .B2(_11987_),
    .Y(_04075_));
 NAND2x1_ASAP7_75t_R _33599_ (.A(_01591_),
    .B(_12013_),
    .Y(_12434_));
 OA21x2_ASAP7_75t_R _33600_ (.A1(net163),
    .A2(_12423_),
    .B(_12434_),
    .Y(_04076_));
 NAND2x1_ASAP7_75t_R _33601_ (.A(_01590_),
    .B(_12013_),
    .Y(_12435_));
 OA21x2_ASAP7_75t_R _33602_ (.A1(net164),
    .A2(_12423_),
    .B(_12435_),
    .Y(_04077_));
 NAND2x1_ASAP7_75t_R _33603_ (.A(_01589_),
    .B(_12013_),
    .Y(_12436_));
 OA21x2_ASAP7_75t_R _33604_ (.A1(net165),
    .A2(_12423_),
    .B(_12436_),
    .Y(_04078_));
 NAND2x1_ASAP7_75t_R _33605_ (.A(_01588_),
    .B(_12013_),
    .Y(_12437_));
 OA21x2_ASAP7_75t_R _33606_ (.A1(net166),
    .A2(_12015_),
    .B(_12437_),
    .Y(_04079_));
 NAND2x1_ASAP7_75t_R _33607_ (.A(_01587_),
    .B(_12013_),
    .Y(_12438_));
 OA21x2_ASAP7_75t_R _33608_ (.A1(net168),
    .A2(_12015_),
    .B(_12438_),
    .Y(_04080_));
 NAND2x1_ASAP7_75t_R _33609_ (.A(_01586_),
    .B(_12013_),
    .Y(_12439_));
 OA21x2_ASAP7_75t_R _33610_ (.A1(net169),
    .A2(_12015_),
    .B(_12439_),
    .Y(_04081_));
 NOR2x1_ASAP7_75t_R _33611_ (.A(_02225_),
    .B(_11974_),
    .Y(_12440_));
 NAND2x1_ASAP7_75t_R _33612_ (.A(_12182_),
    .B(_01645_),
    .Y(_12441_));
 OA21x2_ASAP7_75t_R _33613_ (.A1(net176),
    .A2(_12182_),
    .B(_12441_),
    .Y(_12442_));
 AO32x1_ASAP7_75t_R _33614_ (.A1(_11969_),
    .A2(_11972_),
    .A3(_12440_),
    .B1(_12442_),
    .B2(_11987_),
    .Y(_04082_));
 BUFx4f_ASAP7_75t_R _33615_ (.A(_05469_),
    .Y(_12443_));
 BUFx6f_ASAP7_75t_R _33616_ (.A(_05469_),
    .Y(_12444_));
 NOR2x1_ASAP7_75t_R _33617_ (.A(_12444_),
    .B(_01585_),
    .Y(_12445_));
 AO21x1_ASAP7_75t_R _33618_ (.A1(_12443_),
    .A2(_11698_),
    .B(_12445_),
    .Y(net268));
 OR3x1_ASAP7_75t_R _33619_ (.A(_05507_),
    .B(net140),
    .C(_05512_),
    .Y(_12446_));
 BUFx4f_ASAP7_75t_R _33620_ (.A(_12446_),
    .Y(_12447_));
 BUFx4f_ASAP7_75t_R _33621_ (.A(_12447_),
    .Y(_12448_));
 NAND2x1_ASAP7_75t_R _33622_ (.A(_01585_),
    .B(_12448_),
    .Y(_12449_));
 OA21x2_ASAP7_75t_R _33623_ (.A1(net268),
    .A2(_12448_),
    .B(_12449_),
    .Y(_04083_));
 NOR2x1_ASAP7_75t_R _33624_ (.A(_12444_),
    .B(_01584_),
    .Y(_12450_));
 AO21x1_ASAP7_75t_R _33625_ (.A1(_12443_),
    .A2(_11678_),
    .B(_12450_),
    .Y(net269));
 BUFx4f_ASAP7_75t_R _33626_ (.A(_12447_),
    .Y(_12451_));
 NAND2x1_ASAP7_75t_R _33627_ (.A(_01584_),
    .B(_12448_),
    .Y(_12452_));
 OA21x2_ASAP7_75t_R _33628_ (.A1(_12451_),
    .A2(net269),
    .B(_12452_),
    .Y(_04084_));
 NOR2x1_ASAP7_75t_R _33629_ (.A(_12444_),
    .B(_01583_),
    .Y(_12453_));
 AO21x1_ASAP7_75t_R _33630_ (.A1(_12443_),
    .A2(_11745_),
    .B(_12453_),
    .Y(net270));
 NAND2x1_ASAP7_75t_R _33631_ (.A(_01583_),
    .B(_12448_),
    .Y(_12454_));
 OA21x2_ASAP7_75t_R _33632_ (.A1(_12451_),
    .A2(net270),
    .B(_12454_),
    .Y(_04085_));
 NOR2x1_ASAP7_75t_R _33633_ (.A(_12444_),
    .B(_01582_),
    .Y(_12455_));
 AO21x1_ASAP7_75t_R _33634_ (.A1(_05470_),
    .A2(_11746_),
    .B(_12455_),
    .Y(net271));
 BUFx6f_ASAP7_75t_R _33635_ (.A(_12447_),
    .Y(_12456_));
 NAND2x1_ASAP7_75t_R _33636_ (.A(_01582_),
    .B(_12456_),
    .Y(_12457_));
 OA21x2_ASAP7_75t_R _33637_ (.A1(_12451_),
    .A2(net271),
    .B(_12457_),
    .Y(_04086_));
 NOR2x1_ASAP7_75t_R _33638_ (.A(_12444_),
    .B(_01581_),
    .Y(_12458_));
 AO21x1_ASAP7_75t_R _33639_ (.A1(_05470_),
    .A2(_11721_),
    .B(_12458_),
    .Y(net272));
 NAND2x1_ASAP7_75t_R _33640_ (.A(_01581_),
    .B(_12456_),
    .Y(_12459_));
 OA21x2_ASAP7_75t_R _33641_ (.A1(_12451_),
    .A2(net272),
    .B(_12459_),
    .Y(_04087_));
 NOR2x1_ASAP7_75t_R _33642_ (.A(_12444_),
    .B(_01580_),
    .Y(_12460_));
 AO21x1_ASAP7_75t_R _33643_ (.A1(_05470_),
    .A2(_11749_),
    .B(_12460_),
    .Y(net273));
 NAND2x1_ASAP7_75t_R _33644_ (.A(_01580_),
    .B(_12456_),
    .Y(_12461_));
 OA21x2_ASAP7_75t_R _33645_ (.A1(_12451_),
    .A2(net273),
    .B(_12461_),
    .Y(_04088_));
 NOR2x1_ASAP7_75t_R _33646_ (.A(_12444_),
    .B(_01579_),
    .Y(_12462_));
 AO21x1_ASAP7_75t_R _33647_ (.A1(_05470_),
    .A2(_11744_),
    .B(_12462_),
    .Y(net274));
 NAND2x1_ASAP7_75t_R _33648_ (.A(_01579_),
    .B(_12456_),
    .Y(_12463_));
 OA21x2_ASAP7_75t_R _33649_ (.A1(_12451_),
    .A2(net274),
    .B(_12463_),
    .Y(_04089_));
 BUFx6f_ASAP7_75t_R _33650_ (.A(_05469_),
    .Y(_12464_));
 INVx1_ASAP7_75t_R _33651_ (.A(_01578_),
    .Y(_12465_));
 BUFx6f_ASAP7_75t_R _33652_ (.A(_05469_),
    .Y(_12466_));
 NAND2x1_ASAP7_75t_R _33653_ (.A(_12466_),
    .B(_11758_),
    .Y(_12467_));
 OA21x2_ASAP7_75t_R _33654_ (.A1(_12464_),
    .A2(_12465_),
    .B(_12467_),
    .Y(net275));
 INVx1_ASAP7_75t_R _33655_ (.A(net140),
    .Y(_12468_));
 AND2x2_ASAP7_75t_R _33656_ (.A(_12468_),
    .B(_18773_),
    .Y(_12469_));
 BUFx3_ASAP7_75t_R _33657_ (.A(_12469_),
    .Y(_12470_));
 BUFx4f_ASAP7_75t_R _33658_ (.A(_12447_),
    .Y(_12471_));
 AND2x2_ASAP7_75t_R _33659_ (.A(_12465_),
    .B(_12471_),
    .Y(_12472_));
 AO21x1_ASAP7_75t_R _33660_ (.A1(_12470_),
    .A2(net275),
    .B(_12472_),
    .Y(_04090_));
 AND2x2_ASAP7_75t_R _33661_ (.A(_05507_),
    .B(_01577_),
    .Y(_12473_));
 AOI21x1_ASAP7_75t_R _33662_ (.A1(_12464_),
    .A2(_11766_),
    .B(_12473_),
    .Y(net276));
 NAND2x1_ASAP7_75t_R _33663_ (.A(_01577_),
    .B(_12456_),
    .Y(_12474_));
 OA21x2_ASAP7_75t_R _33664_ (.A1(_12451_),
    .A2(net276),
    .B(_12474_),
    .Y(_04091_));
 INVx1_ASAP7_75t_R _33665_ (.A(_01576_),
    .Y(_12475_));
 NAND2x1_ASAP7_75t_R _33666_ (.A(_12466_),
    .B(_11779_),
    .Y(_12476_));
 OA21x2_ASAP7_75t_R _33667_ (.A1(_12464_),
    .A2(_12475_),
    .B(_12476_),
    .Y(net277));
 AND2x2_ASAP7_75t_R _33668_ (.A(_12475_),
    .B(_12471_),
    .Y(_12477_));
 AO21x1_ASAP7_75t_R _33669_ (.A1(_12470_),
    .A2(net277),
    .B(_12477_),
    .Y(_04092_));
 NOR2x1_ASAP7_75t_R _33670_ (.A(_12444_),
    .B(_01575_),
    .Y(_12478_));
 AO21x1_ASAP7_75t_R _33671_ (.A1(_05470_),
    .A2(_11792_),
    .B(_12478_),
    .Y(net278));
 NAND2x1_ASAP7_75t_R _33672_ (.A(_01575_),
    .B(_12456_),
    .Y(_12479_));
 OA21x2_ASAP7_75t_R _33673_ (.A1(_12451_),
    .A2(net278),
    .B(_12479_),
    .Y(_04093_));
 NOR2x1_ASAP7_75t_R _33674_ (.A(_05469_),
    .B(_01574_),
    .Y(_12480_));
 AO21x1_ASAP7_75t_R _33675_ (.A1(_05470_),
    .A2(_11813_),
    .B(_12480_),
    .Y(net279));
 NAND2x1_ASAP7_75t_R _33676_ (.A(_01574_),
    .B(_12456_),
    .Y(_12481_));
 OA21x2_ASAP7_75t_R _33677_ (.A1(_12451_),
    .A2(net279),
    .B(_12481_),
    .Y(_04094_));
 NOR2x1_ASAP7_75t_R _33678_ (.A(_05469_),
    .B(_01573_),
    .Y(_12482_));
 AO21x1_ASAP7_75t_R _33679_ (.A1(_05470_),
    .A2(_11811_),
    .B(_12482_),
    .Y(net280));
 NAND2x1_ASAP7_75t_R _33680_ (.A(_01573_),
    .B(_12456_),
    .Y(_12483_));
 OA21x2_ASAP7_75t_R _33681_ (.A1(_12451_),
    .A2(net280),
    .B(_12483_),
    .Y(_04095_));
 NOR2x1_ASAP7_75t_R _33682_ (.A(_05469_),
    .B(_01572_),
    .Y(_12484_));
 AO21x1_ASAP7_75t_R _33683_ (.A1(_05470_),
    .A2(_11822_),
    .B(_12484_),
    .Y(net281));
 NAND2x1_ASAP7_75t_R _33684_ (.A(_01572_),
    .B(_12456_),
    .Y(_12485_));
 OA21x2_ASAP7_75t_R _33685_ (.A1(_12448_),
    .A2(net281),
    .B(_12485_),
    .Y(_04096_));
 NOR2x1_ASAP7_75t_R _33686_ (.A(_05469_),
    .B(_01571_),
    .Y(_12486_));
 AO21x1_ASAP7_75t_R _33687_ (.A1(_05470_),
    .A2(_11844_),
    .B(_12486_),
    .Y(net282));
 NAND2x1_ASAP7_75t_R _33688_ (.A(_01571_),
    .B(_12456_),
    .Y(_12487_));
 OA21x2_ASAP7_75t_R _33689_ (.A1(_12448_),
    .A2(net282),
    .B(_12487_),
    .Y(_04097_));
 NAND2x1_ASAP7_75t_R _33690_ (.A(_05507_),
    .B(_01570_),
    .Y(_12488_));
 OA21x2_ASAP7_75t_R _33691_ (.A1(_05507_),
    .A2(_11854_),
    .B(_12488_),
    .Y(net283));
 NAND2x1_ASAP7_75t_R _33692_ (.A(_01570_),
    .B(_12471_),
    .Y(_12489_));
 OA21x2_ASAP7_75t_R _33693_ (.A1(_12448_),
    .A2(net283),
    .B(_12489_),
    .Y(_04098_));
 INVx1_ASAP7_75t_R _33694_ (.A(_01569_),
    .Y(_12490_));
 NAND2x1_ASAP7_75t_R _33695_ (.A(_12466_),
    .B(_11853_),
    .Y(_12491_));
 OA21x2_ASAP7_75t_R _33696_ (.A1(_12464_),
    .A2(_12490_),
    .B(_12491_),
    .Y(net284));
 AND2x2_ASAP7_75t_R _33697_ (.A(_12490_),
    .B(_12471_),
    .Y(_12492_));
 AO21x1_ASAP7_75t_R _33698_ (.A1(_12470_),
    .A2(net284),
    .B(_12492_),
    .Y(_04099_));
 INVx1_ASAP7_75t_R _33699_ (.A(_01568_),
    .Y(_12493_));
 NAND2x1_ASAP7_75t_R _33700_ (.A(_12466_),
    .B(_11867_),
    .Y(_12494_));
 OA21x2_ASAP7_75t_R _33701_ (.A1(_12464_),
    .A2(_12493_),
    .B(_12494_),
    .Y(net285));
 AND2x2_ASAP7_75t_R _33702_ (.A(_12493_),
    .B(_12471_),
    .Y(_12495_));
 AO21x1_ASAP7_75t_R _33703_ (.A1(_12470_),
    .A2(net285),
    .B(_12495_),
    .Y(_04100_));
 INVx1_ASAP7_75t_R _33704_ (.A(_01567_),
    .Y(_12496_));
 NAND2x1_ASAP7_75t_R _33705_ (.A(_12466_),
    .B(_11877_),
    .Y(_12497_));
 OA21x2_ASAP7_75t_R _33706_ (.A1(_12464_),
    .A2(_12496_),
    .B(_12497_),
    .Y(net286));
 AND2x2_ASAP7_75t_R _33707_ (.A(_12496_),
    .B(_12471_),
    .Y(_12498_));
 AO21x1_ASAP7_75t_R _33708_ (.A1(_12470_),
    .A2(net286),
    .B(_12498_),
    .Y(_04101_));
 INVx1_ASAP7_75t_R _33709_ (.A(_01566_),
    .Y(_12499_));
 NAND2x1_ASAP7_75t_R _33710_ (.A(_12466_),
    .B(_11885_),
    .Y(_12500_));
 OA21x2_ASAP7_75t_R _33711_ (.A1(_12443_),
    .A2(_12499_),
    .B(_12500_),
    .Y(net287));
 AND2x2_ASAP7_75t_R _33712_ (.A(_12499_),
    .B(_12471_),
    .Y(_12501_));
 AO21x1_ASAP7_75t_R _33713_ (.A1(_12470_),
    .A2(net287),
    .B(_12501_),
    .Y(_04102_));
 AND2x2_ASAP7_75t_R _33714_ (.A(_05507_),
    .B(_01565_),
    .Y(_12502_));
 AOI21x1_ASAP7_75t_R _33715_ (.A1(_12464_),
    .A2(_05435_),
    .B(_12502_),
    .Y(net288));
 NOR2x1_ASAP7_75t_R _33716_ (.A(_01565_),
    .B(_12469_),
    .Y(_12503_));
 AO21x1_ASAP7_75t_R _33717_ (.A1(_12470_),
    .A2(net288),
    .B(_12503_),
    .Y(_04103_));
 INVx1_ASAP7_75t_R _33718_ (.A(_01564_),
    .Y(_12504_));
 NAND2x1_ASAP7_75t_R _33719_ (.A(_12466_),
    .B(_11896_),
    .Y(_12505_));
 OA21x2_ASAP7_75t_R _33720_ (.A1(_12443_),
    .A2(_12504_),
    .B(_12505_),
    .Y(net289));
 AND2x2_ASAP7_75t_R _33721_ (.A(_12504_),
    .B(_12447_),
    .Y(_12506_));
 AO21x1_ASAP7_75t_R _33722_ (.A1(_12470_),
    .A2(net289),
    .B(_12506_),
    .Y(_04104_));
 INVx1_ASAP7_75t_R _33723_ (.A(_01563_),
    .Y(_12507_));
 NAND2x1_ASAP7_75t_R _33724_ (.A(_11904_),
    .B(_12466_),
    .Y(_12508_));
 OA21x2_ASAP7_75t_R _33725_ (.A1(_12443_),
    .A2(_12507_),
    .B(_12508_),
    .Y(net290));
 AND2x2_ASAP7_75t_R _33726_ (.A(_12507_),
    .B(_12447_),
    .Y(_12509_));
 AO21x1_ASAP7_75t_R _33727_ (.A1(_12470_),
    .A2(net290),
    .B(_12509_),
    .Y(_04105_));
 INVx1_ASAP7_75t_R _33728_ (.A(_01562_),
    .Y(_12510_));
 NAND2x1_ASAP7_75t_R _33729_ (.A(_12466_),
    .B(_05464_),
    .Y(_12511_));
 OA21x2_ASAP7_75t_R _33730_ (.A1(_12443_),
    .A2(_12510_),
    .B(_12511_),
    .Y(net291));
 AND2x2_ASAP7_75t_R _33731_ (.A(_12510_),
    .B(_12447_),
    .Y(_12512_));
 AO21x1_ASAP7_75t_R _33732_ (.A1(_12470_),
    .A2(net291),
    .B(_12512_),
    .Y(_04106_));
 INVx1_ASAP7_75t_R _33733_ (.A(_01561_),
    .Y(_12513_));
 NAND2x1_ASAP7_75t_R _33734_ (.A(_12466_),
    .B(_11641_),
    .Y(_12514_));
 OA21x2_ASAP7_75t_R _33735_ (.A1(_12443_),
    .A2(_12513_),
    .B(_12514_),
    .Y(net292));
 AND2x2_ASAP7_75t_R _33736_ (.A(_12513_),
    .B(_12447_),
    .Y(_12515_));
 AO21x1_ASAP7_75t_R _33737_ (.A1(_12469_),
    .A2(net292),
    .B(_12515_),
    .Y(_04107_));
 INVx1_ASAP7_75t_R _33738_ (.A(_01560_),
    .Y(_12516_));
 NAND2x1_ASAP7_75t_R _33739_ (.A(_12444_),
    .B(_11646_),
    .Y(_12517_));
 OA21x2_ASAP7_75t_R _33740_ (.A1(_12443_),
    .A2(_12516_),
    .B(_12517_),
    .Y(net293));
 AND2x2_ASAP7_75t_R _33741_ (.A(_12516_),
    .B(_12447_),
    .Y(_12518_));
 AO21x1_ASAP7_75t_R _33742_ (.A1(_12469_),
    .A2(net293),
    .B(_12518_),
    .Y(_04108_));
 INVx1_ASAP7_75t_R _33743_ (.A(_01559_),
    .Y(_12519_));
 NAND2x1_ASAP7_75t_R _33744_ (.A(_12444_),
    .B(_11637_),
    .Y(_12520_));
 OA21x2_ASAP7_75t_R _33745_ (.A1(_12443_),
    .A2(_12519_),
    .B(_12520_),
    .Y(net294));
 AND2x2_ASAP7_75t_R _33746_ (.A(_12519_),
    .B(_12447_),
    .Y(_12521_));
 AO21x1_ASAP7_75t_R _33747_ (.A1(_12469_),
    .A2(net294),
    .B(_12521_),
    .Y(_04109_));
 AND2x2_ASAP7_75t_R _33748_ (.A(_05507_),
    .B(_01558_),
    .Y(_12522_));
 AOI21x1_ASAP7_75t_R _33749_ (.A1(_12464_),
    .A2(_11924_),
    .B(_12522_),
    .Y(net295));
 NAND2x1_ASAP7_75t_R _33750_ (.A(_01558_),
    .B(_12471_),
    .Y(_12523_));
 OA21x2_ASAP7_75t_R _33751_ (.A1(_12448_),
    .A2(net295),
    .B(_12523_),
    .Y(_04110_));
 AND2x2_ASAP7_75t_R _33752_ (.A(_05507_),
    .B(_01557_),
    .Y(_12524_));
 AOI21x1_ASAP7_75t_R _33753_ (.A1(_12464_),
    .A2(_11932_),
    .B(_12524_),
    .Y(net296));
 NAND2x1_ASAP7_75t_R _33754_ (.A(_01557_),
    .B(_12471_),
    .Y(_12525_));
 OA21x2_ASAP7_75t_R _33755_ (.A1(_12448_),
    .A2(net296),
    .B(_12525_),
    .Y(_04111_));
 AND2x2_ASAP7_75t_R _33756_ (.A(_05507_),
    .B(_02228_),
    .Y(_12526_));
 AOI21x1_ASAP7_75t_R _33757_ (.A1(_12464_),
    .A2(_11931_),
    .B(_12526_),
    .Y(net297));
 NAND2x1_ASAP7_75t_R _33758_ (.A(_02228_),
    .B(_12471_),
    .Y(_12527_));
 OA21x2_ASAP7_75t_R _33759_ (.A1(_12448_),
    .A2(net297),
    .B(_12527_),
    .Y(_04112_));
 OA21x2_ASAP7_75t_R _33760_ (.A1(_13362_),
    .A2(_05754_),
    .B(_05752_),
    .Y(_12528_));
 AO21x1_ASAP7_75t_R _33761_ (.A1(_01508_),
    .A2(_13358_),
    .B(_13359_),
    .Y(_12529_));
 OA211x2_ASAP7_75t_R _33762_ (.A1(_05751_),
    .A2(_13359_),
    .B(_13357_),
    .C(net104),
    .Y(_12530_));
 AO22x1_ASAP7_75t_R _33763_ (.A1(_05751_),
    .A2(_12529_),
    .B1(_12530_),
    .B2(_04920_),
    .Y(_12531_));
 OAI21x1_ASAP7_75t_R _33764_ (.A1(_13360_),
    .A2(_12528_),
    .B(_12531_),
    .Y(_12532_));
 BUFx6f_ASAP7_75t_R _33765_ (.A(_12532_),
    .Y(_12533_));
 BUFx6f_ASAP7_75t_R _33766_ (.A(_12532_),
    .Y(_12534_));
 NAND2x1_ASAP7_75t_R _33767_ (.A(_01543_),
    .B(_12534_),
    .Y(_12535_));
 OA21x2_ASAP7_75t_R _33768_ (.A1(\alu_adder_result_ex[0] ),
    .A2(_12533_),
    .B(_12535_),
    .Y(_04196_));
 NAND2x1_ASAP7_75t_R _33769_ (.A(_01542_),
    .B(_12534_),
    .Y(_12536_));
 OA21x2_ASAP7_75t_R _33770_ (.A1(\alu_adder_result_ex[10] ),
    .A2(_12533_),
    .B(_12536_),
    .Y(_04197_));
 NAND2x1_ASAP7_75t_R _33771_ (.A(_01541_),
    .B(_12534_),
    .Y(_12537_));
 OA21x2_ASAP7_75t_R _33772_ (.A1(\alu_adder_result_ex[11] ),
    .A2(_12533_),
    .B(_12537_),
    .Y(_04198_));
 NAND2x1_ASAP7_75t_R _33773_ (.A(_01540_),
    .B(_12534_),
    .Y(_12538_));
 OA21x2_ASAP7_75t_R _33774_ (.A1(\alu_adder_result_ex[12] ),
    .A2(_12533_),
    .B(_12538_),
    .Y(_04199_));
 NAND2x1_ASAP7_75t_R _33775_ (.A(_01539_),
    .B(_12534_),
    .Y(_12539_));
 OA21x2_ASAP7_75t_R _33776_ (.A1(\alu_adder_result_ex[13] ),
    .A2(_12533_),
    .B(_12539_),
    .Y(_04200_));
 BUFx4f_ASAP7_75t_R _33777_ (.A(_12532_),
    .Y(_12540_));
 NOR2x1_ASAP7_75t_R _33778_ (.A(_16028_),
    .B(_12532_),
    .Y(_12541_));
 AO21x1_ASAP7_75t_R _33779_ (.A1(_15867_),
    .A2(_12540_),
    .B(_12541_),
    .Y(_04201_));
 NAND2x1_ASAP7_75t_R _33780_ (.A(_01537_),
    .B(_12534_),
    .Y(_12542_));
 OA21x2_ASAP7_75t_R _33781_ (.A1(\alu_adder_result_ex[15] ),
    .A2(_12533_),
    .B(_12542_),
    .Y(_04202_));
 NAND2x1_ASAP7_75t_R _33782_ (.A(_01536_),
    .B(_12534_),
    .Y(_12543_));
 OA21x2_ASAP7_75t_R _33783_ (.A1(\alu_adder_result_ex[16] ),
    .A2(_12533_),
    .B(_12543_),
    .Y(_04203_));
 NAND2x1_ASAP7_75t_R _33784_ (.A(_01535_),
    .B(_12534_),
    .Y(_12544_));
 OA21x2_ASAP7_75t_R _33785_ (.A1(\alu_adder_result_ex[17] ),
    .A2(_12533_),
    .B(_12544_),
    .Y(_04204_));
 BUFx6f_ASAP7_75t_R _33786_ (.A(_12532_),
    .Y(_12545_));
 NAND2x1_ASAP7_75t_R _33787_ (.A(_01534_),
    .B(_12545_),
    .Y(_12546_));
 OA21x2_ASAP7_75t_R _33788_ (.A1(\alu_adder_result_ex[18] ),
    .A2(_12533_),
    .B(_12546_),
    .Y(_04205_));
 NAND2x1_ASAP7_75t_R _33789_ (.A(_01533_),
    .B(_12545_),
    .Y(_12547_));
 OA21x2_ASAP7_75t_R _33790_ (.A1(\alu_adder_result_ex[19] ),
    .A2(_12533_),
    .B(_12547_),
    .Y(_04206_));
 BUFx4f_ASAP7_75t_R _33791_ (.A(_12532_),
    .Y(_12548_));
 NAND2x1_ASAP7_75t_R _33792_ (.A(_01532_),
    .B(_12545_),
    .Y(_12549_));
 OA21x2_ASAP7_75t_R _33793_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_12548_),
    .B(_12549_),
    .Y(_04207_));
 NAND2x1_ASAP7_75t_R _33794_ (.A(_01531_),
    .B(_12545_),
    .Y(_12550_));
 OA21x2_ASAP7_75t_R _33795_ (.A1(\alu_adder_result_ex[20] ),
    .A2(_12548_),
    .B(_12550_),
    .Y(_04208_));
 NAND2x1_ASAP7_75t_R _33796_ (.A(_01530_),
    .B(_12545_),
    .Y(_12551_));
 OA21x2_ASAP7_75t_R _33797_ (.A1(\alu_adder_result_ex[21] ),
    .A2(_12548_),
    .B(_12551_),
    .Y(_04209_));
 NAND2x1_ASAP7_75t_R _33798_ (.A(_01529_),
    .B(_12545_),
    .Y(_12552_));
 OA21x2_ASAP7_75t_R _33799_ (.A1(\alu_adder_result_ex[22] ),
    .A2(_12548_),
    .B(_12552_),
    .Y(_04210_));
 NAND2x1_ASAP7_75t_R _33800_ (.A(_01528_),
    .B(_12545_),
    .Y(_12553_));
 OA21x2_ASAP7_75t_R _33801_ (.A1(\alu_adder_result_ex[23] ),
    .A2(_12548_),
    .B(_12553_),
    .Y(_04211_));
 NOR2x1_ASAP7_75t_R _33802_ (.A(_17257_),
    .B(_12532_),
    .Y(_12554_));
 AO21x1_ASAP7_75t_R _33803_ (.A1(_17125_),
    .A2(_12540_),
    .B(_12554_),
    .Y(_04212_));
 NAND2x1_ASAP7_75t_R _33804_ (.A(_01526_),
    .B(_12545_),
    .Y(_12555_));
 OA21x2_ASAP7_75t_R _33805_ (.A1(\alu_adder_result_ex[25] ),
    .A2(_12548_),
    .B(_12555_),
    .Y(_04213_));
 NOR2x1_ASAP7_75t_R _33806_ (.A(_04414_),
    .B(_12532_),
    .Y(_12556_));
 AO21x1_ASAP7_75t_R _33807_ (.A1(_04283_),
    .A2(_12534_),
    .B(_12556_),
    .Y(_04214_));
 NAND2x1_ASAP7_75t_R _33808_ (.A(_01524_),
    .B(_12545_),
    .Y(_12557_));
 OA21x2_ASAP7_75t_R _33809_ (.A1(\alu_adder_result_ex[27] ),
    .A2(_12548_),
    .B(_12557_),
    .Y(_04215_));
 NAND2x1_ASAP7_75t_R _33810_ (.A(_01523_),
    .B(_12545_),
    .Y(_12558_));
 OA21x2_ASAP7_75t_R _33811_ (.A1(\alu_adder_result_ex[28] ),
    .A2(_12548_),
    .B(_12558_),
    .Y(_04216_));
 BUFx6f_ASAP7_75t_R _33812_ (.A(_12532_),
    .Y(_12559_));
 NAND2x1_ASAP7_75t_R _33813_ (.A(_01522_),
    .B(_12559_),
    .Y(_12560_));
 OA21x2_ASAP7_75t_R _33814_ (.A1(\alu_adder_result_ex[29] ),
    .A2(_12548_),
    .B(_12560_),
    .Y(_04217_));
 NAND2x1_ASAP7_75t_R _33815_ (.A(_01521_),
    .B(_12559_),
    .Y(_12561_));
 OA21x2_ASAP7_75t_R _33816_ (.A1(\alu_adder_result_ex[2] ),
    .A2(_12548_),
    .B(_12561_),
    .Y(_04218_));
 NAND2x1_ASAP7_75t_R _33817_ (.A(_01520_),
    .B(_12559_),
    .Y(_12562_));
 OA21x2_ASAP7_75t_R _33818_ (.A1(\alu_adder_result_ex[30] ),
    .A2(_12540_),
    .B(_12562_),
    .Y(_04219_));
 NAND2x1_ASAP7_75t_R _33819_ (.A(_01519_),
    .B(_12559_),
    .Y(_12563_));
 OA21x2_ASAP7_75t_R _33820_ (.A1(\alu_adder_result_ex[31] ),
    .A2(_12540_),
    .B(_12563_),
    .Y(_04220_));
 NAND2x1_ASAP7_75t_R _33821_ (.A(_01518_),
    .B(_12559_),
    .Y(_12564_));
 OA21x2_ASAP7_75t_R _33822_ (.A1(\alu_adder_result_ex[3] ),
    .A2(_12540_),
    .B(_12564_),
    .Y(_04221_));
 NAND2x1_ASAP7_75t_R _33823_ (.A(_01517_),
    .B(_12559_),
    .Y(_12565_));
 OA21x2_ASAP7_75t_R _33824_ (.A1(\alu_adder_result_ex[4] ),
    .A2(_12540_),
    .B(_12565_),
    .Y(_04222_));
 NAND2x1_ASAP7_75t_R _33825_ (.A(_01516_),
    .B(_12559_),
    .Y(_12566_));
 OA21x2_ASAP7_75t_R _33826_ (.A1(\alu_adder_result_ex[5] ),
    .A2(_12540_),
    .B(_12566_),
    .Y(_04223_));
 NAND2x1_ASAP7_75t_R _33827_ (.A(_01515_),
    .B(_12559_),
    .Y(_12567_));
 OA21x2_ASAP7_75t_R _33828_ (.A1(\alu_adder_result_ex[6] ),
    .A2(_12540_),
    .B(_12567_),
    .Y(_04224_));
 NAND2x1_ASAP7_75t_R _33829_ (.A(_01514_),
    .B(_12559_),
    .Y(_12568_));
 OA21x2_ASAP7_75t_R _33830_ (.A1(\alu_adder_result_ex[7] ),
    .A2(_12540_),
    .B(_12568_),
    .Y(_04225_));
 NOR2x1_ASAP7_75t_R _33831_ (.A(_15417_),
    .B(_12532_),
    .Y(_12569_));
 AO21x1_ASAP7_75t_R _33832_ (.A1(_15338_),
    .A2(_12534_),
    .B(_12569_),
    .Y(_04226_));
 NAND2x1_ASAP7_75t_R _33833_ (.A(_01512_),
    .B(_12559_),
    .Y(_12570_));
 OA21x2_ASAP7_75t_R _33834_ (.A1(\alu_adder_result_ex[9] ),
    .A2(_12540_),
    .B(_12570_),
    .Y(_04227_));
 INVx1_ASAP7_75t_R _33835_ (.A(_01511_),
    .Y(_12571_));
 AND4x1_ASAP7_75t_R _33836_ (.A(_13595_),
    .B(net2013),
    .C(_14026_),
    .D(_05758_),
    .Y(_12572_));
 AO21x1_ASAP7_75t_R _33837_ (.A1(_12571_),
    .A2(_05756_),
    .B(_12572_),
    .Y(_04228_));
 AND3x4_ASAP7_75t_R _33838_ (.A(_13399_),
    .B(_14026_),
    .C(_04928_),
    .Y(net267));
 AND2x2_ASAP7_75t_R _33839_ (.A(_05758_),
    .B(net267),
    .Y(_12573_));
 AO21x1_ASAP7_75t_R _33840_ (.A1(_04924_),
    .A2(_05756_),
    .B(_12573_),
    .Y(_04229_));
 AO21x1_ASAP7_75t_R _33841_ (.A1(net104),
    .A2(_13357_),
    .B(_05752_),
    .Y(_12574_));
 OA21x2_ASAP7_75t_R _33842_ (.A1(_13358_),
    .A2(_05754_),
    .B(_05752_),
    .Y(_12575_));
 AO21x1_ASAP7_75t_R _33843_ (.A1(_13425_),
    .A2(_12574_),
    .B(_12575_),
    .Y(_12576_));
 AND2x2_ASAP7_75t_R _33844_ (.A(_05751_),
    .B(_12576_),
    .Y(_12577_));
 INVx3_ASAP7_75t_R _33845_ (.A(_18762_),
    .Y(_12578_));
 NAND2x2_ASAP7_75t_R _33846_ (.A(_13585_),
    .B(_14026_),
    .Y(_12579_));
 OR3x1_ASAP7_75t_R _33847_ (.A(_13561_),
    .B(_02287_),
    .C(_12579_),
    .Y(_12580_));
 OA21x2_ASAP7_75t_R _33848_ (.A1(_12578_),
    .A2(_05761_),
    .B(_12580_),
    .Y(_12581_));
 INVx1_ASAP7_75t_R _33849_ (.A(net104),
    .Y(_12582_));
 OR3x1_ASAP7_75t_R _33850_ (.A(_05752_),
    .B(_12582_),
    .C(_13358_),
    .Y(_12583_));
 AND2x2_ASAP7_75t_R _33851_ (.A(_05751_),
    .B(_13425_),
    .Y(_12584_));
 AO32x1_ASAP7_75t_R _33852_ (.A1(_13359_),
    .A2(_13357_),
    .A3(_12581_),
    .B1(_12583_),
    .B2(_12584_),
    .Y(_12585_));
 NAND2x1_ASAP7_75t_R _33853_ (.A(_12577_),
    .B(_12585_),
    .Y(_12586_));
 OA21x2_ASAP7_75t_R _33854_ (.A1(_13424_),
    .A2(_12577_),
    .B(_12586_),
    .Y(_04230_));
 INVx1_ASAP7_75t_R _33855_ (.A(_05752_),
    .Y(_12587_));
 AO21x1_ASAP7_75t_R _33856_ (.A1(net104),
    .A2(_13425_),
    .B(_05755_),
    .Y(_12588_));
 AND3x1_ASAP7_75t_R _33857_ (.A(_05751_),
    .B(_12587_),
    .C(_12588_),
    .Y(_04231_));
 INVx1_ASAP7_75t_R _33858_ (.A(_05754_),
    .Y(_12589_));
 OAI21x1_ASAP7_75t_R _33859_ (.A1(_12589_),
    .A2(_12581_),
    .B(_13357_),
    .Y(_12590_));
 AO21x1_ASAP7_75t_R _33860_ (.A1(_13359_),
    .A2(_12590_),
    .B(_12587_),
    .Y(_12591_));
 AND3x1_ASAP7_75t_R _33861_ (.A(_13357_),
    .B(_05754_),
    .C(_12581_),
    .Y(_12592_));
 OR3x1_ASAP7_75t_R _33862_ (.A(_05752_),
    .B(_13425_),
    .C(_12592_),
    .Y(_12593_));
 AND3x1_ASAP7_75t_R _33863_ (.A(_05751_),
    .B(_12591_),
    .C(_12593_),
    .Y(_04232_));
 AND2x2_ASAP7_75t_R _33864_ (.A(_13360_),
    .B(_13359_),
    .Y(_12594_));
 AND3x1_ASAP7_75t_R _33865_ (.A(_05751_),
    .B(_05752_),
    .C(_13425_),
    .Y(_12595_));
 OA211x2_ASAP7_75t_R _33866_ (.A1(_12594_),
    .A2(_12595_),
    .B(_12582_),
    .C(_13357_),
    .Y(_04233_));
 OA211x2_ASAP7_75t_R _33867_ (.A1(_12584_),
    .A2(_12594_),
    .B(net104),
    .C(_13357_),
    .Y(_12596_));
 BUFx4f_ASAP7_75t_R _33868_ (.A(_12596_),
    .Y(_12597_));
 AOI211x1_ASAP7_75t_R _33869_ (.A1(_04922_),
    .A2(_05754_),
    .B(_12597_),
    .C(_01508_),
    .Y(_12598_));
 AO21x1_ASAP7_75t_R _33870_ (.A1(net47),
    .A2(_12597_),
    .B(_12598_),
    .Y(_04234_));
 NAND2x1_ASAP7_75t_R _33871_ (.A(_18769_),
    .B(_05758_),
    .Y(_12599_));
 OA21x2_ASAP7_75t_R _33872_ (.A1(_08908_),
    .A2(_05758_),
    .B(_12599_),
    .Y(_04235_));
 NAND2x1_ASAP7_75t_R _33873_ (.A(_18764_),
    .B(_05758_),
    .Y(_12600_));
 OA21x2_ASAP7_75t_R _33874_ (.A1(_08885_),
    .A2(_05758_),
    .B(_12600_),
    .Y(_04236_));
 NAND2x2_ASAP7_75t_R _33875_ (.A(_01454_),
    .B(_12596_),
    .Y(_12601_));
 BUFx4f_ASAP7_75t_R _33876_ (.A(_12601_),
    .Y(_12602_));
 AO21x1_ASAP7_75t_R _33877_ (.A1(_04919_),
    .A2(_12597_),
    .B(_08569_),
    .Y(_12603_));
 OA21x2_ASAP7_75t_R _33878_ (.A1(net102),
    .A2(_12602_),
    .B(_12603_),
    .Y(_04237_));
 AO21x1_ASAP7_75t_R _33879_ (.A1(_04919_),
    .A2(_12597_),
    .B(_08958_),
    .Y(_12604_));
 OA21x2_ASAP7_75t_R _33880_ (.A1(net80),
    .A2(_12602_),
    .B(_12604_),
    .Y(_04238_));
 AO21x1_ASAP7_75t_R _33881_ (.A1(_04919_),
    .A2(_12597_),
    .B(_09001_),
    .Y(_12605_));
 OA21x2_ASAP7_75t_R _33882_ (.A1(net81),
    .A2(_12602_),
    .B(_12605_),
    .Y(_04239_));
 AO21x1_ASAP7_75t_R _33883_ (.A1(_04919_),
    .A2(_12597_),
    .B(_08602_),
    .Y(_12606_));
 OA21x2_ASAP7_75t_R _33884_ (.A1(net83),
    .A2(_12602_),
    .B(_12606_),
    .Y(_04240_));
 AO21x1_ASAP7_75t_R _33885_ (.A1(_04919_),
    .A2(_12597_),
    .B(_08687_),
    .Y(_12607_));
 OA21x2_ASAP7_75t_R _33886_ (.A1(net84),
    .A2(_12602_),
    .B(_12607_),
    .Y(_04241_));
 AO21x1_ASAP7_75t_R _33887_ (.A1(_04919_),
    .A2(_12597_),
    .B(_08767_),
    .Y(_12608_));
 OA21x2_ASAP7_75t_R _33888_ (.A1(net85),
    .A2(_12602_),
    .B(_12608_),
    .Y(_04242_));
 AO21x1_ASAP7_75t_R _33889_ (.A1(_04919_),
    .A2(_12597_),
    .B(_08813_),
    .Y(_12609_));
 OA21x2_ASAP7_75t_R _33890_ (.A1(net86),
    .A2(_12602_),
    .B(_12609_),
    .Y(_04243_));
 BUFx4f_ASAP7_75t_R _33891_ (.A(_12601_),
    .Y(_12610_));
 NAND2x1_ASAP7_75t_R _33892_ (.A(_01498_),
    .B(_12610_),
    .Y(_12611_));
 OA21x2_ASAP7_75t_R _33893_ (.A1(net87),
    .A2(_12602_),
    .B(_12611_),
    .Y(_04244_));
 BUFx4f_ASAP7_75t_R _33894_ (.A(_12596_),
    .Y(_12612_));
 AND3x1_ASAP7_75t_R _33895_ (.A(_04918_),
    .B(_09446_),
    .C(_12612_),
    .Y(_12613_));
 AOI21x1_ASAP7_75t_R _33896_ (.A1(_01497_),
    .A2(_12602_),
    .B(_12613_),
    .Y(_04245_));
 NAND2x1_ASAP7_75t_R _33897_ (.A(_01496_),
    .B(_12610_),
    .Y(_12614_));
 OA21x2_ASAP7_75t_R _33898_ (.A1(net89),
    .A2(_12602_),
    .B(_12614_),
    .Y(_04246_));
 BUFx4f_ASAP7_75t_R _33899_ (.A(_12601_),
    .Y(_12615_));
 NAND2x1_ASAP7_75t_R _33900_ (.A(_01495_),
    .B(_12610_),
    .Y(_12616_));
 OA21x2_ASAP7_75t_R _33901_ (.A1(net90),
    .A2(_12615_),
    .B(_12616_),
    .Y(_04247_));
 AO21x1_ASAP7_75t_R _33902_ (.A1(_04919_),
    .A2(_12597_),
    .B(_09667_),
    .Y(_12617_));
 OA21x2_ASAP7_75t_R _33903_ (.A1(net103),
    .A2(_12615_),
    .B(_12617_),
    .Y(_04248_));
 NAND2x1_ASAP7_75t_R _33904_ (.A(_01493_),
    .B(_12610_),
    .Y(_12618_));
 OA21x2_ASAP7_75t_R _33905_ (.A1(net91),
    .A2(_12615_),
    .B(_12618_),
    .Y(_04249_));
 NAND2x1_ASAP7_75t_R _33906_ (.A(_01492_),
    .B(_12610_),
    .Y(_12619_));
 OA21x2_ASAP7_75t_R _33907_ (.A1(net92),
    .A2(_12615_),
    .B(_12619_),
    .Y(_04250_));
 AO21x1_ASAP7_75t_R _33908_ (.A1(_04919_),
    .A2(_12612_),
    .B(_09135_),
    .Y(_12620_));
 OA21x2_ASAP7_75t_R _33909_ (.A1(net94),
    .A2(_12615_),
    .B(_12620_),
    .Y(_04251_));
 AO21x1_ASAP7_75t_R _33910_ (.A1(_04918_),
    .A2(_12612_),
    .B(_09410_),
    .Y(_12621_));
 OA21x2_ASAP7_75t_R _33911_ (.A1(net96),
    .A2(_12615_),
    .B(_12621_),
    .Y(_04252_));
 AO21x1_ASAP7_75t_R _33912_ (.A1(_04918_),
    .A2(_12612_),
    .B(_09681_),
    .Y(_12622_));
 OA21x2_ASAP7_75t_R _33913_ (.A1(net49),
    .A2(_12615_),
    .B(_12622_),
    .Y(_04253_));
 AO21x1_ASAP7_75t_R _33914_ (.A1(_04918_),
    .A2(_12612_),
    .B(_09699_),
    .Y(_12623_));
 OA21x2_ASAP7_75t_R _33915_ (.A1(net50),
    .A2(_12615_),
    .B(_12623_),
    .Y(_04254_));
 AO21x1_ASAP7_75t_R _33916_ (.A1(_04918_),
    .A2(_12612_),
    .B(_08605_),
    .Y(_12624_));
 OA21x2_ASAP7_75t_R _33917_ (.A1(net51),
    .A2(_12615_),
    .B(_12624_),
    .Y(_04255_));
 AO21x1_ASAP7_75t_R _33918_ (.A1(_04918_),
    .A2(_12612_),
    .B(_08688_),
    .Y(_12625_));
 OA21x2_ASAP7_75t_R _33919_ (.A1(net75),
    .A2(_12615_),
    .B(_12625_),
    .Y(_04256_));
 AO21x1_ASAP7_75t_R _33920_ (.A1(_04918_),
    .A2(_12612_),
    .B(_08768_),
    .Y(_12626_));
 OA21x2_ASAP7_75t_R _33921_ (.A1(net76),
    .A2(_12610_),
    .B(_12626_),
    .Y(_04257_));
 AO21x1_ASAP7_75t_R _33922_ (.A1(_04918_),
    .A2(_12612_),
    .B(_08814_),
    .Y(_12627_));
 OA21x2_ASAP7_75t_R _33923_ (.A1(net77),
    .A2(_12610_),
    .B(_12627_),
    .Y(_04258_));
 AO21x1_ASAP7_75t_R _33924_ (.A1(_04918_),
    .A2(_12612_),
    .B(_08568_),
    .Y(_12628_));
 OA21x2_ASAP7_75t_R _33925_ (.A1(net78),
    .A2(_12610_),
    .B(_12628_),
    .Y(_04259_));
 NAND2x1_ASAP7_75t_R _33926_ (.A(_01482_),
    .B(_12610_),
    .Y(_12629_));
 OA21x2_ASAP7_75t_R _33927_ (.A1(net79),
    .A2(_12610_),
    .B(_12629_),
    .Y(_04260_));
 NOR2x1_ASAP7_75t_R _33928_ (.A(_04952_),
    .B(_04984_),
    .Y(_12630_));
 AO21x2_ASAP7_75t_R _33929_ (.A1(_12630_),
    .A2(_07764_),
    .B(_07251_),
    .Y(_12631_));
 NOR3x2_ASAP7_75t_R _33930_ (.B(_06475_),
    .C(_07251_),
    .Y(_12632_),
    .A(_05840_));
 AOI21x1_ASAP7_75t_R _33931_ (.A1(_14812_),
    .A2(_07251_),
    .B(_12632_),
    .Y(_12633_));
 NOR2x1_ASAP7_75t_R _33932_ (.A(_02081_),
    .B(_12631_),
    .Y(_12634_));
 AO21x1_ASAP7_75t_R _33933_ (.A1(_12631_),
    .A2(_12633_),
    .B(_12634_),
    .Y(_02491_));
 AOI21x1_ASAP7_75t_R _33934_ (.A1(_05068_),
    .A2(_07251_),
    .B(_12632_),
    .Y(_12635_));
 NOR2x1_ASAP7_75t_R _33935_ (.A(_02078_),
    .B(_12631_),
    .Y(_12636_));
 AO21x1_ASAP7_75t_R _33936_ (.A1(_12631_),
    .A2(_12635_),
    .B(_12636_),
    .Y(_02496_));
 BUFx4f_ASAP7_75t_R _33937_ (.A(_11957_),
    .Y(_12637_));
 BUFx6f_ASAP7_75t_R _33938_ (.A(_12637_),
    .Y(_12638_));
 AND2x2_ASAP7_75t_R _33939_ (.A(net156),
    .B(_07311_),
    .Y(_12639_));
 AO21x1_ASAP7_75t_R _33940_ (.A1(net150),
    .A2(_05484_),
    .B(_12639_),
    .Y(_12640_));
 INVx1_ASAP7_75t_R _33941_ (.A(_01672_),
    .Y(_12641_));
 NAND2x1_ASAP7_75t_R _33942_ (.A(_07311_),
    .B(_01669_),
    .Y(_12642_));
 OA211x2_ASAP7_75t_R _33943_ (.A1(_07311_),
    .A2(_12641_),
    .B(_12642_),
    .C(_05490_),
    .Y(_12643_));
 AOI21x1_ASAP7_75t_R _33944_ (.A1(_05487_),
    .A2(_12640_),
    .B(_12643_),
    .Y(_12644_));
 BUFx4f_ASAP7_75t_R _33945_ (.A(_12644_),
    .Y(_12645_));
 BUFx4f_ASAP7_75t_R _33946_ (.A(_12645_),
    .Y(_12646_));
 AND2x2_ASAP7_75t_R _33947_ (.A(net144),
    .B(_07310_),
    .Y(_12647_));
 AO21x1_ASAP7_75t_R _33948_ (.A1(net165),
    .A2(_05483_),
    .B(_12647_),
    .Y(_12648_));
 INVx1_ASAP7_75t_R _33949_ (.A(_01660_),
    .Y(_12649_));
 NAND2x1_ASAP7_75t_R _33950_ (.A(_07310_),
    .B(_01677_),
    .Y(_12650_));
 OA211x2_ASAP7_75t_R _33951_ (.A1(_07310_),
    .A2(_12649_),
    .B(_12650_),
    .C(_05490_),
    .Y(_12651_));
 AOI21x1_ASAP7_75t_R _33952_ (.A1(_05487_),
    .A2(_12648_),
    .B(_12651_),
    .Y(_12652_));
 BUFx4f_ASAP7_75t_R _33953_ (.A(_12652_),
    .Y(_12653_));
 AND2x2_ASAP7_75t_R _33954_ (.A(net143),
    .B(_05471_),
    .Y(_12654_));
 AO21x1_ASAP7_75t_R _33955_ (.A1(net164),
    .A2(_05472_),
    .B(_12654_),
    .Y(_12655_));
 INVx1_ASAP7_75t_R _33956_ (.A(_01661_),
    .Y(_12656_));
 NAND2x1_ASAP7_75t_R _33957_ (.A(_05471_),
    .B(_01678_),
    .Y(_12657_));
 OA211x2_ASAP7_75t_R _33958_ (.A1(_07308_),
    .A2(_12656_),
    .B(_12657_),
    .C(_05489_),
    .Y(_12658_));
 AO21x2_ASAP7_75t_R _33959_ (.A1(_05473_),
    .A2(_12655_),
    .B(_12658_),
    .Y(_12659_));
 BUFx4f_ASAP7_75t_R _33960_ (.A(_12659_),
    .Y(_12660_));
 AND2x2_ASAP7_75t_R _33961_ (.A(net142),
    .B(_05471_),
    .Y(_12661_));
 AO21x1_ASAP7_75t_R _33962_ (.A1(net163),
    .A2(_05472_),
    .B(_12661_),
    .Y(_12662_));
 INVx1_ASAP7_75t_R _33963_ (.A(_01662_),
    .Y(_12663_));
 NAND2x1_ASAP7_75t_R _33964_ (.A(_05471_),
    .B(_01679_),
    .Y(_12664_));
 OA211x2_ASAP7_75t_R _33965_ (.A1(_07308_),
    .A2(_12663_),
    .B(_12664_),
    .C(_05489_),
    .Y(_12665_));
 AOI21x1_ASAP7_75t_R _33966_ (.A1(_11958_),
    .A2(_12662_),
    .B(_12665_),
    .Y(_12666_));
 AND2x2_ASAP7_75t_R _33967_ (.A(net148),
    .B(_07309_),
    .Y(_12667_));
 AO21x1_ASAP7_75t_R _33968_ (.A1(net169),
    .A2(_05483_),
    .B(_12667_),
    .Y(_12668_));
 BUFx4f_ASAP7_75t_R _33969_ (.A(_07308_),
    .Y(_12669_));
 INVx1_ASAP7_75t_R _33970_ (.A(_01656_),
    .Y(_12670_));
 NAND2x1_ASAP7_75t_R _33971_ (.A(_07309_),
    .B(_01674_),
    .Y(_12671_));
 OA211x2_ASAP7_75t_R _33972_ (.A1(_12669_),
    .A2(_12670_),
    .B(_12671_),
    .C(_05489_),
    .Y(_12672_));
 AOI21x1_ASAP7_75t_R _33973_ (.A1(_05485_),
    .A2(_12668_),
    .B(_12672_),
    .Y(_12673_));
 AND2x2_ASAP7_75t_R _33974_ (.A(net147),
    .B(_07309_),
    .Y(_12674_));
 AO21x1_ASAP7_75t_R _33975_ (.A1(net168),
    .A2(_05483_),
    .B(_12674_),
    .Y(_12675_));
 INVx1_ASAP7_75t_R _33976_ (.A(_01657_),
    .Y(_12676_));
 NAND2x1_ASAP7_75t_R _33977_ (.A(_07309_),
    .B(_01675_),
    .Y(_12677_));
 OA211x2_ASAP7_75t_R _33978_ (.A1(_12669_),
    .A2(_12676_),
    .B(_12677_),
    .C(_05489_),
    .Y(_12678_));
 AO21x2_ASAP7_75t_R _33979_ (.A1(_05485_),
    .A2(_12675_),
    .B(_12678_),
    .Y(_12679_));
 BUFx4f_ASAP7_75t_R _33980_ (.A(_12679_),
    .Y(_12680_));
 AND2x2_ASAP7_75t_R _33981_ (.A(net146),
    .B(_12669_),
    .Y(_12681_));
 AO21x1_ASAP7_75t_R _33982_ (.A1(net166),
    .A2(_05483_),
    .B(_12681_),
    .Y(_12682_));
 INVx1_ASAP7_75t_R _33983_ (.A(_01659_),
    .Y(_12683_));
 NAND2x1_ASAP7_75t_R _33984_ (.A(_12669_),
    .B(_01676_),
    .Y(_12684_));
 OA211x2_ASAP7_75t_R _33985_ (.A1(_12669_),
    .A2(_12683_),
    .B(_12684_),
    .C(_05490_),
    .Y(_12685_));
 AO21x2_ASAP7_75t_R _33986_ (.A1(_05486_),
    .A2(_12682_),
    .B(_12685_),
    .Y(_12686_));
 OR3x4_ASAP7_75t_R _33987_ (.A(_12673_),
    .B(_12680_),
    .C(_12686_),
    .Y(_12687_));
 AO21x1_ASAP7_75t_R _33988_ (.A1(_12660_),
    .A2(_12666_),
    .B(_12687_),
    .Y(_12688_));
 AO21x1_ASAP7_75t_R _33989_ (.A1(_05486_),
    .A2(_12648_),
    .B(_12651_),
    .Y(_12689_));
 BUFx4f_ASAP7_75t_R _33990_ (.A(_12689_),
    .Y(_12690_));
 BUFx4f_ASAP7_75t_R _33991_ (.A(_12690_),
    .Y(_12691_));
 AOI21x1_ASAP7_75t_R _33992_ (.A1(_05485_),
    .A2(_12682_),
    .B(_12685_),
    .Y(_12692_));
 BUFx6f_ASAP7_75t_R _33993_ (.A(_12692_),
    .Y(_12693_));
 BUFx4f_ASAP7_75t_R _33994_ (.A(_12693_),
    .Y(_12694_));
 AND2x2_ASAP7_75t_R _33995_ (.A(_07309_),
    .B(net170),
    .Y(_12695_));
 AO21x1_ASAP7_75t_R _33996_ (.A1(_05483_),
    .A2(net155),
    .B(_12695_),
    .Y(_12696_));
 INVx1_ASAP7_75t_R _33997_ (.A(_01670_),
    .Y(_12697_));
 NAND2x1_ASAP7_75t_R _33998_ (.A(_07309_),
    .B(_01647_),
    .Y(_12698_));
 OA211x2_ASAP7_75t_R _33999_ (.A1(_12669_),
    .A2(_12697_),
    .B(_12698_),
    .C(_05489_),
    .Y(_12699_));
 AO21x1_ASAP7_75t_R _34000_ (.A1(_05485_),
    .A2(_12696_),
    .B(_12699_),
    .Y(_12700_));
 BUFx4f_ASAP7_75t_R _34001_ (.A(_12700_),
    .Y(_12701_));
 AND2x2_ASAP7_75t_R _34002_ (.A(_07308_),
    .B(net173),
    .Y(_12702_));
 AO21x1_ASAP7_75t_R _34003_ (.A1(_05472_),
    .A2(net159),
    .B(_12702_),
    .Y(_12703_));
 INVx1_ASAP7_75t_R _34004_ (.A(_01666_),
    .Y(_12704_));
 NAND2x1_ASAP7_75t_R _34005_ (.A(_07309_),
    .B(_01614_),
    .Y(_12705_));
 OA211x2_ASAP7_75t_R _34006_ (.A1(_07309_),
    .A2(_12704_),
    .B(_12705_),
    .C(_05489_),
    .Y(_12706_));
 AO21x1_ASAP7_75t_R _34007_ (.A1(_05485_),
    .A2(_12703_),
    .B(_12706_),
    .Y(_12707_));
 AND2x2_ASAP7_75t_R _34008_ (.A(_07308_),
    .B(net172),
    .Y(_12708_));
 AO21x1_ASAP7_75t_R _34009_ (.A1(_05472_),
    .A2(net158),
    .B(_12708_),
    .Y(_12709_));
 INVx1_ASAP7_75t_R _34010_ (.A(_01667_),
    .Y(_12710_));
 NAND2x1_ASAP7_75t_R _34011_ (.A(_07308_),
    .B(_01625_),
    .Y(_12711_));
 OA211x2_ASAP7_75t_R _34012_ (.A1(_07309_),
    .A2(_12710_),
    .B(_12711_),
    .C(_05489_),
    .Y(_12712_));
 AO21x1_ASAP7_75t_R _34013_ (.A1(_05473_),
    .A2(_12709_),
    .B(_12712_),
    .Y(_12713_));
 OR2x2_ASAP7_75t_R _34014_ (.A(_12707_),
    .B(_12713_),
    .Y(_12714_));
 AND2x2_ASAP7_75t_R _34015_ (.A(_12669_),
    .B(net167),
    .Y(_12715_));
 AO21x1_ASAP7_75t_R _34016_ (.A1(_05483_),
    .A2(net154),
    .B(_12715_),
    .Y(_12716_));
 INVx1_ASAP7_75t_R _34017_ (.A(_01671_),
    .Y(_12717_));
 NAND2x1_ASAP7_75t_R _34018_ (.A(_12669_),
    .B(_01658_),
    .Y(_12718_));
 OA211x2_ASAP7_75t_R _34019_ (.A1(_07310_),
    .A2(_12717_),
    .B(_12718_),
    .C(_05490_),
    .Y(_12719_));
 AO21x2_ASAP7_75t_R _34020_ (.A1(_05485_),
    .A2(_12716_),
    .B(_12719_),
    .Y(_12720_));
 AND2x2_ASAP7_75t_R _34021_ (.A(_07310_),
    .B(net171),
    .Y(_12721_));
 AO21x1_ASAP7_75t_R _34022_ (.A1(_05483_),
    .A2(net157),
    .B(_12721_),
    .Y(_12722_));
 INVx1_ASAP7_75t_R _34023_ (.A(_01668_),
    .Y(_12723_));
 NAND2x1_ASAP7_75t_R _34024_ (.A(_07310_),
    .B(_01636_),
    .Y(_12724_));
 OA211x2_ASAP7_75t_R _34025_ (.A1(_07310_),
    .A2(_12723_),
    .B(_12724_),
    .C(_05490_),
    .Y(_12725_));
 AO21x1_ASAP7_75t_R _34026_ (.A1(_05486_),
    .A2(_12722_),
    .B(_12725_),
    .Y(_12726_));
 OR4x1_ASAP7_75t_R _34027_ (.A(_12701_),
    .B(_12714_),
    .C(_12720_),
    .D(_12726_),
    .Y(_12727_));
 BUFx4f_ASAP7_75t_R _34028_ (.A(_12727_),
    .Y(_12728_));
 NAND2x2_ASAP7_75t_R _34029_ (.A(_12673_),
    .B(_12679_),
    .Y(_12729_));
 OR4x1_ASAP7_75t_R _34030_ (.A(_12691_),
    .B(_12694_),
    .C(_12728_),
    .D(_12729_),
    .Y(_12730_));
 AND2x2_ASAP7_75t_R _34031_ (.A(net141),
    .B(_07311_),
    .Y(_12731_));
 AO21x1_ASAP7_75t_R _34032_ (.A1(net149),
    .A2(_05483_),
    .B(_12731_),
    .Y(_12732_));
 NAND2x1_ASAP7_75t_R _34033_ (.A(_07311_),
    .B(_01680_),
    .Y(_12733_));
 OA211x2_ASAP7_75t_R _34034_ (.A1(_07311_),
    .A2(_05476_),
    .B(_12733_),
    .C(_05490_),
    .Y(_12734_));
 AO21x2_ASAP7_75t_R _34035_ (.A1(_05487_),
    .A2(_12732_),
    .B(_12734_),
    .Y(_12735_));
 BUFx3_ASAP7_75t_R _34036_ (.A(_12735_),
    .Y(_12736_));
 OA211x2_ASAP7_75t_R _34037_ (.A1(_12653_),
    .A2(_12688_),
    .B(_12730_),
    .C(_12736_),
    .Y(_12737_));
 INVx1_ASAP7_75t_R _34038_ (.A(_12737_),
    .Y(_12738_));
 BUFx3_ASAP7_75t_R _34039_ (.A(_12735_),
    .Y(_12739_));
 AO21x2_ASAP7_75t_R _34040_ (.A1(_05485_),
    .A2(_12668_),
    .B(_12672_),
    .Y(_12740_));
 BUFx4f_ASAP7_75t_R _34041_ (.A(_12740_),
    .Y(_12741_));
 AOI21x1_ASAP7_75t_R _34042_ (.A1(_05485_),
    .A2(_12675_),
    .B(_12678_),
    .Y(_12742_));
 BUFx4f_ASAP7_75t_R _34043_ (.A(_12742_),
    .Y(_12743_));
 BUFx4f_ASAP7_75t_R _34044_ (.A(_12686_),
    .Y(_12744_));
 AO21x2_ASAP7_75t_R _34045_ (.A1(_12741_),
    .A2(_12743_),
    .B(_12744_),
    .Y(_12745_));
 BUFx3_ASAP7_75t_R _34046_ (.A(_12745_),
    .Y(_12746_));
 BUFx4f_ASAP7_75t_R _34047_ (.A(_12680_),
    .Y(_12747_));
 AND2x2_ASAP7_75t_R _34048_ (.A(_12669_),
    .B(net175),
    .Y(_12748_));
 AO21x1_ASAP7_75t_R _34049_ (.A1(_05483_),
    .A2(net161),
    .B(_12748_),
    .Y(_12749_));
 INVx1_ASAP7_75t_R _34050_ (.A(_01664_),
    .Y(_12750_));
 NAND2x1_ASAP7_75t_R _34051_ (.A(_12669_),
    .B(_01592_),
    .Y(_12751_));
 OA211x2_ASAP7_75t_R _34052_ (.A1(_07310_),
    .A2(_12750_),
    .B(_12751_),
    .C(_05490_),
    .Y(_12752_));
 AO21x1_ASAP7_75t_R _34053_ (.A1(_05485_),
    .A2(_12749_),
    .B(_12752_),
    .Y(_12753_));
 BUFx4f_ASAP7_75t_R _34054_ (.A(_12753_),
    .Y(_12754_));
 AND2x2_ASAP7_75t_R _34055_ (.A(_05471_),
    .B(net176),
    .Y(_12755_));
 AO21x1_ASAP7_75t_R _34056_ (.A1(_05472_),
    .A2(net162),
    .B(_12755_),
    .Y(_12756_));
 INVx1_ASAP7_75t_R _34057_ (.A(_01663_),
    .Y(_12757_));
 NAND2x1_ASAP7_75t_R _34058_ (.A(_05471_),
    .B(_02225_),
    .Y(_12758_));
 OA211x2_ASAP7_75t_R _34059_ (.A1(_07308_),
    .A2(_12757_),
    .B(_12758_),
    .C(_05489_),
    .Y(_12759_));
 AO21x2_ASAP7_75t_R _34060_ (.A1(_05473_),
    .A2(_12756_),
    .B(_12759_),
    .Y(_12760_));
 AND2x2_ASAP7_75t_R _34061_ (.A(_05471_),
    .B(net174),
    .Y(_12761_));
 AO21x1_ASAP7_75t_R _34062_ (.A1(_05472_),
    .A2(net160),
    .B(_12761_),
    .Y(_12762_));
 INVx1_ASAP7_75t_R _34063_ (.A(_01665_),
    .Y(_12763_));
 NAND2x1_ASAP7_75t_R _34064_ (.A(_07308_),
    .B(_01603_),
    .Y(_12764_));
 OA211x2_ASAP7_75t_R _34065_ (.A1(_07308_),
    .A2(_12763_),
    .B(_12764_),
    .C(_05489_),
    .Y(_12765_));
 AO21x2_ASAP7_75t_R _34066_ (.A1(_05473_),
    .A2(_12762_),
    .B(_12765_),
    .Y(_12766_));
 AO21x1_ASAP7_75t_R _34067_ (.A1(_05473_),
    .A2(_12662_),
    .B(_12665_),
    .Y(_12767_));
 OR4x1_ASAP7_75t_R _34068_ (.A(_12760_),
    .B(_12766_),
    .C(_12659_),
    .D(_12767_),
    .Y(_12768_));
 OR2x2_ASAP7_75t_R _34069_ (.A(_12754_),
    .B(_12768_),
    .Y(_12769_));
 OR4x1_ASAP7_75t_R _34070_ (.A(_12747_),
    .B(_12691_),
    .C(_12769_),
    .D(_12714_),
    .Y(_12770_));
 INVx1_ASAP7_75t_R _34071_ (.A(_12770_),
    .Y(_12771_));
 OR3x1_ASAP7_75t_R _34072_ (.A(_12739_),
    .B(_12746_),
    .C(_12771_),
    .Y(_12772_));
 BUFx4f_ASAP7_75t_R _34073_ (.A(_05486_),
    .Y(_12773_));
 AOI21x1_ASAP7_75t_R _34074_ (.A1(_12773_),
    .A2(_12732_),
    .B(_12734_),
    .Y(_12774_));
 AO21x2_ASAP7_75t_R _34075_ (.A1(_05487_),
    .A2(_12640_),
    .B(_12643_),
    .Y(_12775_));
 AND2x2_ASAP7_75t_R _34076_ (.A(_12774_),
    .B(_12775_),
    .Y(_12776_));
 BUFx4f_ASAP7_75t_R _34077_ (.A(_12776_),
    .Y(_12777_));
 BUFx4f_ASAP7_75t_R _34078_ (.A(_12673_),
    .Y(_12778_));
 AND2x2_ASAP7_75t_R _34079_ (.A(_12742_),
    .B(_12690_),
    .Y(_12779_));
 INVx1_ASAP7_75t_R _34080_ (.A(_12769_),
    .Y(_12780_));
 INVx1_ASAP7_75t_R _34081_ (.A(_12728_),
    .Y(_12781_));
 BUFx4f_ASAP7_75t_R _34082_ (.A(_12740_),
    .Y(_12782_));
 BUFx4f_ASAP7_75t_R _34083_ (.A(_12743_),
    .Y(_12783_));
 AND3x1_ASAP7_75t_R _34084_ (.A(_12782_),
    .B(_12783_),
    .C(_12653_),
    .Y(_12784_));
 AND2x6_ASAP7_75t_R _34085_ (.A(_12673_),
    .B(_12679_),
    .Y(_12785_));
 AO21x1_ASAP7_75t_R _34086_ (.A1(_12781_),
    .A2(_12784_),
    .B(_12785_),
    .Y(_12786_));
 BUFx4f_ASAP7_75t_R _34087_ (.A(_12744_),
    .Y(_12787_));
 AO221x1_ASAP7_75t_R _34088_ (.A1(_12778_),
    .A2(_12779_),
    .B1(_12780_),
    .B2(_12786_),
    .C(_12787_),
    .Y(_12788_));
 AO32x1_ASAP7_75t_R _34089_ (.A1(_12646_),
    .A2(_12738_),
    .A3(_12772_),
    .B1(_12777_),
    .B2(_12788_),
    .Y(_12789_));
 BUFx4f_ASAP7_75t_R _34090_ (.A(_06859_),
    .Y(_12790_));
 BUFx4f_ASAP7_75t_R _34091_ (.A(_11955_),
    .Y(_12791_));
 AO21x1_ASAP7_75t_R _34092_ (.A1(_12790_),
    .A2(_12791_),
    .B(_14029_),
    .Y(_12792_));
 OA21x2_ASAP7_75t_R _34093_ (.A1(_12638_),
    .A2(_12789_),
    .B(_12792_),
    .Y(_04113_));
 BUFx6f_ASAP7_75t_R _34094_ (.A(_12637_),
    .Y(_12793_));
 OA21x2_ASAP7_75t_R _34095_ (.A1(_05479_),
    .A2(_05477_),
    .B(_05508_),
    .Y(_12794_));
 OAI21x1_ASAP7_75t_R _34096_ (.A1(_07313_),
    .A2(_12794_),
    .B(_05481_),
    .Y(_12795_));
 INVx1_ASAP7_75t_R _34097_ (.A(_01712_),
    .Y(_12796_));
 NOR2x1_ASAP7_75t_R _34098_ (.A(_01711_),
    .B(_05482_),
    .Y(_12797_));
 OR4x1_ASAP7_75t_R _34099_ (.A(_07313_),
    .B(_05508_),
    .C(_12796_),
    .D(_12797_),
    .Y(_12798_));
 AND3x2_ASAP7_75t_R _34100_ (.A(_12075_),
    .B(_12795_),
    .C(_12798_),
    .Y(_12799_));
 AO21x1_ASAP7_75t_R _34101_ (.A1(_05079_),
    .A2(_12793_),
    .B(_12799_),
    .Y(_04114_));
 BUFx6f_ASAP7_75t_R _34102_ (.A(_12080_),
    .Y(_12800_));
 OR3x1_ASAP7_75t_R _34103_ (.A(_11959_),
    .B(_05479_),
    .C(_11979_),
    .Y(_12801_));
 OA21x2_ASAP7_75t_R _34104_ (.A1(_05508_),
    .A2(_01711_),
    .B(_12801_),
    .Y(_12802_));
 OR4x2_ASAP7_75t_R _34105_ (.A(_07313_),
    .B(_12796_),
    .C(_12637_),
    .D(_12802_),
    .Y(_12803_));
 OAI21x1_ASAP7_75t_R _34106_ (.A1(_07787_),
    .A2(_12800_),
    .B(_12803_),
    .Y(_04115_));
 AND2x4_ASAP7_75t_R _34107_ (.A(_12735_),
    .B(_12775_),
    .Y(_12804_));
 NAND2x1_ASAP7_75t_R _34108_ (.A(_12075_),
    .B(_12804_),
    .Y(_12805_));
 OA21x2_ASAP7_75t_R _34109_ (.A1(_07777_),
    .A2(_12800_),
    .B(_12805_),
    .Y(_04116_));
 BUFx4f_ASAP7_75t_R _34110_ (.A(_12774_),
    .Y(_12806_));
 AND2x4_ASAP7_75t_R _34111_ (.A(_12740_),
    .B(_12743_),
    .Y(_12807_));
 AO21x1_ASAP7_75t_R _34112_ (.A1(_12807_),
    .A2(_12646_),
    .B(_12787_),
    .Y(_12808_));
 AND3x1_ASAP7_75t_R _34113_ (.A(_12075_),
    .B(_12806_),
    .C(_12808_),
    .Y(_12809_));
 AOI21x1_ASAP7_75t_R _34114_ (.A1(_13380_),
    .A2(_12638_),
    .B(_12809_),
    .Y(_04117_));
 BUFx4f_ASAP7_75t_R _34115_ (.A(_12074_),
    .Y(_12810_));
 INVx1_ASAP7_75t_R _34116_ (.A(_12777_),
    .Y(_12811_));
 OR3x1_ASAP7_75t_R _34117_ (.A(_12728_),
    .B(_12687_),
    .C(_12811_),
    .Y(_12812_));
 AND3x1_ASAP7_75t_R _34118_ (.A(_12735_),
    .B(_12783_),
    .C(_12644_),
    .Y(_12813_));
 OAI21x1_ASAP7_75t_R _34119_ (.A1(_12666_),
    .A2(_12813_),
    .B(_12787_),
    .Y(_12814_));
 AO21x1_ASAP7_75t_R _34120_ (.A1(_12736_),
    .A2(_12783_),
    .B(_12778_),
    .Y(_12815_));
 BUFx3_ASAP7_75t_R _34121_ (.A(_12782_),
    .Y(_12816_));
 OA21x2_ASAP7_75t_R _34122_ (.A1(_12774_),
    .A2(_12816_),
    .B(_12646_),
    .Y(_12817_));
 BUFx6f_ASAP7_75t_R _34123_ (.A(_12767_),
    .Y(_12818_));
 AO21x1_ASAP7_75t_R _34124_ (.A1(_12815_),
    .A2(_12817_),
    .B(_12818_),
    .Y(_12819_));
 AND4x1_ASAP7_75t_R _34125_ (.A(_12810_),
    .B(_12812_),
    .C(_12814_),
    .D(_12819_),
    .Y(_12820_));
 AO21x1_ASAP7_75t_R _34126_ (.A1(_14303_),
    .A2(_12793_),
    .B(_12820_),
    .Y(_04118_));
 INVx1_ASAP7_75t_R _34127_ (.A(_12660_),
    .Y(_12821_));
 BUFx3_ASAP7_75t_R _34128_ (.A(_12775_),
    .Y(_12822_));
 AND2x2_ASAP7_75t_R _34129_ (.A(_12774_),
    .B(_12693_),
    .Y(_12823_));
 AO221x1_ASAP7_75t_R _34130_ (.A1(_12747_),
    .A2(_12821_),
    .B1(_12781_),
    .B2(_12807_),
    .C(_12645_),
    .Y(_12824_));
 OA211x2_ASAP7_75t_R _34131_ (.A1(_12778_),
    .A2(_12822_),
    .B(_12823_),
    .C(_12824_),
    .Y(_12825_));
 AND3x1_ASAP7_75t_R _34132_ (.A(_12740_),
    .B(_12742_),
    .C(_12692_),
    .Y(_12826_));
 BUFx4f_ASAP7_75t_R _34133_ (.A(_12826_),
    .Y(_12827_));
 AND2x2_ASAP7_75t_R _34134_ (.A(_12659_),
    .B(_12818_),
    .Y(_12828_));
 AND3x4_ASAP7_75t_R _34135_ (.A(_12690_),
    .B(_12827_),
    .C(_12828_),
    .Y(_12829_));
 INVx1_ASAP7_75t_R _34136_ (.A(_12829_),
    .Y(_12830_));
 AND2x4_ASAP7_75t_R _34137_ (.A(_12735_),
    .B(_12644_),
    .Y(_12831_));
 OR3x1_ASAP7_75t_R _34138_ (.A(_12740_),
    .B(_12679_),
    .C(_12686_),
    .Y(_12832_));
 BUFx4f_ASAP7_75t_R _34139_ (.A(_12832_),
    .Y(_12833_));
 AND2x4_ASAP7_75t_R _34140_ (.A(_12831_),
    .B(_12833_),
    .Y(_12834_));
 AND3x1_ASAP7_75t_R _34141_ (.A(_12783_),
    .B(_12830_),
    .C(_12834_),
    .Y(_12835_));
 OR4x1_ASAP7_75t_R _34142_ (.A(_12023_),
    .B(_12821_),
    .C(_12825_),
    .D(_12835_),
    .Y(_12836_));
 OAI21x1_ASAP7_75t_R _34143_ (.A1(_14231_),
    .A2(_12800_),
    .B(_12836_),
    .Y(_04119_));
 BUFx4f_ASAP7_75t_R _34144_ (.A(_12691_),
    .Y(_12837_));
 NAND2x2_ASAP7_75t_R _34145_ (.A(_12659_),
    .B(_12818_),
    .Y(_12838_));
 BUFx4f_ASAP7_75t_R _34146_ (.A(_12707_),
    .Y(_12839_));
 AND2x2_ASAP7_75t_R _34147_ (.A(_12839_),
    .B(_12713_),
    .Y(_12840_));
 BUFx3_ASAP7_75t_R _34148_ (.A(_12694_),
    .Y(_12841_));
 OA21x2_ASAP7_75t_R _34149_ (.A1(_12838_),
    .A2(_12840_),
    .B(_12841_),
    .Y(_12842_));
 OA21x2_ASAP7_75t_R _34150_ (.A1(_12837_),
    .A2(_12842_),
    .B(_12807_),
    .Y(_12843_));
 AO21x1_ASAP7_75t_R _34151_ (.A1(_12782_),
    .A2(_12747_),
    .B(_12779_),
    .Y(_12844_));
 INVx1_ASAP7_75t_R _34152_ (.A(_12768_),
    .Y(_12845_));
 AND2x2_ASAP7_75t_R _34153_ (.A(_12753_),
    .B(_12845_),
    .Y(_12846_));
 NOR3x2_ASAP7_75t_R _34154_ (.B(_12729_),
    .C(_12846_),
    .Y(_12847_),
    .A(_12692_));
 BUFx4f_ASAP7_75t_R _34155_ (.A(_12847_),
    .Y(_12848_));
 BUFx4f_ASAP7_75t_R _34156_ (.A(_12720_),
    .Y(_12849_));
 AO22x1_ASAP7_75t_R _34157_ (.A1(_12787_),
    .A2(_12844_),
    .B1(_12848_),
    .B2(_12849_),
    .Y(_12850_));
 OA21x2_ASAP7_75t_R _34158_ (.A1(_12843_),
    .A2(_12850_),
    .B(_12834_),
    .Y(_12851_));
 AND3x2_ASAP7_75t_R _34159_ (.A(_12673_),
    .B(_12742_),
    .C(_12692_),
    .Y(_12852_));
 BUFx4f_ASAP7_75t_R _34160_ (.A(_12852_),
    .Y(_12853_));
 NAND2x1_ASAP7_75t_R _34161_ (.A(_12736_),
    .B(_12653_),
    .Y(_12854_));
 OA21x2_ASAP7_75t_R _34162_ (.A1(_12736_),
    .A2(_12853_),
    .B(_12854_),
    .Y(_12855_));
 AO32x1_ASAP7_75t_R _34163_ (.A1(_12806_),
    .A2(_12837_),
    .A3(_12808_),
    .B1(_12855_),
    .B2(_12822_),
    .Y(_12856_));
 OR3x2_ASAP7_75t_R _34164_ (.A(_12023_),
    .B(_12851_),
    .C(_12856_),
    .Y(_12857_));
 OA21x2_ASAP7_75t_R _34165_ (.A1(_13573_),
    .A2(_12800_),
    .B(_12857_),
    .Y(_04120_));
 NAND2x2_ASAP7_75t_R _34166_ (.A(_12735_),
    .B(_12644_),
    .Y(_12858_));
 AO21x1_ASAP7_75t_R _34167_ (.A1(_12653_),
    .A2(_12839_),
    .B(_12666_),
    .Y(_12859_));
 AND2x4_ASAP7_75t_R _34168_ (.A(_12742_),
    .B(_12686_),
    .Y(_12860_));
 AO32x1_ASAP7_75t_R _34169_ (.A1(_12660_),
    .A2(_12827_),
    .A3(_12859_),
    .B1(_12860_),
    .B2(_12837_),
    .Y(_12861_));
 AO21x1_ASAP7_75t_R _34170_ (.A1(_12701_),
    .A2(_12848_),
    .B(_12861_),
    .Y(_12862_));
 OA211x2_ASAP7_75t_R _34171_ (.A1(_12736_),
    .A2(_12783_),
    .B(_12841_),
    .C(_12858_),
    .Y(_12863_));
 INVx1_ASAP7_75t_R _34172_ (.A(_12863_),
    .Y(_12864_));
 OA211x2_ASAP7_75t_R _34173_ (.A1(_12858_),
    .A2(_12862_),
    .B(_12864_),
    .C(_12810_),
    .Y(_12865_));
 AO21x1_ASAP7_75t_R _34174_ (.A1(_13563_),
    .A2(_12793_),
    .B(_12865_),
    .Y(_04121_));
 AND2x2_ASAP7_75t_R _34175_ (.A(_12673_),
    .B(_12743_),
    .Y(_12866_));
 NOR2x1_ASAP7_75t_R _34176_ (.A(_12806_),
    .B(_12866_),
    .Y(_12867_));
 BUFx4f_ASAP7_75t_R _34177_ (.A(_12831_),
    .Y(_12868_));
 BUFx4f_ASAP7_75t_R _34178_ (.A(_12726_),
    .Y(_12869_));
 AO21x1_ASAP7_75t_R _34179_ (.A1(_12653_),
    .A2(_12714_),
    .B(_12838_),
    .Y(_12870_));
 AO222x2_ASAP7_75t_R _34180_ (.A1(_12869_),
    .A2(_12848_),
    .B1(_12870_),
    .B2(_12827_),
    .C1(_12860_),
    .C2(_12837_),
    .Y(_12871_));
 AND2x2_ASAP7_75t_R _34181_ (.A(_12747_),
    .B(_12858_),
    .Y(_12872_));
 AO21x1_ASAP7_75t_R _34182_ (.A1(_12868_),
    .A2(_12871_),
    .B(_12872_),
    .Y(_12873_));
 OA211x2_ASAP7_75t_R _34183_ (.A1(_12787_),
    .A2(_12867_),
    .B(_12873_),
    .C(_12810_),
    .Y(_12874_));
 AO21x1_ASAP7_75t_R _34184_ (.A1(_13567_),
    .A2(_12793_),
    .B(_12874_),
    .Y(_04122_));
 BUFx4f_ASAP7_75t_R _34185_ (.A(_12766_),
    .Y(_12875_));
 AND2x2_ASAP7_75t_R _34186_ (.A(_12680_),
    .B(_12693_),
    .Y(_12876_));
 BUFx4f_ASAP7_75t_R _34187_ (.A(_12876_),
    .Y(_12877_));
 AND2x2_ASAP7_75t_R _34188_ (.A(_12774_),
    .B(_12644_),
    .Y(_12878_));
 BUFx3_ASAP7_75t_R _34189_ (.A(_12878_),
    .Y(_12879_));
 NAND2x2_ASAP7_75t_R _34190_ (.A(_12680_),
    .B(_12693_),
    .Y(_12880_));
 AO21x1_ASAP7_75t_R _34191_ (.A1(_12880_),
    .A2(_12878_),
    .B(_12804_),
    .Y(_12881_));
 AO32x1_ASAP7_75t_R _34192_ (.A1(_12875_),
    .A2(_12877_),
    .A3(_12879_),
    .B1(_12881_),
    .B2(_12816_),
    .Y(_12882_));
 BUFx4f_ASAP7_75t_R _34193_ (.A(_12713_),
    .Y(_12883_));
 AND2x2_ASAP7_75t_R _34194_ (.A(_12690_),
    .B(_12686_),
    .Y(_12884_));
 AO21x1_ASAP7_75t_R _34195_ (.A1(_12875_),
    .A2(_12694_),
    .B(_12884_),
    .Y(_12885_));
 AND3x1_ASAP7_75t_R _34196_ (.A(_12743_),
    .B(_12691_),
    .C(_12828_),
    .Y(_12886_));
 AO21x1_ASAP7_75t_R _34197_ (.A1(_12680_),
    .A2(_12875_),
    .B(_12886_),
    .Y(_12887_));
 AO222x2_ASAP7_75t_R _34198_ (.A1(_12883_),
    .A2(_12848_),
    .B1(_12885_),
    .B2(_12783_),
    .C1(_12782_),
    .C2(_12887_),
    .Y(_12888_));
 NAND2x2_ASAP7_75t_R _34199_ (.A(_12652_),
    .B(_12728_),
    .Y(_12889_));
 AO21x1_ASAP7_75t_R _34200_ (.A1(_12875_),
    .A2(_12889_),
    .B(_12778_),
    .Y(_12890_));
 AND2x4_ASAP7_75t_R _34201_ (.A(_12742_),
    .B(_12692_),
    .Y(_12891_));
 AO22x1_ASAP7_75t_R _34202_ (.A1(_12782_),
    .A2(_12744_),
    .B1(_12890_),
    .B2(_12891_),
    .Y(_12892_));
 AO22x1_ASAP7_75t_R _34203_ (.A1(_12868_),
    .A2(_12888_),
    .B1(_12892_),
    .B2(_12777_),
    .Y(_12893_));
 OA21x2_ASAP7_75t_R _34204_ (.A1(_12875_),
    .A2(_12833_),
    .B(_12893_),
    .Y(_12894_));
 OR3x2_ASAP7_75t_R _34205_ (.A(_12023_),
    .B(_12882_),
    .C(_12894_),
    .Y(_12895_));
 OA21x2_ASAP7_75t_R _34206_ (.A1(_13945_),
    .A2(_12800_),
    .B(_12895_),
    .Y(_04123_));
 NAND2x2_ASAP7_75t_R _34207_ (.A(_12774_),
    .B(_12645_),
    .Y(_12896_));
 NOR2x1_ASAP7_75t_R _34208_ (.A(_05487_),
    .B(_01673_),
    .Y(_12897_));
 OA21x2_ASAP7_75t_R _34209_ (.A1(_05474_),
    .A2(_12897_),
    .B(_07312_),
    .Y(_12898_));
 AO21x1_ASAP7_75t_R _34210_ (.A1(_05484_),
    .A2(_12177_),
    .B(_12898_),
    .Y(_12899_));
 AO221x1_ASAP7_75t_R _34211_ (.A1(_12754_),
    .A2(_12877_),
    .B1(_12746_),
    .B2(_12899_),
    .C(_12853_),
    .Y(_12900_));
 AO21x1_ASAP7_75t_R _34212_ (.A1(_12736_),
    .A2(_12899_),
    .B(_12646_),
    .Y(_12901_));
 AO21x1_ASAP7_75t_R _34213_ (.A1(_12754_),
    .A2(_12889_),
    .B(_12687_),
    .Y(_12902_));
 OA211x2_ASAP7_75t_R _34214_ (.A1(_12693_),
    .A2(_12899_),
    .B(_12902_),
    .C(_12776_),
    .Y(_12903_));
 AO21x1_ASAP7_75t_R _34215_ (.A1(_12839_),
    .A2(_12785_),
    .B(_12779_),
    .Y(_12904_));
 AND3x2_ASAP7_75t_R _34216_ (.A(_12686_),
    .B(_12785_),
    .C(_12846_),
    .Y(_12905_));
 AO221x1_ASAP7_75t_R _34217_ (.A1(_12829_),
    .A2(_12899_),
    .B1(_12904_),
    .B2(_12744_),
    .C(_12905_),
    .Y(_12906_));
 OA21x2_ASAP7_75t_R _34218_ (.A1(_12903_),
    .A2(_12906_),
    .B(_12833_),
    .Y(_12907_));
 OR3x2_ASAP7_75t_R _34219_ (.A(_12673_),
    .B(_12652_),
    .C(_12838_),
    .Y(_12908_));
 AO21x1_ASAP7_75t_R _34220_ (.A1(_12693_),
    .A2(_12908_),
    .B(_12680_),
    .Y(_12909_));
 AND2x2_ASAP7_75t_R _34221_ (.A(_12729_),
    .B(_12909_),
    .Y(_12910_));
 OA21x2_ASAP7_75t_R _34222_ (.A1(_12906_),
    .A2(_12910_),
    .B(_12831_),
    .Y(_12911_));
 OA22x2_ASAP7_75t_R _34223_ (.A1(_12754_),
    .A2(_12907_),
    .B1(_12911_),
    .B2(_12903_),
    .Y(_12912_));
 AO21x1_ASAP7_75t_R _34224_ (.A1(_12858_),
    .A2(_12901_),
    .B(_12912_),
    .Y(_12913_));
 OA211x2_ASAP7_75t_R _34225_ (.A1(_12896_),
    .A2(_12900_),
    .B(_12913_),
    .C(_12810_),
    .Y(_12914_));
 AO21x1_ASAP7_75t_R _34226_ (.A1(_13777_),
    .A2(_12793_),
    .B(_12914_),
    .Y(_04124_));
 BUFx6f_ASAP7_75t_R _34227_ (.A(_05484_),
    .Y(_12915_));
 AO21x1_ASAP7_75t_R _34228_ (.A1(_12773_),
    .A2(net150),
    .B(_05475_),
    .Y(_12916_));
 AND2x2_ASAP7_75t_R _34229_ (.A(_07312_),
    .B(_12916_),
    .Y(_12917_));
 AO21x1_ASAP7_75t_R _34230_ (.A1(_12915_),
    .A2(_12216_),
    .B(_12917_),
    .Y(_12918_));
 AO21x1_ASAP7_75t_R _34231_ (.A1(_12746_),
    .A2(_12879_),
    .B(_12804_),
    .Y(_12919_));
 OA21x2_ASAP7_75t_R _34232_ (.A1(_12847_),
    .A2(_12860_),
    .B(_12691_),
    .Y(_12920_));
 AO221x1_ASAP7_75t_R _34233_ (.A1(_12760_),
    .A2(_12910_),
    .B1(_12918_),
    .B2(_12829_),
    .C(_12920_),
    .Y(_12921_));
 AND4x1_ASAP7_75t_R _34234_ (.A(_12760_),
    .B(_12693_),
    .C(_12807_),
    .D(_12889_),
    .Y(_12922_));
 AO21x1_ASAP7_75t_R _34235_ (.A1(_12744_),
    .A2(_12918_),
    .B(_12853_),
    .Y(_12923_));
 OA21x2_ASAP7_75t_R _34236_ (.A1(_12922_),
    .A2(_12923_),
    .B(_12777_),
    .Y(_12924_));
 AO21x1_ASAP7_75t_R _34237_ (.A1(_12868_),
    .A2(_12921_),
    .B(_12924_),
    .Y(_12925_));
 AO21x1_ASAP7_75t_R _34238_ (.A1(_12877_),
    .A2(_12879_),
    .B(_12925_),
    .Y(_12926_));
 AO21x1_ASAP7_75t_R _34239_ (.A1(_12833_),
    .A2(_12925_),
    .B(_12760_),
    .Y(_12927_));
 AO221x2_ASAP7_75t_R _34240_ (.A1(_12918_),
    .A2(_12919_),
    .B1(_12926_),
    .B2(_12927_),
    .C(_12637_),
    .Y(_12928_));
 OA21x2_ASAP7_75t_R _34241_ (.A1(_14732_),
    .A2(_12800_),
    .B(_12928_),
    .Y(_04125_));
 NAND2x1_ASAP7_75t_R _34242_ (.A(_05487_),
    .B(_12331_),
    .Y(_12929_));
 OA211x2_ASAP7_75t_R _34243_ (.A1(_12773_),
    .A2(_12717_),
    .B(_12929_),
    .C(_07312_),
    .Y(_12930_));
 AO21x2_ASAP7_75t_R _34244_ (.A1(_05484_),
    .A2(_12255_),
    .B(_12930_),
    .Y(_12931_));
 AO21x1_ASAP7_75t_R _34245_ (.A1(_12816_),
    .A2(_12931_),
    .B(_12877_),
    .Y(_12932_));
 AOI21x1_ASAP7_75t_R _34246_ (.A1(_12827_),
    .A2(_12889_),
    .B(_12853_),
    .Y(_12933_));
 NOR3x1_ASAP7_75t_R _34247_ (.A(_12666_),
    .B(_12646_),
    .C(_12933_),
    .Y(_12934_));
 AO221x1_ASAP7_75t_R _34248_ (.A1(_12787_),
    .A2(_12931_),
    .B1(_12932_),
    .B2(_12646_),
    .C(_12934_),
    .Y(_12935_));
 INVx1_ASAP7_75t_R _34249_ (.A(_12931_),
    .Y(_12936_));
 OAI21x1_ASAP7_75t_R _34250_ (.A1(_12847_),
    .A2(_12860_),
    .B(_12690_),
    .Y(_12937_));
 OAI21x1_ASAP7_75t_R _34251_ (.A1(_12908_),
    .A2(_12931_),
    .B(_12693_),
    .Y(_12938_));
 AO21x1_ASAP7_75t_R _34252_ (.A1(_12743_),
    .A2(_12938_),
    .B(_12785_),
    .Y(_12939_));
 AO221x1_ASAP7_75t_R _34253_ (.A1(_12666_),
    .A2(_12853_),
    .B1(_12937_),
    .B2(_12939_),
    .C(_12775_),
    .Y(_12940_));
 OA211x2_ASAP7_75t_R _34254_ (.A1(_12646_),
    .A2(_12936_),
    .B(_12940_),
    .C(_12736_),
    .Y(_12941_));
 INVx1_ASAP7_75t_R _34255_ (.A(_12941_),
    .Y(_12942_));
 OA211x2_ASAP7_75t_R _34256_ (.A1(_12739_),
    .A2(_12935_),
    .B(_12942_),
    .C(_12810_),
    .Y(_12943_));
 AO21x1_ASAP7_75t_R _34257_ (.A1(_13857_),
    .A2(_12793_),
    .B(_12943_),
    .Y(_04126_));
 AND2x4_ASAP7_75t_R _34258_ (.A(_12745_),
    .B(_12878_),
    .Y(_12944_));
 NOR2x1_ASAP7_75t_R _34259_ (.A(_12804_),
    .B(_12944_),
    .Y(_12945_));
 NAND2x1_ASAP7_75t_R _34260_ (.A(_05487_),
    .B(_12337_),
    .Y(_12946_));
 OA211x2_ASAP7_75t_R _34261_ (.A1(_12773_),
    .A2(_12697_),
    .B(_12946_),
    .C(_07312_),
    .Y(_12947_));
 AOI21x1_ASAP7_75t_R _34262_ (.A1(_12915_),
    .A2(_12293_),
    .B(_12947_),
    .Y(_12948_));
 OA211x2_ASAP7_75t_R _34263_ (.A1(_12830_),
    .A2(_12948_),
    .B(_12937_),
    .C(_12833_),
    .Y(_12949_));
 OR2x2_ASAP7_75t_R _34264_ (.A(_12858_),
    .B(_12949_),
    .Y(_12950_));
 OR2x2_ASAP7_75t_R _34265_ (.A(_12694_),
    .B(_12948_),
    .Y(_12951_));
 AO21x1_ASAP7_75t_R _34266_ (.A1(_12950_),
    .A2(_12951_),
    .B(_12853_),
    .Y(_12952_));
 AO21x1_ASAP7_75t_R _34267_ (.A1(_12933_),
    .A2(_12951_),
    .B(_12811_),
    .Y(_12953_));
 AO22x1_ASAP7_75t_R _34268_ (.A1(_12821_),
    .A2(_12952_),
    .B1(_12953_),
    .B2(_12950_),
    .Y(_12954_));
 OA211x2_ASAP7_75t_R _34269_ (.A1(_12945_),
    .A2(_12948_),
    .B(_12954_),
    .C(_12080_),
    .Y(_12955_));
 AOI21x1_ASAP7_75t_R _34270_ (.A1(_15025_),
    .A2(_12638_),
    .B(_12955_),
    .Y(_04127_));
 AOI211x1_ASAP7_75t_R _34271_ (.A1(_12868_),
    .A2(_12829_),
    .B(_12944_),
    .C(_12018_),
    .Y(_12956_));
 AO21x1_ASAP7_75t_R _34272_ (.A1(_13555_),
    .A2(_12117_),
    .B(_12956_),
    .Y(_04128_));
 NAND2x1_ASAP7_75t_R _34273_ (.A(_12740_),
    .B(_12743_),
    .Y(_12957_));
 AO21x1_ASAP7_75t_R _34274_ (.A1(_12690_),
    .A2(_12828_),
    .B(_12957_),
    .Y(_12958_));
 NAND2x1_ASAP7_75t_R _34275_ (.A(_12729_),
    .B(_12958_),
    .Y(_12959_));
 NAND2x1_ASAP7_75t_R _34276_ (.A(_12773_),
    .B(_12342_),
    .Y(_12960_));
 OA211x2_ASAP7_75t_R _34277_ (.A1(_11958_),
    .A2(_12723_),
    .B(_12960_),
    .C(_07312_),
    .Y(_12961_));
 AO21x1_ASAP7_75t_R _34278_ (.A1(_12915_),
    .A2(_12330_),
    .B(_12961_),
    .Y(_12962_));
 AO32x1_ASAP7_75t_R _34279_ (.A1(_12694_),
    .A2(_12849_),
    .A3(_12959_),
    .B1(_12962_),
    .B2(_12829_),
    .Y(_12963_));
 OR3x1_ASAP7_75t_R _34280_ (.A(_12853_),
    .B(_12920_),
    .C(_12963_),
    .Y(_12964_));
 OR3x2_ASAP7_75t_R _34281_ (.A(_12652_),
    .B(_12753_),
    .C(_12768_),
    .Y(_12965_));
 INVx1_ASAP7_75t_R _34282_ (.A(_12720_),
    .Y(_12966_));
 OAI21x1_ASAP7_75t_R _34283_ (.A1(_12728_),
    .A2(_12965_),
    .B(_12966_),
    .Y(_12967_));
 AO221x1_ASAP7_75t_R _34284_ (.A1(_12741_),
    .A2(_12849_),
    .B1(_12967_),
    .B2(_12743_),
    .C(_12744_),
    .Y(_12968_));
 OA211x2_ASAP7_75t_R _34285_ (.A1(_12694_),
    .A2(_12962_),
    .B(_12968_),
    .C(_12777_),
    .Y(_12969_));
 AO21x1_ASAP7_75t_R _34286_ (.A1(_12868_),
    .A2(_12964_),
    .B(_12969_),
    .Y(_12970_));
 OA21x2_ASAP7_75t_R _34287_ (.A1(_12849_),
    .A2(_12833_),
    .B(_12970_),
    .Y(_12971_));
 AO32x1_ASAP7_75t_R _34288_ (.A1(_12816_),
    .A2(_12849_),
    .A3(_12877_),
    .B1(_12745_),
    .B2(_12962_),
    .Y(_12972_));
 AO22x1_ASAP7_75t_R _34289_ (.A1(_12804_),
    .A2(_12962_),
    .B1(_12972_),
    .B2(_12879_),
    .Y(_12973_));
 OR3x2_ASAP7_75t_R _34290_ (.A(_12023_),
    .B(_12971_),
    .C(_12973_),
    .Y(_12974_));
 OA21x2_ASAP7_75t_R _34291_ (.A1(net19),
    .A2(_12800_),
    .B(_12974_),
    .Y(_04129_));
 AO21x1_ASAP7_75t_R _34292_ (.A1(_12784_),
    .A2(_12840_),
    .B(_12785_),
    .Y(_12975_));
 AND2x2_ASAP7_75t_R _34293_ (.A(_12826_),
    .B(_12828_),
    .Y(_12976_));
 NAND2x1_ASAP7_75t_R _34294_ (.A(_11959_),
    .B(_12348_),
    .Y(_12977_));
 OA211x2_ASAP7_75t_R _34295_ (.A1(_11959_),
    .A2(_12710_),
    .B(_12977_),
    .C(_07313_),
    .Y(_12978_));
 AO21x1_ASAP7_75t_R _34296_ (.A1(_12915_),
    .A2(_12378_),
    .B(_12978_),
    .Y(_12979_));
 AO21x1_ASAP7_75t_R _34297_ (.A1(_12976_),
    .A2(_12979_),
    .B(_12848_),
    .Y(_12980_));
 AO32x1_ASAP7_75t_R _34298_ (.A1(_12841_),
    .A2(_12701_),
    .A3(_12975_),
    .B1(_12980_),
    .B2(_12837_),
    .Y(_12981_));
 OA21x2_ASAP7_75t_R _34299_ (.A1(_12691_),
    .A2(_12840_),
    .B(_12828_),
    .Y(_12982_));
 AND3x1_ASAP7_75t_R _34300_ (.A(_12741_),
    .B(_12694_),
    .C(_12982_),
    .Y(_12983_));
 INVx1_ASAP7_75t_R _34301_ (.A(_12983_),
    .Y(_12984_));
 AO32x1_ASAP7_75t_R _34302_ (.A1(_12729_),
    .A2(_12775_),
    .A3(_12823_),
    .B1(_12984_),
    .B2(_12813_),
    .Y(_12985_));
 AO32x1_ASAP7_75t_R _34303_ (.A1(_12816_),
    .A2(_12701_),
    .A3(_12877_),
    .B1(_12745_),
    .B2(_12979_),
    .Y(_12986_));
 NOR2x2_ASAP7_75t_R _34304_ (.A(_12644_),
    .B(_12823_),
    .Y(_12987_));
 AO222x2_ASAP7_75t_R _34305_ (.A1(_12701_),
    .A2(_12985_),
    .B1(_12986_),
    .B2(_12879_),
    .C1(_12987_),
    .C2(_12979_),
    .Y(_12988_));
 AO21x1_ASAP7_75t_R _34306_ (.A1(_12834_),
    .A2(_12981_),
    .B(_12988_),
    .Y(_12989_));
 AO21x1_ASAP7_75t_R _34307_ (.A1(_12790_),
    .A2(_12791_),
    .B(_15502_),
    .Y(_12990_));
 OA21x2_ASAP7_75t_R _34308_ (.A1(_12638_),
    .A2(_12989_),
    .B(_12990_),
    .Y(_04130_));
 NAND2x1_ASAP7_75t_R _34309_ (.A(_12673_),
    .B(_12693_),
    .Y(_12991_));
 NAND2x1_ASAP7_75t_R _34310_ (.A(_12880_),
    .B(_12991_),
    .Y(_12992_));
 OR3x1_ASAP7_75t_R _34311_ (.A(_12778_),
    .B(_12783_),
    .C(_12869_),
    .Y(_12993_));
 OA21x2_ASAP7_75t_R _34312_ (.A1(_12782_),
    .A2(_12839_),
    .B(_12645_),
    .Y(_12994_));
 AO21x1_ASAP7_75t_R _34313_ (.A1(_12993_),
    .A2(_12994_),
    .B(_12787_),
    .Y(_12995_));
 NAND2x1_ASAP7_75t_R _34314_ (.A(_11958_),
    .B(_12352_),
    .Y(_12996_));
 OA211x2_ASAP7_75t_R _34315_ (.A1(_11959_),
    .A2(_12704_),
    .B(_12996_),
    .C(_07313_),
    .Y(_12997_));
 AO21x2_ASAP7_75t_R _34316_ (.A1(_12915_),
    .A2(_12403_),
    .B(_12997_),
    .Y(_12998_));
 AO32x1_ASAP7_75t_R _34317_ (.A1(_12992_),
    .A2(_12993_),
    .A3(_12994_),
    .B1(_12995_),
    .B2(_12998_),
    .Y(_12999_));
 AO21x1_ASAP7_75t_R _34318_ (.A1(_12976_),
    .A2(_12998_),
    .B(_12848_),
    .Y(_13000_));
 AND4x1_ASAP7_75t_R _34319_ (.A(_12653_),
    .B(_12869_),
    .C(_12827_),
    .D(_12840_),
    .Y(_13001_));
 AO21x1_ASAP7_75t_R _34320_ (.A1(_12837_),
    .A2(_13000_),
    .B(_13001_),
    .Y(_13002_));
 NAND2x1_ASAP7_75t_R _34321_ (.A(_12694_),
    .B(_12982_),
    .Y(_13003_));
 AO21x1_ASAP7_75t_R _34322_ (.A1(_12778_),
    .A2(_12831_),
    .B(_12777_),
    .Y(_13004_));
 AO32x1_ASAP7_75t_R _34323_ (.A1(_12783_),
    .A2(_12868_),
    .A3(_13003_),
    .B1(_13004_),
    .B2(_12841_),
    .Y(_13005_));
 AO222x2_ASAP7_75t_R _34324_ (.A1(_12804_),
    .A2(_12998_),
    .B1(_13002_),
    .B2(_12834_),
    .C1(_13005_),
    .C2(_12869_),
    .Y(_13006_));
 AO21x1_ASAP7_75t_R _34325_ (.A1(_12806_),
    .A2(_12999_),
    .B(_13006_),
    .Y(_13007_));
 AO21x1_ASAP7_75t_R _34326_ (.A1(_12790_),
    .A2(_12791_),
    .B(_15529_),
    .Y(_13008_));
 OA21x2_ASAP7_75t_R _34327_ (.A1(_12638_),
    .A2(_13007_),
    .B(_13008_),
    .Y(_04131_));
 AO21x1_ASAP7_75t_R _34328_ (.A1(_12807_),
    .A2(_12838_),
    .B(_12785_),
    .Y(_13009_));
 NAND2x1_ASAP7_75t_R _34329_ (.A(_12773_),
    .B(_12356_),
    .Y(_13010_));
 OA211x2_ASAP7_75t_R _34330_ (.A1(_11958_),
    .A2(_12763_),
    .B(_13010_),
    .C(_07312_),
    .Y(_13011_));
 AO21x2_ASAP7_75t_R _34331_ (.A1(_05484_),
    .A2(_12418_),
    .B(_13011_),
    .Y(_13012_));
 OR2x2_ASAP7_75t_R _34332_ (.A(_12653_),
    .B(_13012_),
    .Y(_13013_));
 AO32x1_ASAP7_75t_R _34333_ (.A1(_12841_),
    .A2(_12883_),
    .A3(_13009_),
    .B1(_13013_),
    .B2(_12976_),
    .Y(_13014_));
 AO21x1_ASAP7_75t_R _34334_ (.A1(_12837_),
    .A2(_12848_),
    .B(_13014_),
    .Y(_13015_));
 OR3x1_ASAP7_75t_R _34335_ (.A(_12741_),
    .B(_12818_),
    .C(_12880_),
    .Y(_13016_));
 OA211x2_ASAP7_75t_R _34336_ (.A1(_12992_),
    .A2(_13012_),
    .B(_13016_),
    .C(_12878_),
    .Y(_13017_));
 AND4x1_ASAP7_75t_R _34337_ (.A(_12782_),
    .B(_12883_),
    .C(_12876_),
    .D(_12777_),
    .Y(_13018_));
 AO221x1_ASAP7_75t_R _34338_ (.A1(_12987_),
    .A2(_13012_),
    .B1(_13017_),
    .B2(_12833_),
    .C(_13018_),
    .Y(_13019_));
 AO21x1_ASAP7_75t_R _34339_ (.A1(_12834_),
    .A2(_13015_),
    .B(_13019_),
    .Y(_13020_));
 NAND2x1_ASAP7_75t_R _34340_ (.A(_12782_),
    .B(_12747_),
    .Y(_13021_));
 NAND2x2_ASAP7_75t_R _34341_ (.A(_12741_),
    .B(_12693_),
    .Y(_13022_));
 AO32x1_ASAP7_75t_R _34342_ (.A1(_12775_),
    .A2(_12823_),
    .A3(_13021_),
    .B1(_13022_),
    .B2(_12813_),
    .Y(_13023_));
 OA21x2_ASAP7_75t_R _34343_ (.A1(_13017_),
    .A2(_13023_),
    .B(_12883_),
    .Y(_13024_));
 OR3x2_ASAP7_75t_R _34344_ (.A(_12023_),
    .B(_13020_),
    .C(_13024_),
    .Y(_13025_));
 OA21x2_ASAP7_75t_R _34345_ (.A1(_15499_),
    .A2(_12800_),
    .B(_13025_),
    .Y(_04132_));
 NAND2x1_ASAP7_75t_R _34346_ (.A(_05486_),
    .B(_12360_),
    .Y(_13026_));
 OA211x2_ASAP7_75t_R _34347_ (.A1(_05486_),
    .A2(_12750_),
    .B(_13026_),
    .C(_07311_),
    .Y(_13027_));
 AO21x2_ASAP7_75t_R _34348_ (.A1(_05484_),
    .A2(_12433_),
    .B(_13027_),
    .Y(_13028_));
 AND2x4_ASAP7_75t_R _34349_ (.A(_12673_),
    .B(_12692_),
    .Y(_13029_));
 AO21x1_ASAP7_75t_R _34350_ (.A1(_12827_),
    .A2(_12838_),
    .B(_13029_),
    .Y(_13030_));
 OA21x2_ASAP7_75t_R _34351_ (.A1(_12905_),
    .A2(_13030_),
    .B(_12839_),
    .Y(_13031_));
 AO21x1_ASAP7_75t_R _34352_ (.A1(_12976_),
    .A2(_13028_),
    .B(_12847_),
    .Y(_13032_));
 AO221x1_ASAP7_75t_R _34353_ (.A1(_12660_),
    .A2(_12860_),
    .B1(_13032_),
    .B2(_12690_),
    .C(_12852_),
    .Y(_13033_));
 OA21x2_ASAP7_75t_R _34354_ (.A1(_13031_),
    .A2(_13033_),
    .B(_12831_),
    .Y(_13034_));
 OA21x2_ASAP7_75t_R _34355_ (.A1(_12694_),
    .A2(_13028_),
    .B(_12777_),
    .Y(_13035_));
 OA21x2_ASAP7_75t_R _34356_ (.A1(_12741_),
    .A2(_12680_),
    .B(_13034_),
    .Y(_13036_));
 OR3x1_ASAP7_75t_R _34357_ (.A(_12744_),
    .B(_12839_),
    .C(_13036_),
    .Y(_13037_));
 OA21x2_ASAP7_75t_R _34358_ (.A1(_13034_),
    .A2(_13035_),
    .B(_13037_),
    .Y(_13038_));
 AO21x1_ASAP7_75t_R _34359_ (.A1(_12739_),
    .A2(_13028_),
    .B(_13038_),
    .Y(_13039_));
 AO32x1_ASAP7_75t_R _34360_ (.A1(_12778_),
    .A2(_12660_),
    .A3(_12841_),
    .B1(_12746_),
    .B2(_13028_),
    .Y(_13040_));
 AO22x1_ASAP7_75t_R _34361_ (.A1(_12739_),
    .A2(_13038_),
    .B1(_13040_),
    .B2(_12879_),
    .Y(_13041_));
 AO21x1_ASAP7_75t_R _34362_ (.A1(_12822_),
    .A2(_13039_),
    .B(_13041_),
    .Y(_13042_));
 AO21x1_ASAP7_75t_R _34363_ (.A1(_12790_),
    .A2(_12791_),
    .B(_15745_),
    .Y(_13043_));
 OA21x2_ASAP7_75t_R _34364_ (.A1(_12638_),
    .A2(_13042_),
    .B(_13043_),
    .Y(_04133_));
 NAND2x1_ASAP7_75t_R _34365_ (.A(_12773_),
    .B(_12364_),
    .Y(_13044_));
 OA211x2_ASAP7_75t_R _34366_ (.A1(_11958_),
    .A2(_12757_),
    .B(_13044_),
    .C(_07312_),
    .Y(_13045_));
 AO21x1_ASAP7_75t_R _34367_ (.A1(_12915_),
    .A2(_12442_),
    .B(_13045_),
    .Y(_13046_));
 OR3x1_ASAP7_75t_R _34368_ (.A(_12877_),
    .B(_13029_),
    .C(_13046_),
    .Y(_13047_));
 OA21x2_ASAP7_75t_R _34369_ (.A1(_12837_),
    .A2(_12746_),
    .B(_13047_),
    .Y(_13048_));
 OA21x2_ASAP7_75t_R _34370_ (.A1(_12691_),
    .A2(_12833_),
    .B(_12831_),
    .Y(_13049_));
 OA22x2_ASAP7_75t_R _34371_ (.A1(_12691_),
    .A2(_12852_),
    .B1(_12847_),
    .B2(_13029_),
    .Y(_13050_));
 AND3x2_ASAP7_75t_R _34372_ (.A(_12690_),
    .B(_12660_),
    .C(_12827_),
    .Y(_13051_));
 OA21x2_ASAP7_75t_R _34373_ (.A1(_12666_),
    .A2(_13046_),
    .B(_13051_),
    .Y(_13052_));
 NOR2x2_ASAP7_75t_R _34374_ (.A(_12785_),
    .B(_12891_),
    .Y(_13053_));
 OA21x2_ASAP7_75t_R _34375_ (.A1(_12905_),
    .A2(_13053_),
    .B(_12849_),
    .Y(_13054_));
 OR3x1_ASAP7_75t_R _34376_ (.A(_13050_),
    .B(_13052_),
    .C(_13054_),
    .Y(_13055_));
 AND2x2_ASAP7_75t_R _34377_ (.A(_12680_),
    .B(_12690_),
    .Y(_13056_));
 AO21x1_ASAP7_75t_R _34378_ (.A1(_12841_),
    .A2(_13056_),
    .B(_12645_),
    .Y(_13057_));
 AO222x2_ASAP7_75t_R _34379_ (.A1(_12987_),
    .A2(_13046_),
    .B1(_13049_),
    .B2(_13055_),
    .C1(_13057_),
    .C2(_12806_),
    .Y(_13058_));
 OA211x2_ASAP7_75t_R _34380_ (.A1(_12896_),
    .A2(_13048_),
    .B(_13058_),
    .C(_12810_),
    .Y(_13059_));
 AO21x1_ASAP7_75t_R _34381_ (.A1(_13602_),
    .A2(_12117_),
    .B(_13059_),
    .Y(_04134_));
 AND2x2_ASAP7_75t_R _34382_ (.A(_12680_),
    .B(_12883_),
    .Y(_13060_));
 AO21x1_ASAP7_75t_R _34383_ (.A1(_12875_),
    .A2(_12866_),
    .B(_13060_),
    .Y(_13061_));
 NAND2x1_ASAP7_75t_R _34384_ (.A(_05486_),
    .B(_12368_),
    .Y(_13062_));
 OA211x2_ASAP7_75t_R _34385_ (.A1(_12773_),
    .A2(_12663_),
    .B(_13062_),
    .C(_07311_),
    .Y(_13063_));
 AO21x1_ASAP7_75t_R _34386_ (.A1(_05484_),
    .A2(_12180_),
    .B(_13063_),
    .Y(_13064_));
 AO221x1_ASAP7_75t_R _34387_ (.A1(_12841_),
    .A2(_13061_),
    .B1(_13064_),
    .B2(_12746_),
    .C(_12896_),
    .Y(_13065_));
 AO32x1_ASAP7_75t_R _34388_ (.A1(_12754_),
    .A2(_12845_),
    .A3(_13060_),
    .B1(_12766_),
    .B2(_12743_),
    .Y(_13066_));
 AO32x1_ASAP7_75t_R _34389_ (.A1(_12741_),
    .A2(_12680_),
    .A3(_12883_),
    .B1(_13066_),
    .B2(_12744_),
    .Y(_13067_));
 AND2x2_ASAP7_75t_R _34390_ (.A(_12673_),
    .B(_12720_),
    .Y(_13068_));
 AO21x1_ASAP7_75t_R _34391_ (.A1(_12741_),
    .A2(_12766_),
    .B(_13068_),
    .Y(_13069_));
 AO21x1_ASAP7_75t_R _34392_ (.A1(_12876_),
    .A2(_13069_),
    .B(_12645_),
    .Y(_13070_));
 AO32x1_ASAP7_75t_R _34393_ (.A1(_12831_),
    .A2(_12833_),
    .A3(_13067_),
    .B1(_13070_),
    .B2(_12774_),
    .Y(_13071_));
 OA211x2_ASAP7_75t_R _34394_ (.A1(_12666_),
    .A2(_13064_),
    .B(_12827_),
    .C(_12660_),
    .Y(_13072_));
 OR3x1_ASAP7_75t_R _34395_ (.A(_13029_),
    .B(_12848_),
    .C(_13072_),
    .Y(_13073_));
 AO32x1_ASAP7_75t_R _34396_ (.A1(_12837_),
    .A2(_12645_),
    .A3(_13073_),
    .B1(_13064_),
    .B2(_12987_),
    .Y(_13074_));
 OR2x2_ASAP7_75t_R _34397_ (.A(_13071_),
    .B(_13074_),
    .Y(_13075_));
 AND3x1_ASAP7_75t_R _34398_ (.A(_12075_),
    .B(_13065_),
    .C(_13075_),
    .Y(_13076_));
 AO21x1_ASAP7_75t_R _34399_ (.A1(_14059_),
    .A2(_12117_),
    .B(_13076_),
    .Y(_04135_));
 NAND2x1_ASAP7_75t_R _34400_ (.A(_05487_),
    .B(_12372_),
    .Y(_13077_));
 OA211x2_ASAP7_75t_R _34401_ (.A1(_12773_),
    .A2(_12656_),
    .B(_13077_),
    .C(_07312_),
    .Y(_13078_));
 AO21x1_ASAP7_75t_R _34402_ (.A1(_05484_),
    .A2(_12184_),
    .B(_13078_),
    .Y(_13079_));
 AND2x2_ASAP7_75t_R _34403_ (.A(_12741_),
    .B(_12754_),
    .Y(_13080_));
 AO21x1_ASAP7_75t_R _34404_ (.A1(_12778_),
    .A2(_12701_),
    .B(_13080_),
    .Y(_13081_));
 AO21x1_ASAP7_75t_R _34405_ (.A1(_12877_),
    .A2(_13081_),
    .B(_12645_),
    .Y(_13082_));
 OA21x2_ASAP7_75t_R _34406_ (.A1(_12666_),
    .A2(_13079_),
    .B(_13051_),
    .Y(_13083_));
 AO221x1_ASAP7_75t_R _34407_ (.A1(_12701_),
    .A2(_12905_),
    .B1(_13053_),
    .B2(_12839_),
    .C(_13083_),
    .Y(_13084_));
 OA21x2_ASAP7_75t_R _34408_ (.A1(_13050_),
    .A2(_13084_),
    .B(_13049_),
    .Y(_13085_));
 AO221x1_ASAP7_75t_R _34409_ (.A1(_12987_),
    .A2(_13079_),
    .B1(_13082_),
    .B2(_12806_),
    .C(_13085_),
    .Y(_13086_));
 AO221x1_ASAP7_75t_R _34410_ (.A1(_12754_),
    .A2(_12853_),
    .B1(_13079_),
    .B2(_12746_),
    .C(_12896_),
    .Y(_13087_));
 AND3x2_ASAP7_75t_R _34411_ (.A(_12075_),
    .B(_13086_),
    .C(_13087_),
    .Y(_13088_));
 AO21x1_ASAP7_75t_R _34412_ (.A1(_14487_),
    .A2(_12117_),
    .B(_13088_),
    .Y(_04136_));
 NAND2x1_ASAP7_75t_R _34413_ (.A(_11958_),
    .B(_12379_),
    .Y(_13089_));
 OA211x2_ASAP7_75t_R _34414_ (.A1(_11958_),
    .A2(_12649_),
    .B(_13089_),
    .C(_07313_),
    .Y(_13090_));
 AO21x1_ASAP7_75t_R _34415_ (.A1(_12915_),
    .A2(_12187_),
    .B(_13090_),
    .Y(_13091_));
 AO221x1_ASAP7_75t_R _34416_ (.A1(_12760_),
    .A2(_12853_),
    .B1(_13091_),
    .B2(_12746_),
    .C(_12896_),
    .Y(_13092_));
 OA21x2_ASAP7_75t_R _34417_ (.A1(_12666_),
    .A2(_13091_),
    .B(_13051_),
    .Y(_13093_));
 AO32x1_ASAP7_75t_R _34418_ (.A1(_12743_),
    .A2(_12760_),
    .A3(_12744_),
    .B1(_13056_),
    .B2(_12741_),
    .Y(_13094_));
 AO21x1_ASAP7_75t_R _34419_ (.A1(_12869_),
    .A2(_12905_),
    .B(_13094_),
    .Y(_13095_));
 OR3x1_ASAP7_75t_R _34420_ (.A(_13050_),
    .B(_13093_),
    .C(_13095_),
    .Y(_13096_));
 AO221x1_ASAP7_75t_R _34421_ (.A1(_12987_),
    .A2(_13091_),
    .B1(_13096_),
    .B2(_13049_),
    .C(_12879_),
    .Y(_13097_));
 AND3x1_ASAP7_75t_R _34422_ (.A(_12075_),
    .B(_13092_),
    .C(_13097_),
    .Y(_13098_));
 AO21x1_ASAP7_75t_R _34423_ (.A1(_14546_),
    .A2(_12117_),
    .B(_13098_),
    .Y(_04137_));
 NAND2x1_ASAP7_75t_R _34424_ (.A(_11958_),
    .B(_12383_),
    .Y(_13099_));
 OA211x2_ASAP7_75t_R _34425_ (.A1(_11958_),
    .A2(_12683_),
    .B(_13099_),
    .C(_07313_),
    .Y(_13100_));
 AO21x1_ASAP7_75t_R _34426_ (.A1(_12915_),
    .A2(_12190_),
    .B(_13100_),
    .Y(_13101_));
 AO221x1_ASAP7_75t_R _34427_ (.A1(_12818_),
    .A2(_12853_),
    .B1(_13101_),
    .B2(_12746_),
    .C(_12896_),
    .Y(_13102_));
 OA211x2_ASAP7_75t_R _34428_ (.A1(_12818_),
    .A2(_12694_),
    .B(_13022_),
    .C(_12783_),
    .Y(_13103_));
 OA21x2_ASAP7_75t_R _34429_ (.A1(_12666_),
    .A2(_13101_),
    .B(_13051_),
    .Y(_13104_));
 OR3x1_ASAP7_75t_R _34430_ (.A(_13056_),
    .B(_13103_),
    .C(_13104_),
    .Y(_13105_));
 AO221x1_ASAP7_75t_R _34431_ (.A1(_12987_),
    .A2(_13101_),
    .B1(_13105_),
    .B2(_13049_),
    .C(_12879_),
    .Y(_13106_));
 AND3x1_ASAP7_75t_R _34432_ (.A(_12080_),
    .B(_13102_),
    .C(_13106_),
    .Y(_13107_));
 AO21x1_ASAP7_75t_R _34433_ (.A1(_14604_),
    .A2(_12117_),
    .B(_13107_),
    .Y(_04138_));
 OA21x2_ASAP7_75t_R _34434_ (.A1(_12822_),
    .A2(_12829_),
    .B(_12739_),
    .Y(_13108_));
 OA21x2_ASAP7_75t_R _34435_ (.A1(_12944_),
    .A2(_13108_),
    .B(_12849_),
    .Y(_13109_));
 AO32x1_ASAP7_75t_R _34436_ (.A1(_12781_),
    .A2(_12827_),
    .A3(_12965_),
    .B1(_12849_),
    .B2(_12787_),
    .Y(_13110_));
 OA21x2_ASAP7_75t_R _34437_ (.A1(_12848_),
    .A2(_12860_),
    .B(_12868_),
    .Y(_13111_));
 AO21x1_ASAP7_75t_R _34438_ (.A1(_12777_),
    .A2(_13110_),
    .B(_13111_),
    .Y(_13112_));
 OR3x1_ASAP7_75t_R _34439_ (.A(_12023_),
    .B(_13109_),
    .C(_13112_),
    .Y(_13113_));
 OA21x2_ASAP7_75t_R _34440_ (.A1(_13391_),
    .A2(_12800_),
    .B(_13113_),
    .Y(_04139_));
 NAND2x1_ASAP7_75t_R _34441_ (.A(_05487_),
    .B(_12387_),
    .Y(_13114_));
 OA211x2_ASAP7_75t_R _34442_ (.A1(_12773_),
    .A2(_12676_),
    .B(_13114_),
    .C(_07311_),
    .Y(_13115_));
 AOI21x1_ASAP7_75t_R _34443_ (.A1(_05484_),
    .A2(_12193_),
    .B(_13115_),
    .Y(_13116_));
 NOR2x1_ASAP7_75t_R _34444_ (.A(_12944_),
    .B(_12987_),
    .Y(_13117_));
 AO21x1_ASAP7_75t_R _34445_ (.A1(_12691_),
    .A2(_12660_),
    .B(_12818_),
    .Y(_13118_));
 AND3x1_ASAP7_75t_R _34446_ (.A(_12690_),
    .B(_12818_),
    .C(_13116_),
    .Y(_13119_));
 AO21x1_ASAP7_75t_R _34447_ (.A1(_12653_),
    .A2(_12714_),
    .B(_13119_),
    .Y(_13120_));
 NAND2x1_ASAP7_75t_R _34448_ (.A(_12660_),
    .B(_13120_),
    .Y(_13121_));
 AO21x1_ASAP7_75t_R _34449_ (.A1(_13118_),
    .A2(_13121_),
    .B(_13022_),
    .Y(_13122_));
 OA211x2_ASAP7_75t_R _34450_ (.A1(_12754_),
    .A2(_12841_),
    .B(_13122_),
    .C(_12783_),
    .Y(_13123_));
 OAI21x1_ASAP7_75t_R _34451_ (.A1(_13056_),
    .A2(_13123_),
    .B(_13049_),
    .Y(_13124_));
 OA211x2_ASAP7_75t_R _34452_ (.A1(_13116_),
    .A2(_13117_),
    .B(_13124_),
    .C(_12080_),
    .Y(_13125_));
 AOI21x1_ASAP7_75t_R _34453_ (.A1(_13575_),
    .A2(_12638_),
    .B(_13125_),
    .Y(_04140_));
 NAND2x1_ASAP7_75t_R _34454_ (.A(_11959_),
    .B(_12391_),
    .Y(_13126_));
 OA211x2_ASAP7_75t_R _34455_ (.A1(_11959_),
    .A2(_12670_),
    .B(_13126_),
    .C(_07313_),
    .Y(_13127_));
 AOI21x1_ASAP7_75t_R _34456_ (.A1(_12915_),
    .A2(_12196_),
    .B(_13127_),
    .Y(_13128_));
 AO21x1_ASAP7_75t_R _34457_ (.A1(_12818_),
    .A2(_13128_),
    .B(_12821_),
    .Y(_13129_));
 OR3x1_ASAP7_75t_R _34458_ (.A(_12806_),
    .B(_12653_),
    .C(_12822_),
    .Y(_13130_));
 AO21x1_ASAP7_75t_R _34459_ (.A1(_12827_),
    .A2(_13129_),
    .B(_13130_),
    .Y(_13131_));
 OA211x2_ASAP7_75t_R _34460_ (.A1(_13117_),
    .A2(_13128_),
    .B(_13131_),
    .C(_12080_),
    .Y(_13132_));
 AOI21x1_ASAP7_75t_R _34461_ (.A1(_13576_),
    .A2(_12638_),
    .B(_13132_),
    .Y(_04141_));
 AO221x1_ASAP7_75t_R _34462_ (.A1(_12829_),
    .A2(_12834_),
    .B1(_12879_),
    .B2(_12746_),
    .C(_12987_),
    .Y(_13133_));
 AO221x1_ASAP7_75t_R _34463_ (.A1(_12868_),
    .A2(_12860_),
    .B1(_13133_),
    .B2(_12701_),
    .C(_12637_),
    .Y(_13134_));
 OA21x2_ASAP7_75t_R _34464_ (.A1(_13392_),
    .A2(_12800_),
    .B(_13134_),
    .Y(_04142_));
 INVx1_ASAP7_75t_R _34465_ (.A(_12869_),
    .Y(_13135_));
 AO21x1_ASAP7_75t_R _34466_ (.A1(_12816_),
    .A2(_12645_),
    .B(_12787_),
    .Y(_13136_));
 AND4x1_ASAP7_75t_R _34467_ (.A(_12782_),
    .B(_12841_),
    .C(_12781_),
    .D(_12775_),
    .Y(_13137_));
 AO221x1_ASAP7_75t_R _34468_ (.A1(_13135_),
    .A2(_13136_),
    .B1(_13137_),
    .B2(_12965_),
    .C(_12877_),
    .Y(_13138_));
 OR2x2_ASAP7_75t_R _34469_ (.A(_12785_),
    .B(_12891_),
    .Y(_13139_));
 AO21x1_ASAP7_75t_R _34470_ (.A1(_12645_),
    .A2(_12908_),
    .B(_12869_),
    .Y(_13140_));
 OA211x2_ASAP7_75t_R _34471_ (.A1(_12822_),
    .A2(_13139_),
    .B(_13140_),
    .C(_12739_),
    .Y(_13141_));
 INVx1_ASAP7_75t_R _34472_ (.A(_13141_),
    .Y(_13142_));
 OA211x2_ASAP7_75t_R _34473_ (.A1(_12739_),
    .A2(_13138_),
    .B(_13142_),
    .C(_12080_),
    .Y(_13143_));
 AOI21x1_ASAP7_75t_R _34474_ (.A1(_13569_),
    .A2(_12638_),
    .B(_13143_),
    .Y(_04143_));
 BUFx6f_ASAP7_75t_R _34475_ (.A(_12080_),
    .Y(_13144_));
 OA21x2_ASAP7_75t_R _34476_ (.A1(_12653_),
    .A2(_12883_),
    .B(_12976_),
    .Y(_13145_));
 OR3x1_ASAP7_75t_R _34477_ (.A(_12848_),
    .B(_13053_),
    .C(_13145_),
    .Y(_13146_));
 OR2x2_ASAP7_75t_R _34478_ (.A(_12747_),
    .B(_12883_),
    .Y(_13147_));
 AO21x1_ASAP7_75t_R _34479_ (.A1(_12806_),
    .A2(_13147_),
    .B(_12822_),
    .Y(_13148_));
 OA22x2_ASAP7_75t_R _34480_ (.A1(_12739_),
    .A2(_12991_),
    .B1(_12823_),
    .B2(_12883_),
    .Y(_13149_));
 AO221x1_ASAP7_75t_R _34481_ (.A1(_12834_),
    .A2(_13146_),
    .B1(_13148_),
    .B2(_13149_),
    .C(_12637_),
    .Y(_13150_));
 OA21x2_ASAP7_75t_R _34482_ (.A1(_13399_),
    .A2(_13144_),
    .B(_13150_),
    .Y(_04144_));
 BUFx3_ASAP7_75t_R _34483_ (.A(_12637_),
    .Y(_13151_));
 NOR2x1_ASAP7_75t_R _34484_ (.A(_12728_),
    .B(_12687_),
    .Y(_13152_));
 AO222x2_ASAP7_75t_R _34485_ (.A1(_12777_),
    .A2(_13152_),
    .B1(_12868_),
    .B2(_13053_),
    .C1(_13133_),
    .C2(_12839_),
    .Y(_13153_));
 AO21x1_ASAP7_75t_R _34486_ (.A1(_12790_),
    .A2(_12791_),
    .B(_13375_),
    .Y(_13154_));
 OA21x2_ASAP7_75t_R _34487_ (.A1(_13151_),
    .A2(_13153_),
    .B(_13154_),
    .Y(_04145_));
 AO21x1_ASAP7_75t_R _34488_ (.A1(_12728_),
    .A2(_12807_),
    .B(_13022_),
    .Y(_13155_));
 AND4x1_ASAP7_75t_R _34489_ (.A(_12691_),
    .B(_12769_),
    .C(_13152_),
    .D(_12833_),
    .Y(_13156_));
 AO21x1_ASAP7_75t_R _34490_ (.A1(_12875_),
    .A2(_13155_),
    .B(_13156_),
    .Y(_13157_));
 AO221x1_ASAP7_75t_R _34491_ (.A1(_12849_),
    .A2(_13029_),
    .B1(_12745_),
    .B2(_12875_),
    .C(_12775_),
    .Y(_13158_));
 OA21x2_ASAP7_75t_R _34492_ (.A1(_12646_),
    .A2(_13157_),
    .B(_13158_),
    .Y(_13159_));
 OR3x1_ASAP7_75t_R _34493_ (.A(_12778_),
    .B(_12775_),
    .C(_12891_),
    .Y(_13160_));
 AO22x1_ASAP7_75t_R _34494_ (.A1(_12744_),
    .A2(_12866_),
    .B1(_13056_),
    .B2(_12782_),
    .Y(_13161_));
 AO221x1_ASAP7_75t_R _34495_ (.A1(_12875_),
    .A2(_13160_),
    .B1(_13161_),
    .B2(_12646_),
    .C(_12806_),
    .Y(_13162_));
 OA211x2_ASAP7_75t_R _34496_ (.A1(_12739_),
    .A2(_13159_),
    .B(_13162_),
    .C(_12810_),
    .Y(_13163_));
 AO21x1_ASAP7_75t_R _34497_ (.A1(_08329_),
    .A2(_12117_),
    .B(_13163_),
    .Y(_04146_));
 AND3x1_ASAP7_75t_R _34498_ (.A(_12736_),
    .B(_12816_),
    .C(_12747_),
    .Y(_13164_));
 AO21x1_ASAP7_75t_R _34499_ (.A1(_12806_),
    .A2(_13029_),
    .B(_13164_),
    .Y(_13165_));
 AO21x1_ASAP7_75t_R _34500_ (.A1(_12736_),
    .A2(_13139_),
    .B(_12822_),
    .Y(_13166_));
 OR2x2_ASAP7_75t_R _34501_ (.A(_12736_),
    .B(_13155_),
    .Y(_13167_));
 AO21x1_ASAP7_75t_R _34502_ (.A1(_13166_),
    .A2(_13167_),
    .B(_12944_),
    .Y(_13168_));
 AO32x1_ASAP7_75t_R _34503_ (.A1(_12701_),
    .A2(_12646_),
    .A3(_13165_),
    .B1(_13168_),
    .B2(_12754_),
    .Y(_13169_));
 AO21x1_ASAP7_75t_R _34504_ (.A1(_12790_),
    .A2(_12791_),
    .B(_09773_),
    .Y(_13170_));
 OA21x2_ASAP7_75t_R _34505_ (.A1(_13151_),
    .A2(_13169_),
    .B(_13170_),
    .Y(_04147_));
 AO32x1_ASAP7_75t_R _34506_ (.A1(_12816_),
    .A2(_12747_),
    .A3(_12869_),
    .B1(_12891_),
    .B2(_12760_),
    .Y(_13171_));
 AO32x1_ASAP7_75t_R _34507_ (.A1(_12816_),
    .A2(_12839_),
    .A3(_12877_),
    .B1(_13029_),
    .B2(_12869_),
    .Y(_13172_));
 AO22x1_ASAP7_75t_R _34508_ (.A1(_12868_),
    .A2(_13171_),
    .B1(_13172_),
    .B2(_12879_),
    .Y(_13173_));
 AND3x1_ASAP7_75t_R _34509_ (.A(_12735_),
    .B(_12778_),
    .C(_12747_),
    .Y(_13174_));
 AO21x1_ASAP7_75t_R _34510_ (.A1(_12774_),
    .A2(_12745_),
    .B(_13174_),
    .Y(_13175_));
 OA211x2_ASAP7_75t_R _34511_ (.A1(_12822_),
    .A2(_13175_),
    .B(_12812_),
    .C(_12760_),
    .Y(_13176_));
 OR3x1_ASAP7_75t_R _34512_ (.A(_12023_),
    .B(_13173_),
    .C(_13176_),
    .Y(_13177_));
 OA21x2_ASAP7_75t_R _34513_ (.A1(_14153_),
    .A2(_13144_),
    .B(_13177_),
    .Y(_04148_));
 NAND2x1_ASAP7_75t_R _34514_ (.A(_01545_),
    .B(_12154_),
    .Y(_13178_));
 OA21x2_ASAP7_75t_R _34515_ (.A1(_13151_),
    .A2(_12739_),
    .B(_13178_),
    .Y(_04149_));
 NAND2x1_ASAP7_75t_R _34516_ (.A(_00038_),
    .B(_12154_),
    .Y(_13179_));
 OA21x2_ASAP7_75t_R _34517_ (.A1(_13151_),
    .A2(_12818_),
    .B(_13179_),
    .Y(_04150_));
 NAND2x1_ASAP7_75t_R _34518_ (.A(_00041_),
    .B(_12154_),
    .Y(_13180_));
 OA21x2_ASAP7_75t_R _34519_ (.A1(_13151_),
    .A2(_12660_),
    .B(_13180_),
    .Y(_04151_));
 NAND2x1_ASAP7_75t_R _34520_ (.A(_00043_),
    .B(_12154_),
    .Y(_13181_));
 OA21x2_ASAP7_75t_R _34521_ (.A1(_13151_),
    .A2(_12837_),
    .B(_13181_),
    .Y(_04152_));
 NAND2x1_ASAP7_75t_R _34522_ (.A(_00045_),
    .B(_12154_),
    .Y(_13182_));
 OA21x2_ASAP7_75t_R _34523_ (.A1(_13151_),
    .A2(_12787_),
    .B(_13182_),
    .Y(_04153_));
 NAND2x1_ASAP7_75t_R _34524_ (.A(_00047_),
    .B(_12154_),
    .Y(_13183_));
 OA21x2_ASAP7_75t_R _34525_ (.A1(_13151_),
    .A2(_12747_),
    .B(_13183_),
    .Y(_04154_));
 NAND2x1_ASAP7_75t_R _34526_ (.A(_00049_),
    .B(_12154_),
    .Y(_13184_));
 OA21x2_ASAP7_75t_R _34527_ (.A1(_13151_),
    .A2(_12816_),
    .B(_13184_),
    .Y(_04155_));
 NAND2x1_ASAP7_75t_R _34528_ (.A(_00014_),
    .B(_12154_),
    .Y(_13185_));
 OA21x2_ASAP7_75t_R _34529_ (.A1(_13151_),
    .A2(_12822_),
    .B(_13185_),
    .Y(_04156_));
 BUFx4f_ASAP7_75t_R _34530_ (.A(_12637_),
    .Y(_13186_));
 NAND2x1_ASAP7_75t_R _34531_ (.A(_00016_),
    .B(_12154_),
    .Y(_13187_));
 OA21x2_ASAP7_75t_R _34532_ (.A1(_13186_),
    .A2(_12849_),
    .B(_13187_),
    .Y(_04157_));
 NAND2x1_ASAP7_75t_R _34533_ (.A(_00019_),
    .B(_12018_),
    .Y(_13188_));
 OA21x2_ASAP7_75t_R _34534_ (.A1(_13186_),
    .A2(_12701_),
    .B(_13188_),
    .Y(_04158_));
 NAND2x1_ASAP7_75t_R _34535_ (.A(_00022_),
    .B(_12018_),
    .Y(_13189_));
 OA21x2_ASAP7_75t_R _34536_ (.A1(_13186_),
    .A2(_12869_),
    .B(_13189_),
    .Y(_04159_));
 NAND2x1_ASAP7_75t_R _34537_ (.A(_00025_),
    .B(_12018_),
    .Y(_13190_));
 OA21x2_ASAP7_75t_R _34538_ (.A1(_13186_),
    .A2(_12883_),
    .B(_13190_),
    .Y(_04160_));
 NAND2x1_ASAP7_75t_R _34539_ (.A(_00027_),
    .B(_12018_),
    .Y(_13191_));
 OA21x2_ASAP7_75t_R _34540_ (.A1(_13186_),
    .A2(_12839_),
    .B(_13191_),
    .Y(_04161_));
 NAND2x1_ASAP7_75t_R _34541_ (.A(_00029_),
    .B(_12018_),
    .Y(_13192_));
 OA21x2_ASAP7_75t_R _34542_ (.A1(_13186_),
    .A2(_12875_),
    .B(_13192_),
    .Y(_04162_));
 NAND2x1_ASAP7_75t_R _34543_ (.A(_00032_),
    .B(_12018_),
    .Y(_13193_));
 OA21x2_ASAP7_75t_R _34544_ (.A1(_13186_),
    .A2(_12754_),
    .B(_13193_),
    .Y(_04163_));
 NAND2x1_ASAP7_75t_R _34545_ (.A(_00035_),
    .B(_12018_),
    .Y(_13194_));
 OA21x2_ASAP7_75t_R _34546_ (.A1(_13186_),
    .A2(_12760_),
    .B(_13194_),
    .Y(_04164_));
 BUFx4f_ASAP7_75t_R _34547_ (.A(_12810_),
    .Y(_13195_));
 NAND2x1_ASAP7_75t_R _34548_ (.A(_07255_),
    .B(_13195_),
    .Y(_13196_));
 OA21x2_ASAP7_75t_R _34549_ (.A1(_15464_),
    .A2(_13144_),
    .B(_13196_),
    .Y(_04165_));
 NAND2x1_ASAP7_75t_R _34550_ (.A(_01709_),
    .B(_13195_),
    .Y(_13197_));
 OA21x2_ASAP7_75t_R _34551_ (.A1(_14806_),
    .A2(_13144_),
    .B(_13197_),
    .Y(_04166_));
 BUFx6f_ASAP7_75t_R _34552_ (.A(_12810_),
    .Y(_13198_));
 NAND2x1_ASAP7_75t_R _34553_ (.A(_01708_),
    .B(_13198_),
    .Y(_13199_));
 OA21x2_ASAP7_75t_R _34554_ (.A1(_14014_),
    .A2(_13144_),
    .B(_13199_),
    .Y(_04167_));
 NAND2x1_ASAP7_75t_R _34555_ (.A(_01707_),
    .B(_13198_),
    .Y(_13200_));
 OA21x2_ASAP7_75t_R _34556_ (.A1(_15724_),
    .A2(_13144_),
    .B(_13200_),
    .Y(_04168_));
 NAND2x1_ASAP7_75t_R _34557_ (.A(_07276_),
    .B(_13198_),
    .Y(_13201_));
 OA21x2_ASAP7_75t_R _34558_ (.A1(_15864_),
    .A2(_13144_),
    .B(_13201_),
    .Y(_04169_));
 NAND2x1_ASAP7_75t_R _34559_ (.A(_01705_),
    .B(_13198_),
    .Y(_13202_));
 OA21x2_ASAP7_75t_R _34560_ (.A1(_16003_),
    .A2(_13144_),
    .B(_13202_),
    .Y(_04170_));
 NAND2x1_ASAP7_75t_R _34561_ (.A(_07286_),
    .B(_13198_),
    .Y(_13203_));
 OA21x2_ASAP7_75t_R _34562_ (.A1(_16141_),
    .A2(_13144_),
    .B(_13203_),
    .Y(_04171_));
 AO21x1_ASAP7_75t_R _34563_ (.A1(_12790_),
    .A2(_12791_),
    .B(_16256_),
    .Y(_13204_));
 OA21x2_ASAP7_75t_R _34564_ (.A1(_12064_),
    .A2(_13186_),
    .B(_13204_),
    .Y(_04172_));
 NAND2x1_ASAP7_75t_R _34565_ (.A(_01702_),
    .B(_13198_),
    .Y(_13205_));
 OA21x2_ASAP7_75t_R _34566_ (.A1(_16401_),
    .A2(_13144_),
    .B(_13205_),
    .Y(_04173_));
 BUFx3_ASAP7_75t_R _34567_ (.A(_12080_),
    .Y(_13206_));
 NAND2x1_ASAP7_75t_R _34568_ (.A(_07302_),
    .B(_13198_),
    .Y(_13207_));
 OA21x2_ASAP7_75t_R _34569_ (.A1(_16513_),
    .A2(_13206_),
    .B(_13207_),
    .Y(_04174_));
 OR3x1_ASAP7_75t_R _34570_ (.A(_12915_),
    .B(_11072_),
    .C(_11966_),
    .Y(_13208_));
 OA21x2_ASAP7_75t_R _34571_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(_13206_),
    .B(_13208_),
    .Y(_04175_));
 NAND2x1_ASAP7_75t_R _34572_ (.A(_01700_),
    .B(_13198_),
    .Y(_13209_));
 OA21x2_ASAP7_75t_R _34573_ (.A1(_16642_),
    .A2(_13206_),
    .B(_13209_),
    .Y(_04176_));
 NAND2x1_ASAP7_75t_R _34574_ (.A(_01699_),
    .B(_13198_),
    .Y(_13210_));
 OA21x2_ASAP7_75t_R _34575_ (.A1(_16752_),
    .A2(_13206_),
    .B(_13210_),
    .Y(_04177_));
 NAND2x1_ASAP7_75t_R _34576_ (.A(_01698_),
    .B(_13198_),
    .Y(_13211_));
 OA21x2_ASAP7_75t_R _34577_ (.A1(_16883_),
    .A2(_13206_),
    .B(_13211_),
    .Y(_04178_));
 BUFx6f_ASAP7_75t_R _34578_ (.A(_12810_),
    .Y(_13212_));
 NAND2x1_ASAP7_75t_R _34579_ (.A(_07333_),
    .B(_13212_),
    .Y(_13213_));
 OA21x2_ASAP7_75t_R _34580_ (.A1(_16993_),
    .A2(_13206_),
    .B(_13213_),
    .Y(_04179_));
 NAND2x1_ASAP7_75t_R _34581_ (.A(_01696_),
    .B(_13212_),
    .Y(_13214_));
 OA21x2_ASAP7_75t_R _34582_ (.A1(_17122_),
    .A2(_13206_),
    .B(_13214_),
    .Y(_04180_));
 AO21x1_ASAP7_75t_R _34583_ (.A1(_12790_),
    .A2(_12791_),
    .B(_17231_),
    .Y(_13215_));
 OA21x2_ASAP7_75t_R _34584_ (.A1(_12115_),
    .A2(_13186_),
    .B(_13215_),
    .Y(_04181_));
 NAND2x1_ASAP7_75t_R _34585_ (.A(_01694_),
    .B(_13212_),
    .Y(_13216_));
 OA21x2_ASAP7_75t_R _34586_ (.A1(_04280_),
    .A2(_13206_),
    .B(_13216_),
    .Y(_04182_));
 NAND2x1_ASAP7_75t_R _34587_ (.A(_01693_),
    .B(_13212_),
    .Y(_13217_));
 OA21x2_ASAP7_75t_R _34588_ (.A1(_04389_),
    .A2(_13206_),
    .B(_13217_),
    .Y(_04183_));
 AO21x1_ASAP7_75t_R _34589_ (.A1(_12790_),
    .A2(_12791_),
    .B(_04519_),
    .Y(_13218_));
 OA21x2_ASAP7_75t_R _34590_ (.A1(_12127_),
    .A2(_12793_),
    .B(_13218_),
    .Y(_04184_));
 NAND2x1_ASAP7_75t_R _34591_ (.A(_01691_),
    .B(_13212_),
    .Y(_13219_));
 OA21x2_ASAP7_75t_R _34592_ (.A1(_04629_),
    .A2(_13206_),
    .B(_13219_),
    .Y(_04185_));
 AO21x1_ASAP7_75t_R _34593_ (.A1(_06859_),
    .A2(_12791_),
    .B(\cs_registers_i.pc_id_i[2] ),
    .Y(_13220_));
 OA21x2_ASAP7_75t_R _34594_ (.A1(\cs_registers_i.pc_if_i[2] ),
    .A2(_12793_),
    .B(_13220_),
    .Y(_04186_));
 AO21x1_ASAP7_75t_R _34595_ (.A1(_06859_),
    .A2(_11955_),
    .B(_04743_),
    .Y(_13221_));
 OA21x2_ASAP7_75t_R _34596_ (.A1(_12137_),
    .A2(_12793_),
    .B(_13221_),
    .Y(_04187_));
 NAND2x1_ASAP7_75t_R _34597_ (.A(_01688_),
    .B(_13212_),
    .Y(_13222_));
 OA21x2_ASAP7_75t_R _34598_ (.A1(_04864_),
    .A2(_13195_),
    .B(_13222_),
    .Y(_04188_));
 OR3x1_ASAP7_75t_R _34599_ (.A(_12024_),
    .B(_11072_),
    .C(_11966_),
    .Y(_13223_));
 OA21x2_ASAP7_75t_R _34600_ (.A1(_14979_),
    .A2(_13195_),
    .B(_13223_),
    .Y(_04189_));
 NAND2x1_ASAP7_75t_R _34601_ (.A(_07378_),
    .B(_13212_),
    .Y(_13224_));
 OA21x2_ASAP7_75t_R _34602_ (.A1(_15054_),
    .A2(_13195_),
    .B(_13224_),
    .Y(_04190_));
 NAND2x1_ASAP7_75t_R _34603_ (.A(_07383_),
    .B(_13212_),
    .Y(_13225_));
 OA21x2_ASAP7_75t_R _34604_ (.A1(_15116_),
    .A2(_13195_),
    .B(_13225_),
    .Y(_04191_));
 NAND2x1_ASAP7_75t_R _34605_ (.A(_01685_),
    .B(_13212_),
    .Y(_13226_));
 OA21x2_ASAP7_75t_R _34606_ (.A1(_15180_),
    .A2(_13195_),
    .B(_13226_),
    .Y(_04192_));
 NAND2x1_ASAP7_75t_R _34607_ (.A(_07392_),
    .B(_13212_),
    .Y(_13227_));
 OA21x2_ASAP7_75t_R _34608_ (.A1(_15235_),
    .A2(_13195_),
    .B(_13227_),
    .Y(_04193_));
 NAND2x1_ASAP7_75t_R _34609_ (.A(_07397_),
    .B(_12075_),
    .Y(_13228_));
 OA21x2_ASAP7_75t_R _34610_ (.A1(_15333_),
    .A2(_13195_),
    .B(_13228_),
    .Y(_04194_));
 NAND2x1_ASAP7_75t_R _34611_ (.A(_01682_),
    .B(_12075_),
    .Y(_13229_));
 OA21x2_ASAP7_75t_R _34612_ (.A1(_15391_),
    .A2(_13195_),
    .B(_13229_),
    .Y(_04195_));
 INVx1_ASAP7_75t_R _34613_ (.A(_19026_),
    .Y(_17580_));
 INVx1_ASAP7_75t_R _34614_ (.A(_19008_),
    .Y(_17581_));
 INVx1_ASAP7_75t_R _34615_ (.A(_18466_),
    .Y(_18014_));
 INVx1_ASAP7_75t_R _34616_ (.A(_18517_),
    .Y(_18112_));
 INVx1_ASAP7_75t_R _34617_ (.A(_18498_),
    .Y(_18113_));
 INVx1_ASAP7_75t_R _34618_ (.A(_02242_),
    .Y(_18121_));
 INVx1_ASAP7_75t_R _34619_ (.A(_00251_),
    .Y(_18087_));
 INVx1_ASAP7_75t_R _34620_ (.A(_00147_),
    .Y(_17359_));
 INVx1_ASAP7_75t_R _34621_ (.A(_19047_),
    .Y(_17672_));
 INVx1_ASAP7_75t_R _34622_ (.A(_18350_),
    .Y(_17789_));
 INVx1_ASAP7_75t_R _34623_ (.A(_18326_),
    .Y(_17790_));
 INVx1_ASAP7_75t_R _34624_ (.A(_18321_),
    .Y(_17725_));
 INVx1_ASAP7_75t_R _34625_ (.A(_19065_),
    .Y(_17726_));
 INVx1_ASAP7_75t_R _34626_ (.A(_18351_),
    .Y(_17787_));
 INVx1_ASAP7_75t_R _34627_ (.A(_18325_),
    .Y(_17788_));
 INVx1_ASAP7_75t_R _34628_ (.A(_18324_),
    .Y(_17721_));
 INVx1_ASAP7_75t_R _34629_ (.A(_19064_),
    .Y(_17722_));
 INVx1_ASAP7_75t_R _34630_ (.A(_19063_),
    .Y(_17671_));
 INVx1_ASAP7_75t_R _34631_ (.A(_19061_),
    .Y(_17657_));
 INVx1_ASAP7_75t_R _34632_ (.A(_19042_),
    .Y(_17611_));
 INVx1_ASAP7_75t_R _34633_ (.A(_19043_),
    .Y(_17615_));
 INVx1_ASAP7_75t_R _34634_ (.A(_19022_),
    .Y(_17616_));
 INVx1_ASAP7_75t_R _34635_ (.A(_18374_),
    .Y(_17835_));
 INVx1_ASAP7_75t_R _34636_ (.A(_18349_),
    .Y(_17836_));
 INVx1_ASAP7_75t_R _34637_ (.A(_18346_),
    .Y(_17778_));
 INVx1_ASAP7_75t_R _34638_ (.A(_18320_),
    .Y(_17779_));
 INVx1_ASAP7_75t_R _34639_ (.A(_18355_),
    .Y(_17795_));
 INVx1_ASAP7_75t_R _34640_ (.A(_02339_),
    .Y(_17551_));
 INVx1_ASAP7_75t_R _34641_ (.A(_19083_),
    .Y(_17776_));
 INVx1_ASAP7_75t_R _34642_ (.A(_19080_),
    .Y(_17707_));
 INVx1_ASAP7_75t_R _34643_ (.A(_19058_),
    .Y(_17655_));
 INVx1_ASAP7_75t_R _34644_ (.A(_19041_),
    .Y(_17656_));
 INVx1_ASAP7_75t_R _34645_ (.A(_19082_),
    .Y(_17719_));
 INVx1_ASAP7_75t_R _34646_ (.A(_19062_),
    .Y(_17720_));
 INVx1_ASAP7_75t_R _34647_ (.A(_19059_),
    .Y(_17665_));
 INVx1_ASAP7_75t_R _34648_ (.A(_19044_),
    .Y(_17666_));
 INVx1_ASAP7_75t_R _34649_ (.A(_18370_),
    .Y(_17825_));
 INVx1_ASAP7_75t_R _34650_ (.A(_18345_),
    .Y(_17826_));
 INVx1_ASAP7_75t_R _34651_ (.A(_18338_),
    .Y(_17763_));
 INVx1_ASAP7_75t_R _34652_ (.A(_19077_),
    .Y(_17764_));
 INVx1_ASAP7_75t_R _34653_ (.A(_18362_),
    .Y(_17811_));
 INVx1_ASAP7_75t_R _34654_ (.A(_18337_),
    .Y(_17812_));
 INVx1_ASAP7_75t_R _34655_ (.A(_18333_),
    .Y(_17752_));
 INVx1_ASAP7_75t_R _34656_ (.A(_19073_),
    .Y(_17753_));
 INVx1_ASAP7_75t_R _34657_ (.A(_19072_),
    .Y(_17693_));
 INVx1_ASAP7_75t_R _34658_ (.A(_18367_),
    .Y(_17809_));
 INVx1_ASAP7_75t_R _34659_ (.A(_18336_),
    .Y(_17810_));
 INVx1_ASAP7_75t_R _34660_ (.A(_18344_),
    .Y(_17824_));
 INVx1_ASAP7_75t_R _34661_ (.A(_18342_),
    .Y(_17760_));
 INVx1_ASAP7_75t_R _34662_ (.A(_19076_),
    .Y(_17761_));
 INVx1_ASAP7_75t_R _34663_ (.A(_19075_),
    .Y(_17704_));
 INVx1_ASAP7_75t_R _34664_ (.A(_19057_),
    .Y(_17705_));
 INVx1_ASAP7_75t_R _34665_ (.A(_18335_),
    .Y(_17757_));
 INVx1_ASAP7_75t_R _34666_ (.A(_19074_),
    .Y(_17758_));
 INVx1_ASAP7_75t_R _34667_ (.A(_18597_),
    .Y(_18273_));
 INVx1_ASAP7_75t_R _34668_ (.A(_18588_),
    .Y(_18274_));
 INVx1_ASAP7_75t_R _34669_ (.A(_18584_),
    .Y(_18265_));
 INVx1_ASAP7_75t_R _34670_ (.A(_02244_),
    .Y(_18184_));
 INVx1_ASAP7_75t_R _34671_ (.A(_18343_),
    .Y(_17774_));
 INVx1_ASAP7_75t_R _34672_ (.A(_19081_),
    .Y(_17775_));
 INVx1_ASAP7_75t_R _34673_ (.A(_02243_),
    .Y(_18154_));
 INVx1_ASAP7_75t_R _34674_ (.A(_00254_),
    .Y(_18123_));
 INVx1_ASAP7_75t_R _34675_ (.A(_18445_),
    .Y(_18015_));
 INVx1_ASAP7_75t_R _34676_ (.A(_18927_),
    .Y(_17395_));
 INVx1_ASAP7_75t_R _34677_ (.A(_18330_),
    .Y(_17796_));
 INVx1_ASAP7_75t_R _34678_ (.A(_18334_),
    .Y(_17807_));
 INVx1_ASAP7_75t_R _34679_ (.A(_19034_),
    .Y(_17604_));
 INVx1_ASAP7_75t_R _34680_ (.A(_18969_),
    .Y(_17466_));
 INVx1_ASAP7_75t_R _34681_ (.A(_18955_),
    .Y(_17437_));
 INVx1_ASAP7_75t_R _34682_ (.A(_18939_),
    .Y(_17438_));
 INVx1_ASAP7_75t_R _34683_ (.A(_18966_),
    .Y(_17460_));
 INVx1_ASAP7_75t_R _34684_ (.A(_18954_),
    .Y(_17461_));
 INVx1_ASAP7_75t_R _34685_ (.A(_02338_),
    .Y(_17528_));
 INVx1_ASAP7_75t_R _34686_ (.A(_00190_),
    .Y(_17499_));
 INVx1_ASAP7_75t_R _34687_ (.A(_18463_),
    .Y(_18008_));
 INVx1_ASAP7_75t_R _34688_ (.A(_18441_),
    .Y(_18009_));
 INVx1_ASAP7_75t_R _34689_ (.A(_18437_),
    .Y(_17958_));
 INVx1_ASAP7_75t_R _34690_ (.A(_18417_),
    .Y(_17959_));
 INVx1_ASAP7_75t_R _34691_ (.A(_18416_),
    .Y(_17957_));
 INVx1_ASAP7_75t_R _34692_ (.A(_18389_),
    .Y(_17916_));
 INVx1_ASAP7_75t_R _34693_ (.A(_18415_),
    .Y(_17915_));
 INVx1_ASAP7_75t_R _34694_ (.A(_18917_),
    .Y(_17396_));
 INVx1_ASAP7_75t_R _34695_ (.A(_00220_),
    .Y(_17661_));
 INVx1_ASAP7_75t_R _34696_ (.A(_02346_),
    .Y(_17658_));
 INVx1_ASAP7_75t_R _34697_ (.A(_00212_),
    .Y(_19021_));
 INVx1_ASAP7_75t_R _34698_ (.A(_18390_),
    .Y(_17854_));
 INVx1_ASAP7_75t_R _34699_ (.A(_18360_),
    .Y(_17855_));
 INVx1_ASAP7_75t_R _34700_ (.A(_18520_),
    .Y(_18148_));
 INVx1_ASAP7_75t_R _34701_ (.A(_19050_),
    .Y(_17636_));
 INVx1_ASAP7_75t_R _34702_ (.A(_19030_),
    .Y(_17637_));
 INVx1_ASAP7_75t_R _34703_ (.A(_18519_),
    .Y(_18110_));
 INVx1_ASAP7_75t_R _34704_ (.A(_18496_),
    .Y(_18111_));
 INVx1_ASAP7_75t_R _34705_ (.A(_02344_),
    .Y(_17630_));
 INVx1_ASAP7_75t_R _34706_ (.A(_00208_),
    .Y(_17590_));
 INVx1_ASAP7_75t_R _34707_ (.A(_18388_),
    .Y(_17861_));
 INVx1_ASAP7_75t_R _34708_ (.A(_18363_),
    .Y(_17862_));
 INVx1_ASAP7_75t_R _34709_ (.A(_18409_),
    .Y(_17903_));
 INVx1_ASAP7_75t_R _34710_ (.A(_18385_),
    .Y(_17904_));
 INVx1_ASAP7_75t_R _34711_ (.A(_18949_),
    .Y(_17428_));
 INVx1_ASAP7_75t_R _34712_ (.A(_18933_),
    .Y(_17429_));
 INVx1_ASAP7_75t_R _34713_ (.A(_19068_),
    .Y(_17741_));
 INVx1_ASAP7_75t_R _34714_ (.A(_18327_),
    .Y(_17740_));
 INVx1_ASAP7_75t_R _34715_ (.A(_18493_),
    .Y(_18064_));
 INVx1_ASAP7_75t_R _34716_ (.A(_19027_),
    .Y(_17576_));
 INVx1_ASAP7_75t_R _34717_ (.A(_18468_),
    .Y(_18065_));
 INVx1_ASAP7_75t_R _34718_ (.A(_18495_),
    .Y(_18071_));
 INVx1_ASAP7_75t_R _34719_ (.A(_19006_),
    .Y(_17536_));
 INVx1_ASAP7_75t_R _34720_ (.A(_19029_),
    .Y(_17586_));
 INVx1_ASAP7_75t_R _34721_ (.A(_19010_),
    .Y(_17587_));
 INVx1_ASAP7_75t_R _34722_ (.A(_19009_),
    .Y(_17540_));
 INVx1_ASAP7_75t_R _34723_ (.A(_18995_),
    .Y(_17541_));
 INVx1_ASAP7_75t_R _34724_ (.A(_18471_),
    .Y(_18072_));
 INVx1_ASAP7_75t_R _34725_ (.A(_19048_),
    .Y(_17628_));
 INVx1_ASAP7_75t_R _34726_ (.A(_19028_),
    .Y(_17629_));
 INVx1_ASAP7_75t_R _34727_ (.A(_19045_),
    .Y(_17622_));
 INVx1_ASAP7_75t_R _34728_ (.A(_19025_),
    .Y(_17623_));
 INVx1_ASAP7_75t_R _34729_ (.A(_18366_),
    .Y(_17869_));
 INVx1_ASAP7_75t_R _34730_ (.A(_18391_),
    .Y(_17868_));
 INVx1_ASAP7_75t_R _34731_ (.A(_18442_),
    .Y(_17968_));
 INVx1_ASAP7_75t_R _34732_ (.A(_18421_),
    .Y(_17969_));
 INVx1_ASAP7_75t_R _34733_ (.A(_18393_),
    .Y(_17919_));
 INVx1_ASAP7_75t_R _34734_ (.A(_18392_),
    .Y(_17917_));
 INVx1_ASAP7_75t_R _34735_ (.A(_18395_),
    .Y(_17866_));
 INVx1_ASAP7_75t_R _34736_ (.A(_18365_),
    .Y(_17867_));
 INVx1_ASAP7_75t_R _34737_ (.A(_18386_),
    .Y(_17856_));
 INVx1_ASAP7_75t_R _34738_ (.A(_18361_),
    .Y(_17857_));
 INVx1_ASAP7_75t_R _34739_ (.A(_18357_),
    .Y(_17801_));
 INVx1_ASAP7_75t_R _34740_ (.A(_18332_),
    .Y(_17802_));
 INVx1_ASAP7_75t_R _34741_ (.A(_18492_),
    .Y(_18066_));
 INVx1_ASAP7_75t_R _34742_ (.A(_18469_),
    .Y(_18067_));
 INVx1_ASAP7_75t_R _34743_ (.A(_00154_),
    .Y(_17367_));
 INVx1_ASAP7_75t_R _34744_ (.A(_00148_),
    .Y(_17368_));
 INVx1_ASAP7_75t_R _34745_ (.A(_00152_),
    .Y(_17375_));
 INVx1_ASAP7_75t_R _34746_ (.A(_18564_),
    .Y(_18188_));
 INVx1_ASAP7_75t_R _34747_ (.A(_18545_),
    .Y(_18189_));
 INVx1_ASAP7_75t_R _34748_ (.A(_18906_),
    .Y(_17363_));
 INVx1_ASAP7_75t_R _34749_ (.A(_18540_),
    .Y(_18149_));
 INVx1_ASAP7_75t_R _34750_ (.A(_18522_),
    .Y(_18150_));
 INVx1_ASAP7_75t_R _34751_ (.A(_00273_),
    .Y(_18296_));
 INVx1_ASAP7_75t_R _34752_ (.A(_02249_),
    .Y(_18311_));
 INVx1_ASAP7_75t_R _34753_ (.A(_18918_),
    .Y(_17379_));
 INVx1_ASAP7_75t_R _34754_ (.A(_19079_),
    .Y(_17713_));
 INVx1_ASAP7_75t_R _34755_ (.A(_19060_),
    .Y(_17714_));
 INVx1_ASAP7_75t_R _34756_ (.A(_18368_),
    .Y(_17822_));
 INVx1_ASAP7_75t_R _34757_ (.A(_18341_),
    .Y(_17823_));
 INVx1_ASAP7_75t_R _34758_ (.A(_18905_),
    .Y(_17380_));
 INVx1_ASAP7_75t_R _34759_ (.A(_19078_),
    .Y(_17769_));
 INVx1_ASAP7_75t_R _34760_ (.A(_00142_),
    .Y(_18892_));
 INVx1_ASAP7_75t_R _34761_ (.A(_02324_),
    .Y(_18891_));
 INVx1_ASAP7_75t_R _34762_ (.A(_18485_),
    .Y(_18053_));
 INVx1_ASAP7_75t_R _34763_ (.A(_18462_),
    .Y(_18054_));
 INVx1_ASAP7_75t_R _34764_ (.A(_18459_),
    .Y(_17999_));
 INVx1_ASAP7_75t_R _34765_ (.A(_18438_),
    .Y(_18000_));
 INVx1_ASAP7_75t_R _34766_ (.A(_18433_),
    .Y(_17949_));
 INVx1_ASAP7_75t_R _34767_ (.A(_18410_),
    .Y(_17950_));
 INVx1_ASAP7_75t_R _34768_ (.A(_18405_),
    .Y(_17893_));
 INVx1_ASAP7_75t_R _34769_ (.A(_18380_),
    .Y(_17894_));
 INVx1_ASAP7_75t_R _34770_ (.A(_18379_),
    .Y(_17840_));
 INVx1_ASAP7_75t_R _34771_ (.A(_18354_),
    .Y(_17841_));
 INVx1_ASAP7_75t_R _34772_ (.A(_18436_),
    .Y(_17998_));
 INVx1_ASAP7_75t_R _34773_ (.A(_02237_),
    .Y(_17923_));
 INVx1_ASAP7_75t_R _34774_ (.A(_00236_),
    .Y(_17879_));
 INVx1_ASAP7_75t_R _34775_ (.A(_18413_),
    .Y(_17901_));
 INVx1_ASAP7_75t_R _34776_ (.A(_18384_),
    .Y(_17902_));
 INVx1_ASAP7_75t_R _34777_ (.A(_00209_),
    .Y(_17600_));
 INVx1_ASAP7_75t_R _34778_ (.A(_02345_),
    .Y(_17640_));
 INVx1_ASAP7_75t_R _34779_ (.A(_18358_),
    .Y(_17852_));
 INVx1_ASAP7_75t_R _34780_ (.A(_18514_),
    .Y(_18102_));
 INVx1_ASAP7_75t_R _34781_ (.A(_18516_),
    .Y(_18145_));
 INVx1_ASAP7_75t_R _34782_ (.A(_18539_),
    .Y(_18178_));
 INVx1_ASAP7_75t_R _34783_ (.A(_18467_),
    .Y(_18060_));
 INVx1_ASAP7_75t_R _34784_ (.A(_18489_),
    .Y(_18059_));
 INVx1_ASAP7_75t_R _34785_ (.A(_00224_),
    .Y(_17697_));
 INVx1_ASAP7_75t_R _34786_ (.A(_18491_),
    .Y(_18105_));
 INVx1_ASAP7_75t_R _34787_ (.A(_00195_),
    .Y(_18975_));
 INVx1_ASAP7_75t_R _34788_ (.A(_18536_),
    .Y(_18146_));
 INVx1_ASAP7_75t_R _34789_ (.A(_18541_),
    .Y(_18180_));
 INVx1_ASAP7_75t_R _34790_ (.A(_18583_),
    .Y(_18234_));
 INVx1_ASAP7_75t_R _34791_ (.A(_00159_),
    .Y(_18913_));
 INVx1_ASAP7_75t_R _34792_ (.A(_02331_),
    .Y(_17409_));
 INVx1_ASAP7_75t_R _34793_ (.A(_00163_),
    .Y(_18921_));
 INVx1_ASAP7_75t_R _34794_ (.A(_18563_),
    .Y(_18217_));
 INVx1_ASAP7_75t_R _34795_ (.A(_18579_),
    .Y(_18216_));
 INVx1_ASAP7_75t_R _34796_ (.A(_18429_),
    .Y(_17986_));
 INVx1_ASAP7_75t_R _34797_ (.A(_18451_),
    .Y(_17985_));
 INVx1_ASAP7_75t_R _34798_ (.A(_19066_),
    .Y(_17678_));
 INVx1_ASAP7_75t_R _34799_ (.A(_19049_),
    .Y(_17679_));
 INVx1_ASAP7_75t_R _34800_ (.A(_18560_),
    .Y(_18208_));
 INVx1_ASAP7_75t_R _34801_ (.A(_18589_),
    .Y(_18246_));
 INVx1_ASAP7_75t_R _34802_ (.A(_18494_),
    .Y(_18109_));
 INVx1_ASAP7_75t_R _34803_ (.A(_18490_),
    .Y(_18103_));
 INVx1_ASAP7_75t_R _34804_ (.A(_18538_),
    .Y(_18144_));
 INVx1_ASAP7_75t_R _34805_ (.A(_19067_),
    .Y(_17687_));
 INVx1_ASAP7_75t_R _34806_ (.A(_19053_),
    .Y(_17688_));
 INVx1_ASAP7_75t_R _34807_ (.A(_18041_),
    .Y(_17994_));
 INVx1_ASAP7_75t_R _34808_ (.A(_18512_),
    .Y(_18104_));
 INVx1_ASAP7_75t_R _34809_ (.A(_18572_),
    .Y(_18202_));
 INVx1_ASAP7_75t_R _34810_ (.A(_18518_),
    .Y(_18147_));
 INVx1_ASAP7_75t_R _34811_ (.A(_18559_),
    .Y(_18179_));
 INVx1_ASAP7_75t_R _34812_ (.A(_02246_),
    .Y(_18244_));
 INVx1_ASAP7_75t_R _34813_ (.A(_18233_),
    .Y(_18198_));
 INVx1_ASAP7_75t_R _34814_ (.A(_18455_),
    .Y(_18040_));
 INVx1_ASAP7_75t_R _34815_ (.A(_18478_),
    .Y(_18039_));
 INVx1_ASAP7_75t_R _34816_ (.A(_18480_),
    .Y(_18083_));
 INVx1_ASAP7_75t_R _34817_ (.A(_00196_),
    .Y(_17529_));
 INVx1_ASAP7_75t_R _34818_ (.A(_02340_),
    .Y(_17563_));
 INVx1_ASAP7_75t_R _34819_ (.A(_18550_),
    .Y(_18199_));
 INVx1_ASAP7_75t_R _34820_ (.A(_18940_),
    .Y(_17416_));
 INVx1_ASAP7_75t_R _34821_ (.A(_18382_),
    .Y(_17899_));
 INVx1_ASAP7_75t_R _34822_ (.A(_18999_),
    .Y(_17521_));
 INVx1_ASAP7_75t_R _34823_ (.A(_00219_),
    .Y(_17659_));
 INVx1_ASAP7_75t_R _34824_ (.A(_02349_),
    .Y(_17698_));
 INVx1_ASAP7_75t_R _34825_ (.A(_02232_),
    .Y(_18310_));
 INVx1_ASAP7_75t_R _34826_ (.A(_18515_),
    .Y(_18108_));
 INVx1_ASAP7_75t_R _34827_ (.A(_18926_),
    .Y(_17417_));
 INVx1_ASAP7_75t_R _34828_ (.A(_18383_),
    .Y(_17851_));
 INVx1_ASAP7_75t_R _34829_ (.A(_02350_),
    .Y(_17709_));
 INVx1_ASAP7_75t_R _34830_ (.A(_18381_),
    .Y(_17846_));
 INVx1_ASAP7_75t_R _34831_ (.A(_19016_),
    .Y(_17605_));
 INVx1_ASAP7_75t_R _34832_ (.A(_18981_),
    .Y(_17522_));
 INVx1_ASAP7_75t_R _34833_ (.A(_02327_),
    .Y(_18898_));
 INVx1_ASAP7_75t_R _34834_ (.A(_00149_),
    .Y(_18899_));
 INVx1_ASAP7_75t_R _34835_ (.A(_18359_),
    .Y(_17806_));
 INVx1_ASAP7_75t_R _34836_ (.A(_02348_),
    .Y(_17683_));
 INVx1_ASAP7_75t_R _34837_ (.A(_00214_),
    .Y(_17641_));
 INVx1_ASAP7_75t_R _34838_ (.A(_18434_),
    .Y(_17947_));
 INVx1_ASAP7_75t_R _34839_ (.A(_18408_),
    .Y(_17948_));
 INVx1_ASAP7_75t_R _34840_ (.A(_18407_),
    .Y(_17898_));
 INVx1_ASAP7_75t_R _34841_ (.A(_00194_),
    .Y(_18973_));
 INVx1_ASAP7_75t_R _34842_ (.A(_02240_),
    .Y(_18051_));
 INVx1_ASAP7_75t_R _34843_ (.A(_00245_),
    .Y(_18006_));
 INVx1_ASAP7_75t_R _34844_ (.A(_02241_),
    .Y(_18089_));
 INVx1_ASAP7_75t_R _34845_ (.A(_00248_),
    .Y(_18049_));
 INVx1_ASAP7_75t_R _34846_ (.A(_00143_),
    .Y(_18894_));
 INVx1_ASAP7_75t_R _34847_ (.A(_02325_),
    .Y(_18893_));
 INVx1_ASAP7_75t_R _34848_ (.A(_00150_),
    .Y(_18900_));
 INVx1_ASAP7_75t_R _34849_ (.A(_00277_),
    .Y(_18309_));
 INVx1_ASAP7_75t_R _34850_ (.A(_18435_),
    .Y(_17955_));
 INVx1_ASAP7_75t_R _34851_ (.A(_18414_),
    .Y(_17956_));
 INVx1_ASAP7_75t_R _34852_ (.A(_18412_),
    .Y(_17954_));
 INVx1_ASAP7_75t_R _34853_ (.A(_18411_),
    .Y(_17908_));
 INVx1_ASAP7_75t_R _34854_ (.A(_18387_),
    .Y(_17909_));
 INVx1_ASAP7_75t_R _34855_ (.A(_18506_),
    .Y(_18091_));
 INVx1_ASAP7_75t_R _34856_ (.A(_18484_),
    .Y(_18092_));
 INVx1_ASAP7_75t_R _34857_ (.A(_18481_),
    .Y(_18044_));
 INVx1_ASAP7_75t_R _34858_ (.A(_18458_),
    .Y(_18045_));
 INVx1_ASAP7_75t_R _34859_ (.A(_18454_),
    .Y(_17990_));
 INVx1_ASAP7_75t_R _34860_ (.A(_18432_),
    .Y(_17991_));
 INVx1_ASAP7_75t_R _34861_ (.A(_18428_),
    .Y(_17939_));
 INVx1_ASAP7_75t_R _34862_ (.A(_18404_),
    .Y(_17940_));
 INVx1_ASAP7_75t_R _34863_ (.A(_18402_),
    .Y(_17887_));
 INVx1_ASAP7_75t_R _34864_ (.A(_18378_),
    .Y(_17888_));
 INVx1_ASAP7_75t_R _34865_ (.A(_18457_),
    .Y(_18043_));
 INVx1_ASAP7_75t_R _34866_ (.A(_18456_),
    .Y(_17988_));
 INVx1_ASAP7_75t_R _34867_ (.A(_18431_),
    .Y(_17989_));
 INVx1_ASAP7_75t_R _34868_ (.A(_18430_),
    .Y(_17944_));
 INVx1_ASAP7_75t_R _34869_ (.A(_18406_),
    .Y(_17945_));
 INVx1_ASAP7_75t_R _34870_ (.A(_18525_),
    .Y(_18125_));
 INVx1_ASAP7_75t_R _34871_ (.A(_18505_),
    .Y(_18126_));
 INVx1_ASAP7_75t_R _34872_ (.A(_18502_),
    .Y(_18082_));
 INVx1_ASAP7_75t_R _34873_ (.A(_18475_),
    .Y(_18031_));
 INVx1_ASAP7_75t_R _34874_ (.A(_18453_),
    .Y(_18032_));
 INVx1_ASAP7_75t_R _34875_ (.A(_18449_),
    .Y(_17980_));
 INVx1_ASAP7_75t_R _34876_ (.A(_18427_),
    .Y(_17981_));
 INVx1_ASAP7_75t_R _34877_ (.A(_18426_),
    .Y(_17933_));
 INVx1_ASAP7_75t_R _34878_ (.A(_18403_),
    .Y(_17934_));
 INVx1_ASAP7_75t_R _34879_ (.A(_18479_),
    .Y(_18081_));
 INVx1_ASAP7_75t_R _34880_ (.A(_18934_),
    .Y(_17404_));
 INVx1_ASAP7_75t_R _34881_ (.A(_19005_),
    .Y(_17574_));
 INVx1_ASAP7_75t_R _34882_ (.A(_19023_),
    .Y(_17573_));
 INVx1_ASAP7_75t_R _34883_ (.A(_18569_),
    .Y(_18232_));
 INVx1_ASAP7_75t_R _34884_ (.A(_18575_),
    .Y(_18207_));
 INVx1_ASAP7_75t_R _34885_ (.A(_18573_),
    .Y(_18236_));
 INVx1_ASAP7_75t_R _34886_ (.A(_18554_),
    .Y(_18203_));
 INVx1_ASAP7_75t_R _34887_ (.A(_19071_),
    .Y(_17747_));
 INVx1_ASAP7_75t_R _34888_ (.A(_18331_),
    .Y(_17746_));
 INVx1_ASAP7_75t_R _34889_ (.A(_00170_),
    .Y(_18925_));
 INVx1_ASAP7_75t_R _34890_ (.A(_18339_),
    .Y(_17817_));
 INVx1_ASAP7_75t_R _34891_ (.A(_18364_),
    .Y(_17816_));
 INVx1_ASAP7_75t_R _34892_ (.A(_18418_),
    .Y(_17918_));
 INVx1_ASAP7_75t_R _34893_ (.A(_02329_),
    .Y(_18903_));
 INVx1_ASAP7_75t_R _34894_ (.A(_18571_),
    .Y(_18235_));
 INVx1_ASAP7_75t_R _34895_ (.A(_18578_),
    .Y(_18247_));
 INVx1_ASAP7_75t_R _34896_ (.A(_18567_),
    .Y(_18200_));
 INVx1_ASAP7_75t_R _34897_ (.A(_18552_),
    .Y(_18201_));
 INVx1_ASAP7_75t_R _34898_ (.A(_18556_),
    .Y(_18205_));
 INVx1_ASAP7_75t_R _34899_ (.A(_00160_),
    .Y(_17391_));
 INVx1_ASAP7_75t_R _34900_ (.A(_18998_),
    .Y(_17557_));
 INVx1_ASAP7_75t_R _34901_ (.A(_00156_),
    .Y(_18910_));
 INVx1_ASAP7_75t_R _34902_ (.A(_19013_),
    .Y(_17556_));
 INVx1_ASAP7_75t_R _34903_ (.A(_18570_),
    .Y(_18204_));
 INVx1_ASAP7_75t_R _34904_ (.A(_00263_),
    .Y(_18214_));
 INVx1_ASAP7_75t_R _34905_ (.A(_18452_),
    .Y(_18030_));
 INVx1_ASAP7_75t_R _34906_ (.A(_02333_),
    .Y(_17443_));
 INVx1_ASAP7_75t_R _34907_ (.A(_18356_),
    .Y(_17847_));
 INVx1_ASAP7_75t_R _34908_ (.A(_18340_),
    .Y(_17768_));
 INVx1_ASAP7_75t_R _34909_ (.A(_18558_),
    .Y(_18206_));
 INVx1_ASAP7_75t_R _34910_ (.A(_18977_),
    .Y(_17510_));
 INVx1_ASAP7_75t_R _34911_ (.A(_00177_),
    .Y(_17447_));
 INVx1_ASAP7_75t_R _34912_ (.A(_18477_),
    .Y(_18029_));
 INVx1_ASAP7_75t_R _34913_ (.A(_02330_),
    .Y(_18908_));
 INVx1_ASAP7_75t_R _34914_ (.A(_00155_),
    .Y(_18909_));
 INVx1_ASAP7_75t_R _34915_ (.A(_18593_),
    .Y(_18264_));
 INVx1_ASAP7_75t_R _34916_ (.A(_18574_),
    .Y(_18238_));
 INVx1_ASAP7_75t_R _34917_ (.A(_18585_),
    .Y(_18237_));
 INVx1_ASAP7_75t_R _34918_ (.A(_18994_),
    .Y(_17509_));
 INVx1_ASAP7_75t_R _34919_ (.A(_00174_),
    .Y(_18936_));
 INVx1_ASAP7_75t_R _34920_ (.A(_18996_),
    .Y(_17547_));
 INVx1_ASAP7_75t_R _34921_ (.A(_19011_),
    .Y(_17546_));
 INVx1_ASAP7_75t_R _34922_ (.A(_02239_),
    .Y(_18005_));
 INVx1_ASAP7_75t_R _34923_ (.A(_19002_),
    .Y(_17527_));
 INVx1_ASAP7_75t_R _34924_ (.A(_02247_),
    .Y(_18271_));
 INVx1_ASAP7_75t_R _34925_ (.A(_00180_),
    .Y(_18948_));
 INVx1_ASAP7_75t_R _34926_ (.A(_02336_),
    .Y(_18947_));
 INVx1_ASAP7_75t_R _34927_ (.A(_00182_),
    .Y(_17468_));
 INVx1_ASAP7_75t_R _34928_ (.A(_02337_),
    .Y(_17498_));
 INVx1_ASAP7_75t_R _34929_ (.A(_00188_),
    .Y(_18959_));
 INVx1_ASAP7_75t_R _34930_ (.A(_18447_),
    .Y(_18020_));
 INVx1_ASAP7_75t_R _34931_ (.A(_18472_),
    .Y(_18019_));
 INVx1_ASAP7_75t_R _34932_ (.A(_18450_),
    .Y(_18027_));
 INVx1_ASAP7_75t_R _34933_ (.A(_18473_),
    .Y(_18026_));
 INVx1_ASAP7_75t_R _34934_ (.A(_18474_),
    .Y(_18074_));
 INVx1_ASAP7_75t_R _34935_ (.A(_18499_),
    .Y(_18073_));
 INVx1_ASAP7_75t_R _34936_ (.A(_18500_),
    .Y(_18115_));
 INVx1_ASAP7_75t_R _34937_ (.A(_18425_),
    .Y(_17975_));
 INVx1_ASAP7_75t_R _34938_ (.A(_18446_),
    .Y(_17974_));
 INVx1_ASAP7_75t_R _34939_ (.A(_18448_),
    .Y(_18022_));
 INVx1_ASAP7_75t_R _34940_ (.A(_18470_),
    .Y(_18021_));
 INVx1_ASAP7_75t_R _34941_ (.A(_18476_),
    .Y(_18076_));
 INVx1_ASAP7_75t_R _34942_ (.A(_18497_),
    .Y(_18075_));
 INVx1_ASAP7_75t_R _34943_ (.A(_18501_),
    .Y(_18117_));
 INVx1_ASAP7_75t_R _34944_ (.A(_18521_),
    .Y(_18116_));
 INVx1_ASAP7_75t_R _34945_ (.A(_18526_),
    .Y(_18159_));
 INVx1_ASAP7_75t_R _34946_ (.A(_18544_),
    .Y(_18158_));
 INVx1_ASAP7_75t_R _34947_ (.A(_02238_),
    .Y(_17966_));
 INVx1_ASAP7_75t_R _34948_ (.A(_00141_),
    .Y(_18888_));
 INVx1_ASAP7_75t_R _34949_ (.A(_02323_),
    .Y(_17365_));
 INVx1_ASAP7_75t_R _34950_ (.A(_00213_),
    .Y(_17632_));
 INVx1_ASAP7_75t_R _34951_ (.A(_02347_),
    .Y(_17674_));
 INVx1_ASAP7_75t_R _34952_ (.A(_00144_),
    .Y(_18895_));
 INVx1_ASAP7_75t_R _34953_ (.A(_00260_),
    .Y(_18186_));
 INVx1_ASAP7_75t_R _34954_ (.A(_02245_),
    .Y(_18213_));
 INVx1_ASAP7_75t_R _34955_ (.A(_18978_),
    .Y(_17516_));
 INVx1_ASAP7_75t_R _34956_ (.A(_18997_),
    .Y(_17515_));
 INVx1_ASAP7_75t_R _34957_ (.A(_02351_),
    .Y(_17736_));
 INVx1_ASAP7_75t_R _34958_ (.A(_19012_),
    .Y(_17596_));
 INVx1_ASAP7_75t_R _34959_ (.A(_19031_),
    .Y(_17595_));
 INVx1_ASAP7_75t_R _34960_ (.A(_00203_),
    .Y(_17559_));
 INVx1_ASAP7_75t_R _34961_ (.A(_02343_),
    .Y(_17599_));
 INVx1_ASAP7_75t_R _34962_ (.A(_00207_),
    .Y(_17569_));
 INVx1_ASAP7_75t_R _34963_ (.A(_19035_),
    .Y(_17646_));
 INVx1_ASAP7_75t_R _34964_ (.A(_19054_),
    .Y(_17645_));
 INVx1_ASAP7_75t_R _34965_ (.A(_00269_),
    .Y(_18269_));
 INVx1_ASAP7_75t_R _34966_ (.A(_02248_),
    .Y(_18295_));
 INVx1_ASAP7_75t_R _34967_ (.A(_18596_),
    .Y(_18299_));
 INVx1_ASAP7_75t_R _34968_ (.A(_18603_),
    .Y(_18298_));
 INVx1_ASAP7_75t_R _34969_ (.A(_00145_),
    .Y(_18896_));
 INVx1_ASAP7_75t_R _34970_ (.A(_19046_),
    .Y(_17618_));
 INVx1_ASAP7_75t_R _34971_ (.A(_18965_),
    .Y(_17492_));
 INVx1_ASAP7_75t_R _34972_ (.A(_18982_),
    .Y(_17491_));
 INVx1_ASAP7_75t_R _34973_ (.A(_00175_),
    .Y(_18938_));
 INVx1_ASAP7_75t_R _34974_ (.A(_02334_),
    .Y(_17467_));
 INVx1_ASAP7_75t_R _34975_ (.A(_00164_),
    .Y(_18922_));
 INVx1_ASAP7_75t_R _34976_ (.A(_02326_),
    .Y(_18897_));
 INVx1_ASAP7_75t_R _34977_ (.A(_00161_),
    .Y(_18915_));
 INVx1_ASAP7_75t_R _34978_ (.A(_02332_),
    .Y(_18914_));
 INVx1_ASAP7_75t_R _34979_ (.A(_18985_),
    .Y(_17497_));
 INVx1_ASAP7_75t_R _34980_ (.A(_18369_),
    .Y(_17870_));
 INVx1_ASAP7_75t_R _34981_ (.A(_18371_),
    .Y(_17872_));
 INVx1_ASAP7_75t_R _34982_ (.A(_18394_),
    .Y(_17871_));
 INVx1_ASAP7_75t_R _34983_ (.A(_00183_),
    .Y(_17470_));
 INVx1_ASAP7_75t_R _34984_ (.A(_00184_),
    .Y(_17474_));
 INVx1_ASAP7_75t_R _34985_ (.A(_18510_),
    .Y(_18132_));
 INVx1_ASAP7_75t_R _34986_ (.A(_18530_),
    .Y(_18131_));
 INVx1_ASAP7_75t_R _34987_ (.A(_18529_),
    .Y(_18165_));
 INVx1_ASAP7_75t_R _34988_ (.A(_18548_),
    .Y(_18164_));
 INVx1_ASAP7_75t_R _34989_ (.A(_18531_),
    .Y(_18170_));
 INVx1_ASAP7_75t_R _34990_ (.A(_18553_),
    .Y(_18169_));
 INVx1_ASAP7_75t_R _34991_ (.A(_18532_),
    .Y(_18172_));
 INVx1_ASAP7_75t_R _34992_ (.A(_18551_),
    .Y(_18171_));
 INVx1_ASAP7_75t_R _34993_ (.A(_18961_),
    .Y(_17482_));
 INVx1_ASAP7_75t_R _34994_ (.A(_18976_),
    .Y(_17481_));
 INVx1_ASAP7_75t_R _34995_ (.A(_18511_),
    .Y(_18137_));
 INVx1_ASAP7_75t_R _34996_ (.A(_18534_),
    .Y(_18136_));
 INVx1_ASAP7_75t_R _34997_ (.A(_18535_),
    .Y(_18175_));
 INVx1_ASAP7_75t_R _34998_ (.A(_18557_),
    .Y(_18174_));
 INVx1_ASAP7_75t_R _34999_ (.A(_18488_),
    .Y(_18098_));
 INVx1_ASAP7_75t_R _35000_ (.A(_18509_),
    .Y(_18097_));
 INVx1_ASAP7_75t_R _35001_ (.A(_18513_),
    .Y(_18139_));
 INVx1_ASAP7_75t_R _35002_ (.A(_18533_),
    .Y(_18138_));
 INVx1_ASAP7_75t_R _35003_ (.A(_18537_),
    .Y(_18177_));
 INVx1_ASAP7_75t_R _35004_ (.A(_18555_),
    .Y(_18176_));
 INVx1_ASAP7_75t_R _35005_ (.A(_00176_),
    .Y(_17445_));
 INVx1_ASAP7_75t_R _35006_ (.A(_02335_),
    .Y(_17471_));
 INVx1_ASAP7_75t_R _35007_ (.A(_18979_),
    .Y(_17487_));
 INVx1_ASAP7_75t_R _35008_ (.A(_18230_),
    .Y(_18222_));
 INVx1_ASAP7_75t_R _35009_ (.A(_18549_),
    .Y(_18195_));
 INVx1_ASAP7_75t_R _35010_ (.A(_18231_),
    .Y(_18194_));
 INVx1_ASAP7_75t_R _35011_ (.A(_18568_),
    .Y(_18229_));
 INVx1_ASAP7_75t_R _35012_ (.A(_18259_),
    .Y(_18228_));
 INVx1_ASAP7_75t_R _35013_ (.A(_18582_),
    .Y(_18258_));
 INVx1_ASAP7_75t_R _35014_ (.A(_18290_),
    .Y(_18257_));
 INVx1_ASAP7_75t_R _35015_ (.A(_18289_),
    .Y(_18282_));
 INVx1_ASAP7_75t_R _35016_ (.A(_18592_),
    .Y(_18288_));
 INVx1_ASAP7_75t_R _35017_ (.A(_18600_),
    .Y(_18287_));
 INVx1_ASAP7_75t_R _35018_ (.A(_18602_),
    .Y(_18315_));
 INVx1_ASAP7_75t_R _35019_ (.A(_00200_),
    .Y(_18993_));
 INVx1_ASAP7_75t_R _35020_ (.A(_00201_),
    .Y(_17549_));
 INVx1_ASAP7_75t_R _35021_ (.A(_02342_),
    .Y(_17589_));
 INVx1_ASAP7_75t_R _35022_ (.A(_02322_),
    .Y(_18885_));
 INVx1_ASAP7_75t_R _35023_ (.A(_02318_),
    .Y(_18875_));
 INVx1_ASAP7_75t_R _35024_ (.A(_02319_),
    .Y(_18877_));
 INVx1_ASAP7_75t_R _35025_ (.A(_00139_),
    .Y(_18883_));
 INVx1_ASAP7_75t_R _35026_ (.A(_02321_),
    .Y(_18882_));
 INVx1_ASAP7_75t_R _35027_ (.A(_00138_),
    .Y(_18881_));
 INVx1_ASAP7_75t_R _35028_ (.A(_02320_),
    .Y(_18880_));
 INVx1_ASAP7_75t_R _35029_ (.A(_18375_),
    .Y(_17882_));
 INVx1_ASAP7_75t_R _35030_ (.A(_18399_),
    .Y(_17881_));
 INVx1_ASAP7_75t_R _35031_ (.A(_02236_),
    .Y(_17878_));
 INVx1_ASAP7_75t_R _35032_ (.A(_00153_),
    .Y(_18904_));
 INVx1_ASAP7_75t_R _35033_ (.A(_02341_),
    .Y(_17561_));
 INVx1_ASAP7_75t_R _35034_ (.A(_00162_),
    .Y(_18916_));
 INVx1_ASAP7_75t_R _35035_ (.A(_18950_),
    .Y(_17452_));
 INVx1_ASAP7_75t_R _35036_ (.A(_18960_),
    .Y(_17451_));
 INVx1_ASAP7_75t_R _35037_ (.A(_02235_),
    .Y(_17833_));
 INVx1_ASAP7_75t_R _35038_ (.A(_18398_),
    .Y(_17928_));
 INVx1_ASAP7_75t_R _35039_ (.A(_18422_),
    .Y(_17927_));
 INVx2_ASAP7_75t_R _35040_ (.A(net1997),
    .Y(_17913_));
 INVx1_ASAP7_75t_R _35041_ (.A(_00189_),
    .Y(_18964_));
 INVx1_ASAP7_75t_R _35042_ (.A(_00181_),
    .Y(_18953_));
 AND2x2_ASAP7_75t_R _35043_ (.A(_05469_),
    .B(_05512_),
    .Y(_13230_));
 AND5x1_ASAP7_75t_R _35044_ (.A(_00289_),
    .B(_02227_),
    .C(_04922_),
    .D(_11060_),
    .E(_13230_),
    .Y(_13231_));
 INVx1_ASAP7_75t_R _35045_ (.A(_13231_),
    .Y(core_busy_d));
 AND2x2_ASAP7_75t_R _35046_ (.A(clknet_1_0__leaf_clk_i),
    .B(\core_clock_gate_i.en_latch ),
    .Y(clk));
 INVx1_ASAP7_75t_R _35047_ (.A(_02285_),
    .Y(_13232_));
 OR2x2_ASAP7_75t_R _35048_ (.A(_13561_),
    .B(_02284_),
    .Y(_13233_));
 OA211x2_ASAP7_75t_R _35049_ (.A1(_13573_),
    .A2(_12578_),
    .B(_05761_),
    .C(_13233_),
    .Y(_13234_));
 AO21x2_ASAP7_75t_R _35050_ (.A1(_13232_),
    .A2(_12579_),
    .B(_13234_),
    .Y(net230));
 INVx1_ASAP7_75t_R _35051_ (.A(_02286_),
    .Y(_13235_));
 INVx1_ASAP7_75t_R _35052_ (.A(_00359_),
    .Y(_13236_));
 NAND2x1_ASAP7_75t_R _35053_ (.A(_13573_),
    .B(_00360_),
    .Y(_13237_));
 OA211x2_ASAP7_75t_R _35054_ (.A1(_13573_),
    .A2(_13236_),
    .B(_05761_),
    .C(_13237_),
    .Y(_13238_));
 AO21x2_ASAP7_75t_R _35055_ (.A1(_13235_),
    .A2(_12579_),
    .B(_13238_),
    .Y(net231));
 INVx1_ASAP7_75t_R _35056_ (.A(_00362_),
    .Y(_13239_));
 INVx1_ASAP7_75t_R _35057_ (.A(_00361_),
    .Y(_13240_));
 OR3x1_ASAP7_75t_R _35058_ (.A(_13561_),
    .B(_00363_),
    .C(_12579_),
    .Y(_13241_));
 OA211x2_ASAP7_75t_R _35059_ (.A1(_13240_),
    .A2(_05761_),
    .B(_13241_),
    .C(_18763_),
    .Y(_13242_));
 INVx1_ASAP7_75t_R _35060_ (.A(_13242_),
    .Y(_13243_));
 INVx2_ASAP7_75t_R _35061_ (.A(_02287_),
    .Y(_13244_));
 BUFx4f_ASAP7_75t_R _35062_ (.A(_13244_),
    .Y(_13245_));
 AO21x1_ASAP7_75t_R _35063_ (.A1(_13245_),
    .A2(_12579_),
    .B(_18763_),
    .Y(_13246_));
 AO32x2_ASAP7_75t_R _35064_ (.A1(_13561_),
    .A2(_13239_),
    .A3(_05761_),
    .B1(_13243_),
    .B2(_13246_),
    .Y(net232));
 NAND2x1_ASAP7_75t_R _35065_ (.A(_13573_),
    .B(_00364_),
    .Y(_13247_));
 OA211x2_ASAP7_75t_R _35066_ (.A1(_13573_),
    .A2(_13245_),
    .B(_05761_),
    .C(_13247_),
    .Y(_13248_));
 AO21x2_ASAP7_75t_R _35067_ (.A1(_18763_),
    .A2(_12579_),
    .B(_13248_),
    .Y(net233));
 OA21x2_ASAP7_75t_R _35068_ (.A1(_13362_),
    .A2(_05754_),
    .B(_05751_),
    .Y(net234));
 BUFx6f_ASAP7_75t_R _35069_ (.A(_12578_),
    .Y(_13249_));
 BUFx6f_ASAP7_75t_R _35070_ (.A(_13249_),
    .Y(_13250_));
 BUFx3_ASAP7_75t_R _35071_ (.A(_02288_),
    .Y(_13251_));
 INVx1_ASAP7_75t_R _35072_ (.A(_02289_),
    .Y(_13252_));
 BUFx4f_ASAP7_75t_R _35073_ (.A(_13252_),
    .Y(_13253_));
 AOI22x1_ASAP7_75t_R _35074_ (.A1(_13245_),
    .A2(_05230_),
    .B1(_16094_),
    .B2(_13253_),
    .Y(_13254_));
 BUFx3_ASAP7_75t_R _35075_ (.A(_18762_),
    .Y(_13255_));
 OA211x2_ASAP7_75t_R _35076_ (.A1(_13251_),
    .A2(_17076_),
    .B(_13254_),
    .C(_13255_),
    .Y(_13256_));
 AOI21x1_ASAP7_75t_R _35077_ (.A1(_13250_),
    .A2(_05672_),
    .B(_13256_),
    .Y(net235));
 BUFx4f_ASAP7_75t_R _35078_ (.A(_18762_),
    .Y(_13257_));
 BUFx4f_ASAP7_75t_R _35079_ (.A(_18762_),
    .Y(_13258_));
 INVx1_ASAP7_75t_R _35080_ (.A(_14148_),
    .Y(_13259_));
 BUFx3_ASAP7_75t_R _35081_ (.A(_02289_),
    .Y(_13260_));
 INVx1_ASAP7_75t_R _35082_ (.A(_16354_),
    .Y(_13261_));
 BUFx3_ASAP7_75t_R _35083_ (.A(_02287_),
    .Y(_13262_));
 OA222x2_ASAP7_75t_R _35084_ (.A1(_13251_),
    .A2(_13259_),
    .B1(_17316_),
    .B2(_13260_),
    .C1(_13261_),
    .C2(_13262_),
    .Y(_13263_));
 NAND2x1_ASAP7_75t_R _35085_ (.A(_13258_),
    .B(_13263_),
    .Y(_13264_));
 OA21x2_ASAP7_75t_R _35086_ (.A1(_13257_),
    .A2(_14666_),
    .B(_13264_),
    .Y(net236));
 BUFx4f_ASAP7_75t_R _35087_ (.A(_02289_),
    .Y(_13265_));
 INVx2_ASAP7_75t_R _35088_ (.A(_02288_),
    .Y(_13266_));
 AOI22x1_ASAP7_75t_R _35089_ (.A1(_13266_),
    .A2(_14225_),
    .B1(_16466_),
    .B2(_13244_),
    .Y(_13267_));
 OA211x2_ASAP7_75t_R _35090_ (.A1(_13265_),
    .A2(_04343_),
    .B(_13267_),
    .C(_18762_),
    .Y(_13268_));
 AOI21x1_ASAP7_75t_R _35091_ (.A1(_13250_),
    .A2(_05589_),
    .B(_13268_),
    .Y(net237));
 BUFx4f_ASAP7_75t_R _35092_ (.A(_12578_),
    .Y(_13269_));
 BUFx3_ASAP7_75t_R _35093_ (.A(_02288_),
    .Y(_13270_));
 INVx1_ASAP7_75t_R _35094_ (.A(_14295_),
    .Y(_13271_));
 OA222x2_ASAP7_75t_R _35095_ (.A1(_13270_),
    .A2(_13271_),
    .B1(_04473_),
    .B2(_13260_),
    .C1(_16592_),
    .C2(_13262_),
    .Y(_13272_));
 NOR2x1_ASAP7_75t_R _35096_ (.A(_13249_),
    .B(_13272_),
    .Y(_13273_));
 AO21x2_ASAP7_75t_R _35097_ (.A1(_13269_),
    .A2(_05261_),
    .B(_13273_),
    .Y(net238));
 OA222x2_ASAP7_75t_R _35098_ (.A1(_13270_),
    .A2(_14371_),
    .B1(_04583_),
    .B2(_13260_),
    .C1(_16706_),
    .C2(_13262_),
    .Y(_13274_));
 NOR2x1_ASAP7_75t_R _35099_ (.A(_13249_),
    .B(_13274_),
    .Y(_13275_));
 AO21x2_ASAP7_75t_R _35100_ (.A1(_13269_),
    .A2(_15671_),
    .B(_13275_),
    .Y(net239));
 OA222x2_ASAP7_75t_R _35101_ (.A1(_13270_),
    .A2(_05558_),
    .B1(_04697_),
    .B2(_02289_),
    .C1(_16836_),
    .C2(_02287_),
    .Y(_13276_));
 NOR2x1_ASAP7_75t_R _35102_ (.A(_13249_),
    .B(_13276_),
    .Y(_13277_));
 AO21x2_ASAP7_75t_R _35103_ (.A1(_13269_),
    .A2(_15816_),
    .B(_13277_),
    .Y(net240));
 BUFx3_ASAP7_75t_R _35104_ (.A(_13266_),
    .Y(_13278_));
 AO222x2_ASAP7_75t_R _35105_ (.A1(_13278_),
    .A2(_14486_),
    .B1(_11085_),
    .B2(_13253_),
    .C1(_16946_),
    .C2(_13245_),
    .Y(_13279_));
 AND3x1_ASAP7_75t_R _35106_ (.A(_13249_),
    .B(_15911_),
    .C(_15949_),
    .Y(_13280_));
 AO21x2_ASAP7_75t_R _35107_ (.A1(_13257_),
    .A2(_13279_),
    .B(_13280_),
    .Y(net241));
 BUFx4f_ASAP7_75t_R _35108_ (.A(_02287_),
    .Y(_13281_));
 OAI22x1_ASAP7_75t_R _35109_ (.A1(_13265_),
    .A2(_05672_),
    .B1(_17076_),
    .B2(_13281_),
    .Y(_13282_));
 AO21x1_ASAP7_75t_R _35110_ (.A1(_13278_),
    .A2(_05230_),
    .B(_13282_),
    .Y(_13283_));
 AND3x1_ASAP7_75t_R _35111_ (.A(_13249_),
    .B(_16060_),
    .C(_16093_),
    .Y(_13284_));
 AO21x2_ASAP7_75t_R _35112_ (.A1(_13257_),
    .A2(_13283_),
    .B(_13284_),
    .Y(net242));
 OAI22x1_ASAP7_75t_R _35113_ (.A1(_13265_),
    .A2(_05528_),
    .B1(_17185_),
    .B2(_13281_),
    .Y(_13285_));
 AO21x1_ASAP7_75t_R _35114_ (.A1(_13278_),
    .A2(_14603_),
    .B(_13285_),
    .Y(_13286_));
 AND3x1_ASAP7_75t_R _35115_ (.A(_13249_),
    .B(_16177_),
    .C(_16208_),
    .Y(_13287_));
 AO21x2_ASAP7_75t_R _35116_ (.A1(_13257_),
    .A2(_13286_),
    .B(_13287_),
    .Y(net243));
 INVx1_ASAP7_75t_R _35117_ (.A(_14666_),
    .Y(_13288_));
 OA222x2_ASAP7_75t_R _35118_ (.A1(_13260_),
    .A2(_13259_),
    .B1(_13288_),
    .B2(_13270_),
    .C1(_13262_),
    .C2(_17316_),
    .Y(_13289_));
 NOR2x1_ASAP7_75t_R _35119_ (.A(_13249_),
    .B(_13289_),
    .Y(_13290_));
 AO21x2_ASAP7_75t_R _35120_ (.A1(_13269_),
    .A2(_16354_),
    .B(_13290_),
    .Y(net244));
 INVx1_ASAP7_75t_R _35121_ (.A(_16466_),
    .Y(_13291_));
 AOI22x1_ASAP7_75t_R _35122_ (.A1(_13253_),
    .A2(_14225_),
    .B1(_14723_),
    .B2(_13266_),
    .Y(_13292_));
 OA211x2_ASAP7_75t_R _35123_ (.A1(_13281_),
    .A2(_04343_),
    .B(_13292_),
    .C(_18762_),
    .Y(_13293_));
 AOI21x1_ASAP7_75t_R _35124_ (.A1(_13250_),
    .A2(_13291_),
    .B(_13293_),
    .Y(net245));
 AOI22x1_ASAP7_75t_R _35125_ (.A1(_13245_),
    .A2(_14603_),
    .B1(_16209_),
    .B2(_13253_),
    .Y(_13294_));
 OA211x2_ASAP7_75t_R _35126_ (.A1(_13251_),
    .A2(_17185_),
    .B(_13294_),
    .C(_18762_),
    .Y(_13295_));
 AOI21x1_ASAP7_75t_R _35127_ (.A1(_13269_),
    .A2(_05528_),
    .B(_13295_),
    .Y(net246));
 INVx1_ASAP7_75t_R _35128_ (.A(_05261_),
    .Y(_13296_));
 OA222x2_ASAP7_75t_R _35129_ (.A1(_13265_),
    .A2(_13271_),
    .B1(_13296_),
    .B2(_13251_),
    .C1(_13281_),
    .C2(_04473_),
    .Y(_13297_));
 OR2x2_ASAP7_75t_R _35130_ (.A(_13255_),
    .B(_16592_),
    .Y(_13298_));
 OAI21x1_ASAP7_75t_R _35131_ (.A1(_13250_),
    .A2(_13297_),
    .B(_13298_),
    .Y(net247));
 INVx1_ASAP7_75t_R _35132_ (.A(_15671_),
    .Y(_13299_));
 OA222x2_ASAP7_75t_R _35133_ (.A1(_13265_),
    .A2(_14371_),
    .B1(_13299_),
    .B2(_13251_),
    .C1(_13281_),
    .C2(_04583_),
    .Y(_13300_));
 OR2x2_ASAP7_75t_R _35134_ (.A(_13255_),
    .B(_16706_),
    .Y(_13301_));
 OAI21x1_ASAP7_75t_R _35135_ (.A1(_13250_),
    .A2(_13300_),
    .B(_13301_),
    .Y(net248));
 INVx1_ASAP7_75t_R _35136_ (.A(_15816_),
    .Y(_13302_));
 OA222x2_ASAP7_75t_R _35137_ (.A1(_13265_),
    .A2(_05558_),
    .B1(_13302_),
    .B2(_13251_),
    .C1(_13281_),
    .C2(_04697_),
    .Y(_13303_));
 OR2x2_ASAP7_75t_R _35138_ (.A(_13255_),
    .B(_16836_),
    .Y(_13304_));
 OAI21x1_ASAP7_75t_R _35139_ (.A1(_13250_),
    .A2(_13303_),
    .B(_13304_),
    .Y(net249));
 AO222x2_ASAP7_75t_R _35140_ (.A1(_13253_),
    .A2(_14486_),
    .B1(_15950_),
    .B2(_13278_),
    .C1(_13245_),
    .C2(_11085_),
    .Y(_13305_));
 AND3x1_ASAP7_75t_R _35141_ (.A(_13249_),
    .B(_16914_),
    .C(_16945_),
    .Y(_13306_));
 AO21x2_ASAP7_75t_R _35142_ (.A1(_13258_),
    .A2(_13305_),
    .B(_13306_),
    .Y(net250));
 AO32x1_ASAP7_75t_R _35143_ (.A1(_13244_),
    .A2(_13821_),
    .A3(_13852_),
    .B1(_05230_),
    .B2(_13253_),
    .Y(_13307_));
 AO21x1_ASAP7_75t_R _35144_ (.A1(_13278_),
    .A2(_16094_),
    .B(_13307_),
    .Y(_13308_));
 NAND2x1_ASAP7_75t_R _35145_ (.A(_13269_),
    .B(_17076_),
    .Y(_13309_));
 OA21x2_ASAP7_75t_R _35146_ (.A1(_13269_),
    .A2(_13308_),
    .B(_13309_),
    .Y(net251));
 AO32x1_ASAP7_75t_R _35147_ (.A1(_13244_),
    .A2(_13514_),
    .A3(_13549_),
    .B1(_14603_),
    .B2(_13252_),
    .Y(_13310_));
 AO21x1_ASAP7_75t_R _35148_ (.A1(_13278_),
    .A2(_16209_),
    .B(_13310_),
    .Y(_13311_));
 NAND2x1_ASAP7_75t_R _35149_ (.A(_13269_),
    .B(_17185_),
    .Y(_13312_));
 OA21x2_ASAP7_75t_R _35150_ (.A1(_13269_),
    .A2(_13311_),
    .B(_13312_),
    .Y(net252));
 AO222x2_ASAP7_75t_R _35151_ (.A1(_13245_),
    .A2(_14148_),
    .B1(_14666_),
    .B2(_13253_),
    .C1(_16354_),
    .C2(_13278_),
    .Y(_13313_));
 AND3x1_ASAP7_75t_R _35152_ (.A(_13249_),
    .B(_17284_),
    .C(_17315_),
    .Y(_13314_));
 AO21x2_ASAP7_75t_R _35153_ (.A1(_13258_),
    .A2(_13313_),
    .B(_13314_),
    .Y(net253));
 AO222x2_ASAP7_75t_R _35154_ (.A1(_13245_),
    .A2(_14225_),
    .B1(_14723_),
    .B2(_13253_),
    .C1(_16466_),
    .C2(_13278_),
    .Y(_13315_));
 AND3x1_ASAP7_75t_R _35155_ (.A(_12578_),
    .B(_04311_),
    .C(_04342_),
    .Y(_13316_));
 AO21x2_ASAP7_75t_R _35156_ (.A1(_13258_),
    .A2(_13315_),
    .B(_13316_),
    .Y(net254));
 OA222x2_ASAP7_75t_R _35157_ (.A1(_13281_),
    .A2(_13271_),
    .B1(_13296_),
    .B2(_13265_),
    .C1(_16592_),
    .C2(_13251_),
    .Y(_13317_));
 OR2x2_ASAP7_75t_R _35158_ (.A(_13255_),
    .B(_04473_),
    .Y(_13318_));
 OAI21x1_ASAP7_75t_R _35159_ (.A1(_13250_),
    .A2(_13317_),
    .B(_13318_),
    .Y(net255));
 OA222x2_ASAP7_75t_R _35160_ (.A1(_13281_),
    .A2(_14371_),
    .B1(_13299_),
    .B2(_13265_),
    .C1(_16706_),
    .C2(_13251_),
    .Y(_13319_));
 OR2x2_ASAP7_75t_R _35161_ (.A(_13255_),
    .B(_04583_),
    .Y(_13320_));
 OAI21x1_ASAP7_75t_R _35162_ (.A1(_13250_),
    .A2(_13319_),
    .B(_13320_),
    .Y(net256));
 OA222x2_ASAP7_75t_R _35163_ (.A1(_13262_),
    .A2(_13288_),
    .B1(_13261_),
    .B2(_13260_),
    .C1(_17316_),
    .C2(_13270_),
    .Y(_13321_));
 NAND2x1_ASAP7_75t_R _35164_ (.A(_13258_),
    .B(_13321_),
    .Y(_13322_));
 OA21x2_ASAP7_75t_R _35165_ (.A1(_13257_),
    .A2(_14148_),
    .B(_13322_),
    .Y(net257));
 OA222x2_ASAP7_75t_R _35166_ (.A1(_13281_),
    .A2(_05558_),
    .B1(_13302_),
    .B2(_13265_),
    .C1(_16836_),
    .C2(_13251_),
    .Y(_13323_));
 OR2x2_ASAP7_75t_R _35167_ (.A(_13255_),
    .B(_04697_),
    .Y(_13324_));
 OAI21x1_ASAP7_75t_R _35168_ (.A1(_13250_),
    .A2(_13323_),
    .B(_13324_),
    .Y(net258));
 AO222x2_ASAP7_75t_R _35169_ (.A1(_13245_),
    .A2(_14486_),
    .B1(_15950_),
    .B2(_13253_),
    .C1(_16946_),
    .C2(_13278_),
    .Y(_13325_));
 AO21x1_ASAP7_75t_R _35170_ (.A1(_04875_),
    .A2(_04876_),
    .B(_13255_),
    .Y(_13326_));
 OA21x2_ASAP7_75t_R _35171_ (.A1(_13269_),
    .A2(_13325_),
    .B(_13326_),
    .Y(net259));
 OA222x2_ASAP7_75t_R _35172_ (.A1(_13262_),
    .A2(_05589_),
    .B1(_13291_),
    .B2(_13260_),
    .C1(_04343_),
    .C2(_13270_),
    .Y(_13327_));
 NAND2x1_ASAP7_75t_R _35173_ (.A(_13258_),
    .B(_13327_),
    .Y(_13328_));
 OA21x2_ASAP7_75t_R _35174_ (.A1(_13257_),
    .A2(_14225_),
    .B(_13328_),
    .Y(net260));
 OA222x2_ASAP7_75t_R _35175_ (.A1(_13262_),
    .A2(_13296_),
    .B1(_16592_),
    .B2(_13260_),
    .C1(_04473_),
    .C2(_13270_),
    .Y(_13329_));
 NAND2x1_ASAP7_75t_R _35176_ (.A(_13258_),
    .B(_13329_),
    .Y(_13330_));
 OA21x2_ASAP7_75t_R _35177_ (.A1(_13257_),
    .A2(_14295_),
    .B(_13330_),
    .Y(net261));
 OA222x2_ASAP7_75t_R _35178_ (.A1(_13281_),
    .A2(_13299_),
    .B1(_16706_),
    .B2(_13265_),
    .C1(_04583_),
    .C2(_13251_),
    .Y(_13331_));
 OR2x2_ASAP7_75t_R _35179_ (.A(_13255_),
    .B(_14371_),
    .Y(_13332_));
 OAI21x1_ASAP7_75t_R _35180_ (.A1(_13250_),
    .A2(_13331_),
    .B(_13332_),
    .Y(net262));
 OA222x2_ASAP7_75t_R _35181_ (.A1(_13262_),
    .A2(_13302_),
    .B1(_16836_),
    .B2(_13260_),
    .C1(_04697_),
    .C2(_13270_),
    .Y(_13333_));
 NAND2x1_ASAP7_75t_R _35182_ (.A(_13258_),
    .B(_13333_),
    .Y(_13334_));
 OA21x2_ASAP7_75t_R _35183_ (.A1(_13257_),
    .A2(_14426_),
    .B(_13334_),
    .Y(net263));
 AO222x2_ASAP7_75t_R _35184_ (.A1(_13245_),
    .A2(_15950_),
    .B1(_16946_),
    .B2(_13253_),
    .C1(_11085_),
    .C2(_13278_),
    .Y(_13335_));
 AND2x2_ASAP7_75t_R _35185_ (.A(_12578_),
    .B(_14486_),
    .Y(_13336_));
 AO21x2_ASAP7_75t_R _35186_ (.A1(_13258_),
    .A2(_13335_),
    .B(_13336_),
    .Y(net264));
 INVx1_ASAP7_75t_R _35187_ (.A(_16094_),
    .Y(_13337_));
 OA222x2_ASAP7_75t_R _35188_ (.A1(_13270_),
    .A2(_05672_),
    .B1(_17076_),
    .B2(_13260_),
    .C1(_13337_),
    .C2(_13262_),
    .Y(_13338_));
 NAND2x1_ASAP7_75t_R _35189_ (.A(_13258_),
    .B(_13338_),
    .Y(_13339_));
 OA21x2_ASAP7_75t_R _35190_ (.A1(_13257_),
    .A2(_05230_),
    .B(_13339_),
    .Y(net265));
 OA222x2_ASAP7_75t_R _35191_ (.A1(_13270_),
    .A2(_05528_),
    .B1(_17185_),
    .B2(_13260_),
    .C1(_11114_),
    .C2(_13262_),
    .Y(_13340_));
 NAND2x1_ASAP7_75t_R _35192_ (.A(_13255_),
    .B(_13340_),
    .Y(_13341_));
 OA21x2_ASAP7_75t_R _35193_ (.A1(_13257_),
    .A2(_14603_),
    .B(_13341_),
    .Y(net266));
 OR2x2_ASAP7_75t_R _35194_ (.A(_08347_),
    .B(_08350_),
    .Y(_13342_));
 AND5x1_ASAP7_75t_R _35195_ (.A(_01776_),
    .B(_13570_),
    .C(_04928_),
    .D(_04940_),
    .E(_13342_),
    .Y(\id_stage_i.branch_set_d ));
 OAI21x1_ASAP7_75t_R _35196_ (.A1(net177),
    .A2(_11731_),
    .B(_11946_),
    .Y(_13343_));
 OA21x2_ASAP7_75t_R _35197_ (.A1(_00289_),
    .A2(_05468_),
    .B(_02224_),
    .Y(_13344_));
 AOI22x1_ASAP7_75t_R _35198_ (.A1(_02223_),
    .A2(_13343_),
    .B1(_13344_),
    .B2(_11963_),
    .Y(_13345_));
 AO21x1_ASAP7_75t_R _35199_ (.A1(net140),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .B(_13345_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 NAND3x1_ASAP7_75t_R _35200_ (.A(net140),
    .B(_11946_),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Y(_13346_));
 AOI21x1_ASAP7_75t_R _35201_ (.A1(_13344_),
    .A2(_13346_),
    .B(_11963_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 OA22x2_ASAP7_75t_R _35202_ (.A1(_11964_),
    .A2(_11984_),
    .B1(_11971_),
    .B2(_12637_),
    .Y(_13347_));
 AOI221x1_ASAP7_75t_R _35203_ (.A1(_11950_),
    .A2(_11984_),
    .B1(_13347_),
    .B2(_11959_),
    .C(_11709_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 OA211x2_ASAP7_75t_R _35204_ (.A1(_11962_),
    .A2(_12017_),
    .B(_11947_),
    .C(_05490_),
    .Y(_13348_));
 OR2x2_ASAP7_75t_R _35205_ (.A(_11962_),
    .B(_11947_),
    .Y(_13349_));
 OA21x2_ASAP7_75t_R _35206_ (.A1(_12637_),
    .A2(_13349_),
    .B(_11980_),
    .Y(_13350_));
 OA31x2_ASAP7_75t_R _35207_ (.A1(_12006_),
    .A2(_13348_),
    .A3(_13350_),
    .B1(_11704_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 OA21x2_ASAP7_75t_R _35208_ (.A1(_12263_),
    .A2(_11994_),
    .B(_11889_),
    .Y(_13351_));
 OA21x2_ASAP7_75t_R _35209_ (.A1(_11962_),
    .A2(_12793_),
    .B(_13351_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 INVx1_ASAP7_75t_R _35210_ (.A(_13230_),
    .Y(net298));
 AOI21x1_ASAP7_75t_R _35211_ (.A1(_00289_),
    .A2(net177),
    .B(_02227_),
    .Y(_13352_));
 AO21x1_ASAP7_75t_R _35212_ (.A1(net140),
    .A2(net298),
    .B(_13352_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 OR3x1_ASAP7_75t_R _35213_ (.A(_12468_),
    .B(_02227_),
    .C(_13230_),
    .Y(_13353_));
 AOI21x1_ASAP7_75t_R _35214_ (.A1(_00289_),
    .A2(_13353_),
    .B(_11963_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 AND2x2_ASAP7_75t_R _35215_ (.A(_12468_),
    .B(net298),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 AO21x1_ASAP7_75t_R _35216_ (.A1(_11064_),
    .A2(_11076_),
    .B(_11048_),
    .Y(_13354_));
 AO221x1_ASAP7_75t_R _35217_ (.A1(_05077_),
    .A2(_05335_),
    .B1(_13354_),
    .B2(_04934_),
    .C(_05062_),
    .Y(_13355_));
 OA21x2_ASAP7_75t_R _35218_ (.A1(_05423_),
    .A2(_11045_),
    .B(_12790_),
    .Y(_13356_));
 OAI22x1_ASAP7_75t_R _35219_ (.A1(_11709_),
    .A2(_12638_),
    .B1(_13355_),
    .B2(_13356_),
    .Y(\if_stage_i.instr_valid_id_d ));
 FAx1_ASAP7_75t_R _35220_ (.SN(_18769_),
    .A(_17344_),
    .B(_17345_),
    .CI(_17346_),
    .CON(_02229_));
 FAx1_ASAP7_75t_R _35221_ (.SN(_18876_),
    .A(_17347_),
    .B(_17348_),
    .CI(_17349_),
    .CON(_18878_));
 FAx1_ASAP7_75t_R _35222_ (.SN(_18879_),
    .A(_17350_),
    .B(_17351_),
    .CI(_17352_),
    .CON(_18889_));
 FAx1_ASAP7_75t_R _35223_ (.SN(_18890_),
    .A(_17353_),
    .B(_17354_),
    .CI(_17355_),
    .CON(_17364_));
 FAx1_ASAP7_75t_R _35224_ (.SN(_00147_),
    .A(_17356_),
    .B(_17357_),
    .CI(_17358_),
    .CON(_17381_));
 FAx1_ASAP7_75t_R _35225_ (.SN(_17366_),
    .A(_17360_),
    .B(_17361_),
    .CI(_17362_),
    .CON(_18906_));
 FAx1_ASAP7_75t_R _35226_ (.SN(_00148_),
    .A(_17364_),
    .B(_17365_),
    .CI(_17366_),
    .CON(_00154_));
 FAx1_ASAP7_75t_R _35227_ (.SN(_18901_),
    .A(_17369_),
    .B(_17370_),
    .CI(_17371_),
    .CON(_17387_));
 FAx1_ASAP7_75t_R _35228_ (.SN(_00152_),
    .A(_17372_),
    .B(_17373_),
    .CI(_17374_),
    .CON(_17397_));
 FAx1_ASAP7_75t_R _35229_ (.SN(_18905_),
    .A(_17376_),
    .B(_17377_),
    .CI(_17378_),
    .CON(_18918_));
 FAx1_ASAP7_75t_R _35230_ (.SN(_18907_),
    .A(_17363_),
    .B(_17381_),
    .CI(_17380_),
    .CON(_18919_));
 FAx1_ASAP7_75t_R _35231_ (.SN(_17386_),
    .A(_17382_),
    .B(_17383_),
    .CI(_17384_),
    .CON(_18924_));
 FAx1_ASAP7_75t_R _35232_ (.SN(_00158_),
    .A(_17385_),
    .B(_17386_),
    .CI(_17387_),
    .CON(_00167_));
 FAx1_ASAP7_75t_R _35233_ (.SN(_00160_),
    .A(_17388_),
    .B(_17389_),
    .CI(_17390_),
    .CON(_17418_));
 FAx1_ASAP7_75t_R _35234_ (.SN(_18917_),
    .A(_17392_),
    .B(_17393_),
    .CI(_17394_),
    .CON(_18927_));
 FAx1_ASAP7_75t_R _35235_ (.SN(_18920_),
    .A(_17397_),
    .B(_17396_),
    .CI(_17379_),
    .CON(_18929_));
 FAx1_ASAP7_75t_R _35236_ (.SN(_18923_),
    .A(_17398_),
    .B(_17399_),
    .CI(_17400_),
    .CON(_18932_));
 FAx1_ASAP7_75t_R _35237_ (.SN(_17410_),
    .A(_17401_),
    .B(_17402_),
    .CI(_17403_),
    .CON(_18934_));
 FAx1_ASAP7_75t_R _35238_ (.SN(_00168_),
    .A(_17405_),
    .B(_17406_),
    .CI(_17407_),
    .CON(_17439_));
 FAx1_ASAP7_75t_R _35239_ (.SN(_00169_),
    .A(_17409_),
    .B(_17408_),
    .CI(_17410_),
    .CON(_00173_));
 FAx1_ASAP7_75t_R _35240_ (.SN(_18926_),
    .A(_17413_),
    .B(_17414_),
    .CI(_17415_),
    .CON(_18940_));
 FAx1_ASAP7_75t_R _35241_ (.SN(_18928_),
    .A(_17395_),
    .B(_17418_),
    .CI(_17417_),
    .CON(_18942_));
 FAx1_ASAP7_75t_R _35242_ (.SN(_18930_),
    .A(_17419_),
    .B(_17420_),
    .CI(_17421_),
    .CON(_17444_));
 FAx1_ASAP7_75t_R _35243_ (.SN(_18931_),
    .A(_17422_),
    .B(_17423_),
    .CI(_17424_),
    .CON(_18944_));
 FAx1_ASAP7_75t_R _35244_ (.SN(_18933_),
    .A(_17425_),
    .B(_17426_),
    .CI(_17427_),
    .CON(_18949_));
 FAx1_ASAP7_75t_R _35245_ (.SN(_17433_),
    .A(_17430_),
    .B(_17431_),
    .CI(_17432_),
    .CON(_17462_));
 FAx1_ASAP7_75t_R _35246_ (.SN(_18935_),
    .A(_17433_),
    .B(_17429_),
    .CI(_17404_),
    .CON(_18952_));
 FAx1_ASAP7_75t_R _35247_ (.SN(_18939_),
    .A(_17434_),
    .B(_17435_),
    .CI(_17436_),
    .CON(_18955_));
 FAx1_ASAP7_75t_R _35248_ (.SN(_18941_),
    .A(_17439_),
    .B(_17438_),
    .CI(_17416_),
    .CON(_18957_));
 FAx1_ASAP7_75t_R _35249_ (.SN(_18943_),
    .A(_17440_),
    .B(_17441_),
    .CI(_17442_),
    .CON(_17472_));
 FAx1_ASAP7_75t_R _35250_ (.SN(_00177_),
    .A(_17443_),
    .B(_17444_),
    .CI(_17445_),
    .CON(_00185_));
 FAx1_ASAP7_75t_R _35251_ (.SN(_18950_),
    .A(_17448_),
    .B(_17449_),
    .CI(_17450_),
    .CON(_18960_));
 FAx1_ASAP7_75t_R _35252_ (.SN(_17456_),
    .A(_17453_),
    .B(_17454_),
    .CI(_17455_),
    .CON(_17493_));
 FAx1_ASAP7_75t_R _35253_ (.SN(_18951_),
    .A(_17428_),
    .B(_17456_),
    .CI(_17452_),
    .CON(_18963_));
 FAx1_ASAP7_75t_R _35254_ (.SN(_18954_),
    .A(_17457_),
    .B(_17458_),
    .CI(_17459_),
    .CON(_18966_));
 FAx1_ASAP7_75t_R _35255_ (.SN(_18956_),
    .A(_17462_),
    .B(_17461_),
    .CI(_17437_),
    .CON(_18968_));
 FAx1_ASAP7_75t_R _35256_ (.SN(_17469_),
    .A(_17463_),
    .B(_17464_),
    .CI(_17465_),
    .CON(_18969_));
 FAx1_ASAP7_75t_R _35257_ (.SN(_00183_),
    .A(_17467_),
    .B(_17468_),
    .CI(_17469_),
    .CON(_17502_));
 FAx1_ASAP7_75t_R _35258_ (.SN(_00184_),
    .A(_17471_),
    .B(_17472_),
    .CI(_17470_),
    .CON(_00191_));
 FAx1_ASAP7_75t_R _35259_ (.SN(_18958_),
    .A(_17475_),
    .B(_17476_),
    .CI(_17477_),
    .CON(_18971_));
 FAx1_ASAP7_75t_R _35260_ (.SN(_18961_),
    .A(_17478_),
    .B(_17479_),
    .CI(_17480_),
    .CON(_18976_));
 FAx1_ASAP7_75t_R _35261_ (.SN(_17486_),
    .A(_17483_),
    .B(_17484_),
    .CI(_17485_),
    .CON(_17523_));
 FAx1_ASAP7_75t_R _35262_ (.SN(_18962_),
    .A(_17451_),
    .B(_17486_),
    .CI(_17482_),
    .CON(_18979_));
 FAx1_ASAP7_75t_R _35263_ (.SN(_18965_),
    .A(_17488_),
    .B(_17489_),
    .CI(_17490_),
    .CON(_18982_));
 FAx1_ASAP7_75t_R _35264_ (.SN(_18967_),
    .A(_17493_),
    .B(_17492_),
    .CI(_17460_),
    .CON(_18984_));
 FAx1_ASAP7_75t_R _35265_ (.SN(_17500_),
    .A(_17494_),
    .B(_17495_),
    .CI(_17496_),
    .CON(_18985_));
 FAx1_ASAP7_75t_R _35266_ (.SN(_17501_),
    .A(_17498_),
    .B(_17499_),
    .CI(_17500_),
    .CON(_17532_));
 FAx1_ASAP7_75t_R _35267_ (.SN(_18970_),
    .A(_17501_),
    .B(_17502_),
    .CI(_17466_),
    .CON(_18987_));
 FAx1_ASAP7_75t_R _35268_ (.SN(_18972_),
    .A(_17503_),
    .B(_17504_),
    .CI(_17505_),
    .CON(_18992_));
 FAx1_ASAP7_75t_R _35269_ (.SN(_18977_),
    .A(_17506_),
    .B(_17507_),
    .CI(_17508_),
    .CON(_18994_));
 FAx1_ASAP7_75t_R _35270_ (.SN(_17514_),
    .A(_17511_),
    .B(_17512_),
    .CI(_17513_),
    .CON(_17558_));
 FAx1_ASAP7_75t_R _35271_ (.SN(_18978_),
    .A(_17481_),
    .B(_17514_),
    .CI(_17510_),
    .CON(_18997_));
 FAx1_ASAP7_75t_R _35272_ (.SN(_18980_),
    .A(_17517_),
    .B(_17516_),
    .CI(_17487_),
    .CON(_17560_));
 FAx1_ASAP7_75t_R _35273_ (.SN(_18981_),
    .A(_17518_),
    .B(_17519_),
    .CI(_17520_),
    .CON(_18999_));
 FAx1_ASAP7_75t_R _35274_ (.SN(_18983_),
    .A(_17523_),
    .B(_17522_),
    .CI(_17491_),
    .CON(_19001_));
 FAx1_ASAP7_75t_R _35275_ (.SN(_17530_),
    .A(_17524_),
    .B(_17525_),
    .CI(_17526_),
    .CON(_19002_));
 FAx1_ASAP7_75t_R _35276_ (.SN(_17531_),
    .A(_17528_),
    .B(_17529_),
    .CI(_17530_),
    .CON(_17565_));
 FAx1_ASAP7_75t_R _35277_ (.SN(_18986_),
    .A(_17531_),
    .B(_17532_),
    .CI(_17497_),
    .CON(_19004_));
 FAx1_ASAP7_75t_R _35278_ (.SN(_18991_),
    .A(_17533_),
    .B(_17534_),
    .CI(_17535_),
    .CON(_19006_));
 FAx1_ASAP7_75t_R _35279_ (.SN(_18995_),
    .A(_17537_),
    .B(_17538_),
    .CI(_17539_),
    .CON(_19009_));
 FAx1_ASAP7_75t_R _35280_ (.SN(_17545_),
    .A(_17543_),
    .B(_17542_),
    .CI(_17544_),
    .CON(_17597_));
 FAx1_ASAP7_75t_R _35281_ (.SN(_18996_),
    .A(_17509_),
    .B(_17545_),
    .CI(_17541_),
    .CON(_19011_));
 FAx1_ASAP7_75t_R _35282_ (.SN(_17550_),
    .A(_17547_),
    .B(_17548_),
    .CI(_17515_),
    .CON(_17598_));
 FAx1_ASAP7_75t_R _35283_ (.SN(_00202_),
    .A(_17549_),
    .B(_17551_),
    .CI(_17550_),
    .CON(_17603_));
 FAx1_ASAP7_75t_R _35284_ (.SN(_18998_),
    .A(_17553_),
    .B(_17554_),
    .CI(_17555_),
    .CON(_19013_));
 FAx1_ASAP7_75t_R _35285_ (.SN(_19000_),
    .A(_17558_),
    .B(_17557_),
    .CI(_17521_),
    .CON(_19015_));
 FAx1_ASAP7_75t_R _35286_ (.SN(_00204_),
    .A(_17559_),
    .B(_17560_),
    .CI(_17561_),
    .CON(_17607_));
 FAx1_ASAP7_75t_R _35287_ (.SN(_17564_),
    .A(_17552_),
    .B(_17563_),
    .CI(_17562_),
    .CON(_17606_));
 FAx1_ASAP7_75t_R _35288_ (.SN(_19003_),
    .A(_17564_),
    .B(_17565_),
    .CI(_17527_),
    .CON(_19017_));
 FAx1_ASAP7_75t_R _35289_ (.SN(_00207_),
    .A(_17566_),
    .B(_17567_),
    .CI(_17568_),
    .CON(_17617_));
 FAx1_ASAP7_75t_R _35290_ (.SN(_19005_),
    .A(_17570_),
    .B(_17571_),
    .CI(_17572_),
    .CON(_19023_));
 FAx1_ASAP7_75t_R _35291_ (.SN(_19007_),
    .A(_17575_),
    .B(_17574_),
    .CI(_17536_),
    .CON(_19027_));
 FAx1_ASAP7_75t_R _35292_ (.SN(_19008_),
    .A(_17577_),
    .B(_17578_),
    .CI(_17579_),
    .CON(_19026_));
 FAx1_ASAP7_75t_R _35293_ (.SN(_17585_),
    .A(_17582_),
    .B(_17583_),
    .CI(_17584_),
    .CON(_17638_));
 FAx1_ASAP7_75t_R _35294_ (.SN(_19010_),
    .A(_17581_),
    .B(_17540_),
    .CI(_17585_),
    .CON(_19029_));
 FAx1_ASAP7_75t_R _35295_ (.SN(_17591_),
    .A(_17588_),
    .B(_17587_),
    .CI(_17546_),
    .CON(_17639_));
 FAx1_ASAP7_75t_R _35296_ (.SN(_17601_),
    .A(_17589_),
    .B(_17590_),
    .CI(_17591_),
    .CON(_17644_));
 FAx1_ASAP7_75t_R _35297_ (.SN(_19012_),
    .A(_17592_),
    .B(_17593_),
    .CI(_17594_),
    .CON(_19031_));
 FAx1_ASAP7_75t_R _35298_ (.SN(_19014_),
    .A(_17597_),
    .B(_17596_),
    .CI(_17556_),
    .CON(_19033_));
 FAx1_ASAP7_75t_R _35299_ (.SN(_17602_),
    .A(_17598_),
    .B(_17599_),
    .CI(_17600_),
    .CON(_17647_));
 FAx1_ASAP7_75t_R _35300_ (.SN(_19016_),
    .A(_17601_),
    .B(_17602_),
    .CI(_17603_),
    .CON(_19034_));
 FAx1_ASAP7_75t_R _35301_ (.SN(_19018_),
    .A(_17606_),
    .B(_17607_),
    .CI(_17605_),
    .CON(_19036_));
 FAx1_ASAP7_75t_R _35302_ (.SN(_19019_),
    .A(_17608_),
    .B(_17609_),
    .CI(_17610_),
    .CON(_19042_));
 FAx1_ASAP7_75t_R _35303_ (.SN(_19022_),
    .A(_17612_),
    .B(_17613_),
    .CI(_17614_),
    .CON(_19043_));
 FAx1_ASAP7_75t_R _35304_ (.SN(_19024_),
    .A(_17616_),
    .B(_17573_),
    .CI(_17617_),
    .CON(_19046_));
 FAx1_ASAP7_75t_R _35305_ (.SN(_19025_),
    .A(_17619_),
    .B(_17620_),
    .CI(_17621_),
    .CON(_19045_));
 FAx1_ASAP7_75t_R _35306_ (.SN(_17627_),
    .A(_17624_),
    .B(_17625_),
    .CI(_17626_),
    .CON(_17680_));
 FAx1_ASAP7_75t_R _35307_ (.SN(_19028_),
    .A(_17623_),
    .B(_17580_),
    .CI(_17627_),
    .CON(_19048_));
 FAx1_ASAP7_75t_R _35308_ (.SN(_17631_),
    .A(_17576_),
    .B(_17629_),
    .CI(_17586_),
    .CON(_17682_));
 FAx1_ASAP7_75t_R _35309_ (.SN(_17642_),
    .A(_17630_),
    .B(_17631_),
    .CI(_17632_),
    .CON(_17686_));
 FAx1_ASAP7_75t_R _35310_ (.SN(_19030_),
    .A(_17633_),
    .B(_17634_),
    .CI(_17635_),
    .CON(_19050_));
 FAx1_ASAP7_75t_R _35311_ (.SN(_19032_),
    .A(_17638_),
    .B(_17637_),
    .CI(_17595_),
    .CON(_19052_));
 FAx1_ASAP7_75t_R _35312_ (.SN(_17643_),
    .A(_17639_),
    .B(_17640_),
    .CI(_17641_),
    .CON(_17689_));
 FAx1_ASAP7_75t_R _35313_ (.SN(_19035_),
    .A(_17642_),
    .B(_17643_),
    .CI(_17644_),
    .CON(_19054_));
 FAx1_ASAP7_75t_R _35314_ (.SN(_19037_),
    .A(_17604_),
    .B(_17647_),
    .CI(_17646_),
    .CON(_19056_));
 FAx1_ASAP7_75t_R _35315_ (.SN(_00218_),
    .A(_17648_),
    .B(_17649_),
    .CI(_17650_),
    .CON(_17706_));
 FAx1_ASAP7_75t_R _35316_ (.SN(_19041_),
    .A(_17652_),
    .B(_17653_),
    .CI(_17654_),
    .CON(_19058_));
 FAx1_ASAP7_75t_R _35317_ (.SN(_17660_),
    .A(_17656_),
    .B(_17615_),
    .CI(_17611_),
    .CON(_19061_));
 FAx1_ASAP7_75t_R _35318_ (.SN(_00220_),
    .A(_17658_),
    .B(_17659_),
    .CI(_17660_),
    .CON(_17723_));
 FAx1_ASAP7_75t_R _35319_ (.SN(_19044_),
    .A(_17662_),
    .B(_17663_),
    .CI(_17664_),
    .CON(_19059_));
 FAx1_ASAP7_75t_R _35320_ (.SN(_17670_),
    .A(_17667_),
    .B(_17668_),
    .CI(_17669_),
    .CON(_17730_));
 FAx1_ASAP7_75t_R _35321_ (.SN(_19047_),
    .A(_17670_),
    .B(_17666_),
    .CI(_17622_),
    .CON(_19063_));
 FAx1_ASAP7_75t_R _35322_ (.SN(_17673_),
    .A(_17618_),
    .B(_17672_),
    .CI(_17628_),
    .CON(_17737_));
 FAx1_ASAP7_75t_R _35323_ (.SN(_17684_),
    .A(_17661_),
    .B(_17673_),
    .CI(_17674_),
    .CON(_17738_));
 FAx1_ASAP7_75t_R _35324_ (.SN(_19049_),
    .A(_17675_),
    .B(_17676_),
    .CI(_17677_),
    .CON(_19066_));
 FAx1_ASAP7_75t_R _35325_ (.SN(_19051_),
    .A(_17680_),
    .B(_17679_),
    .CI(_17636_),
    .CON(_17734_));
 FAx1_ASAP7_75t_R _35326_ (.SN(_17685_),
    .A(_17681_),
    .B(_17682_),
    .CI(_17683_),
    .CON(_17742_));
 FAx1_ASAP7_75t_R _35327_ (.SN(_19053_),
    .A(_17684_),
    .B(_17685_),
    .CI(_17686_),
    .CON(_19067_));
 FAx1_ASAP7_75t_R _35328_ (.SN(_19055_),
    .A(_17688_),
    .B(_17645_),
    .CI(_17689_),
    .CON(_19069_));
 FAx1_ASAP7_75t_R _35329_ (.SN(_17699_),
    .A(_17690_),
    .B(_17691_),
    .CI(_17692_),
    .CON(_19072_));
 FAx1_ASAP7_75t_R _35330_ (.SN(_00224_),
    .A(_17694_),
    .B(_17695_),
    .CI(_17696_),
    .CON(_17759_));
 FAx1_ASAP7_75t_R _35331_ (.SN(_00225_),
    .A(_17697_),
    .B(_17698_),
    .CI(_17699_),
    .CON(_17762_));
 FAx1_ASAP7_75t_R _35332_ (.SN(_19057_),
    .A(_17701_),
    .B(_17702_),
    .CI(_17703_),
    .CON(_19075_));
 FAx1_ASAP7_75t_R _35333_ (.SN(_17708_),
    .A(_17705_),
    .B(_17655_),
    .CI(_17706_),
    .CON(_19080_));
 FAx1_ASAP7_75t_R _35334_ (.SN(_17724_),
    .A(_17708_),
    .B(_17709_),
    .CI(_17700_),
    .CON(_17777_));
 FAx1_ASAP7_75t_R _35335_ (.SN(_19060_),
    .A(_17710_),
    .B(_17711_),
    .CI(_17712_),
    .CON(_19079_));
 FAx1_ASAP7_75t_R _35336_ (.SN(_17718_),
    .A(_17715_),
    .B(_17716_),
    .CI(_17717_),
    .CON(_17782_));
 FAx1_ASAP7_75t_R _35337_ (.SN(_19062_),
    .A(_17665_),
    .B(_17718_),
    .CI(_17714_),
    .CON(_19082_));
 FAx1_ASAP7_75t_R _35338_ (.SN(_19064_),
    .A(_17657_),
    .B(_17720_),
    .CI(_17671_),
    .CON(_18324_));
 FAx1_ASAP7_75t_R _35339_ (.SN(_19065_),
    .A(_17723_),
    .B(_17722_),
    .CI(_17724_),
    .CON(_18321_));
 FAx1_ASAP7_75t_R _35340_ (.SN(_17731_),
    .A(_17728_),
    .B(_17727_),
    .CI(_17729_),
    .CON(_17784_));
 FAx1_ASAP7_75t_R _35341_ (.SN(_17733_),
    .A(_17730_),
    .B(_17731_),
    .CI(_17678_),
    .CON(_18323_));
 FAx1_ASAP7_75t_R _35342_ (.SN(_00226_),
    .A(_17733_),
    .B(_17732_),
    .CI(_17734_),
    .CON(_17786_));
 FAx1_ASAP7_75t_R _35343_ (.SN(_17739_),
    .A(_17735_),
    .B(_17737_),
    .CI(_17736_),
    .CON(_17791_));
 FAx1_ASAP7_75t_R _35344_ (.SN(_19068_),
    .A(_17738_),
    .B(_17726_),
    .CI(_17739_),
    .CON(_18327_));
 FAx1_ASAP7_75t_R _35345_ (.SN(_19070_),
    .A(_17741_),
    .B(_17742_),
    .CI(_17687_),
    .CON(_18329_));
 FAx1_ASAP7_75t_R _35346_ (.SN(_19071_),
    .A(_17743_),
    .B(_17744_),
    .CI(_17745_),
    .CON(_18331_));
 FAx1_ASAP7_75t_R _35347_ (.SN(_17751_),
    .A(_17748_),
    .B(_17749_),
    .CI(_17750_),
    .CON(_17808_));
 FAx1_ASAP7_75t_R _35348_ (.SN(_19073_),
    .A(_17747_),
    .B(_17693_),
    .CI(_17751_),
    .CON(_18333_));
 FAx1_ASAP7_75t_R _35349_ (.SN(_19074_),
    .A(_17754_),
    .B(_17755_),
    .CI(_17756_),
    .CON(_18335_));
 FAx1_ASAP7_75t_R _35350_ (.SN(_19076_),
    .A(_17758_),
    .B(_17704_),
    .CI(_17759_),
    .CON(_18342_));
 FAx1_ASAP7_75t_R _35351_ (.SN(_19077_),
    .A(_17761_),
    .B(_17753_),
    .CI(_17762_),
    .CON(_18338_));
 FAx1_ASAP7_75t_R _35352_ (.SN(_19078_),
    .A(_17765_),
    .B(_17766_),
    .CI(_17767_),
    .CON(_18340_));
 FAx1_ASAP7_75t_R _35353_ (.SN(_17773_),
    .A(_17770_),
    .B(_17771_),
    .CI(_17772_),
    .CON(_17828_));
 FAx1_ASAP7_75t_R _35354_ (.SN(_19081_),
    .A(_17769_),
    .B(_17713_),
    .CI(_17773_),
    .CON(_18343_));
 FAx1_ASAP7_75t_R _35355_ (.SN(_19083_),
    .A(_17707_),
    .B(_17775_),
    .CI(_17719_),
    .CON(_17832_));
 FAx1_ASAP7_75t_R _35356_ (.SN(_18320_),
    .A(_17764_),
    .B(_17777_),
    .CI(_17776_),
    .CON(_18346_));
 FAx1_ASAP7_75t_R _35357_ (.SN(_17783_),
    .A(_17780_),
    .B(_17727_),
    .CI(_17781_),
    .CON(_17830_));
 FAx1_ASAP7_75t_R _35358_ (.SN(_18322_),
    .A(_17782_),
    .B(_17783_),
    .CI(_17784_),
    .CON(_18348_));
 FAx1_ASAP7_75t_R _35359_ (.SN(_18325_),
    .A(_17721_),
    .B(_17785_),
    .CI(_17786_),
    .CON(_18351_));
 FAx1_ASAP7_75t_R _35360_ (.SN(_18326_),
    .A(_17779_),
    .B(_17725_),
    .CI(_17788_),
    .CON(_18350_));
 FAx1_ASAP7_75t_R _35361_ (.SN(_18328_),
    .A(_17790_),
    .B(_17740_),
    .CI(_17791_),
    .CON(_18353_));
 FAx1_ASAP7_75t_R _35362_ (.SN(_18330_),
    .A(_17792_),
    .B(_17793_),
    .CI(_17794_),
    .CON(_18355_));
 FAx1_ASAP7_75t_R _35363_ (.SN(_17800_),
    .A(_17797_),
    .B(_17798_),
    .CI(_17799_),
    .CON(_17853_));
 FAx1_ASAP7_75t_R _35364_ (.SN(_18332_),
    .A(_17800_),
    .B(_17796_),
    .CI(_17746_),
    .CON(_18357_));
 FAx1_ASAP7_75t_R _35365_ (.SN(_18334_),
    .A(_17803_),
    .B(_17804_),
    .CI(_17805_),
    .CON(_18359_));
 FAx1_ASAP7_75t_R _35366_ (.SN(_18336_),
    .A(_17807_),
    .B(_17757_),
    .CI(_17808_),
    .CON(_18367_));
 FAx1_ASAP7_75t_R _35367_ (.SN(_18337_),
    .A(_17802_),
    .B(_17752_),
    .CI(_17810_),
    .CON(_18362_));
 FAx1_ASAP7_75t_R _35368_ (.SN(_18339_),
    .A(_17813_),
    .B(_17814_),
    .CI(_17815_),
    .CON(_18364_));
 FAx1_ASAP7_75t_R _35369_ (.SN(_17821_),
    .A(_17818_),
    .B(_17819_),
    .CI(_17820_),
    .CON(_17875_));
 FAx1_ASAP7_75t_R _35370_ (.SN(_18341_),
    .A(_17821_),
    .B(_17817_),
    .CI(_17768_),
    .CON(_18368_));
 FAx1_ASAP7_75t_R _35371_ (.SN(_18344_),
    .A(_17823_),
    .B(_17774_),
    .CI(_17760_),
    .CON(_17877_));
 FAx1_ASAP7_75t_R _35372_ (.SN(_18345_),
    .A(_17812_),
    .B(_17763_),
    .CI(_17824_),
    .CON(_18370_));
 FAx1_ASAP7_75t_R _35373_ (.SN(_17829_),
    .A(_17780_),
    .B(_17827_),
    .CI(_17727_),
    .CON(_17876_));
 FAx1_ASAP7_75t_R _35374_ (.SN(_18347_),
    .A(_17828_),
    .B(_17829_),
    .CI(_17830_),
    .CON(_18373_));
 FAx1_ASAP7_75t_R _35375_ (.SN(_17834_),
    .A(_17831_),
    .B(_17832_),
    .CI(_17833_),
    .CON(_17883_));
 FAx1_ASAP7_75t_R _35376_ (.SN(_18349_),
    .A(_17826_),
    .B(_17834_),
    .CI(_17778_),
    .CON(_18374_));
 FAx1_ASAP7_75t_R _35377_ (.SN(_18352_),
    .A(_17836_),
    .B(_17789_),
    .CI(_17787_),
    .CON(_18376_));
 FAx1_ASAP7_75t_R _35378_ (.SN(_18354_),
    .A(_17837_),
    .B(_17838_),
    .CI(_17839_),
    .CON(_18379_));
 FAx1_ASAP7_75t_R _35379_ (.SN(_17845_),
    .A(_17842_),
    .B(_17843_),
    .CI(_17844_),
    .CON(_17900_));
 FAx1_ASAP7_75t_R _35380_ (.SN(_18356_),
    .A(_17845_),
    .B(_17841_),
    .CI(_17795_),
    .CON(_18381_));
 FAx1_ASAP7_75t_R _35381_ (.SN(_18358_),
    .A(_17848_),
    .B(_17849_),
    .CI(_17850_),
    .CON(_18383_));
 FAx1_ASAP7_75t_R _35382_ (.SN(_18360_),
    .A(_17852_),
    .B(_17806_),
    .CI(_17853_),
    .CON(_18390_));
 FAx1_ASAP7_75t_R _35383_ (.SN(_18361_),
    .A(_17847_),
    .B(_17801_),
    .CI(_17855_),
    .CON(_18386_));
 FAx1_ASAP7_75t_R _35384_ (.SN(_18363_),
    .A(_17858_),
    .B(_17859_),
    .CI(_17860_),
    .CON(_18388_));
 FAx1_ASAP7_75t_R _35385_ (.SN(_18365_),
    .A(_17863_),
    .B(_17864_),
    .CI(_17865_),
    .CON(_18395_));
 FAx1_ASAP7_75t_R _35386_ (.SN(_18366_),
    .A(_17862_),
    .B(_17867_),
    .CI(_17816_),
    .CON(_18391_));
 FAx1_ASAP7_75t_R _35387_ (.SN(_18369_),
    .A(_17869_),
    .B(_17822_),
    .CI(_17809_),
    .CON(_17925_));
 FAx1_ASAP7_75t_R _35388_ (.SN(_18371_),
    .A(_17870_),
    .B(_17857_),
    .CI(_17811_),
    .CON(_18394_));
 FAx1_ASAP7_75t_R _35389_ (.SN(_17874_),
    .A(_17780_),
    .B(_17727_),
    .CI(_17873_),
    .CON(_17921_));
 FAx1_ASAP7_75t_R _35390_ (.SN(_18372_),
    .A(_17874_),
    .B(_17875_),
    .CI(_17876_),
    .CON(_18397_));
 FAx1_ASAP7_75t_R _35391_ (.SN(_17880_),
    .A(_17877_),
    .B(_17878_),
    .CI(_17879_),
    .CON(_17929_));
 FAx1_ASAP7_75t_R _35392_ (.SN(_18375_),
    .A(_17825_),
    .B(_17880_),
    .CI(_17872_),
    .CON(_18399_));
 FAx1_ASAP7_75t_R _35393_ (.SN(_18377_),
    .A(_17835_),
    .B(_17883_),
    .CI(_17882_),
    .CON(_18401_));
 FAx1_ASAP7_75t_R _35394_ (.SN(_18378_),
    .A(_17884_),
    .B(_17885_),
    .CI(_17886_),
    .CON(_18402_));
 FAx1_ASAP7_75t_R _35395_ (.SN(_17892_),
    .A(_17889_),
    .B(_17890_),
    .CI(_17891_),
    .CON(_17946_));
 FAx1_ASAP7_75t_R _35396_ (.SN(_18380_),
    .A(_17888_),
    .B(_17840_),
    .CI(_17892_),
    .CON(_18405_));
 FAx1_ASAP7_75t_R _35397_ (.SN(_18382_),
    .A(_17895_),
    .B(_17896_),
    .CI(_17897_),
    .CON(_18407_));
 FAx1_ASAP7_75t_R _35398_ (.SN(_18384_),
    .A(_17899_),
    .B(_17851_),
    .CI(_17900_),
    .CON(_18413_));
 FAx1_ASAP7_75t_R _35399_ (.SN(_18385_),
    .A(_17902_),
    .B(_17894_),
    .CI(_17846_),
    .CON(_18409_));
 FAx1_ASAP7_75t_R _35400_ (.SN(_18387_),
    .A(_17905_),
    .B(_17906_),
    .CI(_17907_),
    .CON(_18411_));
 FAx1_ASAP7_75t_R _35401_ (.SN(_17914_),
    .A(_17911_),
    .B(_17910_),
    .CI(_17820_),
    .CON(_17962_));
 FAx1_ASAP7_75t_R _35402_ (.SN(_18389_),
    .A(_17909_),
    .B(_17861_),
    .CI(net1999),
    .CON(_18415_));
 FAx1_ASAP7_75t_R _35403_ (.SN(_18392_),
    .A(_17916_),
    .B(_17868_),
    .CI(_17854_),
    .CON(_17965_));
 FAx1_ASAP7_75t_R _35404_ (.SN(_18393_),
    .A(_17904_),
    .B(_17856_),
    .CI(_17917_),
    .CON(_18418_));
 FAx1_ASAP7_75t_R _35405_ (.SN(_17922_),
    .A(_17780_),
    .B(_17920_),
    .CI(_17727_),
    .CON(_17963_));
 FAx1_ASAP7_75t_R _35406_ (.SN(_18396_),
    .A(_17866_),
    .B(_17921_),
    .CI(_17922_),
    .CON(_18420_));
 FAx1_ASAP7_75t_R _35407_ (.SN(_17926_),
    .A(_17923_),
    .B(_17924_),
    .CI(_17925_),
    .CON(_17970_));
 FAx1_ASAP7_75t_R _35408_ (.SN(_18398_),
    .A(_17919_),
    .B(_17871_),
    .CI(_17926_),
    .CON(_18422_));
 FAx1_ASAP7_75t_R _35409_ (.SN(_18400_),
    .A(_17928_),
    .B(_17881_),
    .CI(_17929_),
    .CON(_18424_));
 FAx1_ASAP7_75t_R _35410_ (.SN(_18403_),
    .A(_17930_),
    .B(_17931_),
    .CI(_17932_),
    .CON(_18426_));
 FAx1_ASAP7_75t_R _35411_ (.SN(_17938_),
    .A(_17935_),
    .B(_17936_),
    .CI(_17937_),
    .CON(_17987_));
 FAx1_ASAP7_75t_R _35412_ (.SN(_18404_),
    .A(_17887_),
    .B(_17938_),
    .CI(_17934_),
    .CON(_18428_));
 FAx1_ASAP7_75t_R _35413_ (.SN(_18406_),
    .A(_17941_),
    .B(_17942_),
    .CI(_17943_),
    .CON(_18430_));
 FAx1_ASAP7_75t_R _35414_ (.SN(_18408_),
    .A(_17945_),
    .B(_17898_),
    .CI(_17946_),
    .CON(_18434_));
 FAx1_ASAP7_75t_R _35415_ (.SN(_18410_),
    .A(_17948_),
    .B(_17940_),
    .CI(_17893_),
    .CON(_18433_));
 FAx1_ASAP7_75t_R _35416_ (.SN(_18412_),
    .A(_17951_),
    .B(_17952_),
    .CI(_17953_),
    .CON(_17996_));
 FAx1_ASAP7_75t_R _35417_ (.SN(_18414_),
    .A(_17908_),
    .B(net1999),
    .CI(_17954_),
    .CON(_18435_));
 FAx1_ASAP7_75t_R _35418_ (.SN(_18416_),
    .A(_17901_),
    .B(_17956_),
    .CI(_17915_),
    .CON(_18004_));
 FAx1_ASAP7_75t_R _35419_ (.SN(_18417_),
    .A(_17903_),
    .B(_17957_),
    .CI(_17950_),
    .CON(_18437_));
 FAx1_ASAP7_75t_R _35420_ (.SN(_17961_),
    .A(_17780_),
    .B(_17727_),
    .CI(_17960_),
    .CON(_18002_));
 FAx1_ASAP7_75t_R _35421_ (.SN(_18419_),
    .A(_17961_),
    .B(net1969),
    .CI(_17963_),
    .CON(_18440_));
 FAx1_ASAP7_75t_R _35422_ (.SN(_17967_),
    .A(_17964_),
    .B(_17965_),
    .CI(_17966_),
    .CON(_18010_));
 FAx1_ASAP7_75t_R _35423_ (.SN(_18421_),
    .A(_17959_),
    .B(_17918_),
    .CI(_17967_),
    .CON(_18442_));
 FAx1_ASAP7_75t_R _35424_ (.SN(_18423_),
    .A(_17969_),
    .B(_17927_),
    .CI(_17970_),
    .CON(_18444_));
 FAx1_ASAP7_75t_R _35425_ (.SN(_18425_),
    .A(_17971_),
    .B(_17972_),
    .CI(_17973_),
    .CON(_18446_));
 FAx1_ASAP7_75t_R _35426_ (.SN(_17979_),
    .A(_17976_),
    .B(_17977_),
    .CI(_17978_),
    .CON(_18028_));
 FAx1_ASAP7_75t_R _35427_ (.SN(_18427_),
    .A(_17979_),
    .B(_17975_),
    .CI(_17933_),
    .CON(_18449_));
 FAx1_ASAP7_75t_R _35428_ (.SN(_18429_),
    .A(_17982_),
    .B(_17983_),
    .CI(_17984_),
    .CON(_18451_));
 FAx1_ASAP7_75t_R _35429_ (.SN(_18431_),
    .A(_17986_),
    .B(_17944_),
    .CI(_17987_),
    .CON(_18456_));
 FAx1_ASAP7_75t_R _35430_ (.SN(_18432_),
    .A(_17981_),
    .B(_17939_),
    .CI(_17989_),
    .CON(_18454_));
 FAx1_ASAP7_75t_R _35431_ (.SN(_17995_),
    .A(_17951_),
    .B(_17992_),
    .CI(_17993_),
    .CON(_18041_));
 FAx1_ASAP7_75t_R _35432_ (.SN(_17997_),
    .A(_17913_),
    .B(_17995_),
    .CI(_17996_),
    .CON(_18042_));
 FAx1_ASAP7_75t_R _35433_ (.SN(_18436_),
    .A(_17997_),
    .B(_17955_),
    .CI(_17947_),
    .CON(_18050_));
 FAx1_ASAP7_75t_R _35434_ (.SN(_18438_),
    .A(_17998_),
    .B(_17991_),
    .CI(_17949_),
    .CON(_18459_));
 FAx1_ASAP7_75t_R _35435_ (.SN(_18003_),
    .A(_17780_),
    .B(_18001_),
    .CI(_17727_),
    .CON(_18048_));
 FAx1_ASAP7_75t_R _35436_ (.SN(_18439_),
    .A(_18002_),
    .B(net1969),
    .CI(_18003_),
    .CON(_18461_));
 FAx1_ASAP7_75t_R _35437_ (.SN(_18007_),
    .A(_18004_),
    .B(_18005_),
    .CI(_18006_),
    .CON(_18055_));
 FAx1_ASAP7_75t_R _35438_ (.SN(_18441_),
    .A(_17958_),
    .B(_18000_),
    .CI(_18007_),
    .CON(_18463_));
 FAx1_ASAP7_75t_R _35439_ (.SN(_18443_),
    .A(_18009_),
    .B(_17968_),
    .CI(_18010_),
    .CON(_18465_));
 FAx1_ASAP7_75t_R _35440_ (.SN(_18445_),
    .A(_18011_),
    .B(_18012_),
    .CI(_18013_),
    .CON(_18466_));
 FAx1_ASAP7_75t_R _35441_ (.SN(_18447_),
    .A(_18016_),
    .B(_18017_),
    .CI(_18018_),
    .CON(_18472_));
 FAx1_ASAP7_75t_R _35442_ (.SN(_18448_),
    .A(_18015_),
    .B(_17974_),
    .CI(_18020_),
    .CON(_18470_));
 FAx1_ASAP7_75t_R _35443_ (.SN(_18450_),
    .A(_18023_),
    .B(_18024_),
    .CI(_18025_),
    .CON(_18473_));
 FAx1_ASAP7_75t_R _35444_ (.SN(_18452_),
    .A(_18027_),
    .B(_17985_),
    .CI(_18028_),
    .CON(_18477_));
 FAx1_ASAP7_75t_R _35445_ (.SN(_18453_),
    .A(_18030_),
    .B(_18022_),
    .CI(_17980_),
    .CON(_18475_));
 FAx1_ASAP7_75t_R _35446_ (.SN(_18038_),
    .A(_18033_),
    .B(_18034_),
    .CI(_18035_),
    .CON(_18079_));
 FAx1_ASAP7_75t_R _35447_ (.SN(_18455_),
    .A(net1998),
    .B(_18038_),
    .CI(_17994_),
    .CON(_18478_));
 FAx1_ASAP7_75t_R _35448_ (.SN(_18457_),
    .A(_18040_),
    .B(_18042_),
    .CI(_17988_),
    .CON(_18088_));
 FAx1_ASAP7_75t_R _35449_ (.SN(_18458_),
    .A(_18032_),
    .B(_17990_),
    .CI(_18043_),
    .CON(_18481_));
 FAx1_ASAP7_75t_R _35450_ (.SN(_18047_),
    .A(_17780_),
    .B(_17727_),
    .CI(_18046_),
    .CON(_18086_));
 FAx1_ASAP7_75t_R _35451_ (.SN(_18460_),
    .A(net1970),
    .B(_18047_),
    .CI(_18048_),
    .CON(_18483_));
 FAx1_ASAP7_75t_R _35452_ (.SN(_18052_),
    .A(_18049_),
    .B(_18050_),
    .CI(_18051_),
    .CON(_18093_));
 FAx1_ASAP7_75t_R _35453_ (.SN(_18462_),
    .A(_18045_),
    .B(_18052_),
    .CI(_17999_),
    .CON(_18485_));
 FAx1_ASAP7_75t_R _35454_ (.SN(_18464_),
    .A(_18054_),
    .B(_18008_),
    .CI(_18055_),
    .CON(_18487_));
 FAx1_ASAP7_75t_R _35455_ (.SN(_18467_),
    .A(_18056_),
    .B(_18057_),
    .CI(_18058_),
    .CON(_18489_));
 FAx1_ASAP7_75t_R _35456_ (.SN(_18468_),
    .A(_18061_),
    .B(_18062_),
    .CI(_18063_),
    .CON(_18493_));
 FAx1_ASAP7_75t_R _35457_ (.SN(_18469_),
    .A(_18014_),
    .B(_18065_),
    .CI(_18060_),
    .CON(_18492_));
 FAx1_ASAP7_75t_R _35458_ (.SN(_18471_),
    .A(_18068_),
    .B(_18069_),
    .CI(_18070_),
    .CON(_18495_));
 FAx1_ASAP7_75t_R _35459_ (.SN(_18474_),
    .A(_18072_),
    .B(_18026_),
    .CI(_18019_),
    .CON(_18499_));
 FAx1_ASAP7_75t_R _35460_ (.SN(_18476_),
    .A(_18074_),
    .B(_18067_),
    .CI(_18021_),
    .CON(_18497_));
 FAx1_ASAP7_75t_R _35461_ (.SN(_18080_),
    .A(_17913_),
    .B(_18037_),
    .CI(_18036_),
    .CON(_18114_));
 FAx1_ASAP7_75t_R _35462_ (.SN(_18479_),
    .A(net1963),
    .B(_18029_),
    .CI(_18039_),
    .CON(_18122_));
 FAx1_ASAP7_75t_R _35463_ (.SN(_18480_),
    .A(_18081_),
    .B(_18031_),
    .CI(_18076_),
    .CON(_18502_));
 FAx1_ASAP7_75t_R _35464_ (.SN(_18085_),
    .A(_17780_),
    .B(_17727_),
    .CI(_18084_),
    .CON(_18119_));
 FAx1_ASAP7_75t_R _35465_ (.SN(_18482_),
    .A(_18085_),
    .B(net1970),
    .CI(_18086_),
    .CON(_18503_));
 FAx1_ASAP7_75t_R _35466_ (.SN(_18090_),
    .A(_18087_),
    .B(_18088_),
    .CI(_18089_),
    .CON(_18127_));
 FAx1_ASAP7_75t_R _35467_ (.SN(_18484_),
    .A(_18044_),
    .B(_18090_),
    .CI(_18083_),
    .CON(_18506_));
 FAx1_ASAP7_75t_R _35468_ (.SN(_18486_),
    .A(_18053_),
    .B(_18092_),
    .CI(_18093_),
    .CON(_18508_));
 FAx1_ASAP7_75t_R _35469_ (.SN(_18488_),
    .A(_18094_),
    .B(_18095_),
    .CI(_18096_),
    .CON(_18509_));
 FAx1_ASAP7_75t_R _35470_ (.SN(_18490_),
    .A(_18099_),
    .B(_18100_),
    .CI(_18101_),
    .CON(_18514_));
 FAx1_ASAP7_75t_R _35471_ (.SN(_18491_),
    .A(_18103_),
    .B(_18098_),
    .CI(_18059_),
    .CON(_18512_));
 FAx1_ASAP7_75t_R _35472_ (.SN(_18494_),
    .A(_18106_),
    .B(_18070_),
    .CI(_18107_),
    .CON(_18515_));
 FAx1_ASAP7_75t_R _35473_ (.SN(_18496_),
    .A(_18064_),
    .B(_18109_),
    .CI(_18071_),
    .CON(_18519_));
 FAx1_ASAP7_75t_R _35474_ (.SN(_18498_),
    .A(_18105_),
    .B(_18111_),
    .CI(_18066_),
    .CON(_18517_));
 FAx1_ASAP7_75t_R _35475_ (.SN(_18500_),
    .A(_18073_),
    .B(_18114_),
    .CI(net1964),
    .CON(_18155_));
 FAx1_ASAP7_75t_R _35476_ (.SN(_18501_),
    .A(_18075_),
    .B(_18115_),
    .CI(_18113_),
    .CON(_18521_));
 FAx1_ASAP7_75t_R _35477_ (.SN(_18120_),
    .A(_17780_),
    .B(net2023),
    .CI(_18118_),
    .CON(_18153_));
 FAx1_ASAP7_75t_R _35478_ (.SN(_18504_),
    .A(_18119_),
    .B(net1971),
    .CI(_18120_),
    .CON(_18524_));
 FAx1_ASAP7_75t_R _35479_ (.SN(_18124_),
    .A(_18121_),
    .B(_18122_),
    .CI(_18123_),
    .CON(_18160_));
 FAx1_ASAP7_75t_R _35480_ (.SN(_18505_),
    .A(_18117_),
    .B(_18124_),
    .CI(_18082_),
    .CON(_18525_));
 FAx1_ASAP7_75t_R _35481_ (.SN(_18507_),
    .A(_18126_),
    .B(_18091_),
    .CI(_18127_),
    .CON(_18528_));
 FAx1_ASAP7_75t_R _35482_ (.SN(_18510_),
    .A(_18128_),
    .B(_18129_),
    .CI(_18130_),
    .CON(_18530_));
 FAx1_ASAP7_75t_R _35483_ (.SN(_18511_),
    .A(_18133_),
    .B(_18134_),
    .CI(_18135_),
    .CON(_18534_));
 FAx1_ASAP7_75t_R _35484_ (.SN(_18513_),
    .A(_18137_),
    .B(_18097_),
    .CI(_18132_),
    .CON(_18533_));
 FAx1_ASAP7_75t_R _35485_ (.SN(_18143_),
    .A(_18141_),
    .B(_18140_),
    .CI(_18142_),
    .CON(_18173_));
 FAx1_ASAP7_75t_R _35486_ (.SN(_18516_),
    .A(_18108_),
    .B(_18102_),
    .CI(net2024),
    .CON(_18538_));
 FAx1_ASAP7_75t_R _35487_ (.SN(_18518_),
    .A(_18104_),
    .B(_18139_),
    .CI(_18145_),
    .CON(_18536_));
 FAx1_ASAP7_75t_R _35488_ (.SN(_18520_),
    .A(_18110_),
    .B(net2010),
    .CI(net1965),
    .CON(_18185_));
 FAx1_ASAP7_75t_R _35489_ (.SN(_18522_),
    .A(_18112_),
    .B(_18147_),
    .CI(_18148_),
    .CON(_18540_));
 FAx1_ASAP7_75t_R _35490_ (.SN(_18152_),
    .A(_17780_),
    .B(net2023),
    .CI(_18151_),
    .CON(_18183_));
 FAx1_ASAP7_75t_R _35491_ (.SN(_18523_),
    .A(_18152_),
    .B(net1972),
    .CI(_18153_),
    .CON(_18543_));
 FAx1_ASAP7_75t_R _35492_ (.SN(_18157_),
    .A(_18154_),
    .B(_18155_),
    .CI(_18156_),
    .CON(_18190_));
 FAx1_ASAP7_75t_R _35493_ (.SN(_18526_),
    .A(_18116_),
    .B(_18150_),
    .CI(_18157_),
    .CON(_18544_));
 FAx1_ASAP7_75t_R _35494_ (.SN(_18527_),
    .A(_18125_),
    .B(_18160_),
    .CI(_18159_),
    .CON(_18547_));
 FAx1_ASAP7_75t_R _35495_ (.SN(_18529_),
    .A(_18161_),
    .B(_18162_),
    .CI(_18163_),
    .CON(_18548_));
 FAx1_ASAP7_75t_R _35496_ (.SN(_18531_),
    .A(_18166_),
    .B(_18167_),
    .CI(_18168_),
    .CON(_18553_));
 FAx1_ASAP7_75t_R _35497_ (.SN(_18532_),
    .A(_18165_),
    .B(_18170_),
    .CI(_18131_),
    .CON(_18551_));
 FAx1_ASAP7_75t_R _35498_ (.SN(_18535_),
    .A(_18136_),
    .B(_18173_),
    .CI(net2025),
    .CON(_18557_));
 FAx1_ASAP7_75t_R _35499_ (.SN(_18537_),
    .A(_18175_),
    .B(_18172_),
    .CI(_18138_),
    .CON(_18555_));
 FAx1_ASAP7_75t_R _35500_ (.SN(_18539_),
    .A(net2010),
    .B(_18144_),
    .CI(net1966),
    .CON(_18212_));
 FAx1_ASAP7_75t_R _35501_ (.SN(_18541_),
    .A(_18178_),
    .B(_18146_),
    .CI(_18177_),
    .CON(_18559_));
 FAx1_ASAP7_75t_R _35502_ (.SN(_18182_),
    .A(_17780_),
    .B(net2023),
    .CI(_18181_),
    .CON(_18210_));
 FAx1_ASAP7_75t_R _35503_ (.SN(_18542_),
    .A(_18182_),
    .B(net1972),
    .CI(_18183_),
    .CON(_18562_));
 FAx1_ASAP7_75t_R _35504_ (.SN(_18187_),
    .A(_18184_),
    .B(_18185_),
    .CI(_18186_),
    .CON(_18218_));
 FAx1_ASAP7_75t_R _35505_ (.SN(_18545_),
    .A(_18187_),
    .B(_18149_),
    .CI(_18180_),
    .CON(_18564_));
 FAx1_ASAP7_75t_R _35506_ (.SN(_18546_),
    .A(_18158_),
    .B(_18190_),
    .CI(_18189_),
    .CON(_18566_));
 FAx1_ASAP7_75t_R _35507_ (.SN(_18549_),
    .A(_18191_),
    .B(_18192_),
    .CI(_18193_),
    .CON(_18231_));
 FAx1_ASAP7_75t_R _35508_ (.SN(_18550_),
    .A(_18196_),
    .B(_18197_),
    .CI(_18168_),
    .CON(_18233_));
 FAx1_ASAP7_75t_R _35509_ (.SN(_18552_),
    .A(_18164_),
    .B(_18199_),
    .CI(_18195_),
    .CON(_18567_));
 FAx1_ASAP7_75t_R _35510_ (.SN(_18554_),
    .A(_18173_),
    .B(_18169_),
    .CI(net2026),
    .CON(_18572_));
 FAx1_ASAP7_75t_R _35511_ (.SN(_18556_),
    .A(_18203_),
    .B(_18171_),
    .CI(_18201_),
    .CON(_18570_));
 FAx1_ASAP7_75t_R _35512_ (.SN(_18558_),
    .A(net2011),
    .B(_18174_),
    .CI(net1967),
    .CON(_18243_));
 FAx1_ASAP7_75t_R _35513_ (.SN(_18560_),
    .A(_18206_),
    .B(_18176_),
    .CI(_18205_),
    .CON(_18575_));
 FAx1_ASAP7_75t_R _35514_ (.SN(_18211_),
    .A(_18209_),
    .B(_17780_),
    .CI(net2023),
    .CON(_18241_));
 FAx1_ASAP7_75t_R _35515_ (.SN(_18561_),
    .A(_18210_),
    .B(net1),
    .CI(_18211_),
    .CON(_18577_));
 FAx1_ASAP7_75t_R _35516_ (.SN(_18215_),
    .A(_18212_),
    .B(_18213_),
    .CI(_18214_),
    .CON(_18248_));
 FAx1_ASAP7_75t_R _35517_ (.SN(_18563_),
    .A(_18179_),
    .B(_18208_),
    .CI(_18215_),
    .CON(_18579_));
 FAx1_ASAP7_75t_R _35518_ (.SN(_18565_),
    .A(_18217_),
    .B(_18188_),
    .CI(_18218_),
    .CON(_18581_));
 FAx1_ASAP7_75t_R _35519_ (.SN(_18230_),
    .A(_18219_),
    .B(_18220_),
    .CI(_18221_),
    .CON(_18253_));
 FAx1_ASAP7_75t_R _35520_ (.SN(_18227_),
    .A(_18223_),
    .B(_18224_),
    .CI(_18225_),
    .CON(_18254_));
 FAx1_ASAP7_75t_R _35521_ (.SN(_18568_),
    .A(_18222_),
    .B(_18194_),
    .CI(_18227_),
    .CON(_18259_));
 FAx1_ASAP7_75t_R _35522_ (.SN(_18569_),
    .A(_18173_),
    .B(_18198_),
    .CI(net2027),
    .CON(_18261_));
 FAx1_ASAP7_75t_R _35523_ (.SN(_18571_),
    .A(_18200_),
    .B(_18232_),
    .CI(_18229_),
    .CON(_18583_));
 FAx1_ASAP7_75t_R _35524_ (.SN(_18573_),
    .A(_18202_),
    .B(net2012),
    .CI(net1968),
    .CON(_18270_));
 FAx1_ASAP7_75t_R _35525_ (.SN(_18574_),
    .A(_18204_),
    .B(_18236_),
    .CI(_18235_),
    .CON(_18585_));
 FAx1_ASAP7_75t_R _35526_ (.SN(_18240_),
    .A(_17780_),
    .B(net2023),
    .CI(_18239_),
    .CON(_18268_));
 FAx1_ASAP7_75t_R _35527_ (.SN(_18576_),
    .A(_18240_),
    .B(_18241_),
    .CI(net1),
    .CON(_18587_));
 FAx1_ASAP7_75t_R _35528_ (.SN(_18245_),
    .A(_18242_),
    .B(_18243_),
    .CI(_18244_),
    .CON(_18275_));
 FAx1_ASAP7_75t_R _35529_ (.SN(_18578_),
    .A(_18238_),
    .B(_18245_),
    .CI(_18207_),
    .CON(_18589_));
 FAx1_ASAP7_75t_R _35530_ (.SN(_18580_),
    .A(_18247_),
    .B(_18216_),
    .CI(_18248_),
    .CON(_18591_));
 FAx1_ASAP7_75t_R _35531_ (.SN(_18252_),
    .A(_18249_),
    .B(_18250_),
    .CI(_18251_),
    .CON(_18279_));
 FAx1_ASAP7_75t_R _35532_ (.SN(_18256_),
    .A(_18226_),
    .B(_18252_),
    .CI(_18253_),
    .CON(_18281_));
 FAx1_ASAP7_75t_R _35533_ (.SN(_18260_),
    .A(_18173_),
    .B(_18254_),
    .CI(net2027),
    .CON(_18283_));
 FAx1_ASAP7_75t_R _35534_ (.SN(_18582_),
    .A(_18255_),
    .B(_18256_),
    .CI(_18228_),
    .CON(_18290_));
 FAx1_ASAP7_75t_R _35535_ (.SN(_18263_),
    .A(_18078_),
    .B(_18261_),
    .CI(_18077_),
    .CON(_00272_));
 FAx1_ASAP7_75t_R _35536_ (.SN(_18584_),
    .A(_18258_),
    .B(_18234_),
    .CI(_18263_),
    .CON(_18593_));
 FAx1_ASAP7_75t_R _35537_ (.SN(_18267_),
    .A(_17780_),
    .B(net2023),
    .CI(_18266_),
    .CON(_18294_));
 FAx1_ASAP7_75t_R _35538_ (.SN(_18586_),
    .A(_18267_),
    .B(net1),
    .CI(_18268_),
    .CON(_18594_));
 FAx1_ASAP7_75t_R _35539_ (.SN(_18272_),
    .A(_18269_),
    .B(_18270_),
    .CI(_18271_),
    .CON(_18300_));
 FAx1_ASAP7_75t_R _35540_ (.SN(_18588_),
    .A(_18265_),
    .B(_18272_),
    .CI(_18237_),
    .CON(_18597_));
 FAx1_ASAP7_75t_R _35541_ (.SN(_18590_),
    .A(_18274_),
    .B(_18246_),
    .CI(_18275_),
    .CON(_18599_));
 FAx1_ASAP7_75t_R _35542_ (.SN(_18278_),
    .A(_18276_),
    .B(_18277_),
    .CI(_18251_),
    .CON(_18303_));
 FAx1_ASAP7_75t_R _35543_ (.SN(_18280_),
    .A(_18226_),
    .B(_18278_),
    .CI(_18279_),
    .CON(_18305_));
 FAx1_ASAP7_75t_R _35544_ (.SN(_18289_),
    .A(_18255_),
    .B(_18280_),
    .CI(_18281_),
    .CON(_18307_));
 FAx1_ASAP7_75t_R _35545_ (.SN(_18286_),
    .A(_18283_),
    .B(_18077_),
    .CI(_18078_),
    .CON(_00276_));
 FAx1_ASAP7_75t_R _35546_ (.SN(_18592_),
    .A(_18282_),
    .B(_18257_),
    .CI(_18286_),
    .CON(_18600_));
 FAx1_ASAP7_75t_R _35547_ (.SN(_18293_),
    .A(_18291_),
    .B(_17780_),
    .CI(net2023),
    .CON(_00278_));
 FAx1_ASAP7_75t_R _35548_ (.SN(_18595_),
    .A(_18293_),
    .B(_18294_),
    .CI(net1),
    .CON(_18601_));
 FAx1_ASAP7_75t_R _35549_ (.SN(_18297_),
    .A(_18295_),
    .B(_18262_),
    .CI(_18296_),
    .CON(_18316_));
 FAx1_ASAP7_75t_R _35550_ (.SN(_18596_),
    .A(_18288_),
    .B(_18264_),
    .CI(_18297_),
    .CON(_18603_));
 FAx1_ASAP7_75t_R _35551_ (.SN(_18598_),
    .A(_18300_),
    .B(_18299_),
    .CI(_18273_),
    .CON(_18605_));
 FAx1_ASAP7_75t_R _35552_ (.SN(_18302_),
    .A(_18276_),
    .B(_18301_),
    .CI(_18251_),
    .CON(_02230_));
 FAx1_ASAP7_75t_R _35553_ (.SN(_18304_),
    .A(_18226_),
    .B(_18302_),
    .CI(_18303_),
    .CON(_00282_));
 FAx1_ASAP7_75t_R _35554_ (.SN(_18306_),
    .A(_18255_),
    .B(_18304_),
    .CI(_18305_),
    .CON(_02231_));
 FAx1_ASAP7_75t_R _35555_ (.SN(_18313_),
    .A(_18285_),
    .B(_18306_),
    .CI(_18307_),
    .CON(_00283_));
 FAx1_ASAP7_75t_R _35556_ (.SN(_00277_),
    .A(_17780_),
    .B(net2023),
    .CI(_18308_),
    .CON(_00284_));
 FAx1_ASAP7_75t_R _35557_ (.SN(_02232_),
    .A(_18309_),
    .B(_18292_),
    .CI(_17912_),
    .CON(_00285_));
 FAx1_ASAP7_75t_R _35558_ (.SN(_18314_),
    .A(_18284_),
    .B(_18311_),
    .CI(_18312_),
    .CON(_00286_));
 FAx1_ASAP7_75t_R _35559_ (.SN(_18602_),
    .A(_18313_),
    .B(_18287_),
    .CI(_18314_),
    .CON(_02233_));
 FAx1_ASAP7_75t_R _35560_ (.SN(_18604_),
    .A(_18316_),
    .B(_18315_),
    .CI(_18298_),
    .CON(_02234_));
 FAx1_ASAP7_75t_R _35561_ (.SN(_00293_),
    .A(_18317_),
    .B(_18318_),
    .CI(_18319_),
    .CON(_00295_));
 HAxp5_ASAP7_75t_R _35562_ (.A(_17780_),
    .B(net2023),
    .CON(_17343_),
    .SN(_00229_));
 HAxp5_ASAP7_75t_R _35563_ (.A(_18322_),
    .B(_18323_),
    .CON(_02235_),
    .SN(_17785_));
 HAxp5_ASAP7_75t_R _35564_ (.A(_18328_),
    .B(_18329_),
    .CON(_00235_),
    .SN(_00230_));
 HAxp5_ASAP7_75t_R _35565_ (.A(_18347_),
    .B(_18348_),
    .CON(_02236_),
    .SN(_00233_));
 HAxp5_ASAP7_75t_R _35566_ (.A(_18352_),
    .B(_18353_),
    .CON(_00238_),
    .SN(_00234_));
 HAxp5_ASAP7_75t_R _35567_ (.A(_18372_),
    .B(_18373_),
    .CON(_02237_),
    .SN(_00236_));
 HAxp5_ASAP7_75t_R _35568_ (.A(_18376_),
    .B(_18377_),
    .CON(_00241_),
    .SN(_00237_));
 HAxp5_ASAP7_75t_R _35569_ (.A(_18396_),
    .B(_18397_),
    .CON(_02238_),
    .SN(_00239_));
 HAxp5_ASAP7_75t_R _35570_ (.A(_18400_),
    .B(_18401_),
    .CON(_00244_),
    .SN(_00240_));
 HAxp5_ASAP7_75t_R _35571_ (.A(_18419_),
    .B(_18420_),
    .CON(_02239_),
    .SN(_00242_));
 HAxp5_ASAP7_75t_R _35572_ (.A(_18423_),
    .B(_18424_),
    .CON(_00247_),
    .SN(_00243_));
 HAxp5_ASAP7_75t_R _35573_ (.A(_18439_),
    .B(_18440_),
    .CON(_02240_),
    .SN(_00245_));
 HAxp5_ASAP7_75t_R _35574_ (.A(_18443_),
    .B(_18444_),
    .CON(_00250_),
    .SN(_00246_));
 HAxp5_ASAP7_75t_R _35575_ (.A(_18460_),
    .B(_18461_),
    .CON(_02241_),
    .SN(_00248_));
 HAxp5_ASAP7_75t_R _35576_ (.A(_18464_),
    .B(_18465_),
    .CON(_00253_),
    .SN(_00249_));
 HAxp5_ASAP7_75t_R _35577_ (.A(_18482_),
    .B(_18483_),
    .CON(_02242_),
    .SN(_00251_));
 HAxp5_ASAP7_75t_R _35578_ (.A(_18487_),
    .B(_18486_),
    .CON(_00256_),
    .SN(_00252_));
 HAxp5_ASAP7_75t_R _35579_ (.A(_18503_),
    .B(_18504_),
    .CON(_02243_),
    .SN(_00254_));
 HAxp5_ASAP7_75t_R _35580_ (.A(_18507_),
    .B(_18508_),
    .CON(_00259_),
    .SN(_00255_));
 HAxp5_ASAP7_75t_R _35581_ (.A(_18523_),
    .B(_18524_),
    .CON(_02244_),
    .SN(_00257_));
 HAxp5_ASAP7_75t_R _35582_ (.A(_18527_),
    .B(_18528_),
    .CON(_00262_),
    .SN(_00258_));
 HAxp5_ASAP7_75t_R _35583_ (.A(_18542_),
    .B(_18543_),
    .CON(_02245_),
    .SN(_00260_));
 HAxp5_ASAP7_75t_R _35584_ (.A(_18546_),
    .B(_18547_),
    .CON(_00265_),
    .SN(_00261_));
 HAxp5_ASAP7_75t_R _35585_ (.A(_18561_),
    .B(_18562_),
    .CON(_02246_),
    .SN(_00263_));
 HAxp5_ASAP7_75t_R _35586_ (.A(_18565_),
    .B(_18566_),
    .CON(_00268_),
    .SN(_00264_));
 HAxp5_ASAP7_75t_R _35587_ (.A(_18576_),
    .B(_18577_),
    .CON(_02247_),
    .SN(_00266_));
 HAxp5_ASAP7_75t_R _35588_ (.A(_18580_),
    .B(_18581_),
    .CON(_00271_),
    .SN(_00267_));
 HAxp5_ASAP7_75t_R _35589_ (.A(_18586_),
    .B(_18587_),
    .CON(_02248_),
    .SN(_00269_));
 HAxp5_ASAP7_75t_R _35590_ (.A(_18590_),
    .B(_18591_),
    .CON(_00275_),
    .SN(_00270_));
 HAxp5_ASAP7_75t_R _35591_ (.A(_18594_),
    .B(_18595_),
    .CON(_02249_),
    .SN(_00273_));
 HAxp5_ASAP7_75t_R _35592_ (.A(_18598_),
    .B(_18599_),
    .CON(_00281_),
    .SN(_00274_));
 HAxp5_ASAP7_75t_R _35593_ (.A(_18310_),
    .B(_18601_),
    .CON(_02250_),
    .SN(_00279_));
 HAxp5_ASAP7_75t_R _35594_ (.A(_18604_),
    .B(_18605_),
    .CON(_00287_),
    .SN(_00280_));
 HAxp5_ASAP7_75t_R _35595_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_18606_),
    .CON(_00294_),
    .SN(_00292_));
 HAxp5_ASAP7_75t_R _35596_ (.A(_18607_),
    .B(_18608_),
    .CON(_02251_),
    .SN(_00296_));
 HAxp5_ASAP7_75t_R _35597_ (.A(_18609_),
    .B(_18610_),
    .CON(_02252_),
    .SN(_02253_));
 HAxp5_ASAP7_75t_R _35598_ (.A(_18611_),
    .B(_18608_),
    .CON(_00297_),
    .SN(_18612_));
 HAxp5_ASAP7_75t_R _35599_ (.A(_18613_),
    .B(_18614_),
    .CON(_00299_),
    .SN(_00298_));
 HAxp5_ASAP7_75t_R _35600_ (.A(_18615_),
    .B(_18607_),
    .CON(_02254_),
    .SN(_18616_));
 HAxp5_ASAP7_75t_R _35601_ (.A(_18617_),
    .B(_18618_),
    .CON(_00301_),
    .SN(_00300_));
 HAxp5_ASAP7_75t_R _35602_ (.A(_18619_),
    .B(_18620_),
    .CON(_02255_),
    .SN(_18621_));
 HAxp5_ASAP7_75t_R _35603_ (.A(_18622_),
    .B(_18623_),
    .CON(_00303_),
    .SN(_00302_));
 HAxp5_ASAP7_75t_R _35604_ (.A(_18624_),
    .B(_18625_),
    .CON(_02256_),
    .SN(_18626_));
 HAxp5_ASAP7_75t_R _35605_ (.A(_18627_),
    .B(_18628_),
    .CON(_02257_),
    .SN(_00304_));
 HAxp5_ASAP7_75t_R _35606_ (.A(_18629_),
    .B(_18630_),
    .CON(_00305_),
    .SN(_18631_));
 HAxp5_ASAP7_75t_R _35607_ (.A(_18632_),
    .B(_18633_),
    .CON(_00307_),
    .SN(_00306_));
 HAxp5_ASAP7_75t_R _35608_ (.A(_18634_),
    .B(_18635_),
    .CON(_02258_),
    .SN(_18636_));
 HAxp5_ASAP7_75t_R _35609_ (.A(_18637_),
    .B(_18638_),
    .CON(_00309_),
    .SN(_00308_));
 HAxp5_ASAP7_75t_R _35610_ (.A(_18639_),
    .B(_18640_),
    .CON(_02259_),
    .SN(_18641_));
 HAxp5_ASAP7_75t_R _35611_ (.A(_18642_),
    .B(_18643_),
    .CON(_00311_),
    .SN(_00310_));
 HAxp5_ASAP7_75t_R _35612_ (.A(_18644_),
    .B(_18645_),
    .CON(_02260_),
    .SN(_18646_));
 HAxp5_ASAP7_75t_R _35613_ (.A(_18647_),
    .B(_18648_),
    .CON(_00313_),
    .SN(_00312_));
 HAxp5_ASAP7_75t_R _35614_ (.A(_18649_),
    .B(_18650_),
    .CON(_02261_),
    .SN(_18651_));
 HAxp5_ASAP7_75t_R _35615_ (.A(_18652_),
    .B(_18653_),
    .CON(_00315_),
    .SN(_00314_));
 HAxp5_ASAP7_75t_R _35616_ (.A(_18654_),
    .B(_18655_),
    .CON(_02262_),
    .SN(_18656_));
 HAxp5_ASAP7_75t_R _35617_ (.A(_18657_),
    .B(_18658_),
    .CON(_00317_),
    .SN(_00316_));
 HAxp5_ASAP7_75t_R _35618_ (.A(_18659_),
    .B(_18660_),
    .CON(_02263_),
    .SN(_18661_));
 HAxp5_ASAP7_75t_R _35619_ (.A(_18662_),
    .B(_18663_),
    .CON(_00319_),
    .SN(_00318_));
 HAxp5_ASAP7_75t_R _35620_ (.A(_18664_),
    .B(_18665_),
    .CON(_02264_),
    .SN(_18666_));
 HAxp5_ASAP7_75t_R _35621_ (.A(_18667_),
    .B(_18668_),
    .CON(_00321_),
    .SN(_00320_));
 HAxp5_ASAP7_75t_R _35622_ (.A(_18669_),
    .B(_18670_),
    .CON(_02265_),
    .SN(_18671_));
 HAxp5_ASAP7_75t_R _35623_ (.A(_18672_),
    .B(_18673_),
    .CON(_00323_),
    .SN(_00322_));
 HAxp5_ASAP7_75t_R _35624_ (.A(_18674_),
    .B(_18675_),
    .CON(_02266_),
    .SN(_18676_));
 HAxp5_ASAP7_75t_R _35625_ (.A(_18677_),
    .B(_18678_),
    .CON(_02267_),
    .SN(_00324_));
 HAxp5_ASAP7_75t_R _35626_ (.A(_18679_),
    .B(_18680_),
    .CON(_00325_),
    .SN(_18681_));
 HAxp5_ASAP7_75t_R _35627_ (.A(_18682_),
    .B(_18683_),
    .CON(_02268_),
    .SN(_00326_));
 HAxp5_ASAP7_75t_R _35628_ (.A(_18684_),
    .B(_18685_),
    .CON(_00327_),
    .SN(_18686_));
 HAxp5_ASAP7_75t_R _35629_ (.A(_18687_),
    .B(_18688_),
    .CON(_00329_),
    .SN(_00328_));
 HAxp5_ASAP7_75t_R _35630_ (.A(_18689_),
    .B(_18690_),
    .CON(_02269_),
    .SN(_18691_));
 HAxp5_ASAP7_75t_R _35631_ (.A(_18692_),
    .B(_18693_),
    .CON(_00331_),
    .SN(_00330_));
 HAxp5_ASAP7_75t_R _35632_ (.A(_18694_),
    .B(_18695_),
    .CON(_02270_),
    .SN(_18696_));
 HAxp5_ASAP7_75t_R _35633_ (.A(_18697_),
    .B(_18698_),
    .CON(_00333_),
    .SN(_00332_));
 HAxp5_ASAP7_75t_R _35634_ (.A(_18699_),
    .B(_18700_),
    .CON(_02271_),
    .SN(_18701_));
 HAxp5_ASAP7_75t_R _35635_ (.A(_18702_),
    .B(_18703_),
    .CON(_00335_),
    .SN(_00334_));
 HAxp5_ASAP7_75t_R _35636_ (.A(_18704_),
    .B(_18705_),
    .CON(_02272_),
    .SN(_18706_));
 HAxp5_ASAP7_75t_R _35637_ (.A(_18707_),
    .B(_18708_),
    .CON(_00337_),
    .SN(_00336_));
 HAxp5_ASAP7_75t_R _35638_ (.A(_18709_),
    .B(_18710_),
    .CON(_02273_),
    .SN(_18711_));
 HAxp5_ASAP7_75t_R _35639_ (.A(_18712_),
    .B(_18713_),
    .CON(_02274_),
    .SN(_00338_));
 HAxp5_ASAP7_75t_R _35640_ (.A(_18714_),
    .B(_18715_),
    .CON(_00339_),
    .SN(_18716_));
 HAxp5_ASAP7_75t_R _35641_ (.A(_18717_),
    .B(_18718_),
    .CON(_00341_),
    .SN(_00340_));
 HAxp5_ASAP7_75t_R _35642_ (.A(_18719_),
    .B(_18720_),
    .CON(_02275_),
    .SN(_18721_));
 HAxp5_ASAP7_75t_R _35643_ (.A(_18722_),
    .B(_18723_),
    .CON(_02276_),
    .SN(_00342_));
 HAxp5_ASAP7_75t_R _35644_ (.A(_18724_),
    .B(_18725_),
    .CON(_00343_),
    .SN(_18726_));
 HAxp5_ASAP7_75t_R _35645_ (.A(_18727_),
    .B(_18728_),
    .CON(_02277_),
    .SN(_00344_));
 HAxp5_ASAP7_75t_R _35646_ (.A(_18729_),
    .B(_18730_),
    .CON(_00345_),
    .SN(_18731_));
 HAxp5_ASAP7_75t_R _35647_ (.A(_18732_),
    .B(_18733_),
    .CON(_00347_),
    .SN(_00346_));
 HAxp5_ASAP7_75t_R _35648_ (.A(_18734_),
    .B(_18735_),
    .CON(_02278_),
    .SN(_18736_));
 HAxp5_ASAP7_75t_R _35649_ (.A(_18737_),
    .B(_18738_),
    .CON(_02279_),
    .SN(_00348_));
 HAxp5_ASAP7_75t_R _35650_ (.A(_18739_),
    .B(_18740_),
    .CON(_00349_),
    .SN(_18741_));
 HAxp5_ASAP7_75t_R _35651_ (.A(_18742_),
    .B(_18743_),
    .CON(_00351_),
    .SN(_00350_));
 HAxp5_ASAP7_75t_R _35652_ (.A(_18744_),
    .B(_18745_),
    .CON(_02280_),
    .SN(_18746_));
 HAxp5_ASAP7_75t_R _35653_ (.A(_18747_),
    .B(_18748_),
    .CON(_00353_),
    .SN(_00352_));
 HAxp5_ASAP7_75t_R _35654_ (.A(_18749_),
    .B(_18750_),
    .CON(_02281_),
    .SN(_18751_));
 HAxp5_ASAP7_75t_R _35655_ (.A(_18752_),
    .B(_18753_),
    .CON(_00355_),
    .SN(_00354_));
 HAxp5_ASAP7_75t_R _35656_ (.A(_18754_),
    .B(_18755_),
    .CON(_02282_),
    .SN(_18756_));
 HAxp5_ASAP7_75t_R _35657_ (.A(_18757_),
    .B(_18758_),
    .CON(_02283_),
    .SN(_00356_));
 HAxp5_ASAP7_75t_R _35658_ (.A(_18759_),
    .B(_18760_),
    .CON(_00357_),
    .SN(_18761_));
 HAxp5_ASAP7_75t_R _35659_ (.A(_18762_),
    .B(_18763_),
    .CON(_02284_),
    .SN(_02285_));
 HAxp5_ASAP7_75t_R _35660_ (.A(\alu_adder_result_ex[1] ),
    .B(_18763_),
    .CON(_00364_),
    .SN(_02286_));
 HAxp5_ASAP7_75t_R _35661_ (.A(_18764_),
    .B(_18763_),
    .CON(_00360_),
    .SN(_18765_));
 HAxp5_ASAP7_75t_R _35662_ (.A(\alu_adder_result_ex[0] ),
    .B(\alu_adder_result_ex[1] ),
    .CON(_00361_),
    .SN(_00363_));
 HAxp5_ASAP7_75t_R _35663_ (.A(\alu_adder_result_ex[0] ),
    .B(\alu_adder_result_ex[1] ),
    .CON(_02287_),
    .SN(_18766_));
 HAxp5_ASAP7_75t_R _35664_ (.A(\alu_adder_result_ex[0] ),
    .B(_18764_),
    .CON(_00359_),
    .SN(_18767_));
 HAxp5_ASAP7_75t_R _35665_ (.A(\alu_adder_result_ex[0] ),
    .B(_18764_),
    .CON(_02288_),
    .SN(_18768_));
 HAxp5_ASAP7_75t_R _35666_ (.A(net52),
    .B(\alu_adder_result_ex[1] ),
    .CON(_00362_),
    .SN(_18770_));
 HAxp5_ASAP7_75t_R _35667_ (.A(net52),
    .B(\alu_adder_result_ex[1] ),
    .CON(_02289_),
    .SN(_18771_));
 HAxp5_ASAP7_75t_R _35668_ (.A(net52),
    .B(_18764_),
    .CON(_18762_),
    .SN(_18772_));
 HAxp5_ASAP7_75t_R _35669_ (.A(_18773_),
    .B(_18774_),
    .CON(_02290_),
    .SN(_02291_));
 HAxp5_ASAP7_75t_R _35670_ (.A(_18775_),
    .B(_18776_),
    .CON(_02292_),
    .SN(_02293_));
 HAxp5_ASAP7_75t_R _35671_ (.A(_18778_),
    .B(net2002),
    .CON(_01450_),
    .SN(_02294_));
 HAxp5_ASAP7_75t_R _35672_ (.A(net2002),
    .B(_18779_),
    .CON(_02295_),
    .SN(_18780_));
 HAxp5_ASAP7_75t_R _35673_ (.A(_18778_),
    .B(_18781_),
    .CON(_02296_),
    .SN(_18782_));
 HAxp5_ASAP7_75t_R _35674_ (.A(_18781_),
    .B(_18779_),
    .CON(_00406_),
    .SN(_18783_));
 HAxp5_ASAP7_75t_R _35675_ (.A(_18784_),
    .B(_18785_),
    .CON(_00794_),
    .SN(_00415_));
 HAxp5_ASAP7_75t_R _35676_ (.A(_17345_),
    .B(_17346_),
    .CON(_00448_),
    .SN(_02297_));
 HAxp5_ASAP7_75t_R _35677_ (.A(_18787_),
    .B(_18786_),
    .CON(_00797_),
    .SN(_00793_));
 HAxp5_ASAP7_75t_R _35678_ (.A(_18788_),
    .B(_18789_),
    .CON(_00800_),
    .SN(_00796_));
 HAxp5_ASAP7_75t_R _35679_ (.A(_18790_),
    .B(_18791_),
    .CON(_00803_),
    .SN(_00799_));
 HAxp5_ASAP7_75t_R _35680_ (.A(_18792_),
    .B(_18793_),
    .CON(_00806_),
    .SN(_00802_));
 HAxp5_ASAP7_75t_R _35681_ (.A(_18794_),
    .B(_18795_),
    .CON(_00808_),
    .SN(_00805_));
 HAxp5_ASAP7_75t_R _35682_ (.A(_18796_),
    .B(_18797_),
    .CON(_00811_),
    .SN(_02298_));
 HAxp5_ASAP7_75t_R _35683_ (.A(_18799_),
    .B(_18798_),
    .CON(_00814_),
    .SN(_00810_));
 HAxp5_ASAP7_75t_R _35684_ (.A(_18801_),
    .B(_18800_),
    .CON(_00817_),
    .SN(_00813_));
 HAxp5_ASAP7_75t_R _35685_ (.A(_18802_),
    .B(_18803_),
    .CON(_00820_),
    .SN(_00816_));
 HAxp5_ASAP7_75t_R _35686_ (.A(_18804_),
    .B(_18805_),
    .CON(_00823_),
    .SN(_00819_));
 HAxp5_ASAP7_75t_R _35687_ (.A(_18807_),
    .B(_18806_),
    .CON(_00856_),
    .SN(_00822_));
 HAxp5_ASAP7_75t_R _35688_ (.A(_18809_),
    .B(_18808_),
    .CON(_00889_),
    .SN(_00855_));
 HAxp5_ASAP7_75t_R _35689_ (.A(_18810_),
    .B(_18811_),
    .CON(_00922_),
    .SN(_00888_));
 HAxp5_ASAP7_75t_R _35690_ (.A(_18813_),
    .B(_18812_),
    .CON(_00955_),
    .SN(_00921_));
 HAxp5_ASAP7_75t_R _35691_ (.A(_18814_),
    .B(_18815_),
    .CON(_00988_),
    .SN(_00954_));
 HAxp5_ASAP7_75t_R _35692_ (.A(_18816_),
    .B(_18817_),
    .CON(_01021_),
    .SN(_00987_));
 HAxp5_ASAP7_75t_R _35693_ (.A(_18818_),
    .B(_18819_),
    .CON(_01054_),
    .SN(_01020_));
 HAxp5_ASAP7_75t_R _35694_ (.A(_18820_),
    .B(_18821_),
    .CON(_01087_),
    .SN(_01053_));
 HAxp5_ASAP7_75t_R _35695_ (.A(_18822_),
    .B(_18823_),
    .CON(_01120_),
    .SN(_01086_));
 HAxp5_ASAP7_75t_R _35696_ (.A(_18824_),
    .B(_18825_),
    .CON(_01153_),
    .SN(_01119_));
 HAxp5_ASAP7_75t_R _35697_ (.A(_18826_),
    .B(_18827_),
    .CON(_01186_),
    .SN(_01152_));
 HAxp5_ASAP7_75t_R _35698_ (.A(_18828_),
    .B(_18829_),
    .CON(_01219_),
    .SN(_01185_));
 HAxp5_ASAP7_75t_R _35699_ (.A(_18830_),
    .B(_18831_),
    .CON(_01252_),
    .SN(_01218_));
 HAxp5_ASAP7_75t_R _35700_ (.A(_18832_),
    .B(_18833_),
    .CON(_01285_),
    .SN(_01251_));
 HAxp5_ASAP7_75t_R _35701_ (.A(_18834_),
    .B(_18835_),
    .CON(_01318_),
    .SN(_01284_));
 HAxp5_ASAP7_75t_R _35702_ (.A(_18836_),
    .B(_18837_),
    .CON(_01351_),
    .SN(_01317_));
 HAxp5_ASAP7_75t_R _35703_ (.A(_18838_),
    .B(_18839_),
    .CON(_01384_),
    .SN(_01350_));
 HAxp5_ASAP7_75t_R _35704_ (.A(_18840_),
    .B(_18841_),
    .CON(_01417_),
    .SN(_01383_));
 HAxp5_ASAP7_75t_R _35705_ (.A(_18842_),
    .B(_18843_),
    .CON(_01449_),
    .SN(_01416_));
 HAxp5_ASAP7_75t_R _35706_ (.A(_18844_),
    .B(_18845_),
    .CON(_02299_),
    .SN(_01451_));
 HAxp5_ASAP7_75t_R _35707_ (.A(_18846_),
    .B(_18847_),
    .CON(_00358_),
    .SN(_18848_));
 HAxp5_ASAP7_75t_R _35708_ (.A(_18849_),
    .B(_18850_),
    .CON(_02300_),
    .SN(_02301_));
 HAxp5_ASAP7_75t_R _35709_ (.A(_18851_),
    .B(\cs_registers_i.priv_lvl_q[0] ),
    .CON(_02302_),
    .SN(_01452_));
 HAxp5_ASAP7_75t_R _35710_ (.A(_18852_),
    .B(_18853_),
    .CON(_02303_),
    .SN(_02304_));
 HAxp5_ASAP7_75t_R _35711_ (.A(_18854_),
    .B(_18855_),
    .CON(_00571_),
    .SN(_02305_));
 HAxp5_ASAP7_75t_R _35712_ (.A(_18854_),
    .B(_18856_),
    .CON(_02306_),
    .SN(_18857_));
 HAxp5_ASAP7_75t_R _35713_ (.A(_18858_),
    .B(_18855_),
    .CON(_00572_),
    .SN(_18859_));
 HAxp5_ASAP7_75t_R _35714_ (.A(_18858_),
    .B(_18856_),
    .CON(_00479_),
    .SN(_18860_));
 HAxp5_ASAP7_75t_R _35715_ (.A(_18861_),
    .B(_18862_),
    .CON(_02307_),
    .SN(_02308_));
 HAxp5_ASAP7_75t_R _35716_ (.A(_18861_),
    .B(_18863_),
    .CON(_02309_),
    .SN(_18864_));
 HAxp5_ASAP7_75t_R _35717_ (.A(_18865_),
    .B(_18862_),
    .CON(_02310_),
    .SN(_18866_));
 HAxp5_ASAP7_75t_R _35718_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(\cs_registers_i.mhpmcounter[2][1] ),
    .CON(_02311_),
    .SN(_02312_));
 HAxp5_ASAP7_75t_R _35719_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .CON(_02313_),
    .SN(_02314_));
 HAxp5_ASAP7_75t_R _35720_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CON(_02315_),
    .SN(_00017_));
 HAxp5_ASAP7_75t_R _35721_ (.A(_18867_),
    .B(_18868_),
    .CON(_00068_),
    .SN(_02316_));
 HAxp5_ASAP7_75t_R _35722_ (.A(_18867_),
    .B(_18868_),
    .CON(_02317_),
    .SN(_18869_));
 HAxp5_ASAP7_75t_R _35723_ (.A(_18867_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_00074_),
    .SN(_18870_));
 HAxp5_ASAP7_75t_R _35724_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_18868_),
    .CON(_01458_),
    .SN(_18871_));
 HAxp5_ASAP7_75t_R _35725_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_00067_),
    .SN(_18872_));
 HAxp5_ASAP7_75t_R _35726_ (.A(_18873_),
    .B(_18874_),
    .CON(_02318_),
    .SN(_00104_));
 HAxp5_ASAP7_75t_R _35727_ (.A(_18876_),
    .B(_18875_),
    .CON(_02319_),
    .SN(_00137_));
 HAxp5_ASAP7_75t_R _35728_ (.A(_18878_),
    .B(_18879_),
    .CON(_02320_),
    .SN(_00138_));
 HAxp5_ASAP7_75t_R _35729_ (.A(_18881_),
    .B(_18877_),
    .CON(_02321_),
    .SN(_00139_));
 HAxp5_ASAP7_75t_R _35730_ (.A(_18883_),
    .B(_18884_),
    .CON(_02322_),
    .SN(_00140_));
 HAxp5_ASAP7_75t_R _35731_ (.A(_18886_),
    .B(_18887_),
    .CON(_02323_),
    .SN(_00141_));
 HAxp5_ASAP7_75t_R _35732_ (.A(_18889_),
    .B(_18890_),
    .CON(_02324_),
    .SN(_00142_));
 HAxp5_ASAP7_75t_R _35733_ (.A(_18880_),
    .B(_18892_),
    .CON(_02325_),
    .SN(_00143_));
 HAxp5_ASAP7_75t_R _35734_ (.A(_18894_),
    .B(_18882_),
    .CON(_17371_),
    .SN(_00144_));
 HAxp5_ASAP7_75t_R _35735_ (.A(_18895_),
    .B(_18888_),
    .CON(_17369_),
    .SN(_00145_));
 HAxp5_ASAP7_75t_R _35736_ (.A(_18896_),
    .B(_18885_),
    .CON(_02326_),
    .SN(_00146_));
 HAxp5_ASAP7_75t_R _35737_ (.A(_17368_),
    .B(_18891_),
    .CON(_02327_),
    .SN(_00149_));
 HAxp5_ASAP7_75t_R _35738_ (.A(_18893_),
    .B(_18899_),
    .CON(_17383_),
    .SN(_00150_));
 HAxp5_ASAP7_75t_R _35739_ (.A(_17359_),
    .B(_18900_),
    .CON(_17384_),
    .SN(_17370_));
 HAxp5_ASAP7_75t_R _35740_ (.A(_18901_),
    .B(_18897_),
    .CON(_02328_),
    .SN(_00151_));
 HAxp5_ASAP7_75t_R _35741_ (.A(_17375_),
    .B(_18902_),
    .CON(_02329_),
    .SN(_00153_));
 HAxp5_ASAP7_75t_R _35742_ (.A(_17367_),
    .B(_18907_),
    .CON(_02330_),
    .SN(_00155_));
 HAxp5_ASAP7_75t_R _35743_ (.A(_18909_),
    .B(_18898_),
    .CON(_17400_),
    .SN(_00156_));
 HAxp5_ASAP7_75t_R _35744_ (.A(_18910_),
    .B(_18904_),
    .CON(_17398_),
    .SN(_17382_));
 HAxp5_ASAP7_75t_R _35745_ (.A(_17386_),
    .B(_17387_),
    .CON(_00166_),
    .SN(_00157_));
 HAxp5_ASAP7_75t_R _35746_ (.A(_18911_),
    .B(_18912_),
    .CON(_02331_),
    .SN(_00159_));
 HAxp5_ASAP7_75t_R _35747_ (.A(_18913_),
    .B(_17391_),
    .CON(_02332_),
    .SN(_00161_));
 HAxp5_ASAP7_75t_R _35748_ (.A(_18915_),
    .B(_18903_),
    .CON(_17420_),
    .SN(_00162_));
 HAxp5_ASAP7_75t_R _35749_ (.A(_18919_),
    .B(_18920_),
    .CON(_17421_),
    .SN(_00163_));
 HAxp5_ASAP7_75t_R _35750_ (.A(_18908_),
    .B(_18921_),
    .CON(_17423_),
    .SN(_00164_));
 HAxp5_ASAP7_75t_R _35751_ (.A(_18922_),
    .B(_18916_),
    .CON(_17424_),
    .SN(_17399_));
 HAxp5_ASAP7_75t_R _35752_ (.A(_18923_),
    .B(_18924_),
    .CON(_00172_),
    .SN(_00165_));
 HAxp5_ASAP7_75t_R _35753_ (.A(_17412_),
    .B(_18914_),
    .CON(_17440_),
    .SN(_00170_));
 HAxp5_ASAP7_75t_R _35754_ (.A(_18928_),
    .B(_18929_),
    .CON(_17441_),
    .SN(_17419_));
 HAxp5_ASAP7_75t_R _35755_ (.A(_18925_),
    .B(_18930_),
    .CON(_02333_),
    .SN(_17422_));
 HAxp5_ASAP7_75t_R _35756_ (.A(_18931_),
    .B(_18932_),
    .CON(_00179_),
    .SN(_00171_));
 HAxp5_ASAP7_75t_R _35757_ (.A(_17411_),
    .B(_18935_),
    .CON(_17465_),
    .SN(_00174_));
 HAxp5_ASAP7_75t_R _35758_ (.A(_18937_),
    .B(_18936_),
    .CON(_02334_),
    .SN(_00175_));
 HAxp5_ASAP7_75t_R _35759_ (.A(_18941_),
    .B(_18942_),
    .CON(_17463_),
    .SN(_17442_));
 HAxp5_ASAP7_75t_R _35760_ (.A(_18943_),
    .B(_18938_),
    .CON(_02335_),
    .SN(_00176_));
 HAxp5_ASAP7_75t_R _35761_ (.A(_17447_),
    .B(_18944_),
    .CON(_00187_),
    .SN(_00178_));
 HAxp5_ASAP7_75t_R _35762_ (.A(_18945_),
    .B(_18946_),
    .CON(_02336_),
    .SN(_00180_));
 HAxp5_ASAP7_75t_R _35763_ (.A(_18951_),
    .B(_18952_),
    .CON(_17496_),
    .SN(_00181_));
 HAxp5_ASAP7_75t_R _35764_ (.A(_18953_),
    .B(_18948_),
    .CON(_02337_),
    .SN(_00182_));
 HAxp5_ASAP7_75t_R _35765_ (.A(_18956_),
    .B(_18957_),
    .CON(_17494_),
    .SN(_17464_));
 HAxp5_ASAP7_75t_R _35766_ (.A(_17474_),
    .B(_17446_),
    .CON(_00193_),
    .SN(_00186_));
 HAxp5_ASAP7_75t_R _35767_ (.A(_18947_),
    .B(_18958_),
    .CON(_17517_),
    .SN(_00188_));
 HAxp5_ASAP7_75t_R _35768_ (.A(_18962_),
    .B(_18963_),
    .CON(_17526_),
    .SN(_00189_));
 HAxp5_ASAP7_75t_R _35769_ (.A(_18964_),
    .B(_18959_),
    .CON(_02338_),
    .SN(_00190_));
 HAxp5_ASAP7_75t_R _35770_ (.A(_18967_),
    .B(_18968_),
    .CON(_17524_),
    .SN(_17495_));
 HAxp5_ASAP7_75t_R _35771_ (.A(_18970_),
    .B(_17473_),
    .CON(_00198_),
    .SN(_00192_));
 HAxp5_ASAP7_75t_R _35772_ (.A(_18971_),
    .B(_18972_),
    .CON(_17548_),
    .SN(_00194_));
 HAxp5_ASAP7_75t_R _35773_ (.A(_18974_),
    .B(_18973_),
    .CON(_02339_),
    .SN(_00195_));
 HAxp5_ASAP7_75t_R _35774_ (.A(_18980_),
    .B(_18975_),
    .CON(_02340_),
    .SN(_00196_));
 HAxp5_ASAP7_75t_R _35775_ (.A(_18983_),
    .B(_18984_),
    .CON(_02341_),
    .SN(_17525_));
 HAxp5_ASAP7_75t_R _35776_ (.A(_18986_),
    .B(_18987_),
    .CON(_00206_),
    .SN(_00197_));
 HAxp5_ASAP7_75t_R _35777_ (.A(_18988_),
    .B(_18989_),
    .CON(_17575_),
    .SN(_00199_));
 HAxp5_ASAP7_75t_R _35778_ (.A(_18991_),
    .B(_18992_),
    .CON(_17588_),
    .SN(_00200_));
 HAxp5_ASAP7_75t_R _35779_ (.A(_18993_),
    .B(_18990_),
    .CON(_02342_),
    .SN(_00201_));
 HAxp5_ASAP7_75t_R _35780_ (.A(_19000_),
    .B(_19001_),
    .CON(_02343_),
    .SN(_00203_));
 HAxp5_ASAP7_75t_R _35781_ (.A(_19003_),
    .B(_19004_),
    .CON(_00211_),
    .SN(_00205_));
 HAxp5_ASAP7_75t_R _35782_ (.A(_17569_),
    .B(_19007_),
    .CON(_02344_),
    .SN(_00208_));
 HAxp5_ASAP7_75t_R _35783_ (.A(_19014_),
    .B(_19015_),
    .CON(_02345_),
    .SN(_00209_));
 HAxp5_ASAP7_75t_R _35784_ (.A(_19018_),
    .B(_19017_),
    .CON(_00216_),
    .SN(_00210_));
 HAxp5_ASAP7_75t_R _35785_ (.A(_19019_),
    .B(_19020_),
    .CON(_02346_),
    .SN(_00212_));
 HAxp5_ASAP7_75t_R _35786_ (.A(_19021_),
    .B(_19024_),
    .CON(_02347_),
    .SN(_00213_));
 HAxp5_ASAP7_75t_R _35787_ (.A(_19032_),
    .B(_19033_),
    .CON(_02348_),
    .SN(_00214_));
 HAxp5_ASAP7_75t_R _35788_ (.A(_19036_),
    .B(_19037_),
    .CON(_00223_),
    .SN(_00215_));
 HAxp5_ASAP7_75t_R _35789_ (.A(_19038_),
    .B(_19039_),
    .CON(_02349_),
    .SN(_00217_));
 HAxp5_ASAP7_75t_R _35790_ (.A(_19040_),
    .B(_17651_),
    .CON(_02350_),
    .SN(_00219_));
 HAxp5_ASAP7_75t_R _35791_ (.A(_19051_),
    .B(_19052_),
    .CON(_02351_),
    .SN(_00221_));
 HAxp5_ASAP7_75t_R _35792_ (.A(_19055_),
    .B(_19056_),
    .CON(_00228_),
    .SN(_00222_));
 HAxp5_ASAP7_75t_R _35793_ (.A(_19069_),
    .B(_19070_),
    .CON(_00231_),
    .SN(_00227_));
 DFFASRHQNx1_ASAP7_75t_R _35794_ (.CLK(clknet_leaf_44_clk),
    .D(_02352_),
    .QN(_02214_),
    .RESETN(net305),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R _35795_ (.CLK(clknet_leaf_44_clk),
    .D(_02353_),
    .QN(_02213_),
    .RESETN(net306),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R _35796_ (.CLK(clknet_leaf_39_clk),
    .D(_02354_),
    .QN(_00408_),
    .RESETN(net307),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R _35797_ (.CLK(clknet_leaf_39_clk),
    .D(_02355_),
    .QN(_02212_),
    .RESETN(net308),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R _35798_ (.CLK(clknet_leaf_39_clk),
    .D(_02356_),
    .QN(_02211_),
    .RESETN(net74),
    .SETN(net309));
 DFFASRHQNx1_ASAP7_75t_R _35799_ (.CLK(clknet_leaf_8_clk),
    .D(_02357_),
    .QN(_02210_),
    .RESETN(net310),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R _35800_ (.CLK(clknet_leaf_8_clk),
    .D(_02358_),
    .QN(_02215_),
    .RESETN(net311),
    .SETN(net67));
 BUFx16f_ASAP7_75t_R clkbuf_regs_0_core_clock (.A(clk_i),
    .Y(delaynet_0_core_clock));
 TIEHIx1_ASAP7_75t_R _35794__255 (.H(net305));
 BUFx2_ASAP7_75t_R _35803_ (.A(net299),
    .Y(alert_major_o));
 BUFx2_ASAP7_75t_R _35804_ (.A(net300),
    .Y(alert_minor_o));
 BUFx2_ASAP7_75t_R _35805_ (.A(net301),
    .Y(data_addr_o[0]));
 BUFx2_ASAP7_75t_R _35806_ (.A(net302),
    .Y(data_addr_o[1]));
 BUFx2_ASAP7_75t_R _35807_ (.A(\alu_adder_result_ex[2] ),
    .Y(net220));
 BUFx2_ASAP7_75t_R _35808_ (.A(\alu_adder_result_ex[3] ),
    .Y(net223));
 BUFx2_ASAP7_75t_R _35809_ (.A(\alu_adder_result_ex[4] ),
    .Y(net224));
 BUFx4f_ASAP7_75t_R _35810_ (.A(\alu_adder_result_ex[5] ),
    .Y(net225));
 BUFx2_ASAP7_75t_R _35811_ (.A(\alu_adder_result_ex[6] ),
    .Y(net226));
 BUFx3_ASAP7_75t_R _35812_ (.A(\alu_adder_result_ex[7] ),
    .Y(net227));
 BUFx2_ASAP7_75t_R _35813_ (.A(\alu_adder_result_ex[8] ),
    .Y(net228));
 BUFx2_ASAP7_75t_R _35814_ (.A(\alu_adder_result_ex[9] ),
    .Y(net229));
 BUFx2_ASAP7_75t_R _35815_ (.A(\alu_adder_result_ex[10] ),
    .Y(net200));
 BUFx2_ASAP7_75t_R _35816_ (.A(\alu_adder_result_ex[11] ),
    .Y(net201));
 BUFx2_ASAP7_75t_R _35817_ (.A(\alu_adder_result_ex[12] ),
    .Y(net202));
 BUFx3_ASAP7_75t_R _35818_ (.A(\alu_adder_result_ex[13] ),
    .Y(net203));
 BUFx3_ASAP7_75t_R _35819_ (.A(\alu_adder_result_ex[14] ),
    .Y(net204));
 BUFx3_ASAP7_75t_R _35820_ (.A(\alu_adder_result_ex[15] ),
    .Y(net205));
 BUFx2_ASAP7_75t_R _35821_ (.A(\alu_adder_result_ex[16] ),
    .Y(net206));
 BUFx3_ASAP7_75t_R _35822_ (.A(\alu_adder_result_ex[17] ),
    .Y(net207));
 BUFx3_ASAP7_75t_R _35823_ (.A(\alu_adder_result_ex[18] ),
    .Y(net208));
 BUFx3_ASAP7_75t_R _35824_ (.A(\alu_adder_result_ex[19] ),
    .Y(net209));
 BUFx2_ASAP7_75t_R _35825_ (.A(\alu_adder_result_ex[20] ),
    .Y(net210));
 BUFx2_ASAP7_75t_R _35826_ (.A(\alu_adder_result_ex[21] ),
    .Y(net211));
 BUFx2_ASAP7_75t_R _35827_ (.A(\alu_adder_result_ex[22] ),
    .Y(net212));
 BUFx3_ASAP7_75t_R _35828_ (.A(\alu_adder_result_ex[23] ),
    .Y(net213));
 BUFx2_ASAP7_75t_R _35829_ (.A(\alu_adder_result_ex[24] ),
    .Y(net214));
 BUFx4f_ASAP7_75t_R _35830_ (.A(\alu_adder_result_ex[25] ),
    .Y(net215));
 BUFx2_ASAP7_75t_R _35831_ (.A(\alu_adder_result_ex[26] ),
    .Y(net216));
 BUFx4f_ASAP7_75t_R _35832_ (.A(\alu_adder_result_ex[27] ),
    .Y(net217));
 BUFx4f_ASAP7_75t_R _35833_ (.A(\alu_adder_result_ex[28] ),
    .Y(net218));
 BUFx4f_ASAP7_75t_R _35834_ (.A(\alu_adder_result_ex[29] ),
    .Y(net219));
 BUFx3_ASAP7_75t_R _35835_ (.A(\alu_adder_result_ex[30] ),
    .Y(net221));
 BUFx3_ASAP7_75t_R _35836_ (.A(\alu_adder_result_ex[31] ),
    .Y(net222));
 BUFx2_ASAP7_75t_R _35837_ (.A(net303),
    .Y(instr_addr_o[0]));
 BUFx2_ASAP7_75t_R _35838_ (.A(net304),
    .Y(instr_addr_o[1]));
 DFFASRHQNx1_ASAP7_75t_R \core_busy_q$_DFF_PN0_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(core_busy_d),
    .QN(_02209_),
    .RESETN(net312),
    .SETN(net67));
 DLLx1_ASAP7_75t_R \core_clock_gate_i.en_latch$_DLATCH_N_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_00006_),
    .Q(\core_clock_gate_i.en_latch ));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02359_),
    .QN(_00788_),
    .RESETN(net313),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02360_),
    .QN(_01453_),
    .RESETN(net314),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02361_),
    .QN(_00786_),
    .RESETN(net315),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02362_),
    .QN(_02208_),
    .RESETN(net316),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02363_),
    .QN(_02207_),
    .RESETN(net317),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02364_),
    .QN(_02206_),
    .RESETN(net318),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02365_),
    .QN(_02205_),
    .RESETN(net319),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02366_),
    .QN(_02204_),
    .RESETN(net320),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02367_),
    .QN(_02203_),
    .RESETN(net321),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02368_),
    .QN(_02202_),
    .RESETN(net322),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02369_),
    .QN(_02201_),
    .RESETN(net323),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02370_),
    .QN(_02200_),
    .RESETN(net324),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02371_),
    .QN(_02199_),
    .RESETN(net325),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02372_),
    .QN(_02198_),
    .RESETN(net326),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02373_),
    .QN(_02197_),
    .RESETN(net327),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02374_),
    .QN(_02196_),
    .RESETN(net328),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02375_),
    .QN(_02195_),
    .RESETN(net329),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02376_),
    .QN(_02194_),
    .RESETN(net330),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02377_),
    .QN(_02193_),
    .RESETN(net331),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02378_),
    .QN(_02192_),
    .RESETN(net332),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02379_),
    .QN(_02191_),
    .RESETN(net333),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02380_),
    .QN(_02190_),
    .RESETN(net334),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02381_),
    .QN(_02189_),
    .RESETN(net335),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02382_),
    .QN(_02188_),
    .RESETN(net336),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02383_),
    .QN(_02187_),
    .RESETN(net337),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02384_),
    .QN(_02186_),
    .RESETN(net338),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02385_),
    .QN(_02185_),
    .RESETN(net339),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[32]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02386_),
    .QN(_02184_),
    .RESETN(net340),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[33]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02387_),
    .QN(_02183_),
    .RESETN(net341),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02388_),
    .QN(_02182_),
    .RESETN(net342),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02389_),
    .QN(_02181_),
    .RESETN(net343),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02390_),
    .QN(_02180_),
    .RESETN(net344),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_02391_),
    .QN(_02179_),
    .RESETN(net345),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02392_),
    .QN(_02178_),
    .RESETN(net346),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02393_),
    .QN(_02177_),
    .RESETN(net347),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02394_),
    .QN(_02176_),
    .RESETN(net348),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02395_),
    .QN(_02175_),
    .RESETN(net349),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02396_),
    .QN(_02174_),
    .RESETN(net350),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02397_),
    .QN(_02173_),
    .RESETN(net351),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02398_),
    .QN(_02172_),
    .RESETN(net352),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02399_),
    .QN(_02171_),
    .RESETN(net353),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02400_),
    .QN(_02170_),
    .RESETN(net354),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02401_),
    .QN(_02169_),
    .RESETN(net355),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02402_),
    .QN(_02168_),
    .RESETN(net356),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02403_),
    .QN(_02167_),
    .RESETN(net357),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02404_),
    .QN(_02166_),
    .RESETN(net358),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02405_),
    .QN(_02165_),
    .RESETN(net359),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02406_),
    .QN(_02164_),
    .RESETN(net360),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02407_),
    .QN(_02163_),
    .RESETN(net361),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02408_),
    .QN(_02162_),
    .RESETN(net362),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02409_),
    .QN(_02161_),
    .RESETN(net363),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02410_),
    .QN(_02160_),
    .RESETN(net364),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02411_),
    .QN(_02159_),
    .RESETN(net365),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02412_),
    .QN(_02158_),
    .RESETN(net366),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02413_),
    .QN(_02157_),
    .RESETN(net367),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02414_),
    .QN(_02156_),
    .RESETN(net368),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02415_),
    .QN(_02155_),
    .RESETN(net369),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02416_),
    .QN(_02154_),
    .RESETN(net370),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02417_),
    .QN(_02153_),
    .RESETN(net371),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02418_),
    .QN(_02152_),
    .RESETN(net372),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02419_),
    .QN(_02151_),
    .RESETN(net373),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .D(_02420_),
    .QN(_02150_),
    .RESETN(net374),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02421_),
    .QN(_02149_),
    .RESETN(net375),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02422_),
    .QN(_02148_),
    .RESETN(net376),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02423_),
    .QN(_02147_),
    .RESETN(net377),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02424_),
    .QN(_02146_),
    .RESETN(net378),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02425_),
    .QN(_00787_),
    .RESETN(net379),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02426_),
    .QN(_02145_),
    .RESETN(net380),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02427_),
    .QN(_02144_),
    .RESETN(net381),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02428_),
    .QN(_02143_),
    .RESETN(net382),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02429_),
    .QN(_02142_),
    .RESETN(net383),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02430_),
    .QN(_02141_),
    .RESETN(net384),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02431_),
    .QN(_02140_),
    .RESETN(net385),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02432_),
    .QN(_02139_),
    .RESETN(net386),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02433_),
    .QN(_02138_),
    .RESETN(net387),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02434_),
    .QN(_02137_),
    .RESETN(net388),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02435_),
    .QN(_02136_),
    .RESETN(net389),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02436_),
    .QN(_02135_),
    .RESETN(net390),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02437_),
    .QN(_02134_),
    .RESETN(net391),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02438_),
    .QN(_02133_),
    .RESETN(net392),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02439_),
    .QN(_02132_),
    .RESETN(net393),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02440_),
    .QN(_02131_),
    .RESETN(net394),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02441_),
    .QN(_02130_),
    .RESETN(net395),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02442_),
    .QN(_02129_),
    .RESETN(net396),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02443_),
    .QN(_02128_),
    .RESETN(net397),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02444_),
    .QN(_02127_),
    .RESETN(net398),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02445_),
    .QN(_02126_),
    .RESETN(net399),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02446_),
    .QN(_02125_),
    .RESETN(net400),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02447_),
    .QN(_02124_),
    .RESETN(net401),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02448_),
    .QN(_02123_),
    .RESETN(net402),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02449_),
    .QN(_02122_),
    .RESETN(net403),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[32]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02450_),
    .QN(_02121_),
    .RESETN(net404),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[33]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02451_),
    .QN(_02120_),
    .RESETN(net405),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02452_),
    .QN(_02119_),
    .RESETN(net406),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02453_),
    .QN(_02118_),
    .RESETN(net407),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02454_),
    .QN(_02117_),
    .RESETN(net408),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02455_),
    .QN(_02116_),
    .RESETN(net409),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02456_),
    .QN(_02115_),
    .RESETN(net410),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02457_),
    .QN(_02114_),
    .RESETN(net411),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02458_),
    .QN(_02113_),
    .RESETN(net412),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02459_),
    .QN(_02112_),
    .RESETN(net413),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .D(_02460_),
    .QN(_02111_),
    .RESETN(net414),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02461_),
    .QN(_02110_),
    .RESETN(net415),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02462_),
    .QN(_02109_),
    .RESETN(net416),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02463_),
    .QN(_02108_),
    .RESETN(net417),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02464_),
    .QN(_02107_),
    .RESETN(net418),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02465_),
    .QN(_02106_),
    .RESETN(net419),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02466_),
    .QN(_02105_),
    .RESETN(net420),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02467_),
    .QN(_02104_),
    .RESETN(net421),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02468_),
    .QN(_02103_),
    .RESETN(net422),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02469_),
    .QN(_02102_),
    .RESETN(net423),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02470_),
    .QN(_02101_),
    .RESETN(net424),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02471_),
    .QN(_02100_),
    .RESETN(net425),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02472_),
    .QN(_02099_),
    .RESETN(net426),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02473_),
    .QN(_02098_),
    .RESETN(net427),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02474_),
    .QN(_02097_),
    .RESETN(net428),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .D(_02475_),
    .QN(_02096_),
    .RESETN(net429),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02476_),
    .QN(_02095_),
    .RESETN(net430),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02477_),
    .QN(_02094_),
    .RESETN(net431),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02478_),
    .QN(_02093_),
    .RESETN(net432),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02479_),
    .QN(_02092_),
    .RESETN(net433),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02480_),
    .QN(_02091_),
    .RESETN(net434),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02481_),
    .QN(_02090_),
    .RESETN(net435),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02482_),
    .QN(_02089_),
    .RESETN(net436),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02483_),
    .QN(_02088_),
    .RESETN(net437),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .D(_02484_),
    .QN(_02087_),
    .RESETN(net438),
    .SETN(net73));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02485_),
    .QN(_02086_),
    .RESETN(net439),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02486_),
    .QN(_02085_),
    .RESETN(net440),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02487_),
    .QN(_02084_),
    .RESETN(net441),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02488_),
    .QN(_02083_),
    .RESETN(net442),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.priv_lvl_q[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_31_clk),
    .D(_02489_),
    .QN(_02082_),
    .RESETN(net72),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.priv_lvl_q[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_31_clk),
    .D(_02490_),
    .QN(_18850_),
    .RESETN(net72),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[0]$_DFFE_PN1N_  (.CLK(clknet_leaf_31_clk),
    .D(_02491_),
    .QN(_02081_),
    .RESETN(net72),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02492_),
    .QN(_02080_),
    .RESETN(net446),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .D(_02493_),
    .QN(_00783_),
    .RESETN(net447),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02494_),
    .QN(_02079_),
    .RESETN(net448),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02495_),
    .QN(_00790_),
    .RESETN(net449),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[1]$_DFFE_PN1N_  (.CLK(clknet_leaf_31_clk),
    .D(_02496_),
    .QN(_02078_),
    .RESETN(net72),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02497_),
    .QN(_01460_),
    .RESETN(net451),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_02498_),
    .QN(_02077_),
    .RESETN(net452),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_02499_),
    .QN(_02076_),
    .RESETN(net453),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_02500_),
    .QN(_02075_),
    .RESETN(net454),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02501_),
    .QN(_02074_),
    .RESETN(net455),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02502_),
    .QN(_02073_),
    .RESETN(net456),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02503_),
    .QN(_02072_),
    .RESETN(net457),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02504_),
    .QN(_02071_),
    .RESETN(net458),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02505_),
    .QN(_02070_),
    .RESETN(net459),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02506_),
    .QN(_02069_),
    .RESETN(net460),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02507_),
    .QN(_02068_),
    .RESETN(net461),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02508_),
    .QN(_02067_),
    .RESETN(net462),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02509_),
    .QN(_02066_),
    .RESETN(net463),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02510_),
    .QN(_02065_),
    .RESETN(net464),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02511_),
    .QN(_00789_),
    .RESETN(net465),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02512_),
    .QN(_02064_),
    .RESETN(net466),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02513_),
    .QN(_02063_),
    .RESETN(net467),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02514_),
    .QN(_02062_),
    .RESETN(net468),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02515_),
    .QN(_02061_),
    .RESETN(net469),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02516_),
    .QN(_02060_),
    .RESETN(net470),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02517_),
    .QN(_02059_),
    .RESETN(net471),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02518_),
    .QN(_02058_),
    .RESETN(net472),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02519_),
    .QN(_02057_),
    .RESETN(net473),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02520_),
    .QN(_02056_),
    .RESETN(net474),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02521_),
    .QN(_02055_),
    .RESETN(net475),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02522_),
    .QN(_02054_),
    .RESETN(net476),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02523_),
    .QN(_02053_),
    .RESETN(net477),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02524_),
    .QN(_02052_),
    .RESETN(net478),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02525_),
    .QN(_01461_),
    .RESETN(net479),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02526_),
    .QN(_01462_),
    .RESETN(net480),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02527_),
    .QN(_01463_),
    .RESETN(net481),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02528_),
    .QN(_01464_),
    .RESETN(net482),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02529_),
    .QN(_02051_),
    .RESETN(net483),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02530_),
    .QN(_02050_),
    .RESETN(net484),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02531_),
    .QN(_02049_),
    .RESETN(net485),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02532_),
    .QN(_02048_),
    .RESETN(net486),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02533_),
    .QN(_02047_),
    .RESETN(net487),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02534_),
    .QN(_02046_),
    .RESETN(net488),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02535_),
    .QN(_02045_),
    .RESETN(net489),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02536_),
    .QN(_02044_),
    .RESETN(net490),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02537_),
    .QN(_02043_),
    .RESETN(net491),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02538_),
    .QN(_02042_),
    .RESETN(net492),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02539_),
    .QN(_02041_),
    .RESETN(net493),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02540_),
    .QN(_02040_),
    .RESETN(net494),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02541_),
    .QN(_02039_),
    .RESETN(net495),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02542_),
    .QN(_02038_),
    .RESETN(net496),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02543_),
    .QN(_02037_),
    .RESETN(net497),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02544_),
    .QN(_02036_),
    .RESETN(net498),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02545_),
    .QN(_02035_),
    .RESETN(net499),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02546_),
    .QN(_02034_),
    .RESETN(net500),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02547_),
    .QN(_02033_),
    .RESETN(net501),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02548_),
    .QN(_02032_),
    .RESETN(net502),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02549_),
    .QN(_02031_),
    .RESETN(net503),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02550_),
    .QN(_02030_),
    .RESETN(net504),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02551_),
    .QN(_02029_),
    .RESETN(net505),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02552_),
    .QN(_02028_),
    .RESETN(net506),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02553_),
    .QN(_02027_),
    .RESETN(net507),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02554_),
    .QN(_02026_),
    .RESETN(net508),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02555_),
    .QN(_02025_),
    .RESETN(net509),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02556_),
    .QN(_02024_),
    .RESETN(net510),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02557_),
    .QN(_02023_),
    .RESETN(net511),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02558_),
    .QN(_02022_),
    .RESETN(net512),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02559_),
    .QN(_02021_),
    .RESETN(net513),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02560_),
    .QN(_02020_),
    .RESETN(net514),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02561_),
    .QN(_02019_),
    .RESETN(net515),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02562_),
    .QN(_02018_),
    .RESETN(net516),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02563_),
    .QN(_02017_),
    .RESETN(net517),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02564_),
    .QN(_02016_),
    .RESETN(net518),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02565_),
    .QN(_02015_),
    .RESETN(net519),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02566_),
    .QN(_02014_),
    .RESETN(net520),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02567_),
    .QN(_02013_),
    .RESETN(net521),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02568_),
    .QN(_02012_),
    .RESETN(net522),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02569_),
    .QN(_02011_),
    .RESETN(net523),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02570_),
    .QN(_02010_),
    .RESETN(net524),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02571_),
    .QN(_02009_),
    .RESETN(net525),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02572_),
    .QN(_02008_),
    .RESETN(net526),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02573_),
    .QN(_02007_),
    .RESETN(net527),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02574_),
    .QN(_02006_),
    .RESETN(net528),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02575_),
    .QN(_02005_),
    .RESETN(net529),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02576_),
    .QN(_02004_),
    .RESETN(net530),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02577_),
    .QN(_02003_),
    .RESETN(net531),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02578_),
    .QN(_02002_),
    .RESETN(net532),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02579_),
    .QN(_02001_),
    .RESETN(net533),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02580_),
    .QN(_02000_),
    .RESETN(net534),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02581_),
    .QN(_01999_),
    .RESETN(net535),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02582_),
    .QN(_01998_),
    .RESETN(net536),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02583_),
    .QN(_01997_),
    .RESETN(net537),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02584_),
    .QN(_01996_),
    .RESETN(net538),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02585_),
    .QN(_01995_),
    .RESETN(net539),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02586_),
    .QN(_01994_),
    .RESETN(net540),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02587_),
    .QN(_01993_),
    .RESETN(net541),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02588_),
    .QN(_01992_),
    .RESETN(net542),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02589_),
    .QN(_01991_),
    .RESETN(net543),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02590_),
    .QN(_01990_),
    .RESETN(net544),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02591_),
    .QN(_01989_),
    .RESETN(net545),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02592_),
    .QN(_01988_),
    .RESETN(net546),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02593_),
    .QN(_01987_),
    .RESETN(net547),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02594_),
    .QN(_01986_),
    .RESETN(net548),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02595_),
    .QN(_01985_),
    .RESETN(net549),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_02596_),
    .QN(_01984_),
    .RESETN(net550),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02597_),
    .QN(_01983_),
    .RESETN(net551),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02598_),
    .QN(_01982_),
    .RESETN(net552),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02599_),
    .QN(_01981_),
    .RESETN(net553),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02600_),
    .QN(_01980_),
    .RESETN(net554),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02601_),
    .QN(_01979_),
    .RESETN(net555),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02602_),
    .QN(_01978_),
    .RESETN(net556),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02603_),
    .QN(_01977_),
    .RESETN(net557),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02604_),
    .QN(_01976_),
    .RESETN(net558),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02605_),
    .QN(_01975_),
    .RESETN(net559),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02606_),
    .QN(_01974_),
    .RESETN(net560),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02607_),
    .QN(_01973_),
    .RESETN(net561),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02608_),
    .QN(_01972_),
    .RESETN(net562),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02609_),
    .QN(_01971_),
    .RESETN(net563),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02610_),
    .QN(_01970_),
    .RESETN(net564),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02611_),
    .QN(_01969_),
    .RESETN(net565),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02612_),
    .QN(_01968_),
    .RESETN(net566),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02613_),
    .QN(_01967_),
    .RESETN(net567),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02614_),
    .QN(_01966_),
    .RESETN(net568),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02615_),
    .QN(_01965_),
    .RESETN(net569),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02616_),
    .QN(_01964_),
    .RESETN(net570),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02617_),
    .QN(_01963_),
    .RESETN(net571),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02618_),
    .QN(_01962_),
    .RESETN(net572),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02619_),
    .QN(_01961_),
    .RESETN(net573),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02620_),
    .QN(_01960_),
    .RESETN(net574),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02621_),
    .QN(_01959_),
    .RESETN(net575),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02622_),
    .QN(_01958_),
    .RESETN(net576),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02623_),
    .QN(_01957_),
    .RESETN(net577),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02624_),
    .QN(_01956_),
    .RESETN(net578),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02625_),
    .QN(_01955_),
    .RESETN(net579),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02626_),
    .QN(_01954_),
    .RESETN(net580),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02627_),
    .QN(_01953_),
    .RESETN(net581),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02628_),
    .QN(_01952_),
    .RESETN(net582),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02629_),
    .QN(_01951_),
    .RESETN(net583),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02630_),
    .QN(_01950_),
    .RESETN(net584),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02631_),
    .QN(_01949_),
    .RESETN(net585),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02632_),
    .QN(_01948_),
    .RESETN(net586),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02633_),
    .QN(_01947_),
    .RESETN(net587),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02634_),
    .QN(_01946_),
    .RESETN(net588),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02635_),
    .QN(_01945_),
    .RESETN(net589),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02636_),
    .QN(_01944_),
    .RESETN(net590),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02637_),
    .QN(_01943_),
    .RESETN(net591),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02638_),
    .QN(_01942_),
    .RESETN(net592),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02639_),
    .QN(_01941_),
    .RESETN(net593),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02640_),
    .QN(_01940_),
    .RESETN(net594),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02641_),
    .QN(_01939_),
    .RESETN(net595),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02642_),
    .QN(_01938_),
    .RESETN(net596),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02643_),
    .QN(_01937_),
    .RESETN(net597),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02644_),
    .QN(_01936_),
    .RESETN(net598),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02645_),
    .QN(_01935_),
    .RESETN(net599),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02646_),
    .QN(_01934_),
    .RESETN(net600),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02647_),
    .QN(_01933_),
    .RESETN(net601),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02648_),
    .QN(_01932_),
    .RESETN(net602),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02649_),
    .QN(_01931_),
    .RESETN(net603),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02650_),
    .QN(_01930_),
    .RESETN(net604),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02651_),
    .QN(_01929_),
    .RESETN(net605),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02652_),
    .QN(_01928_),
    .RESETN(net606),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02653_),
    .QN(_01927_),
    .RESETN(net607),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02654_),
    .QN(_01926_),
    .RESETN(net608),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02655_),
    .QN(_01925_),
    .RESETN(net609),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02656_),
    .QN(_01924_),
    .RESETN(net610),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02657_),
    .QN(_01923_),
    .RESETN(net611),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02658_),
    .QN(_01922_),
    .RESETN(net612),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02659_),
    .QN(_01921_),
    .RESETN(net613),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02660_),
    .QN(_01920_),
    .RESETN(net614),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02661_),
    .QN(_01919_),
    .RESETN(net615),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02662_),
    .QN(_01918_),
    .RESETN(net616),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02663_),
    .QN(_01917_),
    .RESETN(net617),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02664_),
    .QN(_01916_),
    .RESETN(net618),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02665_),
    .QN(_01915_),
    .RESETN(net619),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02666_),
    .QN(_01914_),
    .RESETN(net620),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02667_),
    .QN(_01913_),
    .RESETN(net621),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02668_),
    .QN(_01912_),
    .RESETN(net622),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_02669_),
    .QN(_01911_),
    .RESETN(net623),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02670_),
    .QN(_01910_),
    .RESETN(net624),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_02671_),
    .QN(_01909_),
    .RESETN(net625),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02672_),
    .QN(_01908_),
    .RESETN(net626),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02673_),
    .QN(_01907_),
    .RESETN(net627),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_02674_),
    .QN(_01906_),
    .RESETN(net628),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02675_),
    .QN(_01905_),
    .RESETN(net629),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02676_),
    .QN(_01904_),
    .RESETN(net630),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02677_),
    .QN(_01903_),
    .RESETN(net631),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02678_),
    .QN(_01902_),
    .RESETN(net632),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_02679_),
    .QN(_01901_),
    .RESETN(net633),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02680_),
    .QN(_01900_),
    .RESETN(net634),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02681_),
    .QN(_01899_),
    .RESETN(net635),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02682_),
    .QN(_01898_),
    .RESETN(net636),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_02683_),
    .QN(_01897_),
    .RESETN(net637),
    .SETN(net71));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_02684_),
    .QN(_01896_),
    .RESETN(net638),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02685_),
    .QN(_01895_),
    .RESETN(net639),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02686_),
    .QN(_01894_),
    .RESETN(net640),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02687_),
    .QN(_01893_),
    .RESETN(net641),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02688_),
    .QN(_01892_),
    .RESETN(net642),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02689_),
    .QN(_01891_),
    .RESETN(net643),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_02690_),
    .QN(_01890_),
    .RESETN(net644),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02691_),
    .QN(_01889_),
    .RESETN(net645),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rdata_q[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .D(_02692_),
    .QN(_01888_),
    .RESETN(net72),
    .SETN(net646));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02693_),
    .QN(_01887_),
    .RESETN(net647),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02694_),
    .QN(_01886_),
    .RESETN(net648),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02695_),
    .QN(_01885_),
    .RESETN(net649),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02696_),
    .QN(_01884_),
    .RESETN(net650),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02697_),
    .QN(_01883_),
    .RESETN(net651),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02698_),
    .QN(_01882_),
    .RESETN(net652),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02699_),
    .QN(_01881_),
    .RESETN(net653),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02700_),
    .QN(_01880_),
    .RESETN(net654),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02701_),
    .QN(_01879_),
    .RESETN(net655),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02702_),
    .QN(_01878_),
    .RESETN(net656),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02703_),
    .QN(_01877_),
    .RESETN(net657),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02704_),
    .QN(_01876_),
    .RESETN(net658),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02705_),
    .QN(_01875_),
    .RESETN(net659),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02706_),
    .QN(_01874_),
    .RESETN(net660),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02707_),
    .QN(_01873_),
    .RESETN(net661),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_02708_),
    .QN(_01872_),
    .RESETN(net662),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02709_),
    .QN(_01871_),
    .RESETN(net663),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02710_),
    .QN(_01870_),
    .RESETN(net664),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02711_),
    .QN(_01869_),
    .RESETN(net665),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02712_),
    .QN(_01868_),
    .RESETN(net666),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02713_),
    .QN(_01867_),
    .RESETN(net667),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02714_),
    .QN(_01866_),
    .RESETN(net668),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02715_),
    .QN(_01865_),
    .RESETN(net669),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02716_),
    .QN(_01864_),
    .RESETN(net670),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02717_),
    .QN(_01863_),
    .RESETN(net671),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02718_),
    .QN(_01862_),
    .RESETN(net672),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02719_),
    .QN(_01861_),
    .RESETN(net673),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_02720_),
    .QN(_01860_),
    .RESETN(net674),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02721_),
    .QN(_01859_),
    .RESETN(net675),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02722_),
    .QN(_01858_),
    .RESETN(net676),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02723_),
    .QN(_01857_),
    .RESETN(net677),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02724_),
    .QN(_01856_),
    .RESETN(net678),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02725_),
    .QN(_01855_),
    .RESETN(net679),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02726_),
    .QN(_01854_),
    .RESETN(net680),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_02727_),
    .QN(_01853_),
    .RESETN(net681),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02728_),
    .QN(_01852_),
    .RESETN(net682),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .D(_02729_),
    .QN(_01851_),
    .RESETN(net72),
    .SETN(net683));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02730_),
    .QN(_01850_),
    .RESETN(net684),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02731_),
    .QN(_01849_),
    .RESETN(net685),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02732_),
    .QN(_01848_),
    .RESETN(net686),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02733_),
    .QN(_01847_),
    .RESETN(net687),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02734_),
    .QN(_01846_),
    .RESETN(net688),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_02735_),
    .QN(_01845_),
    .RESETN(net689),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02736_),
    .QN(_01844_),
    .RESETN(net690),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02737_),
    .QN(_01843_),
    .RESETN(net691),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02738_),
    .QN(_01842_),
    .RESETN(net692),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02739_),
    .QN(_01841_),
    .RESETN(net693),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02740_),
    .QN(_01840_),
    .RESETN(net694),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02741_),
    .QN(_01839_),
    .RESETN(net695),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02742_),
    .QN(_01838_),
    .RESETN(net696),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02743_),
    .QN(_01837_),
    .RESETN(net697),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02744_),
    .QN(_01836_),
    .RESETN(net698),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02745_),
    .QN(_01835_),
    .RESETN(net699),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02746_),
    .QN(_01834_),
    .RESETN(net700),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02747_),
    .QN(_01833_),
    .RESETN(net701),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02748_),
    .QN(_01832_),
    .RESETN(net702),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02749_),
    .QN(_01831_),
    .RESETN(net703),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02750_),
    .QN(_01830_),
    .RESETN(net704),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02751_),
    .QN(_01829_),
    .RESETN(net705),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02752_),
    .QN(_01828_),
    .RESETN(net706),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02753_),
    .QN(_01827_),
    .RESETN(net707),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02754_),
    .QN(_01826_),
    .RESETN(net708),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02755_),
    .QN(_01825_),
    .RESETN(net709),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02756_),
    .QN(_01824_),
    .RESETN(net710),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02757_),
    .QN(_01823_),
    .RESETN(net711),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02758_),
    .QN(_01822_),
    .RESETN(net712),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02759_),
    .QN(_01821_),
    .RESETN(net713),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02760_),
    .QN(_01820_),
    .RESETN(net714),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02761_),
    .QN(_01819_),
    .RESETN(net715),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_02762_),
    .QN(_01818_),
    .RESETN(net716),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02763_),
    .QN(_01467_),
    .RESETN(net717),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02764_),
    .QN(_00785_),
    .RESETN(net718),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02765_),
    .QN(_00784_),
    .RESETN(net719),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02766_),
    .QN(_01468_),
    .RESETN(net720),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02767_),
    .QN(_01469_),
    .RESETN(net721),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02768_),
    .QN(_01470_),
    .RESETN(net722),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02769_),
    .QN(_01471_),
    .RESETN(net723),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02770_),
    .QN(_01472_),
    .RESETN(net724),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02771_),
    .QN(_01473_),
    .RESETN(net725),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02772_),
    .QN(_01474_),
    .RESETN(net726),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_02773_),
    .QN(_01475_),
    .RESETN(net727),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02774_),
    .QN(_01476_),
    .RESETN(net728),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_02775_),
    .QN(_01477_),
    .RESETN(net729),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02776_),
    .QN(_01478_),
    .RESETN(net730),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02777_),
    .QN(_01479_),
    .RESETN(net731),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02778_),
    .QN(_01480_),
    .RESETN(net732),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02779_),
    .QN(_01481_),
    .RESETN(net733),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02780_),
    .QN(_00007_),
    .RESETN(net734),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_02781_),
    .QN(_00008_),
    .RESETN(net735),
    .SETN(net68));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02782_),
    .QN(_00009_),
    .RESETN(net736),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_02783_),
    .QN(_00010_),
    .RESETN(net737),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_02784_),
    .QN(_00011_),
    .RESETN(net738),
    .SETN(net69));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_02785_),
    .QN(_01465_),
    .RESETN(net739),
    .SETN(net70));
 DFFASRHQNx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .D(_02786_),
    .QN(_01466_),
    .RESETN(net740),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02787_),
    .QN(_01817_),
    .RESETN(net741),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02788_),
    .QN(_18867_),
    .RESETN(net742),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02789_),
    .QN(_18868_),
    .RESETN(net743),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02790_),
    .QN(_00069_),
    .RESETN(net744),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02791_),
    .QN(_00070_),
    .RESETN(net745),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02792_),
    .QN(_01457_),
    .RESETN(net746),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.CLK(clknet_leaf_44_clk),
    .D(_00000_),
    .QN(_02216_),
    .RESETN(net74),
    .SETN(net747));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .D(_00001_),
    .QN(_01459_),
    .RESETN(net748),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .D(_00002_),
    .QN(_02217_),
    .RESETN(net749),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .D(_00003_),
    .QN(_02218_),
    .RESETN(net750),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .D(_00004_),
    .QN(_00407_),
    .RESETN(net751),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .D(_00005_),
    .QN(_01816_),
    .RESETN(net752),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02793_),
    .QN(_00106_),
    .RESETN(net753),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02794_),
    .QN(_00116_),
    .RESETN(net754),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02795_),
    .QN(_00115_),
    .RESETN(net755),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02796_),
    .QN(_00118_),
    .RESETN(net756),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02797_),
    .QN(_00117_),
    .RESETN(net757),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02798_),
    .QN(_00120_),
    .RESETN(net758),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02799_),
    .QN(_00119_),
    .RESETN(net759),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02800_),
    .QN(_00122_),
    .RESETN(net760),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02801_),
    .QN(_00121_),
    .RESETN(net761),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02802_),
    .QN(_00124_),
    .RESETN(net762),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02803_),
    .QN(_00123_),
    .RESETN(net763),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02804_),
    .QN(_00105_),
    .RESETN(net764),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02805_),
    .QN(_00126_),
    .RESETN(net765),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02806_),
    .QN(_00125_),
    .RESETN(net766),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02807_),
    .QN(_00128_),
    .RESETN(net767),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02808_),
    .QN(_00127_),
    .RESETN(net768),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02809_),
    .QN(_00130_),
    .RESETN(net769),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02810_),
    .QN(_00129_),
    .RESETN(net770),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02811_),
    .QN(_00132_),
    .RESETN(net771),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02812_),
    .QN(_00131_),
    .RESETN(net772),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02813_),
    .QN(_00134_),
    .RESETN(net773),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02814_),
    .QN(_00133_),
    .RESETN(net774),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02815_),
    .QN(_00108_),
    .RESETN(net775),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02816_),
    .QN(_00136_),
    .RESETN(net776),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02817_),
    .QN(_00135_),
    .RESETN(net777),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02818_),
    .QN(_00107_),
    .RESETN(net778),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02819_),
    .QN(_00110_),
    .RESETN(net779),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02820_),
    .QN(_00109_),
    .RESETN(net780),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02821_),
    .QN(_00112_),
    .RESETN(net781),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02822_),
    .QN(_00111_),
    .RESETN(net782),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02823_),
    .QN(_00114_),
    .RESETN(net783),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .D(_02824_),
    .QN(_00113_),
    .RESETN(net784),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02825_),
    .QN(_00071_),
    .RESETN(net785),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02826_),
    .QN(_00082_),
    .RESETN(net786),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02827_),
    .QN(_00083_),
    .RESETN(net787),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02828_),
    .QN(_00084_),
    .RESETN(net788),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02829_),
    .QN(_00085_),
    .RESETN(net789),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02830_),
    .QN(_00086_),
    .RESETN(net790),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02831_),
    .QN(_00087_),
    .RESETN(net791),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02832_),
    .QN(_00088_),
    .RESETN(net792),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02833_),
    .QN(_00089_),
    .RESETN(net793),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02834_),
    .QN(_00090_),
    .RESETN(net794),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02835_),
    .QN(_00091_),
    .RESETN(net795),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02836_),
    .QN(_00072_),
    .RESETN(net796),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02837_),
    .QN(_00092_),
    .RESETN(net797),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02838_),
    .QN(_00093_),
    .RESETN(net798),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02839_),
    .QN(_00094_),
    .RESETN(net799),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02840_),
    .QN(_00095_),
    .RESETN(net800),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02841_),
    .QN(_00096_),
    .RESETN(net801),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02842_),
    .QN(_00097_),
    .RESETN(net802),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02843_),
    .QN(_00098_),
    .RESETN(net803),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02844_),
    .QN(_00099_),
    .RESETN(net804),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02845_),
    .QN(_00100_),
    .RESETN(net805),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02846_),
    .QN(_00101_),
    .RESETN(net806),
    .SETN(net197));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02847_),
    .QN(_00073_),
    .RESETN(net807),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02848_),
    .QN(_00102_),
    .RESETN(net808),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02849_),
    .QN(_00103_),
    .RESETN(net809),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .D(_02850_),
    .QN(_00075_),
    .RESETN(net810),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02851_),
    .QN(_00076_),
    .RESETN(net811),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02852_),
    .QN(_00077_),
    .RESETN(net812),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02853_),
    .QN(_00078_),
    .RESETN(net813),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02854_),
    .QN(_00079_),
    .RESETN(net814),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_02855_),
    .QN(_00080_),
    .RESETN(net815),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .D(_02856_),
    .QN(_00081_),
    .RESETN(net816),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \fetch_enable_q$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_02857_),
    .QN(_01815_),
    .RESETN(net817),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_02858_),
    .QN(_01814_),
    .RESETN(net818),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[100]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02859_),
    .QN(_00543_),
    .RESETN(net819),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[101]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02860_),
    .QN(_00575_),
    .RESETN(net820),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[102]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02861_),
    .QN(_00605_),
    .RESETN(net821),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[103]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02862_),
    .QN(_00635_),
    .RESETN(net822),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[104]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02863_),
    .QN(_00665_),
    .RESETN(net823),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[105]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02864_),
    .QN(_00695_),
    .RESETN(net824),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[106]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02865_),
    .QN(_00725_),
    .RESETN(net825),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[107]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02866_),
    .QN(_00755_),
    .RESETN(net826),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[108]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02867_),
    .QN(_00451_),
    .RESETN(net827),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[109]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02868_),
    .QN(_00826_),
    .RESETN(net828),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02869_),
    .QN(_01813_),
    .RESETN(net829),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[110]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02870_),
    .QN(_00859_),
    .RESETN(net830),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[111]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02871_),
    .QN(_00892_),
    .RESETN(net831),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[112]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_02872_),
    .QN(_00925_),
    .RESETN(net832),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[113]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02873_),
    .QN(_00958_),
    .RESETN(net833),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[114]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02874_),
    .QN(_00991_),
    .RESETN(net834),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[115]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02875_),
    .QN(_01024_),
    .RESETN(net835),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[116]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02876_),
    .QN(_01057_),
    .RESETN(net836),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[117]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02877_),
    .QN(_01090_),
    .RESETN(net837),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[118]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02878_),
    .QN(_01123_),
    .RESETN(net838),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[119]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02879_),
    .QN(_01156_),
    .RESETN(net839),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_02880_),
    .QN(_01812_),
    .RESETN(net840),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[120]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02881_),
    .QN(_01189_),
    .RESETN(net841),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[121]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02882_),
    .QN(_01222_),
    .RESETN(net842),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[122]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02883_),
    .QN(_01255_),
    .RESETN(net843),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[123]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02884_),
    .QN(_01288_),
    .RESETN(net844),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[124]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_02885_),
    .QN(_01321_),
    .RESETN(net845),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[125]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02886_),
    .QN(_01354_),
    .RESETN(net846),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[126]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_02887_),
    .QN(_01387_),
    .RESETN(net847),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[127]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_02888_),
    .QN(_01420_),
    .RESETN(net848),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[128]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_02889_),
    .QN(_00419_),
    .RESETN(net849),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[129]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02890_),
    .QN(_00372_),
    .RESETN(net850),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_02891_),
    .QN(_01811_),
    .RESETN(net851),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[130]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02892_),
    .QN(_00483_),
    .RESETN(net852),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[131]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02893_),
    .QN(_00514_),
    .RESETN(net853),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[132]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02894_),
    .QN(_00544_),
    .RESETN(net854),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[133]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02895_),
    .QN(_00576_),
    .RESETN(net855),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[134]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02896_),
    .QN(_00606_),
    .RESETN(net856),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[135]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02897_),
    .QN(_00636_),
    .RESETN(net857),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[136]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02898_),
    .QN(_00666_),
    .RESETN(net858),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[137]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_02899_),
    .QN(_00696_),
    .RESETN(net859),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[138]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02900_),
    .QN(_00726_),
    .RESETN(net860),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[139]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_02901_),
    .QN(_00756_),
    .RESETN(net861),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_02902_),
    .QN(_01810_),
    .RESETN(net862),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[140]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_02903_),
    .QN(_00452_),
    .RESETN(net863),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[141]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02904_),
    .QN(_00827_),
    .RESETN(net864),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[142]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02905_),
    .QN(_00860_),
    .RESETN(net865),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[143]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02906_),
    .QN(_00893_),
    .RESETN(net866),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[144]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_02907_),
    .QN(_00926_),
    .RESETN(net867),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[145]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02908_),
    .QN(_00959_),
    .RESETN(net868),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[146]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02909_),
    .QN(_00992_),
    .RESETN(net869),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[147]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02910_),
    .QN(_01025_),
    .RESETN(net870),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[148]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_02911_),
    .QN(_01058_),
    .RESETN(net871),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[149]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02912_),
    .QN(_01091_),
    .RESETN(net872),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_02913_),
    .QN(_01809_),
    .RESETN(net873),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[150]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02914_),
    .QN(_01124_),
    .RESETN(net874),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[151]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02915_),
    .QN(_01157_),
    .RESETN(net875),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[152]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02916_),
    .QN(_01190_),
    .RESETN(net876),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[153]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02917_),
    .QN(_01223_),
    .RESETN(net877),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[154]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02918_),
    .QN(_01256_),
    .RESETN(net878),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[155]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02919_),
    .QN(_01289_),
    .RESETN(net879),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[156]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02920_),
    .QN(_01322_),
    .RESETN(net880),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[157]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_02921_),
    .QN(_01355_),
    .RESETN(net881),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[158]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02922_),
    .QN(_01388_),
    .RESETN(net882),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[159]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_02923_),
    .QN(_01421_),
    .RESETN(net883),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_02924_),
    .QN(_01808_),
    .RESETN(net884),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[160]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02925_),
    .QN(_00420_),
    .RESETN(net885),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[161]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_02926_),
    .QN(_00373_),
    .RESETN(net886),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[162]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02927_),
    .QN(_00484_),
    .RESETN(net887),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[163]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02928_),
    .QN(_00515_),
    .RESETN(net888),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[164]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_02929_),
    .QN(_00545_),
    .RESETN(net889),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[165]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02930_),
    .QN(_00577_),
    .RESETN(net890),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[166]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_02931_),
    .QN(_00607_),
    .RESETN(net891),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[167]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02932_),
    .QN(_00637_),
    .RESETN(net892),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[168]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02933_),
    .QN(_00667_),
    .RESETN(net893),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[169]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02934_),
    .QN(_00697_),
    .RESETN(net894),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_02935_),
    .QN(_01807_),
    .RESETN(net895),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[170]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02936_),
    .QN(_00727_),
    .RESETN(net896),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[171]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02937_),
    .QN(_00757_),
    .RESETN(net897),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[172]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_02938_),
    .QN(_00453_),
    .RESETN(net898),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[173]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02939_),
    .QN(_00828_),
    .RESETN(net899),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[174]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02940_),
    .QN(_00861_),
    .RESETN(net900),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[175]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_02941_),
    .QN(_00894_),
    .RESETN(net901),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[176]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02942_),
    .QN(_00927_),
    .RESETN(net902),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[177]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_02943_),
    .QN(_00960_),
    .RESETN(net903),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[178]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02944_),
    .QN(_00993_),
    .RESETN(net904),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[179]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02945_),
    .QN(_01026_),
    .RESETN(net905),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_02946_),
    .QN(_01806_),
    .RESETN(net906),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[180]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_02947_),
    .QN(_01059_),
    .RESETN(net907),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[181]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_02948_),
    .QN(_01092_),
    .RESETN(net908),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[182]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_02949_),
    .QN(_01125_),
    .RESETN(net909),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[183]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02950_),
    .QN(_01158_),
    .RESETN(net910),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[184]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02951_),
    .QN(_01191_),
    .RESETN(net911),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[185]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02952_),
    .QN(_01224_),
    .RESETN(net912),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[186]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02953_),
    .QN(_01257_),
    .RESETN(net913),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[187]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02954_),
    .QN(_01290_),
    .RESETN(net914),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[188]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02955_),
    .QN(_01323_),
    .RESETN(net915),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[189]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02956_),
    .QN(_01356_),
    .RESETN(net916),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_02957_),
    .QN(_01805_),
    .RESETN(net917),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[190]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02958_),
    .QN(_01389_),
    .RESETN(net918),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[191]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_02959_),
    .QN(_01422_),
    .RESETN(net919),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[192]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02960_),
    .QN(_00421_),
    .RESETN(net920),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[193]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02961_),
    .QN(_00374_),
    .RESETN(net921),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[194]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02962_),
    .QN(_00485_),
    .RESETN(net922),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[195]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02963_),
    .QN(_00516_),
    .RESETN(net923),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[196]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02964_),
    .QN(_00546_),
    .RESETN(net924),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[197]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_02965_),
    .QN(_00578_),
    .RESETN(net925),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[198]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02966_),
    .QN(_00608_),
    .RESETN(net926),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[199]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02967_),
    .QN(_00638_),
    .RESETN(net927),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_02968_),
    .QN(_01804_),
    .RESETN(net928),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_02969_),
    .QN(_01803_),
    .RESETN(net929),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[200]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02970_),
    .QN(_00668_),
    .RESETN(net930),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[201]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02971_),
    .QN(_00698_),
    .RESETN(net931),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[202]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02972_),
    .QN(_00728_),
    .RESETN(net932),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[203]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02973_),
    .QN(_00758_),
    .RESETN(net933),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[204]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_02974_),
    .QN(_00454_),
    .RESETN(net934),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[205]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02975_),
    .QN(_00829_),
    .RESETN(net935),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[206]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02976_),
    .QN(_00862_),
    .RESETN(net936),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[207]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02977_),
    .QN(_00895_),
    .RESETN(net937),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[208]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02978_),
    .QN(_00928_),
    .RESETN(net938),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[209]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_02979_),
    .QN(_00961_),
    .RESETN(net939),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_02980_),
    .QN(_01802_),
    .RESETN(net940),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[210]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_02981_),
    .QN(_00994_),
    .RESETN(net941),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[211]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02982_),
    .QN(_01027_),
    .RESETN(net942),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[212]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02983_),
    .QN(_01060_),
    .RESETN(net943),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[213]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02984_),
    .QN(_01093_),
    .RESETN(net944),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[214]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_02985_),
    .QN(_01126_),
    .RESETN(net945),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[215]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_02986_),
    .QN(_01159_),
    .RESETN(net946),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[216]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02987_),
    .QN(_01192_),
    .RESETN(net947),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[217]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_02988_),
    .QN(_01225_),
    .RESETN(net948),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[218]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02989_),
    .QN(_01258_),
    .RESETN(net949),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[219]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02990_),
    .QN(_01291_),
    .RESETN(net950),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_02991_),
    .QN(_01801_),
    .RESETN(net951),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[220]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02992_),
    .QN(_01324_),
    .RESETN(net952),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[221]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_02993_),
    .QN(_01357_),
    .RESETN(net953),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[222]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_02994_),
    .QN(_01390_),
    .RESETN(net954),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[223]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_02995_),
    .QN(_01423_),
    .RESETN(net955),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[224]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_02996_),
    .QN(_00422_),
    .RESETN(net956),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[225]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_02997_),
    .QN(_00375_),
    .RESETN(net957),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[226]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_02998_),
    .QN(_00486_),
    .RESETN(net958),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[227]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_02999_),
    .QN(_00517_),
    .RESETN(net959),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[228]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03000_),
    .QN(_00547_),
    .RESETN(net960),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[229]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03001_),
    .QN(_00579_),
    .RESETN(net961),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03002_),
    .QN(_01800_),
    .RESETN(net962),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[230]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03003_),
    .QN(_00609_),
    .RESETN(net963),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[231]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03004_),
    .QN(_00639_),
    .RESETN(net964),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[232]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03005_),
    .QN(_00669_),
    .RESETN(net965),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[233]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03006_),
    .QN(_00699_),
    .RESETN(net966),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[234]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03007_),
    .QN(_00729_),
    .RESETN(net967),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[235]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03008_),
    .QN(_00759_),
    .RESETN(net968),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[236]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03009_),
    .QN(_00455_),
    .RESETN(net969),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[237]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03010_),
    .QN(_00830_),
    .RESETN(net970),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[238]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03011_),
    .QN(_00863_),
    .RESETN(net971),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[239]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03012_),
    .QN(_00896_),
    .RESETN(net972),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03013_),
    .QN(_01799_),
    .RESETN(net973),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[240]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03014_),
    .QN(_00929_),
    .RESETN(net974),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[241]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03015_),
    .QN(_00962_),
    .RESETN(net975),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[242]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03016_),
    .QN(_00995_),
    .RESETN(net976),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[243]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03017_),
    .QN(_01028_),
    .RESETN(net977),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[244]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03018_),
    .QN(_01061_),
    .RESETN(net978),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[245]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03019_),
    .QN(_01094_),
    .RESETN(net979),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[246]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03020_),
    .QN(_01127_),
    .RESETN(net980),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[247]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03021_),
    .QN(_01160_),
    .RESETN(net981),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[248]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03022_),
    .QN(_01193_),
    .RESETN(net982),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[249]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03023_),
    .QN(_01226_),
    .RESETN(net983),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03024_),
    .QN(_01798_),
    .RESETN(net984),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[250]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03025_),
    .QN(_01259_),
    .RESETN(net985),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[251]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03026_),
    .QN(_01292_),
    .RESETN(net986),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[252]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03027_),
    .QN(_01325_),
    .RESETN(net987),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[253]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03028_),
    .QN(_01358_),
    .RESETN(net988),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[254]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03029_),
    .QN(_01391_),
    .RESETN(net989),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[255]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03030_),
    .QN(_01424_),
    .RESETN(net990),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[256]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03031_),
    .QN(_00423_),
    .RESETN(net991),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[257]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03032_),
    .QN(_00376_),
    .RESETN(net992),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[258]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03033_),
    .QN(_00487_),
    .RESETN(net993),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[259]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03034_),
    .QN(_00518_),
    .RESETN(net994),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03035_),
    .QN(_01797_),
    .RESETN(net995),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[260]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03036_),
    .QN(_00548_),
    .RESETN(net996),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[261]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03037_),
    .QN(_00580_),
    .RESETN(net997),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[262]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03038_),
    .QN(_00610_),
    .RESETN(net998),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[263]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03039_),
    .QN(_00640_),
    .RESETN(net999),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[264]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03040_),
    .QN(_00670_),
    .RESETN(net1000),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[265]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03041_),
    .QN(_00700_),
    .RESETN(net1001),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[266]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03042_),
    .QN(_00730_),
    .RESETN(net1002),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[267]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03043_),
    .QN(_00760_),
    .RESETN(net1003),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[268]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03044_),
    .QN(_00456_),
    .RESETN(net1004),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[269]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03045_),
    .QN(_00831_),
    .RESETN(net1005),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03046_),
    .QN(_01796_),
    .RESETN(net1006),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[270]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03047_),
    .QN(_00864_),
    .RESETN(net1007),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[271]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03048_),
    .QN(_00897_),
    .RESETN(net1008),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[272]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03049_),
    .QN(_00930_),
    .RESETN(net1009),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[273]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03050_),
    .QN(_00963_),
    .RESETN(net1010),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[274]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03051_),
    .QN(_00996_),
    .RESETN(net1011),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[275]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03052_),
    .QN(_01029_),
    .RESETN(net1012),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[276]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03053_),
    .QN(_01062_),
    .RESETN(net1013),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[277]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03054_),
    .QN(_01095_),
    .RESETN(net1014),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[278]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03055_),
    .QN(_01128_),
    .RESETN(net1015),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[279]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03056_),
    .QN(_01161_),
    .RESETN(net1016),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03057_),
    .QN(_01795_),
    .RESETN(net1017),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[280]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03058_),
    .QN(_01194_),
    .RESETN(net1018),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[281]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03059_),
    .QN(_01227_),
    .RESETN(net1019),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[282]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03060_),
    .QN(_01260_),
    .RESETN(net1020),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[283]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03061_),
    .QN(_01293_),
    .RESETN(net1021),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[284]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03062_),
    .QN(_01326_),
    .RESETN(net1022),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[285]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03063_),
    .QN(_01359_),
    .RESETN(net1023),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[286]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03064_),
    .QN(_01392_),
    .RESETN(net1024),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[287]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03065_),
    .QN(_01425_),
    .RESETN(net1025),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[288]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03066_),
    .QN(_00424_),
    .RESETN(net1026),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[289]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03067_),
    .QN(_00377_),
    .RESETN(net1027),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03068_),
    .QN(_01794_),
    .RESETN(net1028),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[290]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03069_),
    .QN(_00488_),
    .RESETN(net1029),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[291]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03070_),
    .QN(_00519_),
    .RESETN(net1030),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[292]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03071_),
    .QN(_00549_),
    .RESETN(net1031),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[293]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03072_),
    .QN(_00581_),
    .RESETN(net1032),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[294]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03073_),
    .QN(_00611_),
    .RESETN(net1033),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[295]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03074_),
    .QN(_00641_),
    .RESETN(net1034),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[296]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03075_),
    .QN(_00671_),
    .RESETN(net1035),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[297]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03076_),
    .QN(_00701_),
    .RESETN(net1036),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[298]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03077_),
    .QN(_00731_),
    .RESETN(net1037),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[299]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03078_),
    .QN(_00761_),
    .RESETN(net1038),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03079_),
    .QN(_01793_),
    .RESETN(net1039),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03080_),
    .QN(_01792_),
    .RESETN(net1040),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[300]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03081_),
    .QN(_00457_),
    .RESETN(net1041),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[301]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03082_),
    .QN(_00832_),
    .RESETN(net1042),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[302]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03083_),
    .QN(_00865_),
    .RESETN(net1043),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[303]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03084_),
    .QN(_00898_),
    .RESETN(net1044),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[304]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03085_),
    .QN(_00931_),
    .RESETN(net1045),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[305]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03086_),
    .QN(_00964_),
    .RESETN(net1046),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[306]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03087_),
    .QN(_00997_),
    .RESETN(net1047),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[307]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03088_),
    .QN(_01030_),
    .RESETN(net1048),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[308]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03089_),
    .QN(_01063_),
    .RESETN(net1049),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[309]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03090_),
    .QN(_01096_),
    .RESETN(net1050),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03091_),
    .QN(_01791_),
    .RESETN(net1051),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[310]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03092_),
    .QN(_01129_),
    .RESETN(net1052),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[311]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03093_),
    .QN(_01162_),
    .RESETN(net1053),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[312]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03094_),
    .QN(_01195_),
    .RESETN(net1054),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[313]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03095_),
    .QN(_01228_),
    .RESETN(net1055),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[314]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03096_),
    .QN(_01261_),
    .RESETN(net1056),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[315]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03097_),
    .QN(_01294_),
    .RESETN(net1057),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[316]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03098_),
    .QN(_01327_),
    .RESETN(net1058),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[317]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03099_),
    .QN(_01360_),
    .RESETN(net1059),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[318]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03100_),
    .QN(_01393_),
    .RESETN(net1060),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[319]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03101_),
    .QN(_01426_),
    .RESETN(net1061),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03102_),
    .QN(_01790_),
    .RESETN(net1062),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[320]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03103_),
    .QN(_00425_),
    .RESETN(net1063),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[321]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03104_),
    .QN(_00378_),
    .RESETN(net1064),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[322]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03105_),
    .QN(_00489_),
    .RESETN(net1065),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[323]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03106_),
    .QN(_00520_),
    .RESETN(net1066),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[324]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03107_),
    .QN(_00550_),
    .RESETN(net1067),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[325]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03108_),
    .QN(_00582_),
    .RESETN(net1068),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[326]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03109_),
    .QN(_00612_),
    .RESETN(net1069),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[327]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03110_),
    .QN(_00642_),
    .RESETN(net1070),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[328]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03111_),
    .QN(_00672_),
    .RESETN(net1071),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[329]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03112_),
    .QN(_00702_),
    .RESETN(net1072),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[32]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03113_),
    .QN(_00416_),
    .RESETN(net1073),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[330]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03114_),
    .QN(_00732_),
    .RESETN(net1074),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[331]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03115_),
    .QN(_00762_),
    .RESETN(net1075),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[332]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03116_),
    .QN(_00458_),
    .RESETN(net1076),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[333]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03117_),
    .QN(_00833_),
    .RESETN(net1077),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[334]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03118_),
    .QN(_00866_),
    .RESETN(net1078),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[335]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03119_),
    .QN(_00899_),
    .RESETN(net1079),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[336]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03120_),
    .QN(_00932_),
    .RESETN(net1080),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[337]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03121_),
    .QN(_00965_),
    .RESETN(net1081),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[338]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03122_),
    .QN(_00998_),
    .RESETN(net1082),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[339]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03123_),
    .QN(_01031_),
    .RESETN(net1083),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[33]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03124_),
    .QN(_00369_),
    .RESETN(net1084),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[340]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03125_),
    .QN(_01064_),
    .RESETN(net1085),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[341]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03126_),
    .QN(_01097_),
    .RESETN(net1086),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[342]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03127_),
    .QN(_01130_),
    .RESETN(net1087),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[343]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03128_),
    .QN(_01163_),
    .RESETN(net1088),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[344]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03129_),
    .QN(_01196_),
    .RESETN(net1089),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[345]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03130_),
    .QN(_01229_),
    .RESETN(net1090),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[346]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03131_),
    .QN(_01262_),
    .RESETN(net1091),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[347]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03132_),
    .QN(_01295_),
    .RESETN(net1092),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[348]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03133_),
    .QN(_01328_),
    .RESETN(net1093),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[349]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03134_),
    .QN(_01361_),
    .RESETN(net1094),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03135_),
    .QN(_00480_),
    .RESETN(net1095),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[350]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03136_),
    .QN(_01394_),
    .RESETN(net1096),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[351]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03137_),
    .QN(_01427_),
    .RESETN(net1097),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[352]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03138_),
    .QN(_00426_),
    .RESETN(net1098),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[353]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03139_),
    .QN(_00379_),
    .RESETN(net1099),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[354]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03140_),
    .QN(_00490_),
    .RESETN(net1100),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[355]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03141_),
    .QN(_00521_),
    .RESETN(net1101),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[356]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03142_),
    .QN(_00551_),
    .RESETN(net1102),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[357]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03143_),
    .QN(_00583_),
    .RESETN(net1103),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[358]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03144_),
    .QN(_00613_),
    .RESETN(net1104),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[359]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03145_),
    .QN(_00643_),
    .RESETN(net1105),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_03146_),
    .QN(_00511_),
    .RESETN(net1106),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[360]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03147_),
    .QN(_00673_),
    .RESETN(net1107),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[361]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03148_),
    .QN(_00703_),
    .RESETN(net1108),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[362]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03149_),
    .QN(_00733_),
    .RESETN(net1109),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[363]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03150_),
    .QN(_00763_),
    .RESETN(net1110),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[364]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03151_),
    .QN(_00459_),
    .RESETN(net1111),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[365]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03152_),
    .QN(_00834_),
    .RESETN(net1112),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[366]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03153_),
    .QN(_00867_),
    .RESETN(net1113),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[367]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03154_),
    .QN(_00900_),
    .RESETN(net1114),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[368]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03155_),
    .QN(_00933_),
    .RESETN(net1115),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[369]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03156_),
    .QN(_00966_),
    .RESETN(net1116),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03157_),
    .QN(_00541_),
    .RESETN(net1117),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[370]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03158_),
    .QN(_00999_),
    .RESETN(net1118),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[371]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03159_),
    .QN(_01032_),
    .RESETN(net1119),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[372]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03160_),
    .QN(_01065_),
    .RESETN(net1120),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[373]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03161_),
    .QN(_01098_),
    .RESETN(net1121),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[374]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03162_),
    .QN(_01131_),
    .RESETN(net1122),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[375]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03163_),
    .QN(_01164_),
    .RESETN(net1123),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[376]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03164_),
    .QN(_01197_),
    .RESETN(net1124),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[377]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03165_),
    .QN(_01230_),
    .RESETN(net1125),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[378]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03166_),
    .QN(_01263_),
    .RESETN(net1126),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[379]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03167_),
    .QN(_01296_),
    .RESETN(net1127),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03168_),
    .QN(_00573_),
    .RESETN(net1128),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[380]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03169_),
    .QN(_01329_),
    .RESETN(net1129),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[381]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03170_),
    .QN(_01362_),
    .RESETN(net1130),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[382]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03171_),
    .QN(_01395_),
    .RESETN(net1131),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[383]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03172_),
    .QN(_01428_),
    .RESETN(net1132),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[384]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03173_),
    .QN(_00427_),
    .RESETN(net1133),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[385]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03174_),
    .QN(_00380_),
    .RESETN(net1134),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[386]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03175_),
    .QN(_00491_),
    .RESETN(net1135),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[387]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03176_),
    .QN(_00522_),
    .RESETN(net1136),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[388]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03177_),
    .QN(_00552_),
    .RESETN(net1137),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[389]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03178_),
    .QN(_00584_),
    .RESETN(net1138),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03179_),
    .QN(_00603_),
    .RESETN(net1139),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[390]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03180_),
    .QN(_00614_),
    .RESETN(net1140),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[391]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03181_),
    .QN(_00644_),
    .RESETN(net1141),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[392]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03182_),
    .QN(_00674_),
    .RESETN(net1142),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[393]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03183_),
    .QN(_00704_),
    .RESETN(net1143),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[394]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03184_),
    .QN(_00734_),
    .RESETN(net1144),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[395]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03185_),
    .QN(_00764_),
    .RESETN(net1145),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[396]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03186_),
    .QN(_00460_),
    .RESETN(net1146),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[397]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03187_),
    .QN(_00835_),
    .RESETN(net1147),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[398]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03188_),
    .QN(_00868_),
    .RESETN(net1148),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[399]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03189_),
    .QN(_00901_),
    .RESETN(net1149),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03190_),
    .QN(_00633_),
    .RESETN(net1150),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_03191_),
    .QN(_01789_),
    .RESETN(net1151),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[400]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03192_),
    .QN(_00934_),
    .RESETN(net1152),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[401]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03193_),
    .QN(_00967_),
    .RESETN(net1153),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[402]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03194_),
    .QN(_01000_),
    .RESETN(net1154),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[403]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03195_),
    .QN(_01033_),
    .RESETN(net1155),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[404]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03196_),
    .QN(_01066_),
    .RESETN(net1156),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[405]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03197_),
    .QN(_01099_),
    .RESETN(net1157),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[406]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03198_),
    .QN(_01132_),
    .RESETN(net1158),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[407]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03199_),
    .QN(_01165_),
    .RESETN(net1159),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[408]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03200_),
    .QN(_01198_),
    .RESETN(net1160),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[409]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03201_),
    .QN(_01231_),
    .RESETN(net1161),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03202_),
    .QN(_00663_),
    .RESETN(net1162),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[410]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03203_),
    .QN(_01264_),
    .RESETN(net1163),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[411]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03204_),
    .QN(_01297_),
    .RESETN(net1164),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[412]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03205_),
    .QN(_01330_),
    .RESETN(net1165),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[413]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03206_),
    .QN(_01363_),
    .RESETN(net1166),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[414]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03207_),
    .QN(_01396_),
    .RESETN(net1167),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[415]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03208_),
    .QN(_01429_),
    .RESETN(net1168),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[416]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03209_),
    .QN(_00428_),
    .RESETN(net1169),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[417]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03210_),
    .QN(_00381_),
    .RESETN(net1170),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[418]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03211_),
    .QN(_00492_),
    .RESETN(net1171),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[419]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03212_),
    .QN(_00523_),
    .RESETN(net1172),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03213_),
    .QN(_00693_),
    .RESETN(net1173),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[420]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03214_),
    .QN(_00553_),
    .RESETN(net1174),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[421]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03215_),
    .QN(_00585_),
    .RESETN(net1175),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[422]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03216_),
    .QN(_00615_),
    .RESETN(net1176),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[423]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03217_),
    .QN(_00645_),
    .RESETN(net1177),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[424]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03218_),
    .QN(_00675_),
    .RESETN(net1178),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[425]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03219_),
    .QN(_00705_),
    .RESETN(net1179),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[426]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk_i_regs),
    .D(_03220_),
    .QN(_00735_),
    .RESETN(net1180),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[427]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03221_),
    .QN(_00765_),
    .RESETN(net1181),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[428]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03222_),
    .QN(_00461_),
    .RESETN(net1182),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[429]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03223_),
    .QN(_00836_),
    .RESETN(net1183),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03224_),
    .QN(_00723_),
    .RESETN(net1184),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[430]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03225_),
    .QN(_00869_),
    .RESETN(net1185),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[431]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03226_),
    .QN(_00902_),
    .RESETN(net1186),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[432]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03227_),
    .QN(_00935_),
    .RESETN(net1187),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[433]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03228_),
    .QN(_00968_),
    .RESETN(net1188),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[434]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03229_),
    .QN(_01001_),
    .RESETN(net1189),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[435]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03230_),
    .QN(_01034_),
    .RESETN(net1190),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[436]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03231_),
    .QN(_01067_),
    .RESETN(net1191),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[437]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03232_),
    .QN(_01100_),
    .RESETN(net1192),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[438]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03233_),
    .QN(_01133_),
    .RESETN(net1193),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[439]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk_i_regs),
    .D(_03234_),
    .QN(_01166_),
    .RESETN(net1194),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03235_),
    .QN(_00753_),
    .RESETN(net1195),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[440]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03236_),
    .QN(_01199_),
    .RESETN(net1196),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[441]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03237_),
    .QN(_01232_),
    .RESETN(net1197),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[442]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03238_),
    .QN(_01265_),
    .RESETN(net1198),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[443]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03239_),
    .QN(_01298_),
    .RESETN(net1199),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[444]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk_i_regs),
    .D(_03240_),
    .QN(_01331_),
    .RESETN(net1200),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[445]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03241_),
    .QN(_01364_),
    .RESETN(net1201),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[446]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03242_),
    .QN(_01397_),
    .RESETN(net1202),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[447]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03243_),
    .QN(_01430_),
    .RESETN(net1203),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[448]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03244_),
    .QN(_00429_),
    .RESETN(net1204),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[449]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk_i_regs),
    .D(_03245_),
    .QN(_00382_),
    .RESETN(net1205),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03246_),
    .QN(_00449_),
    .RESETN(net1206),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[450]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03247_),
    .QN(_00493_),
    .RESETN(net1207),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[451]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03248_),
    .QN(_00524_),
    .RESETN(net1208),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[452]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03249_),
    .QN(_00554_),
    .RESETN(net1209),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[453]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03250_),
    .QN(_00586_),
    .RESETN(net1210),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[454]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03251_),
    .QN(_00616_),
    .RESETN(net1211),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[455]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03252_),
    .QN(_00646_),
    .RESETN(net1212),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[456]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03253_),
    .QN(_00676_),
    .RESETN(net1213),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[457]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03254_),
    .QN(_00706_),
    .RESETN(net1214),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[458]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03255_),
    .QN(_00736_),
    .RESETN(net1215),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[459]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk_i_regs),
    .D(_03256_),
    .QN(_00766_),
    .RESETN(net1216),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03257_),
    .QN(_00824_),
    .RESETN(net1217),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[460]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03258_),
    .QN(_00462_),
    .RESETN(net1218),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[461]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03259_),
    .QN(_00837_),
    .RESETN(net1219),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[462]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03260_),
    .QN(_00870_),
    .RESETN(net1220),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[463]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03261_),
    .QN(_00903_),
    .RESETN(net1221),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[464]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03262_),
    .QN(_00936_),
    .RESETN(net1222),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[465]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03263_),
    .QN(_00969_),
    .RESETN(net1223),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[466]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03264_),
    .QN(_01002_),
    .RESETN(net1224),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[467]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03265_),
    .QN(_01035_),
    .RESETN(net1225),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[468]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03266_),
    .QN(_01068_),
    .RESETN(net1226),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[469]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03267_),
    .QN(_01101_),
    .RESETN(net1227),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03268_),
    .QN(_00857_),
    .RESETN(net1228),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[470]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03269_),
    .QN(_01134_),
    .RESETN(net1229),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[471]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk_i_regs),
    .D(_03270_),
    .QN(_01167_),
    .RESETN(net1230),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[472]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03271_),
    .QN(_01200_),
    .RESETN(net1231),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[473]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk_i_regs),
    .D(_03272_),
    .QN(_01233_),
    .RESETN(net1232),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[474]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03273_),
    .QN(_01266_),
    .RESETN(net1233),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[475]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk_i_regs),
    .D(_03274_),
    .QN(_01299_),
    .RESETN(net1234),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[476]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03275_),
    .QN(_01332_),
    .RESETN(net1235),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[477]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03276_),
    .QN(_01365_),
    .RESETN(net1236),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[478]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03277_),
    .QN(_01398_),
    .RESETN(net1237),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[479]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03278_),
    .QN(_01431_),
    .RESETN(net1238),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03279_),
    .QN(_00890_),
    .RESETN(net1239),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[480]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03280_),
    .QN(_00430_),
    .RESETN(net1240),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[481]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03281_),
    .QN(_00383_),
    .RESETN(net1241),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[482]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03282_),
    .QN(_00494_),
    .RESETN(net1242),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[483]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03283_),
    .QN(_00525_),
    .RESETN(net1243),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[484]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_03284_),
    .QN(_00555_),
    .RESETN(net1244),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[485]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03285_),
    .QN(_00587_),
    .RESETN(net1245),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[486]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03286_),
    .QN(_00617_),
    .RESETN(net1246),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[487]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03287_),
    .QN(_00647_),
    .RESETN(net1247),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[488]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03288_),
    .QN(_00677_),
    .RESETN(net1248),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[489]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03289_),
    .QN(_00707_),
    .RESETN(net1249),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03290_),
    .QN(_00923_),
    .RESETN(net1250),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[490]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03291_),
    .QN(_00737_),
    .RESETN(net1251),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[491]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03292_),
    .QN(_00767_),
    .RESETN(net1252),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[492]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03293_),
    .QN(_00463_),
    .RESETN(net1253),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[493]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03294_),
    .QN(_00838_),
    .RESETN(net1254),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[494]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03295_),
    .QN(_00871_),
    .RESETN(net1255),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[495]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03296_),
    .QN(_00904_),
    .RESETN(net1256),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[496]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03297_),
    .QN(_00937_),
    .RESETN(net1257),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[497]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03298_),
    .QN(_00970_),
    .RESETN(net1258),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[498]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03299_),
    .QN(_01003_),
    .RESETN(net1259),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[499]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03300_),
    .QN(_01036_),
    .RESETN(net1260),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03301_),
    .QN(_00956_),
    .RESETN(net1261),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03302_),
    .QN(_01788_),
    .RESETN(net1262),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[500]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03303_),
    .QN(_01069_),
    .RESETN(net1263),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[501]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03304_),
    .QN(_01102_),
    .RESETN(net1264),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[502]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03305_),
    .QN(_01135_),
    .RESETN(net1265),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[503]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03306_),
    .QN(_01168_),
    .RESETN(net1266),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[504]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03307_),
    .QN(_01201_),
    .RESETN(net1267),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[505]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03308_),
    .QN(_01234_),
    .RESETN(net1268),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[506]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03309_),
    .QN(_01267_),
    .RESETN(net1269),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[507]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03310_),
    .QN(_01300_),
    .RESETN(net1270),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[508]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03311_),
    .QN(_01333_),
    .RESETN(net1271),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[509]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03312_),
    .QN(_01366_),
    .RESETN(net1272),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03313_),
    .QN(_00989_),
    .RESETN(net1273),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[510]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03314_),
    .QN(_01399_),
    .RESETN(net1274),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[511]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03315_),
    .QN(_01432_),
    .RESETN(net1275),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[512]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03316_),
    .QN(_00431_),
    .RESETN(net1276),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[513]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03317_),
    .QN(_00384_),
    .RESETN(net1277),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[514]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03318_),
    .QN(_00495_),
    .RESETN(net1278),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[515]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03319_),
    .QN(_00526_),
    .RESETN(net1279),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[516]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_03320_),
    .QN(_00556_),
    .RESETN(net1280),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[517]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03321_),
    .QN(_00588_),
    .RESETN(net1281),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[518]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03322_),
    .QN(_00618_),
    .RESETN(net1282),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[519]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03323_),
    .QN(_00648_),
    .RESETN(net1283),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03324_),
    .QN(_01022_),
    .RESETN(net1284),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[520]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03325_),
    .QN(_00678_),
    .RESETN(net1285),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[521]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03326_),
    .QN(_00708_),
    .RESETN(net1286),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[522]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03327_),
    .QN(_00738_),
    .RESETN(net1287),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[523]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03328_),
    .QN(_00768_),
    .RESETN(net1288),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[524]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03329_),
    .QN(_00464_),
    .RESETN(net1289),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[525]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk_i_regs),
    .D(_03330_),
    .QN(_00839_),
    .RESETN(net1290),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[526]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03331_),
    .QN(_00872_),
    .RESETN(net1291),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[527]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03332_),
    .QN(_00905_),
    .RESETN(net1292),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[528]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03333_),
    .QN(_00938_),
    .RESETN(net1293),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[529]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03334_),
    .QN(_00971_),
    .RESETN(net1294),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03335_),
    .QN(_01055_),
    .RESETN(net1295),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[530]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk_i_regs),
    .D(_03336_),
    .QN(_01004_),
    .RESETN(net1296),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[531]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03337_),
    .QN(_01037_),
    .RESETN(net1297),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[532]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03338_),
    .QN(_01070_),
    .RESETN(net1298),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[533]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03339_),
    .QN(_01103_),
    .RESETN(net1299),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[534]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03340_),
    .QN(_01136_),
    .RESETN(net1300),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[535]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03341_),
    .QN(_01169_),
    .RESETN(net1301),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[536]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03342_),
    .QN(_01202_),
    .RESETN(net1302),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[537]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk_i_regs),
    .D(_03343_),
    .QN(_01235_),
    .RESETN(net1303),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[538]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03344_),
    .QN(_01268_),
    .RESETN(net1304),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[539]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03345_),
    .QN(_01301_),
    .RESETN(net1305),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03346_),
    .QN(_01088_),
    .RESETN(net1306),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[540]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03347_),
    .QN(_01334_),
    .RESETN(net1307),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[541]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03348_),
    .QN(_01367_),
    .RESETN(net1308),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[542]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03349_),
    .QN(_01400_),
    .RESETN(net1309),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[543]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03350_),
    .QN(_01433_),
    .RESETN(net1310),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[544]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03351_),
    .QN(_00432_),
    .RESETN(net1311),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[545]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03352_),
    .QN(_00385_),
    .RESETN(net1312),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[546]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03353_),
    .QN(_00496_),
    .RESETN(net1313),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[547]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03354_),
    .QN(_00527_),
    .RESETN(net1314),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[548]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03355_),
    .QN(_00557_),
    .RESETN(net1315),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[549]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03356_),
    .QN(_00589_),
    .RESETN(net1316),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03357_),
    .QN(_01121_),
    .RESETN(net1317),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[550]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03358_),
    .QN(_00619_),
    .RESETN(net1318),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[551]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03359_),
    .QN(_00649_),
    .RESETN(net1319),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[552]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03360_),
    .QN(_00679_),
    .RESETN(net1320),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[553]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03361_),
    .QN(_00709_),
    .RESETN(net1321),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[554]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03362_),
    .QN(_00739_),
    .RESETN(net1322),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[555]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03363_),
    .QN(_00769_),
    .RESETN(net1323),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[556]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03364_),
    .QN(_00465_),
    .RESETN(net1324),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[557]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03365_),
    .QN(_00840_),
    .RESETN(net1325),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[558]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03366_),
    .QN(_00873_),
    .RESETN(net1326),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[559]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03367_),
    .QN(_00906_),
    .RESETN(net1327),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03368_),
    .QN(_01154_),
    .RESETN(net1328),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[560]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03369_),
    .QN(_00939_),
    .RESETN(net1329),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[561]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03370_),
    .QN(_00972_),
    .RESETN(net1330),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[562]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03371_),
    .QN(_01005_),
    .RESETN(net1331),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[563]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03372_),
    .QN(_01038_),
    .RESETN(net1332),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[564]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03373_),
    .QN(_01071_),
    .RESETN(net1333),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[565]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03374_),
    .QN(_01104_),
    .RESETN(net1334),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[566]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03375_),
    .QN(_01137_),
    .RESETN(net1335),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[567]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03376_),
    .QN(_01170_),
    .RESETN(net1336),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[568]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03377_),
    .QN(_01203_),
    .RESETN(net1337),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[569]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03378_),
    .QN(_01236_),
    .RESETN(net1338),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03379_),
    .QN(_01187_),
    .RESETN(net1339),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[570]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03380_),
    .QN(_01269_),
    .RESETN(net1340),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[571]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03381_),
    .QN(_01302_),
    .RESETN(net1341),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[572]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03382_),
    .QN(_01335_),
    .RESETN(net1342),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[573]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03383_),
    .QN(_01368_),
    .RESETN(net1343),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[574]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03384_),
    .QN(_01401_),
    .RESETN(net1344),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[575]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03385_),
    .QN(_01434_),
    .RESETN(net1345),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[576]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03386_),
    .QN(_00433_),
    .RESETN(net1346),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[577]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03387_),
    .QN(_00386_),
    .RESETN(net1347),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[578]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03388_),
    .QN(_00497_),
    .RESETN(net1348),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[579]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03389_),
    .QN(_00528_),
    .RESETN(net1349),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03390_),
    .QN(_01220_),
    .RESETN(net1350),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[580]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03391_),
    .QN(_00558_),
    .RESETN(net1351),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[581]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03392_),
    .QN(_00590_),
    .RESETN(net1352),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[582]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03393_),
    .QN(_00620_),
    .RESETN(net1353),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[583]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03394_),
    .QN(_00650_),
    .RESETN(net1354),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[584]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03395_),
    .QN(_00680_),
    .RESETN(net1355),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[585]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03396_),
    .QN(_00710_),
    .RESETN(net1356),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[586]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03397_),
    .QN(_00740_),
    .RESETN(net1357),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[587]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03398_),
    .QN(_00770_),
    .RESETN(net1358),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[588]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03399_),
    .QN(_00466_),
    .RESETN(net1359),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[589]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03400_),
    .QN(_00841_),
    .RESETN(net1360),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03401_),
    .QN(_01253_),
    .RESETN(net1361),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[590]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03402_),
    .QN(_00874_),
    .RESETN(net1362),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[591]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03403_),
    .QN(_00907_),
    .RESETN(net1363),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[592]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03404_),
    .QN(_00940_),
    .RESETN(net1364),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[593]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03405_),
    .QN(_00973_),
    .RESETN(net1365),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[594]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03406_),
    .QN(_01006_),
    .RESETN(net1366),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[595]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03407_),
    .QN(_01039_),
    .RESETN(net1367),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[596]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03408_),
    .QN(_01072_),
    .RESETN(net1368),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[597]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03409_),
    .QN(_01105_),
    .RESETN(net1369),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[598]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03410_),
    .QN(_01138_),
    .RESETN(net1370),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[599]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03411_),
    .QN(_01171_),
    .RESETN(net1371),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03412_),
    .QN(_01286_),
    .RESETN(net1372),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03413_),
    .QN(_01787_),
    .RESETN(net1373),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[600]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03414_),
    .QN(_01204_),
    .RESETN(net1374),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[601]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03415_),
    .QN(_01237_),
    .RESETN(net1375),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[602]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03416_),
    .QN(_01270_),
    .RESETN(net1376),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[603]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03417_),
    .QN(_01303_),
    .RESETN(net1377),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[604]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03418_),
    .QN(_01336_),
    .RESETN(net1378),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[605]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03419_),
    .QN(_01369_),
    .RESETN(net1379),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[606]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03420_),
    .QN(_01402_),
    .RESETN(net1380),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[607]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03421_),
    .QN(_01435_),
    .RESETN(net1381),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[608]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03422_),
    .QN(_00434_),
    .RESETN(net1382),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[609]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03423_),
    .QN(_00387_),
    .RESETN(net1383),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03424_),
    .QN(_01319_),
    .RESETN(net1384),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[610]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03425_),
    .QN(_00498_),
    .RESETN(net1385),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[611]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03426_),
    .QN(_00529_),
    .RESETN(net1386),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[612]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03427_),
    .QN(_00559_),
    .RESETN(net1387),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[613]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03428_),
    .QN(_00591_),
    .RESETN(net1388),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[614]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03429_),
    .QN(_00621_),
    .RESETN(net1389),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[615]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03430_),
    .QN(_00651_),
    .RESETN(net1390),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[616]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03431_),
    .QN(_00681_),
    .RESETN(net1391),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[617]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03432_),
    .QN(_00711_),
    .RESETN(net1392),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[618]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03433_),
    .QN(_00741_),
    .RESETN(net1393),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[619]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03434_),
    .QN(_00771_),
    .RESETN(net1394),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03435_),
    .QN(_01352_),
    .RESETN(net1395),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[620]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03436_),
    .QN(_00467_),
    .RESETN(net1396),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[621]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03437_),
    .QN(_00842_),
    .RESETN(net1397),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[622]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03438_),
    .QN(_00875_),
    .RESETN(net1398),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[623]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03439_),
    .QN(_00908_),
    .RESETN(net1399),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[624]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03440_),
    .QN(_00941_),
    .RESETN(net1400),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[625]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03441_),
    .QN(_00974_),
    .RESETN(net1401),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[626]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03442_),
    .QN(_01007_),
    .RESETN(net1402),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[627]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03443_),
    .QN(_01040_),
    .RESETN(net1403),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[628]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03444_),
    .QN(_01073_),
    .RESETN(net1404),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[629]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03445_),
    .QN(_01106_),
    .RESETN(net1405),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03446_),
    .QN(_01385_),
    .RESETN(net1406),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[630]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03447_),
    .QN(_01139_),
    .RESETN(net1407),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[631]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03448_),
    .QN(_01172_),
    .RESETN(net1408),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[632]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03449_),
    .QN(_01205_),
    .RESETN(net1409),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[633]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03450_),
    .QN(_01238_),
    .RESETN(net1410),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[634]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03451_),
    .QN(_01271_),
    .RESETN(net1411),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[635]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03452_),
    .QN(_01304_),
    .RESETN(net1412),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[636]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03453_),
    .QN(_01337_),
    .RESETN(net1413),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[637]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03454_),
    .QN(_01370_),
    .RESETN(net1414),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[638]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03455_),
    .QN(_01403_),
    .RESETN(net1415),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[639]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03456_),
    .QN(_01436_),
    .RESETN(net1416),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03457_),
    .QN(_01418_),
    .RESETN(net1417),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[640]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03458_),
    .QN(_00435_),
    .RESETN(net1418),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[641]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03459_),
    .QN(_00388_),
    .RESETN(net1419),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[642]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03460_),
    .QN(_00499_),
    .RESETN(net1420),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[643]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03461_),
    .QN(_00530_),
    .RESETN(net1421),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[644]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03462_),
    .QN(_00560_),
    .RESETN(net1422),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[645]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03463_),
    .QN(_00592_),
    .RESETN(net1423),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[646]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03464_),
    .QN(_00622_),
    .RESETN(net1424),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[647]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03465_),
    .QN(_00652_),
    .RESETN(net1425),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[648]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03466_),
    .QN(_00682_),
    .RESETN(net1426),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[649]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03467_),
    .QN(_00712_),
    .RESETN(net1427),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[64]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03468_),
    .QN(_00417_),
    .RESETN(net1428),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[650]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03469_),
    .QN(_00742_),
    .RESETN(net1429),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[651]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03470_),
    .QN(_00772_),
    .RESETN(net1430),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[652]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03471_),
    .QN(_00468_),
    .RESETN(net1431),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[653]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03472_),
    .QN(_00843_),
    .RESETN(net1432),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[654]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03473_),
    .QN(_00876_),
    .RESETN(net1433),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[655]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03474_),
    .QN(_00909_),
    .RESETN(net1434),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[656]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03475_),
    .QN(_00942_),
    .RESETN(net1435),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[657]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03476_),
    .QN(_00975_),
    .RESETN(net1436),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[658]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03477_),
    .QN(_01008_),
    .RESETN(net1437),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[659]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03478_),
    .QN(_01041_),
    .RESETN(net1438),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[65]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03479_),
    .QN(_00370_),
    .RESETN(net1439),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[660]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03480_),
    .QN(_01074_),
    .RESETN(net1440),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[661]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03481_),
    .QN(_01107_),
    .RESETN(net1441),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[662]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03482_),
    .QN(_01140_),
    .RESETN(net1442),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[663]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03483_),
    .QN(_01173_),
    .RESETN(net1443),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[664]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03484_),
    .QN(_01206_),
    .RESETN(net1444),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[665]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03485_),
    .QN(_01239_),
    .RESETN(net1445),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[666]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03486_),
    .QN(_01272_),
    .RESETN(net1446),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[667]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03487_),
    .QN(_01305_),
    .RESETN(net1447),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[668]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03488_),
    .QN(_01338_),
    .RESETN(net1448),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[669]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03489_),
    .QN(_01371_),
    .RESETN(net1449),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[66]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03490_),
    .QN(_00481_),
    .RESETN(net1450),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[670]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03491_),
    .QN(_01404_),
    .RESETN(net1451),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[671]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03492_),
    .QN(_01437_),
    .RESETN(net1452),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[672]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03493_),
    .QN(_00436_),
    .RESETN(net1453),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[673]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03494_),
    .QN(_00389_),
    .RESETN(net1454),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[674]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03495_),
    .QN(_00500_),
    .RESETN(net1455),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[675]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03496_),
    .QN(_00531_),
    .RESETN(net1456),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[676]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03497_),
    .QN(_00561_),
    .RESETN(net1457),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[677]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk_i_regs),
    .D(_03498_),
    .QN(_00593_),
    .RESETN(net1458),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[678]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03499_),
    .QN(_00623_),
    .RESETN(net1459),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[679]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03500_),
    .QN(_00653_),
    .RESETN(net1460),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[67]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03501_),
    .QN(_00512_),
    .RESETN(net1461),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[680]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03502_),
    .QN(_00683_),
    .RESETN(net1462),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[681]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03503_),
    .QN(_00713_),
    .RESETN(net1463),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[682]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03504_),
    .QN(_00743_),
    .RESETN(net1464),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[683]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03505_),
    .QN(_00773_),
    .RESETN(net1465),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[684]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03506_),
    .QN(_00469_),
    .RESETN(net1466),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[685]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03507_),
    .QN(_00844_),
    .RESETN(net1467),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[686]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03508_),
    .QN(_00877_),
    .RESETN(net1468),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[687]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03509_),
    .QN(_00910_),
    .RESETN(net1469),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[688]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03510_),
    .QN(_00943_),
    .RESETN(net1470),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[689]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03511_),
    .QN(_00976_),
    .RESETN(net1471),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[68]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03512_),
    .QN(_00542_),
    .RESETN(net1472),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[690]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03513_),
    .QN(_01009_),
    .RESETN(net1473),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[691]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03514_),
    .QN(_01042_),
    .RESETN(net1474),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[692]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03515_),
    .QN(_01075_),
    .RESETN(net1475),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[693]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03516_),
    .QN(_01108_),
    .RESETN(net1476),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[694]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03517_),
    .QN(_01141_),
    .RESETN(net1477),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[695]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03518_),
    .QN(_01174_),
    .RESETN(net1478),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[696]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03519_),
    .QN(_01207_),
    .RESETN(net1479),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[697]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03520_),
    .QN(_01240_),
    .RESETN(net1480),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[698]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03521_),
    .QN(_01273_),
    .RESETN(net1481),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[699]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03522_),
    .QN(_01306_),
    .RESETN(net1482),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[69]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03523_),
    .QN(_00574_),
    .RESETN(net1483),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03524_),
    .QN(_01786_),
    .RESETN(net1484),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[700]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03525_),
    .QN(_01339_),
    .RESETN(net1485),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[701]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03526_),
    .QN(_01372_),
    .RESETN(net1486),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[702]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03527_),
    .QN(_01405_),
    .RESETN(net1487),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[703]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03528_),
    .QN(_01438_),
    .RESETN(net1488),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[704]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03529_),
    .QN(_00437_),
    .RESETN(net1489),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[705]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03530_),
    .QN(_00390_),
    .RESETN(net1490),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[706]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03531_),
    .QN(_00501_),
    .RESETN(net1491),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[707]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03532_),
    .QN(_00532_),
    .RESETN(net1492),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[708]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03533_),
    .QN(_00562_),
    .RESETN(net1493),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[709]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03534_),
    .QN(_00594_),
    .RESETN(net1494),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[70]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03535_),
    .QN(_00604_),
    .RESETN(net1495),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[710]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03536_),
    .QN(_00624_),
    .RESETN(net1496),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[711]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03537_),
    .QN(_00654_),
    .RESETN(net1497),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[712]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03538_),
    .QN(_00684_),
    .RESETN(net1498),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[713]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03539_),
    .QN(_00714_),
    .RESETN(net1499),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[714]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03540_),
    .QN(_00744_),
    .RESETN(net1500),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[715]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03541_),
    .QN(_00774_),
    .RESETN(net1501),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[716]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03542_),
    .QN(_00470_),
    .RESETN(net1502),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[717]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03543_),
    .QN(_00845_),
    .RESETN(net1503),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[718]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03544_),
    .QN(_00878_),
    .RESETN(net1504),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[719]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk_i_regs),
    .D(_03545_),
    .QN(_00911_),
    .RESETN(net1505),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[71]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03546_),
    .QN(_00634_),
    .RESETN(net1506),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[720]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03547_),
    .QN(_00944_),
    .RESETN(net1507),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[721]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03548_),
    .QN(_00977_),
    .RESETN(net1508),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[722]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03549_),
    .QN(_01010_),
    .RESETN(net1509),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[723]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03550_),
    .QN(_01043_),
    .RESETN(net1510),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[724]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03551_),
    .QN(_01076_),
    .RESETN(net1511),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[725]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03552_),
    .QN(_01109_),
    .RESETN(net1512),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[726]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03553_),
    .QN(_01142_),
    .RESETN(net1513),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[727]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03554_),
    .QN(_01175_),
    .RESETN(net1514),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[728]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03555_),
    .QN(_01208_),
    .RESETN(net1515),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[729]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03556_),
    .QN(_01241_),
    .RESETN(net1516),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[72]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03557_),
    .QN(_00664_),
    .RESETN(net1517),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[730]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03558_),
    .QN(_01274_),
    .RESETN(net1518),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[731]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03559_),
    .QN(_01307_),
    .RESETN(net1519),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[732]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03560_),
    .QN(_01340_),
    .RESETN(net1520),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[733]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03561_),
    .QN(_01373_),
    .RESETN(net1521),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[734]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03562_),
    .QN(_01406_),
    .RESETN(net1522),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[735]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03563_),
    .QN(_01439_),
    .RESETN(net1523),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[736]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03564_),
    .QN(_00438_),
    .RESETN(net1524),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[737]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03565_),
    .QN(_00391_),
    .RESETN(net1525),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[738]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03566_),
    .QN(_00502_),
    .RESETN(net1526),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[739]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03567_),
    .QN(_00533_),
    .RESETN(net1527),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[73]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03568_),
    .QN(_00694_),
    .RESETN(net1528),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[740]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03569_),
    .QN(_00563_),
    .RESETN(net1529),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[741]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03570_),
    .QN(_00595_),
    .RESETN(net1530),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[742]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03571_),
    .QN(_00625_),
    .RESETN(net1531),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[743]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03572_),
    .QN(_00655_),
    .RESETN(net1532),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[744]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03573_),
    .QN(_00685_),
    .RESETN(net1533),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[745]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03574_),
    .QN(_00715_),
    .RESETN(net1534),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[746]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03575_),
    .QN(_00745_),
    .RESETN(net1535),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[747]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03576_),
    .QN(_00775_),
    .RESETN(net1536),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[748]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03577_),
    .QN(_00471_),
    .RESETN(net1537),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[749]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03578_),
    .QN(_00846_),
    .RESETN(net1538),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[74]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03579_),
    .QN(_00724_),
    .RESETN(net1539),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[750]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03580_),
    .QN(_00879_),
    .RESETN(net1540),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[751]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03581_),
    .QN(_00912_),
    .RESETN(net1541),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[752]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03582_),
    .QN(_00945_),
    .RESETN(net1542),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[753]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03583_),
    .QN(_00978_),
    .RESETN(net1543),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[754]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03584_),
    .QN(_01011_),
    .RESETN(net1544),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[755]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03585_),
    .QN(_01044_),
    .RESETN(net1545),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[756]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03586_),
    .QN(_01077_),
    .RESETN(net1546),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[757]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03587_),
    .QN(_01110_),
    .RESETN(net1547),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[758]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03588_),
    .QN(_01143_),
    .RESETN(net1548),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[759]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03589_),
    .QN(_01176_),
    .RESETN(net1549),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[75]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03590_),
    .QN(_00754_),
    .RESETN(net1550),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[760]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03591_),
    .QN(_01209_),
    .RESETN(net1551),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[761]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03592_),
    .QN(_01242_),
    .RESETN(net1552),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[762]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03593_),
    .QN(_01275_),
    .RESETN(net1553),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[763]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03594_),
    .QN(_01308_),
    .RESETN(net1554),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[764]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03595_),
    .QN(_01341_),
    .RESETN(net1555),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[765]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03596_),
    .QN(_01374_),
    .RESETN(net1556),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[766]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03597_),
    .QN(_01407_),
    .RESETN(net1557),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[767]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03598_),
    .QN(_01440_),
    .RESETN(net1558),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[768]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03599_),
    .QN(_00439_),
    .RESETN(net1559),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[769]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03600_),
    .QN(_00392_),
    .RESETN(net1560),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[76]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03601_),
    .QN(_00450_),
    .RESETN(net1561),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[770]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03602_),
    .QN(_00503_),
    .RESETN(net1562),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[771]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03603_),
    .QN(_00534_),
    .RESETN(net1563),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[772]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03604_),
    .QN(_00564_),
    .RESETN(net1564),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[773]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03605_),
    .QN(_00596_),
    .RESETN(net1565),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[774]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03606_),
    .QN(_00626_),
    .RESETN(net1566),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[775]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03607_),
    .QN(_00656_),
    .RESETN(net1567),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[776]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_03608_),
    .QN(_00686_),
    .RESETN(net1568),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[777]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03609_),
    .QN(_00716_),
    .RESETN(net1569),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[778]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03610_),
    .QN(_00746_),
    .RESETN(net1570),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[779]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03611_),
    .QN(_00776_),
    .RESETN(net1571),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[77]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03612_),
    .QN(_00825_),
    .RESETN(net1572),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[780]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03613_),
    .QN(_00472_),
    .RESETN(net1573),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[781]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03614_),
    .QN(_00847_),
    .RESETN(net1574),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[782]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03615_),
    .QN(_00880_),
    .RESETN(net1575),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[783]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03616_),
    .QN(_00913_),
    .RESETN(net1576),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[784]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03617_),
    .QN(_00946_),
    .RESETN(net1577),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[785]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03618_),
    .QN(_00979_),
    .RESETN(net1578),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[786]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03619_),
    .QN(_01012_),
    .RESETN(net1579),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[787]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03620_),
    .QN(_01045_),
    .RESETN(net1580),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[788]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03621_),
    .QN(_01078_),
    .RESETN(net1581),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[789]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03622_),
    .QN(_01111_),
    .RESETN(net1582),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[78]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03623_),
    .QN(_00858_),
    .RESETN(net1583),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[790]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03624_),
    .QN(_01144_),
    .RESETN(net1584),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[791]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03625_),
    .QN(_01177_),
    .RESETN(net1585),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[792]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03626_),
    .QN(_01210_),
    .RESETN(net1586),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[793]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03627_),
    .QN(_01243_),
    .RESETN(net1587),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[794]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03628_),
    .QN(_01276_),
    .RESETN(net1588),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[795]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03629_),
    .QN(_01309_),
    .RESETN(net1589),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[796]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03630_),
    .QN(_01342_),
    .RESETN(net1590),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[797]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03631_),
    .QN(_01375_),
    .RESETN(net1591),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[798]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03632_),
    .QN(_01408_),
    .RESETN(net1592),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[799]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03633_),
    .QN(_01441_),
    .RESETN(net1593),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[79]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03634_),
    .QN(_00891_),
    .RESETN(net1594),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03635_),
    .QN(_01785_),
    .RESETN(net1595),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[800]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03636_),
    .QN(_00440_),
    .RESETN(net1596),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[801]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03637_),
    .QN(_00393_),
    .RESETN(net1597),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[802]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03638_),
    .QN(_00504_),
    .RESETN(net1598),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[803]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03639_),
    .QN(_00535_),
    .RESETN(net1599),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[804]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03640_),
    .QN(_00565_),
    .RESETN(net1600),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[805]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03641_),
    .QN(_00597_),
    .RESETN(net1601),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[806]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03642_),
    .QN(_00627_),
    .RESETN(net1602),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[807]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03643_),
    .QN(_00657_),
    .RESETN(net1603),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[808]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03644_),
    .QN(_00687_),
    .RESETN(net1604),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[809]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03645_),
    .QN(_00717_),
    .RESETN(net1605),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[80]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03646_),
    .QN(_00924_),
    .RESETN(net1606),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[810]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03647_),
    .QN(_00747_),
    .RESETN(net1607),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[811]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03648_),
    .QN(_00777_),
    .RESETN(net1608),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[812]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03649_),
    .QN(_00473_),
    .RESETN(net1609),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[813]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03650_),
    .QN(_00848_),
    .RESETN(net1610),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[814]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03651_),
    .QN(_00881_),
    .RESETN(net1611),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[815]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03652_),
    .QN(_00914_),
    .RESETN(net1612),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[816]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03653_),
    .QN(_00947_),
    .RESETN(net1613),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[817]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03654_),
    .QN(_00980_),
    .RESETN(net1614),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[818]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03655_),
    .QN(_01013_),
    .RESETN(net1615),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[819]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03656_),
    .QN(_01046_),
    .RESETN(net1616),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[81]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03657_),
    .QN(_00957_),
    .RESETN(net1617),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[820]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03658_),
    .QN(_01079_),
    .RESETN(net1618),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[821]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03659_),
    .QN(_01112_),
    .RESETN(net1619),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[822]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03660_),
    .QN(_01145_),
    .RESETN(net1620),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[823]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03661_),
    .QN(_01178_),
    .RESETN(net1621),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[824]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03662_),
    .QN(_01211_),
    .RESETN(net1622),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[825]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03663_),
    .QN(_01244_),
    .RESETN(net1623),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[826]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03664_),
    .QN(_01277_),
    .RESETN(net1624),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[827]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03665_),
    .QN(_01310_),
    .RESETN(net1625),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[828]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03666_),
    .QN(_01343_),
    .RESETN(net1626),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[829]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03667_),
    .QN(_01376_),
    .RESETN(net1627),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[82]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03668_),
    .QN(_00990_),
    .RESETN(net1628),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[830]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03669_),
    .QN(_01409_),
    .RESETN(net1629),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[831]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03670_),
    .QN(_01442_),
    .RESETN(net1630),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[832]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03671_),
    .QN(_00441_),
    .RESETN(net1631),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[833]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03672_),
    .QN(_00394_),
    .RESETN(net1632),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[834]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03673_),
    .QN(_00505_),
    .RESETN(net1633),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[835]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03674_),
    .QN(_00536_),
    .RESETN(net1634),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[836]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03675_),
    .QN(_00566_),
    .RESETN(net1635),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[837]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk_i_regs),
    .D(_03676_),
    .QN(_00598_),
    .RESETN(net1636),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[838]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03677_),
    .QN(_00628_),
    .RESETN(net1637),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[839]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03678_),
    .QN(_00658_),
    .RESETN(net1638),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[83]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03679_),
    .QN(_01023_),
    .RESETN(net1639),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[840]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03680_),
    .QN(_00688_),
    .RESETN(net1640),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[841]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03681_),
    .QN(_00718_),
    .RESETN(net1641),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[842]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03682_),
    .QN(_00748_),
    .RESETN(net1642),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[843]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03683_),
    .QN(_00778_),
    .RESETN(net1643),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[844]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03684_),
    .QN(_00474_),
    .RESETN(net1644),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[845]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03685_),
    .QN(_00849_),
    .RESETN(net1645),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[846]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03686_),
    .QN(_00882_),
    .RESETN(net1646),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[847]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03687_),
    .QN(_00915_),
    .RESETN(net1647),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[848]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03688_),
    .QN(_00948_),
    .RESETN(net1648),
    .SETN(net59));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[849]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03689_),
    .QN(_00981_),
    .RESETN(net1649),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[84]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03690_),
    .QN(_01056_),
    .RESETN(net1650),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[850]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03691_),
    .QN(_01014_),
    .RESETN(net1651),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[851]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03692_),
    .QN(_01047_),
    .RESETN(net1652),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[852]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03693_),
    .QN(_01080_),
    .RESETN(net1653),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[853]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03694_),
    .QN(_01113_),
    .RESETN(net1654),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[854]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03695_),
    .QN(_01146_),
    .RESETN(net1655),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[855]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03696_),
    .QN(_01179_),
    .RESETN(net1656),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[856]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03697_),
    .QN(_01212_),
    .RESETN(net1657),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[857]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03698_),
    .QN(_01245_),
    .RESETN(net1658),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[858]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03699_),
    .QN(_01278_),
    .RESETN(net1659),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[859]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03700_),
    .QN(_01311_),
    .RESETN(net1660),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[85]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03701_),
    .QN(_01089_),
    .RESETN(net1661),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[860]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03702_),
    .QN(_01344_),
    .RESETN(net1662),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[861]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03703_),
    .QN(_01377_),
    .RESETN(net1663),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[862]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03704_),
    .QN(_01410_),
    .RESETN(net1664),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[863]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03705_),
    .QN(_01443_),
    .RESETN(net1665),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[864]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03706_),
    .QN(_00442_),
    .RESETN(net1666),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[865]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03707_),
    .QN(_00395_),
    .RESETN(net1667),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[866]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03708_),
    .QN(_00506_),
    .RESETN(net1668),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[867]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03709_),
    .QN(_00537_),
    .RESETN(net1669),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[868]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03710_),
    .QN(_00567_),
    .RESETN(net1670),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[869]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03711_),
    .QN(_00599_),
    .RESETN(net1671),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[86]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03712_),
    .QN(_01122_),
    .RESETN(net1672),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[870]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03713_),
    .QN(_00629_),
    .RESETN(net1673),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[871]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03714_),
    .QN(_00659_),
    .RESETN(net1674),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[872]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03715_),
    .QN(_00689_),
    .RESETN(net1675),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[873]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk_i_regs),
    .D(_03716_),
    .QN(_00719_),
    .RESETN(net1676),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[874]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03717_),
    .QN(_00749_),
    .RESETN(net1677),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[875]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03718_),
    .QN(_00779_),
    .RESETN(net1678),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[876]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03719_),
    .QN(_00475_),
    .RESETN(net1679),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[877]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03720_),
    .QN(_00850_),
    .RESETN(net1680),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[878]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03721_),
    .QN(_00883_),
    .RESETN(net1681),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[879]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03722_),
    .QN(_00916_),
    .RESETN(net1682),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[87]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03723_),
    .QN(_01155_),
    .RESETN(net1683),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[880]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03724_),
    .QN(_00949_),
    .RESETN(net1684),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[881]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk_i_regs),
    .D(_03725_),
    .QN(_00982_),
    .RESETN(net1685),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[882]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03726_),
    .QN(_01015_),
    .RESETN(net1686),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[883]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03727_),
    .QN(_01048_),
    .RESETN(net1687),
    .SETN(net2021));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[884]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03728_),
    .QN(_01081_),
    .RESETN(net1688),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[885]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03729_),
    .QN(_01114_),
    .RESETN(net1689),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[886]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03730_),
    .QN(_01147_),
    .RESETN(net1690),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[887]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03731_),
    .QN(_01180_),
    .RESETN(net1691),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[888]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03732_),
    .QN(_01213_),
    .RESETN(net1692),
    .SETN(net57));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[889]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03733_),
    .QN(_01246_),
    .RESETN(net1693),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[88]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03734_),
    .QN(_01188_),
    .RESETN(net1694),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[890]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03735_),
    .QN(_01279_),
    .RESETN(net1695),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[891]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03736_),
    .QN(_01312_),
    .RESETN(net1696),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[892]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03737_),
    .QN(_01345_),
    .RESETN(net1697),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[893]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03738_),
    .QN(_01378_),
    .RESETN(net1698),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[894]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03739_),
    .QN(_01411_),
    .RESETN(net1699),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[895]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03740_),
    .QN(_01444_),
    .RESETN(net1700),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[896]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03741_),
    .QN(_00443_),
    .RESETN(net1701),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[897]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk_i_regs),
    .D(_03742_),
    .QN(_00396_),
    .RESETN(net1702),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[898]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03743_),
    .QN(_00507_),
    .RESETN(net1703),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[899]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03744_),
    .QN(_00538_),
    .RESETN(net1704),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[89]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03745_),
    .QN(_01221_),
    .RESETN(net1705),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03746_),
    .QN(_01784_),
    .RESETN(net1706),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[900]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03747_),
    .QN(_00568_),
    .RESETN(net1707),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[901]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03748_),
    .QN(_00600_),
    .RESETN(net1708),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[902]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03749_),
    .QN(_00630_),
    .RESETN(net1709),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[903]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03750_),
    .QN(_00660_),
    .RESETN(net1710),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[904]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03751_),
    .QN(_00690_),
    .RESETN(net1711),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[905]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03752_),
    .QN(_00720_),
    .RESETN(net1712),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[906]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03753_),
    .QN(_00750_),
    .RESETN(net1713),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[907]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03754_),
    .QN(_00780_),
    .RESETN(net1714),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[908]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03755_),
    .QN(_00476_),
    .RESETN(net1715),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[909]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk_i_regs),
    .D(_03756_),
    .QN(_00851_),
    .RESETN(net1716),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[90]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03757_),
    .QN(_01254_),
    .RESETN(net1717),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[910]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03758_),
    .QN(_00884_),
    .RESETN(net1718),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[911]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03759_),
    .QN(_00917_),
    .RESETN(net1719),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[912]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03760_),
    .QN(_00950_),
    .RESETN(net1720),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[913]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03761_),
    .QN(_00983_),
    .RESETN(net1721),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[914]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03762_),
    .QN(_01016_),
    .RESETN(net1722),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[915]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03763_),
    .QN(_01049_),
    .RESETN(net1723),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[916]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03764_),
    .QN(_01082_),
    .RESETN(net1724),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[917]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03765_),
    .QN(_01115_),
    .RESETN(net1725),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[918]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03766_),
    .QN(_01148_),
    .RESETN(net1726),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[919]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03767_),
    .QN(_01181_),
    .RESETN(net1727),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[91]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03768_),
    .QN(_01287_),
    .RESETN(net1728),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[920]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03769_),
    .QN(_01214_),
    .RESETN(net1729),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[921]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk_i_regs),
    .D(_03770_),
    .QN(_01247_),
    .RESETN(net1730),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[922]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03771_),
    .QN(_01280_),
    .RESETN(net1731),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[923]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03772_),
    .QN(_01313_),
    .RESETN(net1732),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[924]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03773_),
    .QN(_01346_),
    .RESETN(net1733),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[925]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03774_),
    .QN(_01379_),
    .RESETN(net1734),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[926]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03775_),
    .QN(_01412_),
    .RESETN(net1735),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[927]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03776_),
    .QN(_01445_),
    .RESETN(net1736),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[928]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03777_),
    .QN(_00444_),
    .RESETN(net1737),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[929]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03778_),
    .QN(_00397_),
    .RESETN(net1738),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[92]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03779_),
    .QN(_01320_),
    .RESETN(net1739),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[930]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03780_),
    .QN(_00508_),
    .RESETN(net1740),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[931]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03781_),
    .QN(_00539_),
    .RESETN(net1741),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[932]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk_i_regs),
    .D(_03782_),
    .QN(_00569_),
    .RESETN(net1742),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[933]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03783_),
    .QN(_00601_),
    .RESETN(net1743),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[934]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03784_),
    .QN(_00631_),
    .RESETN(net1744),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[935]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03785_),
    .QN(_00661_),
    .RESETN(net1745),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[936]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk_i_regs),
    .D(_03786_),
    .QN(_00691_),
    .RESETN(net1746),
    .SETN(net53));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[937]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk_i_regs),
    .D(_03787_),
    .QN(_00721_),
    .RESETN(net1747),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[938]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03788_),
    .QN(_00751_),
    .RESETN(net1748),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[939]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk_i_regs),
    .D(_03789_),
    .QN(_00781_),
    .RESETN(net1749),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[93]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk_i_regs),
    .D(_03790_),
    .QN(_01353_),
    .RESETN(net1750),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[940]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk_i_regs),
    .D(_03791_),
    .QN(_00477_),
    .RESETN(net1751),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[941]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03792_),
    .QN(_00852_),
    .RESETN(net1752),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[942]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03793_),
    .QN(_00885_),
    .RESETN(net1753),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[943]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03794_),
    .QN(_00918_),
    .RESETN(net1754),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[944]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03795_),
    .QN(_00951_),
    .RESETN(net1755),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[945]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03796_),
    .QN(_00984_),
    .RESETN(net1756),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[946]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03797_),
    .QN(_01017_),
    .RESETN(net1757),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[947]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03798_),
    .QN(_01050_),
    .RESETN(net1758),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[948]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk_i_regs),
    .D(_03799_),
    .QN(_01083_),
    .RESETN(net1759),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[949]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03800_),
    .QN(_01116_),
    .RESETN(net1760),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[94]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03801_),
    .QN(_01386_),
    .RESETN(net1761),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[950]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk_i_regs),
    .D(_03802_),
    .QN(_01149_),
    .RESETN(net1762),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[951]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk_i_regs),
    .D(_03803_),
    .QN(_01182_),
    .RESETN(net1763),
    .SETN(net56));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[952]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03804_),
    .QN(_01215_),
    .RESETN(net1764),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[953]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03805_),
    .QN(_01248_),
    .RESETN(net1765),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[954]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03806_),
    .QN(_01281_),
    .RESETN(net1766),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[955]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk_i_regs),
    .D(_03807_),
    .QN(_01314_),
    .RESETN(net1767),
    .SETN(net58));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[956]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03808_),
    .QN(_01347_),
    .RESETN(net1768),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[957]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk_i_regs),
    .D(_03809_),
    .QN(_01380_),
    .RESETN(net1769),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[958]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk_i_regs),
    .D(_03810_),
    .QN(_01413_),
    .RESETN(net1770),
    .SETN(net65));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[959]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03811_),
    .QN(_01446_),
    .RESETN(net1771),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[95]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03812_),
    .QN(_01419_),
    .RESETN(net1772),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[960]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03813_),
    .QN(_00445_),
    .RESETN(net1773),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[961]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03814_),
    .QN(_00398_),
    .RESETN(net1774),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[962]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03815_),
    .QN(_00509_),
    .RESETN(net1775),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[963]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03816_),
    .QN(_00540_),
    .RESETN(net1776),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[964]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk_i_regs),
    .D(_03817_),
    .QN(_00570_),
    .RESETN(net1777),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[965]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk_i_regs),
    .D(_03818_),
    .QN(_00602_),
    .RESETN(net1778),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[966]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03819_),
    .QN(_00632_),
    .RESETN(net1779),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[967]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03820_),
    .QN(_00662_),
    .RESETN(net1780),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[968]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_03821_),
    .QN(_00692_),
    .RESETN(net1781),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[969]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03822_),
    .QN(_00722_),
    .RESETN(net1782),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[96]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03823_),
    .QN(_00418_),
    .RESETN(net1783),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[970]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03824_),
    .QN(_00752_),
    .RESETN(net1784),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[971]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk_i_regs),
    .D(_03825_),
    .QN(_00782_),
    .RESETN(net1785),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[972]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk_i_regs),
    .D(_03826_),
    .QN(_00478_),
    .RESETN(net1786),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[973]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03827_),
    .QN(_00853_),
    .RESETN(net1787),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[974]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03828_),
    .QN(_00886_),
    .RESETN(net1788),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[975]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03829_),
    .QN(_00919_),
    .RESETN(net1789),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[976]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03830_),
    .QN(_00952_),
    .RESETN(net1790),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[977]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk_i_regs),
    .D(_03831_),
    .QN(_00985_),
    .RESETN(net1791),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[978]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03832_),
    .QN(_01018_),
    .RESETN(net1792),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[979]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03833_),
    .QN(_01051_),
    .RESETN(net1793),
    .SETN(net60));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[97]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk_i_regs),
    .D(_03834_),
    .QN(_00371_),
    .RESETN(net1794),
    .SETN(net63));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[980]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk_i_regs),
    .D(_03835_),
    .QN(_01084_),
    .RESETN(net1795),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[981]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03836_),
    .QN(_01117_),
    .RESETN(net1796),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[982]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03837_),
    .QN(_01150_),
    .RESETN(net1797),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[983]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk_i_regs),
    .D(_03838_),
    .QN(_01183_),
    .RESETN(net1798),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[984]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03839_),
    .QN(_01216_),
    .RESETN(net1799),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[985]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03840_),
    .QN(_01249_),
    .RESETN(net1800),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[986]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03841_),
    .QN(_01282_),
    .RESETN(net1801),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[987]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03842_),
    .QN(_01315_),
    .RESETN(net1802),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[988]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk_i_regs),
    .D(_03843_),
    .QN(_01348_),
    .RESETN(net1803),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[989]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk_i_regs),
    .D(_03844_),
    .QN(_01381_),
    .RESETN(net1804),
    .SETN(net62));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[98]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk_i_regs),
    .D(_03845_),
    .QN(_00482_),
    .RESETN(net1805),
    .SETN(net64));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[990]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03846_),
    .QN(_01414_),
    .RESETN(net1806),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[991]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk_i_regs),
    .D(_03847_),
    .QN(_01447_),
    .RESETN(net1807),
    .SETN(net55));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[99]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk_i_regs),
    .D(_03848_),
    .QN(_00513_),
    .RESETN(net1808),
    .SETN(net61));
 DFFASRHQNx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk_i_regs),
    .D(_03849_),
    .QN(_01783_),
    .RESETN(net1809),
    .SETN(net54));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_03850_),
    .QN(_01782_),
    .RESETN(net1810),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_03851_),
    .QN(_01781_),
    .RESETN(net1811),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_03852_),
    .QN(_01780_),
    .RESETN(net1812),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_03853_),
    .QN(_01779_),
    .RESETN(net1813),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.debug_mode_q$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .D(_03854_),
    .QN(_01455_),
    .RESETN(net1814),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .D(\id_stage_i.controller_i.exc_req_d ),
    .QN(_02219_),
    .RESETN(net1815),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .D(\id_stage_i.controller_i.illegal_insn_d ),
    .QN(_00791_),
    .RESETN(net1816),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .D(\id_stage_i.controller_i.load_err_d ),
    .QN(_01778_),
    .RESETN(net1817),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.nmi_mode_q$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .D(_03855_),
    .QN(_02220_),
    .RESETN(net1818),
    .SETN(net72));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .D(\id_stage_i.controller_i.store_err_d ),
    .QN(_02221_),
    .RESETN(net1819),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.g_branch_set_flop.branch_set_q$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .D(\id_stage_i.branch_set_d ),
    .QN(_01777_),
    .RESETN(net1820),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_03856_),
    .QN(_01776_),
    .RESETN(net1821),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03857_),
    .QN(_01775_),
    .RESETN(net1822),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_03858_),
    .QN(_01774_),
    .RESETN(net1823),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03859_),
    .QN(_01773_),
    .RESETN(net1824),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_03860_),
    .QN(_01772_),
    .RESETN(net1825),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_03861_),
    .QN(_01771_),
    .RESETN(net1826),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03862_),
    .QN(_01770_),
    .RESETN(net1827),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_03863_),
    .QN(_01769_),
    .RESETN(net1828),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_03864_),
    .QN(_01768_),
    .RESETN(net1829),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03865_),
    .QN(_01767_),
    .RESETN(net1830),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_03866_),
    .QN(_01766_),
    .RESETN(net1831),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03867_),
    .QN(_01765_),
    .RESETN(net1832),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03868_),
    .QN(_01764_),
    .RESETN(net1833),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03869_),
    .QN(_01763_),
    .RESETN(net1834),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03870_),
    .QN(_01762_),
    .RESETN(net1835),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03871_),
    .QN(_01761_),
    .RESETN(net1836),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03872_),
    .QN(_01760_),
    .RESETN(net1837),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03873_),
    .QN(_01759_),
    .RESETN(net1838),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03874_),
    .QN(_01758_),
    .RESETN(net1839),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03875_),
    .QN(_01757_),
    .RESETN(net1840),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03876_),
    .QN(_01756_),
    .RESETN(net1841),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03877_),
    .QN(_01755_),
    .RESETN(net1842),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03878_),
    .QN(_01754_),
    .RESETN(net1843),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03879_),
    .QN(_01753_),
    .RESETN(net1844),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03880_),
    .QN(_01752_),
    .RESETN(net1845),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03881_),
    .QN(_01751_),
    .RESETN(net1846),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[34]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03882_),
    .QN(_00447_),
    .RESETN(net1847),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[35]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03883_),
    .QN(_00414_),
    .RESETN(net1848),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[36]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03884_),
    .QN(_00792_),
    .RESETN(net1849),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[37]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03885_),
    .QN(_00795_),
    .RESETN(net1850),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[38]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03886_),
    .QN(_00798_),
    .RESETN(net1851),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[39]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03887_),
    .QN(_00801_),
    .RESETN(net1852),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_03888_),
    .QN(_01750_),
    .RESETN(net1853),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[40]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03889_),
    .QN(_00804_),
    .RESETN(net1854),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[41]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03890_),
    .QN(_00807_),
    .RESETN(net1855),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[42]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03891_),
    .QN(_00809_),
    .RESETN(net1856),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[43]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03892_),
    .QN(_00812_),
    .RESETN(net1857),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[44]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03893_),
    .QN(_00815_),
    .RESETN(net1858),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[45]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03894_),
    .QN(_00818_),
    .RESETN(net1859),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[46]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_03895_),
    .QN(_00821_),
    .RESETN(net1860),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[47]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03896_),
    .QN(_00854_),
    .RESETN(net1861),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[48]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03897_),
    .QN(_00887_),
    .RESETN(net1862),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[49]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03898_),
    .QN(_00920_),
    .RESETN(net1863),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .D(_03899_),
    .QN(_01749_),
    .RESETN(net1864),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[50]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03900_),
    .QN(_00953_),
    .RESETN(net1865),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[51]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03901_),
    .QN(_00986_),
    .RESETN(net1866),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[52]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03902_),
    .QN(_01019_),
    .RESETN(net1867),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[53]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03903_),
    .QN(_01052_),
    .RESETN(net1868),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[54]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03904_),
    .QN(_01085_),
    .RESETN(net1869),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[55]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_03905_),
    .QN(_01118_),
    .RESETN(net1870),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[56]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_03906_),
    .QN(_01151_),
    .RESETN(net1871),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[57]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_03907_),
    .QN(_01184_),
    .RESETN(net1872),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[58]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_03908_),
    .QN(_01217_),
    .RESETN(net1873),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[59]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03909_),
    .QN(_01250_),
    .RESETN(net1874),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03910_),
    .QN(_01748_),
    .RESETN(net1875),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[60]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .D(_03911_),
    .QN(_01283_),
    .RESETN(net1876),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[61]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03912_),
    .QN(_01316_),
    .RESETN(net1877),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[62]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03913_),
    .QN(_01349_),
    .RESETN(net1878),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[63]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03914_),
    .QN(_01382_),
    .RESETN(net1879),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[64]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03915_),
    .QN(_01415_),
    .RESETN(net1880),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[65]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03916_),
    .QN(_01448_),
    .RESETN(net1881),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[66]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03917_),
    .QN(_01747_),
    .RESETN(net1882),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[67]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .D(_03918_),
    .QN(_00232_),
    .RESETN(net1883),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03919_),
    .QN(_01746_),
    .RESETN(net1884),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03920_),
    .QN(_01745_),
    .RESETN(net1885),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03921_),
    .QN(_01744_),
    .RESETN(net1886),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \id_stage_i.imd_val_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .D(_03922_),
    .QN(_02222_),
    .RESETN(net1887),
    .SETN(net74));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .QN(_02223_),
    .RESETN(net1888),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .QN(_02224_),
    .RESETN(net1889),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .QN(_01743_),
    .RESETN(net1890),
    .SETN(net67));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03923_),
    .QN(_01742_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03924_),
    .QN(_01741_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03925_),
    .QN(_01740_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03926_),
    .QN(_01739_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_03927_),
    .QN(_01738_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03928_),
    .QN(_01737_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_03929_),
    .QN(_01736_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_03930_),
    .QN(_01735_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_03931_),
    .QN(_01734_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03932_),
    .QN(_01733_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03933_),
    .QN(_01732_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03934_),
    .QN(_01731_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03935_),
    .QN(_01730_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03936_),
    .QN(_01729_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03937_),
    .QN(_01728_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03938_),
    .QN(_01727_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03939_),
    .QN(_01726_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_03940_),
    .QN(_01725_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_03941_),
    .QN(_01724_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_03942_),
    .QN(_01723_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03943_),
    .QN(_01722_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03944_),
    .QN(_01721_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_03945_),
    .QN(_01720_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03946_),
    .QN(_01719_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03947_),
    .QN(_01718_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03948_),
    .QN(_01717_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03949_),
    .QN(_01716_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03950_),
    .QN(_01715_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03951_),
    .QN(_01714_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03952_),
    .QN(_01713_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_03953_),
    .QN(_01712_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_03954_),
    .QN(_01711_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_03955_),
    .QN(_01710_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_03956_),
    .QN(_00365_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03957_),
    .QN(_01709_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_03958_),
    .QN(_01708_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03959_),
    .QN(_01707_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03960_),
    .QN(_01706_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03961_),
    .QN(_01705_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_03962_),
    .QN(_01704_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03963_),
    .QN(_01703_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_03964_),
    .QN(_01702_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03965_),
    .QN(_01701_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03966_),
    .QN(_01700_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03967_),
    .QN(_18317_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03968_),
    .QN(_01699_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03969_),
    .QN(_01698_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03970_),
    .QN(_01697_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03971_),
    .QN(_01696_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_03972_),
    .QN(_01695_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03973_),
    .QN(_01694_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03974_),
    .QN(_01693_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_03975_),
    .QN(_01692_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_03976_),
    .QN(_01691_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_03977_),
    .QN(_01690_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_03978_),
    .QN(_01689_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03979_),
    .QN(_01688_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03980_),
    .QN(_01687_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03981_),
    .QN(_01686_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_03982_),
    .QN(_01685_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03983_),
    .QN(_01684_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_03984_),
    .QN(_01683_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_03985_),
    .QN(_01682_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_03986_),
    .QN(_01681_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_03987_),
    .QN(_01680_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_03988_),
    .QN(_01679_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_03989_),
    .QN(_01678_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_03990_),
    .QN(_01677_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_03991_),
    .QN(_01676_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_03992_),
    .QN(_01675_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_03993_),
    .QN(_01674_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_03994_),
    .QN(_01673_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_03995_),
    .QN(_01672_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_03996_),
    .QN(_01671_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_03997_),
    .QN(_01670_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_03998_),
    .QN(_01669_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_03999_),
    .QN(_01668_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04000_),
    .QN(_01667_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04001_),
    .QN(_01666_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04002_),
    .QN(_01665_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04003_),
    .QN(_01664_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04004_),
    .QN(_01663_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04005_),
    .QN(_01662_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04006_),
    .QN(_01661_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04007_),
    .QN(_01660_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04008_),
    .QN(_01659_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04009_),
    .QN(_01658_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04010_),
    .QN(_01657_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04011_),
    .QN(_01656_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04012_),
    .QN(_01655_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04013_),
    .QN(_01654_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04014_),
    .QN(_01653_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04015_),
    .QN(_01652_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04016_),
    .QN(_01651_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04017_),
    .QN(_01650_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_04018_),
    .QN(_01649_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04019_),
    .QN(_01648_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04020_),
    .QN(_01647_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04021_),
    .QN(_01646_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04022_),
    .QN(_01645_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04023_),
    .QN(_01644_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04024_),
    .QN(_01643_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04025_),
    .QN(_01642_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04026_),
    .QN(_01641_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04027_),
    .QN(_01640_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04028_),
    .QN(_01639_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04029_),
    .QN(_01638_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04030_),
    .QN(_01637_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04031_),
    .QN(_01636_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04032_),
    .QN(_01635_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04033_),
    .QN(_01634_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04034_),
    .QN(_01633_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04035_),
    .QN(_01632_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04036_),
    .QN(_01631_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04037_),
    .QN(_01630_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04038_),
    .QN(_01629_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04039_),
    .QN(_01628_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04040_),
    .QN(_01627_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04041_),
    .QN(_01626_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04042_),
    .QN(_01625_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04043_),
    .QN(_01624_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04044_),
    .QN(_01623_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04045_),
    .QN(_01622_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04046_),
    .QN(_01621_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04047_),
    .QN(_01620_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_04048_),
    .QN(_01619_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04049_),
    .QN(_01618_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04050_),
    .QN(_01617_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04051_),
    .QN(_01616_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04052_),
    .QN(_01615_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04053_),
    .QN(_01614_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_04054_),
    .QN(_01613_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04055_),
    .QN(_01612_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_04056_),
    .QN(_01611_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04057_),
    .QN(_01610_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04058_),
    .QN(_01609_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04059_),
    .QN(_01608_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04060_),
    .QN(_01607_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04061_),
    .QN(_01606_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_04062_),
    .QN(_01605_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04063_),
    .QN(_01604_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04064_),
    .QN(_01603_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04065_),
    .QN(_01602_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_04066_),
    .QN(_01601_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04067_),
    .QN(_01600_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04068_),
    .QN(_01599_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04069_),
    .QN(_01598_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04070_),
    .QN(_01597_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04071_),
    .QN(_01596_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04072_),
    .QN(_01595_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04073_),
    .QN(_01594_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04074_),
    .QN(_01593_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04075_),
    .QN(_01592_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04076_),
    .QN(_01591_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04077_),
    .QN(_01590_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_04078_),
    .QN(_01589_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04079_),
    .QN(_01588_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04080_),
    .QN(_01587_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_04081_),
    .QN(_01586_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04082_),
    .QN(_02225_));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .QN(_00291_),
    .RESETN(net1891),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .QN(_00290_),
    .RESETN(net1892),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .QN(_02226_),
    .RESETN(net1893),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .QN(_02227_),
    .RESETN(net1894),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .QN(_00289_),
    .RESETN(net1895),
    .SETN(net67));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04083_),
    .QN(_01585_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04084_),
    .QN(_01584_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04085_),
    .QN(_01583_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04086_),
    .QN(_01582_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04087_),
    .QN(_01581_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_04088_),
    .QN(_01580_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_04089_),
    .QN(_01579_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_04090_),
    .QN(_01578_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_04091_),
    .QN(_01577_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_04092_),
    .QN(_01576_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04093_),
    .QN(_01575_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04094_),
    .QN(_01574_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04095_),
    .QN(_01573_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04096_),
    .QN(_01572_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04097_),
    .QN(_01571_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04098_),
    .QN(_01570_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_04099_),
    .QN(_01569_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_04100_),
    .QN(_01568_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_04101_),
    .QN(_01567_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04102_),
    .QN(_01566_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04103_),
    .QN(_01565_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04104_),
    .QN(_01564_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04105_),
    .QN(_01563_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04106_),
    .QN(_01562_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04107_),
    .QN(_01561_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04108_),
    .QN(_01560_));
 DFFHQNx3_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_04109_),
    .QN(_01559_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04110_),
    .QN(_01558_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04111_),
    .QN(_01557_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_04112_),
    .QN(_02228_));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .QN(_00288_),
    .RESETN(net1896),
    .SETN(net67));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04113_),
    .QN(_01556_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04114_),
    .QN(_01555_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.CLK(clknet_leaf_7_clk),
    .D(_04115_),
    .QN(_01554_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04116_),
    .QN(_00510_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[0]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04117_),
    .QN(_01553_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[10]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04118_),
    .QN(_00037_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[11]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .D(_04119_),
    .QN(_00040_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[12]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04120_),
    .QN(_00404_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[13]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04121_),
    .QN(_00403_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[14]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04122_),
    .QN(_00401_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[15]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04123_),
    .QN(_00413_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[16]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04124_),
    .QN(_00412_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[17]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04125_),
    .QN(_00411_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[18]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04126_),
    .QN(_00410_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[19]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04127_),
    .QN(_00409_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[1]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04128_),
    .QN(_00013_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[20]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .D(_04129_),
    .QN(_00368_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[21]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .D(_04130_),
    .QN(_01552_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[22]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .D(_04131_),
    .QN(_01551_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[23]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .D(_04132_),
    .QN(_00367_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[24]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .D(_04133_),
    .QN(_00366_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[25]$_DFFE_PN_  (.CLK(clknet_leaf_9_clk),
    .D(_04134_),
    .QN(_01550_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[26]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04135_),
    .QN(_00405_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[27]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04136_),
    .QN(_01549_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[28]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04137_),
    .QN(_01548_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[29]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04138_),
    .QN(_01547_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[2]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04139_),
    .QN(_00015_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[30]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04140_),
    .QN(_01546_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[31]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04141_),
    .QN(_00402_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[3]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04142_),
    .QN(_00018_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[4]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04143_),
    .QN(_00021_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[5]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04144_),
    .QN(_00024_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[6]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04145_),
    .QN(_00400_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[7]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04146_),
    .QN(_00446_));
 DFFHQNx1_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[8]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04147_),
    .QN(_00031_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_alu_id_o[9]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .D(_04148_),
    .QN(_00034_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04149_),
    .QN(_01545_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04150_),
    .QN(_00038_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04151_),
    .QN(_00041_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04152_),
    .QN(_00043_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04153_),
    .QN(_00045_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04154_),
    .QN(_00047_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04155_),
    .QN(_00049_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04156_),
    .QN(_00014_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04157_),
    .QN(_00016_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04158_),
    .QN(_00019_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .D(_04159_),
    .QN(_00022_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04160_),
    .QN(_00025_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04161_),
    .QN(_00027_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04162_),
    .QN(_00029_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04163_),
    .QN(_00032_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .D(_04164_),
    .QN(_00035_));
 DFFASRHQNx1_ASAP7_75t_R \if_stage_i.instr_valid_id_q$_DFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .D(\if_stage_i.instr_valid_id_d ),
    .QN(_01456_),
    .RESETN(net1897),
    .SETN(net67));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04165_),
    .QN(_00039_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04166_),
    .QN(_00042_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04167_),
    .QN(_00044_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04168_),
    .QN(_00046_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04169_),
    .QN(_00048_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04170_),
    .QN(_00050_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04171_),
    .QN(_00051_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04172_),
    .QN(_00052_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04173_),
    .QN(_00053_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .D(_04174_),
    .QN(_00054_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04175_),
    .QN(_01544_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04176_),
    .QN(_00055_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04177_),
    .QN(_00056_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04178_),
    .QN(_00057_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04179_),
    .QN(_00058_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04180_),
    .QN(_00059_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04181_),
    .QN(_00060_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04182_),
    .QN(_00061_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04183_),
    .QN(_00062_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04184_),
    .QN(_00063_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04185_),
    .QN(_00064_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04186_),
    .QN(_00012_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .D(_04187_),
    .QN(_00065_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04188_),
    .QN(_00066_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04189_),
    .QN(_00020_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04190_),
    .QN(_00023_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04191_),
    .QN(_00026_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04192_),
    .QN(_00028_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .D(_04193_),
    .QN(_00030_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04194_),
    .QN(_00033_));
 DFFHQNx2_ASAP7_75t_R \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.CLK(clknet_leaf_10_clk),
    .D(_04195_),
    .QN(_00036_));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04196_),
    .QN(_01543_),
    .RESETN(net1898),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .D(_04197_),
    .QN(_01542_),
    .RESETN(net1899),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04198_),
    .QN(_01541_),
    .RESETN(net1900),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04199_),
    .QN(_01540_),
    .RESETN(net1901),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04200_),
    .QN(_01539_),
    .RESETN(net1902),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04201_),
    .QN(_01538_),
    .RESETN(net1903),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04202_),
    .QN(_01537_),
    .RESETN(net1904),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04203_),
    .QN(_01536_),
    .RESETN(net1905),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04204_),
    .QN(_01535_),
    .RESETN(net1906),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04205_),
    .QN(_01534_),
    .RESETN(net1907),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04206_),
    .QN(_01533_),
    .RESETN(net1908),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04207_),
    .QN(_01532_),
    .RESETN(net1909),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04208_),
    .QN(_01531_),
    .RESETN(net1910),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04209_),
    .QN(_01530_),
    .RESETN(net1911),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04210_),
    .QN(_01529_),
    .RESETN(net1912),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .D(_04211_),
    .QN(_01528_),
    .RESETN(net1913),
    .SETN(net66));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04212_),
    .QN(_01527_),
    .RESETN(net1914),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04213_),
    .QN(_01526_),
    .RESETN(net1915),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04214_),
    .QN(_01525_),
    .RESETN(net1916),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04215_),
    .QN(_01524_),
    .RESETN(net1917),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04216_),
    .QN(_01523_),
    .RESETN(net1918),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04217_),
    .QN(_01522_),
    .RESETN(net1919),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04218_),
    .QN(_01521_),
    .RESETN(net1920),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04219_),
    .QN(_01520_),
    .RESETN(net1921),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04220_),
    .QN(_01519_),
    .RESETN(net1922),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04221_),
    .QN(_01518_),
    .RESETN(net1923),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04222_),
    .QN(_01517_),
    .RESETN(net1924),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04223_),
    .QN(_01516_),
    .RESETN(net1925),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04224_),
    .QN(_01515_),
    .RESETN(net1926),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04225_),
    .QN(_01514_),
    .RESETN(net1927),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_04226_),
    .QN(_01513_),
    .RESETN(net1928),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_04227_),
    .QN(_01512_),
    .RESETN(net1929),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04228_),
    .QN(_01511_),
    .RESETN(net1930),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04229_),
    .QN(_01454_),
    .RESETN(net1931),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04230_),
    .QN(_18763_),
    .RESETN(net1932),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04231_),
    .QN(_01510_),
    .RESETN(net1933),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04232_),
    .QN(_01509_),
    .RESETN(net1934),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04233_),
    .QN(_00399_),
    .RESETN(net1935),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04234_),
    .QN(_01508_),
    .RESETN(net1936),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04235_),
    .QN(_01507_),
    .RESETN(net1937),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_04236_),
    .QN(_01506_),
    .RESETN(net1938),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04237_),
    .QN(_01505_),
    .RESETN(net1939),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04238_),
    .QN(_01504_),
    .RESETN(net1940),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04239_),
    .QN(_01503_),
    .RESETN(net1941),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04240_),
    .QN(_01502_),
    .RESETN(net1942),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04241_),
    .QN(_01501_),
    .RESETN(net1943),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04242_),
    .QN(_01500_),
    .RESETN(net1944),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04243_),
    .QN(_01499_),
    .RESETN(net1945),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04244_),
    .QN(_01498_),
    .RESETN(net1946),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04245_),
    .QN(_01497_),
    .RESETN(net1947),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04246_),
    .QN(_01496_),
    .RESETN(net1948),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_04247_),
    .QN(_01495_),
    .RESETN(net1949),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04248_),
    .QN(_01494_),
    .RESETN(net1950),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04249_),
    .QN(_01493_),
    .RESETN(net1951),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04250_),
    .QN(_01492_),
    .RESETN(net1952),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04251_),
    .QN(_01491_),
    .RESETN(net1953),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .D(_04252_),
    .QN(_01490_),
    .RESETN(net1954),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04253_),
    .QN(_01489_),
    .RESETN(net1955),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04254_),
    .QN(_01488_),
    .RESETN(net1956),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04255_),
    .QN(_01487_),
    .RESETN(net1957),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04256_),
    .QN(_01486_),
    .RESETN(net1958),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04257_),
    .QN(_01485_),
    .RESETN(net1959),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_04258_),
    .QN(_01484_),
    .RESETN(net1960),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_04259_),
    .QN(_01483_),
    .RESETN(net1961),
    .SETN(net67));
 DFFASRHQNx1_ASAP7_75t_R \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_04260_),
    .QN(_01482_),
    .RESETN(net1962),
    .SETN(net67));
 BUFx6f_ASAP7_75t_R split1 (.A(net1972),
    .Y(net1));
 BUFx2_ASAP7_75t_R clone4 (.A(_00368_),
    .Y(net4));
 BUFx3_ASAP7_75t_R clone9 (.A(_09647_),
    .Y(net9));
 BUFx6f_ASAP7_75t_R clone10 (.A(_13470_),
    .Y(net10));
 BUFx3_ASAP7_75t_R clone11 (.A(net16),
    .Y(net11));
 BUFx6f_ASAP7_75t_R clone12 (.A(_13457_),
    .Y(net12));
 BUFx3_ASAP7_75t_R clone13 (.A(_09580_),
    .Y(net13));
 BUFx3_ASAP7_75t_R clone14 (.A(_13469_),
    .Y(net14));
 BUFx3_ASAP7_75t_R clone15 (.A(_13458_),
    .Y(net15));
 BUFx2_ASAP7_75t_R clone16 (.A(_13467_),
    .Y(net16));
 BUFx2_ASAP7_75t_R clone17 (.A(_13457_),
    .Y(net17));
 BUFx3_ASAP7_75t_R clone18 (.A(_15518_),
    .Y(net18));
 BUFx4f_ASAP7_75t_R clone19 (.A(net18),
    .Y(net19));
 BUFx3_ASAP7_75t_R clone20 (.A(_13456_),
    .Y(net20));
 BUFx2_ASAP7_75t_R clone21 (.A(_15537_),
    .Y(net21));
 BUFx3_ASAP7_75t_R clone22 (.A(_15537_),
    .Y(net22));
 BUFx3_ASAP7_75t_R clone95 (.A(_09543_),
    .Y(net95));
 BUFx2_ASAP7_75t_R clone145 (.A(_15537_),
    .Y(net145));
 BUFx3_ASAP7_75t_R clone151 (.A(_09621_),
    .Y(net151));
 BUFx3_ASAP7_75t_R clone152 (.A(_09621_),
    .Y(net152));
 BUFx3_ASAP7_75t_R clone153 (.A(_09621_),
    .Y(net153));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_Right_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_Right_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_Right_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_Right_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_Right_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_Right_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_Right_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_Right_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_Right_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_Right_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_Right_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_Right_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_Right_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_Right_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_Right_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_Right_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_Right_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_Right_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_Right_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_Right_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_Right_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_Right_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_Right_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_Right_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Left_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Left_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Left_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Left_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Left_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Left_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Left_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Left_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Left_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Left_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Left_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Left_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Left_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Left_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Left_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Left_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Left_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Left_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Left_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Left_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Left_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Left_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Left_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Left_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Left_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Left_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Left_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Left_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Left_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Left_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Left_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Left_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Left_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Left_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Left_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Left_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Left_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Left_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Left_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Left_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Left_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Left_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Left_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Left_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Left_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Left_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Left_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Left_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Left_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Left_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Left_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Left_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Left_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Left_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Left_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Left_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Left_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Left_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Left_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Left_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Left_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Left_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Left_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Left_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Left_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Left_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Left_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Left_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Left_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Left_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Left_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Left_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Left_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Left_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Left_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Left_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Left_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Left_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Left_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Left_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Left_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Left_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Left_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Left_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Left_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Left_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Left_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Left_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Left_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Left_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Left_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Left_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Left_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Left_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Left_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Left_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Left_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Left_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Left_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Left_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Left_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Left_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Left_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Left_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Left_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Left_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Left_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Left_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Left_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Left_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Left_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Left_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_Left_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_Left_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_Left_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_Left_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_Left_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_Left_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_Left_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_Left_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_Left_479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_Left_480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_Left_481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_Left_482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_Left_483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_Left_484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_Left_485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_Left_486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_Left_487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_Left_488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_Left_489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_Left_490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_Left_491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_Left_492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_Left_493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_Left_494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_Left_495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_Left_496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_Left_497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_Left_498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_Left_499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_Left_500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_Left_501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_Left_502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_Left_503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_Left_504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_Left_505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_Left_506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_Left_507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_Left_508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_Left_509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_Left_510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_Left_511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_Left_512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_Left_513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_Left_514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_Left_515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_Left_516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_Left_517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_Left_518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_Left_519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_Left_520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_Left_521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_Left_522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Left_523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Left_524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_Left_525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_Left_526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_Left_527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_Left_528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_Left_529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_Left_530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_Left_531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_Left_532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_Left_533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_Left_534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_Left_535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_Left_536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_Left_537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_Left_538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_Left_539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_Left_540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_Left_541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_Left_542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_Left_543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_Left_544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_Left_545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_Left_546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_Left_547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_Left_548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_Left_549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_Left_550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_Left_551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_Left_552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_Left_553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_Left_554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_Left_555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_Left_556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_Left_557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_Left_558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_Left_559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_Left_560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_Left_561 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_562 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_563 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_564 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_565 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_566 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_567 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_568 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_569 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_570 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_571 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_572 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_573 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_574 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_575 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_576 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_577 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_578 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_579 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_580 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_581 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_582 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_583 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_584 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_585 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_15_586 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_587 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_588 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_17_589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_19_592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_21_595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_23_598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_25_601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_27_604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_29_607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_31_610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_33_613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_35_616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_37_619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_39_622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_41_625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_43_628 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_629 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_630 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_45_631 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_632 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_633 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_47_634 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_635 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_636 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_49_637 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_638 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_639 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_51_640 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_641 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_642 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_53_643 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_644 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_645 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_55_646 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_647 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_648 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_57_649 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_650 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_651 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_59_652 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_653 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_654 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_61_655 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_656 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_657 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_63_658 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_659 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_660 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_65_661 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_662 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_663 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_67_664 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_665 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_666 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_69_667 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_668 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_669 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_71_670 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_671 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_672 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_73_673 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_674 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_675 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_75_676 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_677 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_678 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_77_679 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_680 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_681 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_79_682 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_683 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_684 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_81_685 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_686 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_687 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_83_688 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_689 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_690 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_85_691 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_692 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_693 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_87_694 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_695 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_696 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_89_697 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_698 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_699 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_91_700 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_701 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_702 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_703 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_704 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_705 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_95_706 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_707 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_708 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_97_709 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_710 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_711 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_99_712 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_713 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_714 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_101_715 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_716 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_717 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_103_718 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_719 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_720 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_105_721 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_722 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_723 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_107_724 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_725 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_726 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_109_727 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_728 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_729 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_111_730 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_731 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_732 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_113_733 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_734 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_735 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_115_736 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_737 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_738 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_117_739 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_740 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_741 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_119_742 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_743 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_744 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_121_745 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_746 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_747 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_123_748 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_749 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_750 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_125_751 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_752 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_753 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_127_754 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_755 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_756 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_129_757 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_758 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_759 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_131_760 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_761 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_762 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_133_763 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_764 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_765 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_135_766 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_767 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_768 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_137_769 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_770 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_771 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_139_772 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_773 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_774 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_141_775 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_776 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_777 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_143_778 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_779 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_780 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_145_781 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_782 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_783 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_147_784 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_785 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_786 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_149_787 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_788 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_789 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_151_790 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_152_791 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_152_792 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_153_793 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_154_794 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_154_795 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_155_796 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_156_797 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_156_798 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_157_799 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_158_800 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_158_801 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_159_802 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_160_803 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_160_804 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_161_805 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_806 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_807 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_163_808 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_809 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_810 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_165_811 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_812 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_813 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_167_814 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_815 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_816 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_169_817 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_818 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_819 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_171_820 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_821 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_822 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_823 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_174_824 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_174_825 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_175_826 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_176_827 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_176_828 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_177_829 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_830 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_831 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_832 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_833 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_834 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_835 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_836 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_837 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_838 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_839 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_840 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_841 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_842 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_843 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_844 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_845 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_846 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_847 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_190_848 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_190_849 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_191_850 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_192_851 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_192_852 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_193_853 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_194_854 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_194_855 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_195_856 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_196_857 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_196_858 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_197_859 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_198_860 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_198_861 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_199_862 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_200_863 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_200_864 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_201_865 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_202_866 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_202_867 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_203_868 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_204_869 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_204_870 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_205_871 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_206_872 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_206_873 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_207_874 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_208_875 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_208_876 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_209_877 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_210_878 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_210_879 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_211_880 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_212_881 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_212_882 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_213_883 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_214_884 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_214_885 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_215_886 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_216_887 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_216_888 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_217_889 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_218_890 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_218_891 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_219_892 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_220_893 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_220_894 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_221_895 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_222_896 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_222_897 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_223_898 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_224_899 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_224_900 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_225_901 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_226_902 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_226_903 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_227_904 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_228_905 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_228_906 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_229_907 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_230_908 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_230_909 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_231_910 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_232_911 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_232_912 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_233_913 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_234_914 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_234_915 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_235_916 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_236_917 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_236_918 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_237_919 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_238_920 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_238_921 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_239_922 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_240_923 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_240_924 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_241_925 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_926 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_927 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_243_928 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_244_929 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_244_930 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_245_931 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_246_932 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_246_933 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_247_934 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_248_935 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_248_936 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_249_937 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_250_938 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_250_939 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_251_940 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_252_941 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_252_942 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_253_943 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_254_944 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_254_945 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_255_946 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_256_947 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_256_948 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_257_949 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_258_950 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_258_951 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_259_952 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_260_953 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_260_954 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_261_955 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_262_956 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_262_957 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_263_958 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_264_959 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_264_960 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_265_961 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_266_962 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_266_963 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_267_964 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_268_965 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_268_966 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_269_967 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_270_968 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_270_969 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_271_970 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_272_971 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_272_972 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_273_973 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_274_974 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_274_975 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_275_976 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_276_977 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_276_978 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_277_979 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_278_980 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_278_981 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_279_982 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_280_983 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_280_984 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_280_985 ();
 BUFx6f_ASAP7_75t_R load_slew30 (.A(_18769_),
    .Y(net52));
 BUFx16f_ASAP7_75t_R load_slew31 (.A(net54),
    .Y(net53));
 BUFx16f_ASAP7_75t_R load_slew32 (.A(net55),
    .Y(net54));
 BUFx16f_ASAP7_75t_R load_slew33 (.A(net66),
    .Y(net55));
 BUFx16f_ASAP7_75t_R load_slew34 (.A(net60),
    .Y(net56));
 BUFx16f_ASAP7_75t_R load_slew35 (.A(net58),
    .Y(net57));
 BUFx16f_ASAP7_75t_R load_slew36 (.A(net2021),
    .Y(net58));
 BUFx10_ASAP7_75t_R load_slew37 (.A(net66),
    .Y(net59));
 BUFx16f_ASAP7_75t_R load_slew38 (.A(net66),
    .Y(net60));
 BUFx16f_ASAP7_75t_R load_slew39 (.A(net63),
    .Y(net61));
 BUFx16f_ASAP7_75t_R load_slew40 (.A(net63),
    .Y(net62));
 BUFx16f_ASAP7_75t_R load_slew41 (.A(net64),
    .Y(net63));
 BUFx24_ASAP7_75t_R load_slew42 (.A(net65),
    .Y(net64));
 BUFx16f_ASAP7_75t_R load_slew43 (.A(net66),
    .Y(net65));
 BUFx24_ASAP7_75t_R load_slew44 (.A(net74),
    .Y(net66));
 BUFx16f_ASAP7_75t_R load_slew45 (.A(net72),
    .Y(net67));
 BUFx16f_ASAP7_75t_R load_slew46 (.A(net70),
    .Y(net68));
 BUFx16f_ASAP7_75t_R load_slew47 (.A(net70),
    .Y(net69));
 BUFx16f_ASAP7_75t_R load_slew48 (.A(net72),
    .Y(net70));
 BUFx16f_ASAP7_75t_R load_slew49 (.A(net72),
    .Y(net71));
 BUFx16f_ASAP7_75t_R load_slew50 (.A(net73),
    .Y(net72));
 BUFx16f_ASAP7_75t_R load_slew51 (.A(net197),
    .Y(net73));
 BUFx24_ASAP7_75t_R load_slew52 (.A(net197),
    .Y(net74));
 BUFx2_ASAP7_75t_R input1 (.A(boot_addr_i[10]),
    .Y(net23));
 BUFx2_ASAP7_75t_R input2 (.A(boot_addr_i[11]),
    .Y(net24));
 BUFx2_ASAP7_75t_R input3 (.A(boot_addr_i[12]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input4 (.A(boot_addr_i[13]),
    .Y(net26));
 BUFx2_ASAP7_75t_R input5 (.A(boot_addr_i[14]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input6 (.A(boot_addr_i[15]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input7 (.A(boot_addr_i[16]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input8 (.A(boot_addr_i[17]),
    .Y(net30));
 BUFx2_ASAP7_75t_R input9 (.A(boot_addr_i[18]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input10 (.A(boot_addr_i[19]),
    .Y(net32));
 BUFx2_ASAP7_75t_R input11 (.A(boot_addr_i[20]),
    .Y(net33));
 BUFx2_ASAP7_75t_R input12 (.A(boot_addr_i[21]),
    .Y(net34));
 BUFx2_ASAP7_75t_R input13 (.A(boot_addr_i[22]),
    .Y(net35));
 BUFx2_ASAP7_75t_R input14 (.A(boot_addr_i[23]),
    .Y(net36));
 BUFx2_ASAP7_75t_R input15 (.A(boot_addr_i[24]),
    .Y(net37));
 BUFx2_ASAP7_75t_R input16 (.A(boot_addr_i[25]),
    .Y(net38));
 BUFx2_ASAP7_75t_R input17 (.A(boot_addr_i[26]),
    .Y(net39));
 BUFx2_ASAP7_75t_R input18 (.A(boot_addr_i[27]),
    .Y(net40));
 BUFx2_ASAP7_75t_R input19 (.A(boot_addr_i[28]),
    .Y(net41));
 BUFx2_ASAP7_75t_R input20 (.A(boot_addr_i[29]),
    .Y(net42));
 BUFx2_ASAP7_75t_R input21 (.A(boot_addr_i[30]),
    .Y(net43));
 BUFx2_ASAP7_75t_R input22 (.A(boot_addr_i[31]),
    .Y(net44));
 BUFx2_ASAP7_75t_R input23 (.A(boot_addr_i[8]),
    .Y(net45));
 BUFx2_ASAP7_75t_R input24 (.A(boot_addr_i[9]),
    .Y(net46));
 BUFx2_ASAP7_75t_R input25 (.A(data_err_i),
    .Y(net47));
 BUFx2_ASAP7_75t_R input26 (.A(data_rdata_i[0]),
    .Y(net48));
 BUFx2_ASAP7_75t_R input27 (.A(data_rdata_i[10]),
    .Y(net49));
 BUFx2_ASAP7_75t_R input28 (.A(data_rdata_i[11]),
    .Y(net50));
 BUFx2_ASAP7_75t_R input29 (.A(data_rdata_i[12]),
    .Y(net51));
 BUFx3_ASAP7_75t_R input30 (.A(data_rdata_i[13]),
    .Y(net75));
 BUFx3_ASAP7_75t_R input31 (.A(data_rdata_i[14]),
    .Y(net76));
 BUFx3_ASAP7_75t_R input32 (.A(data_rdata_i[15]),
    .Y(net77));
 BUFx2_ASAP7_75t_R input33 (.A(data_rdata_i[16]),
    .Y(net78));
 BUFx3_ASAP7_75t_R input34 (.A(data_rdata_i[17]),
    .Y(net79));
 BUFx3_ASAP7_75t_R input35 (.A(data_rdata_i[18]),
    .Y(net80));
 BUFx3_ASAP7_75t_R input36 (.A(data_rdata_i[19]),
    .Y(net81));
 BUFx4f_ASAP7_75t_R input37 (.A(data_rdata_i[1]),
    .Y(net82));
 BUFx3_ASAP7_75t_R input38 (.A(data_rdata_i[20]),
    .Y(net83));
 BUFx3_ASAP7_75t_R input39 (.A(data_rdata_i[21]),
    .Y(net84));
 BUFx2_ASAP7_75t_R input40 (.A(data_rdata_i[22]),
    .Y(net85));
 BUFx2_ASAP7_75t_R input41 (.A(data_rdata_i[23]),
    .Y(net86));
 BUFx2_ASAP7_75t_R input42 (.A(data_rdata_i[24]),
    .Y(net87));
 BUFx2_ASAP7_75t_R input43 (.A(data_rdata_i[25]),
    .Y(net88));
 BUFx2_ASAP7_75t_R input44 (.A(data_rdata_i[26]),
    .Y(net89));
 BUFx2_ASAP7_75t_R input45 (.A(data_rdata_i[27]),
    .Y(net90));
 BUFx2_ASAP7_75t_R input46 (.A(data_rdata_i[28]),
    .Y(net91));
 BUFx2_ASAP7_75t_R input47 (.A(data_rdata_i[29]),
    .Y(net92));
 BUFx3_ASAP7_75t_R input48 (.A(data_rdata_i[2]),
    .Y(net93));
 BUFx2_ASAP7_75t_R input49 (.A(data_rdata_i[30]),
    .Y(net94));
 BUFx4f_ASAP7_75t_R input50 (.A(data_rdata_i[31]),
    .Y(net96));
 BUFx2_ASAP7_75t_R input51 (.A(data_rdata_i[3]),
    .Y(net97));
 BUFx2_ASAP7_75t_R input52 (.A(data_rdata_i[4]),
    .Y(net98));
 BUFx2_ASAP7_75t_R input53 (.A(data_rdata_i[5]),
    .Y(net99));
 BUFx2_ASAP7_75t_R input54 (.A(data_rdata_i[6]),
    .Y(net100));
 BUFx2_ASAP7_75t_R input55 (.A(data_rdata_i[7]),
    .Y(net101));
 BUFx2_ASAP7_75t_R input56 (.A(data_rdata_i[8]),
    .Y(net102));
 BUFx2_ASAP7_75t_R input57 (.A(data_rdata_i[9]),
    .Y(net103));
 BUFx3_ASAP7_75t_R input58 (.A(data_rvalid_i),
    .Y(net104));
 BUFx4f_ASAP7_75t_R input59 (.A(debug_req_i),
    .Y(net105));
 BUFx2_ASAP7_75t_R input60 (.A(fetch_enable_i),
    .Y(net106));
 BUFx2_ASAP7_75t_R input61 (.A(hart_id_i[0]),
    .Y(net107));
 BUFx2_ASAP7_75t_R input62 (.A(hart_id_i[10]),
    .Y(net108));
 BUFx2_ASAP7_75t_R input63 (.A(hart_id_i[11]),
    .Y(net109));
 BUFx2_ASAP7_75t_R input64 (.A(hart_id_i[12]),
    .Y(net110));
 BUFx2_ASAP7_75t_R input65 (.A(hart_id_i[13]),
    .Y(net111));
 BUFx2_ASAP7_75t_R input66 (.A(hart_id_i[14]),
    .Y(net112));
 BUFx2_ASAP7_75t_R input67 (.A(hart_id_i[15]),
    .Y(net113));
 BUFx2_ASAP7_75t_R input68 (.A(hart_id_i[16]),
    .Y(net114));
 BUFx2_ASAP7_75t_R input69 (.A(hart_id_i[17]),
    .Y(net115));
 BUFx2_ASAP7_75t_R input70 (.A(hart_id_i[18]),
    .Y(net116));
 BUFx2_ASAP7_75t_R input71 (.A(hart_id_i[19]),
    .Y(net117));
 BUFx2_ASAP7_75t_R input72 (.A(hart_id_i[1]),
    .Y(net118));
 BUFx2_ASAP7_75t_R input73 (.A(hart_id_i[20]),
    .Y(net119));
 BUFx2_ASAP7_75t_R input74 (.A(hart_id_i[21]),
    .Y(net120));
 BUFx2_ASAP7_75t_R input75 (.A(hart_id_i[22]),
    .Y(net121));
 BUFx2_ASAP7_75t_R input76 (.A(hart_id_i[23]),
    .Y(net122));
 BUFx2_ASAP7_75t_R input77 (.A(hart_id_i[24]),
    .Y(net123));
 BUFx2_ASAP7_75t_R input78 (.A(hart_id_i[25]),
    .Y(net124));
 BUFx2_ASAP7_75t_R input79 (.A(hart_id_i[26]),
    .Y(net125));
 BUFx2_ASAP7_75t_R input80 (.A(hart_id_i[27]),
    .Y(net126));
 BUFx2_ASAP7_75t_R input81 (.A(hart_id_i[28]),
    .Y(net127));
 BUFx2_ASAP7_75t_R input82 (.A(hart_id_i[29]),
    .Y(net128));
 BUFx2_ASAP7_75t_R input83 (.A(hart_id_i[2]),
    .Y(net129));
 BUFx2_ASAP7_75t_R input84 (.A(hart_id_i[30]),
    .Y(net130));
 BUFx2_ASAP7_75t_R input85 (.A(hart_id_i[31]),
    .Y(net131));
 BUFx2_ASAP7_75t_R input86 (.A(hart_id_i[3]),
    .Y(net132));
 BUFx2_ASAP7_75t_R input87 (.A(hart_id_i[4]),
    .Y(net133));
 BUFx2_ASAP7_75t_R input88 (.A(hart_id_i[5]),
    .Y(net134));
 BUFx2_ASAP7_75t_R input89 (.A(hart_id_i[6]),
    .Y(net135));
 BUFx2_ASAP7_75t_R input90 (.A(hart_id_i[7]),
    .Y(net136));
 BUFx2_ASAP7_75t_R input91 (.A(hart_id_i[8]),
    .Y(net137));
 BUFx2_ASAP7_75t_R input92 (.A(hart_id_i[9]),
    .Y(net138));
 BUFx2_ASAP7_75t_R input93 (.A(instr_err_i),
    .Y(net139));
 BUFx2_ASAP7_75t_R input94 (.A(instr_gnt_i),
    .Y(net140));
 BUFx3_ASAP7_75t_R input95 (.A(instr_rdata_i[0]),
    .Y(net141));
 BUFx2_ASAP7_75t_R input96 (.A(instr_rdata_i[10]),
    .Y(net142));
 BUFx2_ASAP7_75t_R input97 (.A(instr_rdata_i[11]),
    .Y(net143));
 BUFx2_ASAP7_75t_R input98 (.A(instr_rdata_i[12]),
    .Y(net144));
 BUFx2_ASAP7_75t_R input99 (.A(instr_rdata_i[13]),
    .Y(net146));
 BUFx2_ASAP7_75t_R input100 (.A(instr_rdata_i[14]),
    .Y(net147));
 BUFx2_ASAP7_75t_R input101 (.A(instr_rdata_i[15]),
    .Y(net148));
 BUFx3_ASAP7_75t_R input102 (.A(instr_rdata_i[16]),
    .Y(net149));
 BUFx3_ASAP7_75t_R input103 (.A(instr_rdata_i[17]),
    .Y(net150));
 BUFx2_ASAP7_75t_R input104 (.A(instr_rdata_i[18]),
    .Y(net154));
 BUFx2_ASAP7_75t_R input105 (.A(instr_rdata_i[19]),
    .Y(net155));
 BUFx3_ASAP7_75t_R input106 (.A(instr_rdata_i[1]),
    .Y(net156));
 BUFx2_ASAP7_75t_R input107 (.A(instr_rdata_i[20]),
    .Y(net157));
 BUFx2_ASAP7_75t_R input108 (.A(instr_rdata_i[21]),
    .Y(net158));
 BUFx2_ASAP7_75t_R input109 (.A(instr_rdata_i[22]),
    .Y(net159));
 BUFx2_ASAP7_75t_R input110 (.A(instr_rdata_i[23]),
    .Y(net160));
 BUFx2_ASAP7_75t_R input111 (.A(instr_rdata_i[24]),
    .Y(net161));
 BUFx2_ASAP7_75t_R input112 (.A(instr_rdata_i[25]),
    .Y(net162));
 BUFx2_ASAP7_75t_R input113 (.A(instr_rdata_i[26]),
    .Y(net163));
 BUFx2_ASAP7_75t_R input114 (.A(instr_rdata_i[27]),
    .Y(net164));
 BUFx2_ASAP7_75t_R input115 (.A(instr_rdata_i[28]),
    .Y(net165));
 BUFx2_ASAP7_75t_R input116 (.A(instr_rdata_i[29]),
    .Y(net166));
 BUFx2_ASAP7_75t_R input117 (.A(instr_rdata_i[2]),
    .Y(net167));
 BUFx2_ASAP7_75t_R input118 (.A(instr_rdata_i[30]),
    .Y(net168));
 BUFx2_ASAP7_75t_R input119 (.A(instr_rdata_i[31]),
    .Y(net169));
 BUFx2_ASAP7_75t_R input120 (.A(instr_rdata_i[3]),
    .Y(net170));
 BUFx2_ASAP7_75t_R input121 (.A(instr_rdata_i[4]),
    .Y(net171));
 BUFx2_ASAP7_75t_R input122 (.A(instr_rdata_i[5]),
    .Y(net172));
 BUFx2_ASAP7_75t_R input123 (.A(instr_rdata_i[6]),
    .Y(net173));
 BUFx3_ASAP7_75t_R input124 (.A(instr_rdata_i[7]),
    .Y(net174));
 BUFx2_ASAP7_75t_R input125 (.A(instr_rdata_i[8]),
    .Y(net175));
 BUFx3_ASAP7_75t_R input126 (.A(instr_rdata_i[9]),
    .Y(net176));
 BUFx2_ASAP7_75t_R input127 (.A(instr_rvalid_i),
    .Y(net177));
 BUFx2_ASAP7_75t_R input128 (.A(irq_external_i),
    .Y(net178));
 BUFx2_ASAP7_75t_R input129 (.A(irq_fast_i[0]),
    .Y(net179));
 BUFx2_ASAP7_75t_R input130 (.A(irq_fast_i[10]),
    .Y(net180));
 BUFx2_ASAP7_75t_R input131 (.A(irq_fast_i[11]),
    .Y(net181));
 BUFx2_ASAP7_75t_R input132 (.A(irq_fast_i[12]),
    .Y(net182));
 BUFx2_ASAP7_75t_R input133 (.A(irq_fast_i[13]),
    .Y(net183));
 BUFx2_ASAP7_75t_R input134 (.A(irq_fast_i[14]),
    .Y(net184));
 BUFx2_ASAP7_75t_R input135 (.A(irq_fast_i[1]),
    .Y(net185));
 BUFx2_ASAP7_75t_R input136 (.A(irq_fast_i[2]),
    .Y(net186));
 BUFx2_ASAP7_75t_R input137 (.A(irq_fast_i[3]),
    .Y(net187));
 BUFx2_ASAP7_75t_R input138 (.A(irq_fast_i[4]),
    .Y(net188));
 BUFx2_ASAP7_75t_R input139 (.A(irq_fast_i[5]),
    .Y(net189));
 BUFx2_ASAP7_75t_R input140 (.A(irq_fast_i[6]),
    .Y(net190));
 BUFx2_ASAP7_75t_R input141 (.A(irq_fast_i[7]),
    .Y(net191));
 BUFx2_ASAP7_75t_R input142 (.A(irq_fast_i[8]),
    .Y(net192));
 BUFx2_ASAP7_75t_R input143 (.A(irq_fast_i[9]),
    .Y(net193));
 BUFx3_ASAP7_75t_R input144 (.A(irq_nm_i),
    .Y(net194));
 BUFx2_ASAP7_75t_R input145 (.A(irq_software_i),
    .Y(net195));
 BUFx2_ASAP7_75t_R input146 (.A(irq_timer_i),
    .Y(net196));
 BUFx8_ASAP7_75t_R input147 (.A(rst_ni),
    .Y(net197));
 BUFx2_ASAP7_75t_R input148 (.A(test_en_i),
    .Y(net198));
 BUFx2_ASAP7_75t_R output149 (.A(net199),
    .Y(core_sleep_o));
 BUFx2_ASAP7_75t_R output150 (.A(net200),
    .Y(data_addr_o[10]));
 BUFx2_ASAP7_75t_R output151 (.A(net201),
    .Y(data_addr_o[11]));
 BUFx2_ASAP7_75t_R output152 (.A(net202),
    .Y(data_addr_o[12]));
 BUFx2_ASAP7_75t_R output153 (.A(net203),
    .Y(data_addr_o[13]));
 BUFx2_ASAP7_75t_R output154 (.A(net204),
    .Y(data_addr_o[14]));
 BUFx2_ASAP7_75t_R output155 (.A(net205),
    .Y(data_addr_o[15]));
 BUFx2_ASAP7_75t_R output156 (.A(net206),
    .Y(data_addr_o[16]));
 BUFx2_ASAP7_75t_R output157 (.A(net207),
    .Y(data_addr_o[17]));
 BUFx2_ASAP7_75t_R output158 (.A(net208),
    .Y(data_addr_o[18]));
 BUFx2_ASAP7_75t_R output159 (.A(net209),
    .Y(data_addr_o[19]));
 BUFx2_ASAP7_75t_R output160 (.A(net210),
    .Y(data_addr_o[20]));
 BUFx2_ASAP7_75t_R output161 (.A(net211),
    .Y(data_addr_o[21]));
 BUFx2_ASAP7_75t_R output162 (.A(net212),
    .Y(data_addr_o[22]));
 BUFx2_ASAP7_75t_R output163 (.A(net213),
    .Y(data_addr_o[23]));
 BUFx2_ASAP7_75t_R output164 (.A(net214),
    .Y(data_addr_o[24]));
 BUFx2_ASAP7_75t_R output165 (.A(net215),
    .Y(data_addr_o[25]));
 BUFx2_ASAP7_75t_R output166 (.A(net216),
    .Y(data_addr_o[26]));
 BUFx2_ASAP7_75t_R output167 (.A(net217),
    .Y(data_addr_o[27]));
 BUFx2_ASAP7_75t_R output168 (.A(net218),
    .Y(data_addr_o[28]));
 BUFx2_ASAP7_75t_R output169 (.A(net219),
    .Y(data_addr_o[29]));
 BUFx2_ASAP7_75t_R output170 (.A(net220),
    .Y(data_addr_o[2]));
 BUFx2_ASAP7_75t_R output171 (.A(net221),
    .Y(data_addr_o[30]));
 BUFx2_ASAP7_75t_R output172 (.A(net222),
    .Y(data_addr_o[31]));
 BUFx2_ASAP7_75t_R output173 (.A(net223),
    .Y(data_addr_o[3]));
 BUFx2_ASAP7_75t_R output174 (.A(net224),
    .Y(data_addr_o[4]));
 BUFx2_ASAP7_75t_R output175 (.A(net225),
    .Y(data_addr_o[5]));
 BUFx2_ASAP7_75t_R output176 (.A(net226),
    .Y(data_addr_o[6]));
 BUFx2_ASAP7_75t_R output177 (.A(net227),
    .Y(data_addr_o[7]));
 BUFx2_ASAP7_75t_R output178 (.A(net228),
    .Y(data_addr_o[8]));
 BUFx2_ASAP7_75t_R output179 (.A(net229),
    .Y(data_addr_o[9]));
 BUFx2_ASAP7_75t_R output180 (.A(net230),
    .Y(data_be_o[0]));
 BUFx2_ASAP7_75t_R output181 (.A(net231),
    .Y(data_be_o[1]));
 BUFx2_ASAP7_75t_R output182 (.A(net232),
    .Y(data_be_o[2]));
 BUFx2_ASAP7_75t_R output183 (.A(net233),
    .Y(data_be_o[3]));
 BUFx2_ASAP7_75t_R output184 (.A(net234),
    .Y(data_req_o));
 BUFx2_ASAP7_75t_R output185 (.A(net235),
    .Y(data_wdata_o[0]));
 BUFx2_ASAP7_75t_R output186 (.A(net236),
    .Y(data_wdata_o[10]));
 BUFx2_ASAP7_75t_R output187 (.A(net237),
    .Y(data_wdata_o[11]));
 BUFx2_ASAP7_75t_R output188 (.A(net238),
    .Y(data_wdata_o[12]));
 BUFx2_ASAP7_75t_R output189 (.A(net239),
    .Y(data_wdata_o[13]));
 BUFx2_ASAP7_75t_R output190 (.A(net240),
    .Y(data_wdata_o[14]));
 BUFx2_ASAP7_75t_R output191 (.A(net241),
    .Y(data_wdata_o[15]));
 BUFx2_ASAP7_75t_R output192 (.A(net242),
    .Y(data_wdata_o[16]));
 BUFx2_ASAP7_75t_R output193 (.A(net243),
    .Y(data_wdata_o[17]));
 BUFx2_ASAP7_75t_R output194 (.A(net244),
    .Y(data_wdata_o[18]));
 BUFx2_ASAP7_75t_R output195 (.A(net245),
    .Y(data_wdata_o[19]));
 BUFx2_ASAP7_75t_R output196 (.A(net246),
    .Y(data_wdata_o[1]));
 BUFx2_ASAP7_75t_R output197 (.A(net247),
    .Y(data_wdata_o[20]));
 BUFx2_ASAP7_75t_R output198 (.A(net248),
    .Y(data_wdata_o[21]));
 BUFx2_ASAP7_75t_R output199 (.A(net249),
    .Y(data_wdata_o[22]));
 BUFx2_ASAP7_75t_R output200 (.A(net250),
    .Y(data_wdata_o[23]));
 BUFx2_ASAP7_75t_R output201 (.A(net251),
    .Y(data_wdata_o[24]));
 BUFx2_ASAP7_75t_R output202 (.A(net252),
    .Y(data_wdata_o[25]));
 BUFx2_ASAP7_75t_R output203 (.A(net253),
    .Y(data_wdata_o[26]));
 BUFx2_ASAP7_75t_R output204 (.A(net254),
    .Y(data_wdata_o[27]));
 BUFx2_ASAP7_75t_R output205 (.A(net255),
    .Y(data_wdata_o[28]));
 BUFx2_ASAP7_75t_R output206 (.A(net256),
    .Y(data_wdata_o[29]));
 BUFx2_ASAP7_75t_R output207 (.A(net257),
    .Y(data_wdata_o[2]));
 BUFx2_ASAP7_75t_R output208 (.A(net258),
    .Y(data_wdata_o[30]));
 BUFx2_ASAP7_75t_R output209 (.A(net259),
    .Y(data_wdata_o[31]));
 BUFx2_ASAP7_75t_R output210 (.A(net260),
    .Y(data_wdata_o[3]));
 BUFx2_ASAP7_75t_R output211 (.A(net261),
    .Y(data_wdata_o[4]));
 BUFx2_ASAP7_75t_R output212 (.A(net262),
    .Y(data_wdata_o[5]));
 BUFx2_ASAP7_75t_R output213 (.A(net263),
    .Y(data_wdata_o[6]));
 BUFx2_ASAP7_75t_R output214 (.A(net264),
    .Y(data_wdata_o[7]));
 BUFx2_ASAP7_75t_R output215 (.A(net265),
    .Y(data_wdata_o[8]));
 BUFx2_ASAP7_75t_R output216 (.A(net266),
    .Y(data_wdata_o[9]));
 BUFx2_ASAP7_75t_R output217 (.A(net267),
    .Y(data_we_o));
 BUFx2_ASAP7_75t_R output218 (.A(net268),
    .Y(instr_addr_o[10]));
 BUFx2_ASAP7_75t_R output219 (.A(net269),
    .Y(instr_addr_o[11]));
 BUFx2_ASAP7_75t_R output220 (.A(net270),
    .Y(instr_addr_o[12]));
 BUFx2_ASAP7_75t_R output221 (.A(net271),
    .Y(instr_addr_o[13]));
 BUFx2_ASAP7_75t_R output222 (.A(net272),
    .Y(instr_addr_o[14]));
 BUFx2_ASAP7_75t_R output223 (.A(net273),
    .Y(instr_addr_o[15]));
 BUFx2_ASAP7_75t_R output224 (.A(net274),
    .Y(instr_addr_o[16]));
 BUFx2_ASAP7_75t_R output225 (.A(net275),
    .Y(instr_addr_o[17]));
 BUFx2_ASAP7_75t_R output226 (.A(net276),
    .Y(instr_addr_o[18]));
 BUFx2_ASAP7_75t_R output227 (.A(net277),
    .Y(instr_addr_o[19]));
 BUFx2_ASAP7_75t_R output228 (.A(net278),
    .Y(instr_addr_o[20]));
 BUFx2_ASAP7_75t_R output229 (.A(net279),
    .Y(instr_addr_o[21]));
 BUFx2_ASAP7_75t_R output230 (.A(net280),
    .Y(instr_addr_o[22]));
 BUFx2_ASAP7_75t_R output231 (.A(net281),
    .Y(instr_addr_o[23]));
 BUFx2_ASAP7_75t_R output232 (.A(net282),
    .Y(instr_addr_o[24]));
 BUFx2_ASAP7_75t_R output233 (.A(net283),
    .Y(instr_addr_o[25]));
 BUFx2_ASAP7_75t_R output234 (.A(net284),
    .Y(instr_addr_o[26]));
 BUFx2_ASAP7_75t_R output235 (.A(net285),
    .Y(instr_addr_o[27]));
 BUFx2_ASAP7_75t_R output236 (.A(net286),
    .Y(instr_addr_o[28]));
 BUFx2_ASAP7_75t_R output237 (.A(net287),
    .Y(instr_addr_o[29]));
 BUFx2_ASAP7_75t_R output238 (.A(net288),
    .Y(instr_addr_o[2]));
 BUFx2_ASAP7_75t_R output239 (.A(net289),
    .Y(instr_addr_o[30]));
 BUFx3_ASAP7_75t_R output240 (.A(net290),
    .Y(instr_addr_o[31]));
 BUFx2_ASAP7_75t_R output241 (.A(net291),
    .Y(instr_addr_o[3]));
 BUFx2_ASAP7_75t_R output242 (.A(net292),
    .Y(instr_addr_o[4]));
 BUFx2_ASAP7_75t_R output243 (.A(net293),
    .Y(instr_addr_o[5]));
 BUFx2_ASAP7_75t_R output244 (.A(net294),
    .Y(instr_addr_o[6]));
 BUFx2_ASAP7_75t_R output245 (.A(net295),
    .Y(instr_addr_o[7]));
 BUFx2_ASAP7_75t_R output246 (.A(net296),
    .Y(instr_addr_o[8]));
 BUFx2_ASAP7_75t_R output247 (.A(net297),
    .Y(instr_addr_o[9]));
 BUFx2_ASAP7_75t_R output248 (.A(net298),
    .Y(instr_req_o));
 TIELOx1_ASAP7_75t_R _35803__249 (.L(net299));
 TIELOx1_ASAP7_75t_R _35804__250 (.L(net300));
 TIELOx1_ASAP7_75t_R _35805__251 (.L(net301));
 TIELOx1_ASAP7_75t_R _35806__252 (.L(net302));
 TIELOx1_ASAP7_75t_R _35837__253 (.L(net303));
 TIELOx1_ASAP7_75t_R _35838__254 (.L(net304));
 TIEHIx1_ASAP7_75t_R _35795__256 (.H(net306));
 TIEHIx1_ASAP7_75t_R _35796__257 (.H(net307));
 TIEHIx1_ASAP7_75t_R _35797__258 (.H(net308));
 TIEHIx1_ASAP7_75t_R _35798__259 (.H(net309));
 TIEHIx1_ASAP7_75t_R _35799__260 (.H(net310));
 TIEHIx1_ASAP7_75t_R _35800__261 (.H(net311));
 TIEHIx1_ASAP7_75t_R \core_busy_q$_DFF_PN0__262  (.H(net312));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P__263  (.H(net313));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P__264  (.H(net314));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[0]$_DFFE_PN0P__265  (.H(net315));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[10]$_DFFE_PN0P__266  (.H(net316));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[11]$_DFFE_PN0P__267  (.H(net317));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[12]$_DFFE_PN0P__268  (.H(net318));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[13]$_DFFE_PN0P__269  (.H(net319));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[14]$_DFFE_PN0P__270  (.H(net320));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[15]$_DFFE_PN0P__271  (.H(net321));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[16]$_DFFE_PN0P__272  (.H(net322));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[17]$_DFFE_PN0P__273  (.H(net323));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[18]$_DFFE_PN0P__274  (.H(net324));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[19]$_DFFE_PN0P__275  (.H(net325));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[1]$_DFFE_PN0P__276  (.H(net326));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[20]$_DFFE_PN0P__277  (.H(net327));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[21]$_DFFE_PN0P__278  (.H(net328));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[22]$_DFFE_PN0P__279  (.H(net329));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[23]$_DFFE_PN0P__280  (.H(net330));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[24]$_DFFE_PN0P__281  (.H(net331));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[25]$_DFFE_PN0P__282  (.H(net332));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[26]$_DFFE_PN0P__283  (.H(net333));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[27]$_DFFE_PN0P__284  (.H(net334));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[28]$_DFFE_PN0P__285  (.H(net335));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[29]$_DFFE_PN0P__286  (.H(net336));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[2]$_DFFE_PN0P__287  (.H(net337));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[30]$_DFFE_PN0P__288  (.H(net338));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[31]$_DFFE_PN0P__289  (.H(net339));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[32]$_DFFE_PN0P__290  (.H(net340));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[33]$_DFFE_PN0P__291  (.H(net341));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[34]$_DFFE_PN0P__292  (.H(net342));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[35]$_DFFE_PN0P__293  (.H(net343));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[36]$_DFFE_PN0P__294  (.H(net344));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[37]$_DFFE_PN0P__295  (.H(net345));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[38]$_DFFE_PN0P__296  (.H(net346));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[39]$_DFFE_PN0P__297  (.H(net347));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[3]$_DFFE_PN0P__298  (.H(net348));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[40]$_DFFE_PN0P__299  (.H(net349));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[41]$_DFFE_PN0P__300  (.H(net350));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[42]$_DFFE_PN0P__301  (.H(net351));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[43]$_DFFE_PN0P__302  (.H(net352));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[44]$_DFFE_PN0P__303  (.H(net353));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[45]$_DFFE_PN0P__304  (.H(net354));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[46]$_DFFE_PN0P__305  (.H(net355));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[47]$_DFFE_PN0P__306  (.H(net356));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[48]$_DFFE_PN0P__307  (.H(net357));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[49]$_DFFE_PN0P__308  (.H(net358));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[4]$_DFFE_PN0P__309  (.H(net359));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[50]$_DFFE_PN0P__310  (.H(net360));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[51]$_DFFE_PN0P__311  (.H(net361));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[52]$_DFFE_PN0P__312  (.H(net362));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[53]$_DFFE_PN0P__313  (.H(net363));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[54]$_DFFE_PN0P__314  (.H(net364));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[55]$_DFFE_PN0P__315  (.H(net365));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[56]$_DFFE_PN0P__316  (.H(net366));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[57]$_DFFE_PN0P__317  (.H(net367));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[58]$_DFFE_PN0P__318  (.H(net368));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[59]$_DFFE_PN0P__319  (.H(net369));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[5]$_DFFE_PN0P__320  (.H(net370));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[60]$_DFFE_PN0P__321  (.H(net371));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[61]$_DFFE_PN0P__322  (.H(net372));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[62]$_DFFE_PN0P__323  (.H(net373));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[63]$_DFFE_PN0P__324  (.H(net374));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[6]$_DFFE_PN0P__325  (.H(net375));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[7]$_DFFE_PN0P__326  (.H(net376));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[8]$_DFFE_PN0P__327  (.H(net377));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.mcycle_counter_i.counter_q[9]$_DFFE_PN0P__328  (.H(net378));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[0]$_DFFE_PN0P__329  (.H(net379));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[10]$_DFFE_PN0P__330  (.H(net380));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[11]$_DFFE_PN0P__331  (.H(net381));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[12]$_DFFE_PN0P__332  (.H(net382));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[13]$_DFFE_PN0P__333  (.H(net383));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[14]$_DFFE_PN0P__334  (.H(net384));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[15]$_DFFE_PN0P__335  (.H(net385));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[16]$_DFFE_PN0P__336  (.H(net386));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[17]$_DFFE_PN0P__337  (.H(net387));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[18]$_DFFE_PN0P__338  (.H(net388));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[19]$_DFFE_PN0P__339  (.H(net389));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[1]$_DFFE_PN0P__340  (.H(net390));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[20]$_DFFE_PN0P__341  (.H(net391));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[21]$_DFFE_PN0P__342  (.H(net392));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[22]$_DFFE_PN0P__343  (.H(net393));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[23]$_DFFE_PN0P__344  (.H(net394));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[24]$_DFFE_PN0P__345  (.H(net395));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[25]$_DFFE_PN0P__346  (.H(net396));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[26]$_DFFE_PN0P__347  (.H(net397));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[27]$_DFFE_PN0P__348  (.H(net398));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[28]$_DFFE_PN0P__349  (.H(net399));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[29]$_DFFE_PN0P__350  (.H(net400));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[2]$_DFFE_PN0P__351  (.H(net401));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[30]$_DFFE_PN0P__352  (.H(net402));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[31]$_DFFE_PN0P__353  (.H(net403));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[32]$_DFFE_PN0P__354  (.H(net404));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[33]$_DFFE_PN0P__355  (.H(net405));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[34]$_DFFE_PN0P__356  (.H(net406));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[35]$_DFFE_PN0P__357  (.H(net407));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[36]$_DFFE_PN0P__358  (.H(net408));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[37]$_DFFE_PN0P__359  (.H(net409));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[38]$_DFFE_PN0P__360  (.H(net410));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[39]$_DFFE_PN0P__361  (.H(net411));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[3]$_DFFE_PN0P__362  (.H(net412));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[40]$_DFFE_PN0P__363  (.H(net413));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[41]$_DFFE_PN0P__364  (.H(net414));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[42]$_DFFE_PN0P__365  (.H(net415));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[43]$_DFFE_PN0P__366  (.H(net416));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[44]$_DFFE_PN0P__367  (.H(net417));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[45]$_DFFE_PN0P__368  (.H(net418));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[46]$_DFFE_PN0P__369  (.H(net419));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[47]$_DFFE_PN0P__370  (.H(net420));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[48]$_DFFE_PN0P__371  (.H(net421));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[49]$_DFFE_PN0P__372  (.H(net422));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[4]$_DFFE_PN0P__373  (.H(net423));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[50]$_DFFE_PN0P__374  (.H(net424));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[51]$_DFFE_PN0P__375  (.H(net425));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[52]$_DFFE_PN0P__376  (.H(net426));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[53]$_DFFE_PN0P__377  (.H(net427));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[54]$_DFFE_PN0P__378  (.H(net428));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[55]$_DFFE_PN0P__379  (.H(net429));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[56]$_DFFE_PN0P__380  (.H(net430));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[57]$_DFFE_PN0P__381  (.H(net431));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[58]$_DFFE_PN0P__382  (.H(net432));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[59]$_DFFE_PN0P__383  (.H(net433));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[5]$_DFFE_PN0P__384  (.H(net434));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[60]$_DFFE_PN0P__385  (.H(net435));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[61]$_DFFE_PN0P__386  (.H(net436));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[62]$_DFFE_PN0P__387  (.H(net437));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[63]$_DFFE_PN0P__388  (.H(net438));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[6]$_DFFE_PN0P__389  (.H(net439));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[7]$_DFFE_PN0P__390  (.H(net440));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[8]$_DFFE_PN0P__391  (.H(net441));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.minstret_counter_i.counter_q[9]$_DFFE_PN0P__392  (.H(net442));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.priv_lvl_q[0]$_DFFE_PN1P__393  (.H(net443));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.priv_lvl_q[1]$_DFFE_PN1P__394  (.H(net444));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[0]$_DFFE_PN1N__395  (.H(net445));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[11]$_DFFE_PN0P__396  (.H(net446));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[12]$_DFFE_PN0P__397  (.H(net447));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[13]$_DFFE_PN0P__398  (.H(net448));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[15]$_DFFE_PN0P__399  (.H(net449));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[1]$_DFFE_PN1N__400  (.H(net450));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[2]$_DFFE_PN0P__401  (.H(net451));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[6]$_DFFE_PN0P__402  (.H(net452));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[7]$_DFFE_PN0P__403  (.H(net453));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dcsr_csr.rdata_q[8]$_DFFE_PN0P__404  (.H(net454));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[10]$_DFFE_PN0P__405  (.H(net455));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[11]$_DFFE_PN0P__406  (.H(net456));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[12]$_DFFE_PN0P__407  (.H(net457));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[13]$_DFFE_PN0P__408  (.H(net458));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[14]$_DFFE_PN0P__409  (.H(net459));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[15]$_DFFE_PN0P__410  (.H(net460));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[16]$_DFFE_PN0P__411  (.H(net461));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[17]$_DFFE_PN0P__412  (.H(net462));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[18]$_DFFE_PN0P__413  (.H(net463));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[19]$_DFFE_PN0P__414  (.H(net464));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[1]$_DFFE_PN0P__415  (.H(net465));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[20]$_DFFE_PN0P__416  (.H(net466));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[21]$_DFFE_PN0P__417  (.H(net467));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[22]$_DFFE_PN0P__418  (.H(net468));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[23]$_DFFE_PN0P__419  (.H(net469));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[24]$_DFFE_PN0P__420  (.H(net470));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[25]$_DFFE_PN0P__421  (.H(net471));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[26]$_DFFE_PN0P__422  (.H(net472));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[27]$_DFFE_PN0P__423  (.H(net473));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[28]$_DFFE_PN0P__424  (.H(net474));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[29]$_DFFE_PN0P__425  (.H(net475));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[2]$_DFFE_PN0P__426  (.H(net476));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[30]$_DFFE_PN0P__427  (.H(net477));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[31]$_DFFE_PN0P__428  (.H(net478));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[3]$_DFFE_PN0P__429  (.H(net479));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[4]$_DFFE_PN0P__430  (.H(net480));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[5]$_DFFE_PN0P__431  (.H(net481));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[6]$_DFFE_PN0P__432  (.H(net482));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[7]$_DFFE_PN0P__433  (.H(net483));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[8]$_DFFE_PN0P__434  (.H(net484));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_depc_csr.rdata_q[9]$_DFFE_PN0P__435  (.H(net485));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[0]$_DFFE_PN0P__436  (.H(net486));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[10]$_DFFE_PN0P__437  (.H(net487));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[11]$_DFFE_PN0P__438  (.H(net488));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[12]$_DFFE_PN0P__439  (.H(net489));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[13]$_DFFE_PN0P__440  (.H(net490));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[14]$_DFFE_PN0P__441  (.H(net491));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[15]$_DFFE_PN0P__442  (.H(net492));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[16]$_DFFE_PN0P__443  (.H(net493));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[17]$_DFFE_PN0P__444  (.H(net494));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[18]$_DFFE_PN0P__445  (.H(net495));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[19]$_DFFE_PN0P__446  (.H(net496));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[1]$_DFFE_PN0P__447  (.H(net497));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[20]$_DFFE_PN0P__448  (.H(net498));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[21]$_DFFE_PN0P__449  (.H(net499));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[22]$_DFFE_PN0P__450  (.H(net500));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[23]$_DFFE_PN0P__451  (.H(net501));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[24]$_DFFE_PN0P__452  (.H(net502));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[25]$_DFFE_PN0P__453  (.H(net503));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[26]$_DFFE_PN0P__454  (.H(net504));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[27]$_DFFE_PN0P__455  (.H(net505));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[28]$_DFFE_PN0P__456  (.H(net506));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[29]$_DFFE_PN0P__457  (.H(net507));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[2]$_DFFE_PN0P__458  (.H(net508));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[30]$_DFFE_PN0P__459  (.H(net509));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[31]$_DFFE_PN0P__460  (.H(net510));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[3]$_DFFE_PN0P__461  (.H(net511));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[4]$_DFFE_PN0P__462  (.H(net512));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[5]$_DFFE_PN0P__463  (.H(net513));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[6]$_DFFE_PN0P__464  (.H(net514));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[7]$_DFFE_PN0P__465  (.H(net515));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[8]$_DFFE_PN0P__466  (.H(net516));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch0_csr.rdata_q[9]$_DFFE_PN0P__467  (.H(net517));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[0]$_DFFE_PN0P__468  (.H(net518));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[10]$_DFFE_PN0P__469  (.H(net519));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[11]$_DFFE_PN0P__470  (.H(net520));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[12]$_DFFE_PN0P__471  (.H(net521));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[13]$_DFFE_PN0P__472  (.H(net522));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[14]$_DFFE_PN0P__473  (.H(net523));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[15]$_DFFE_PN0P__474  (.H(net524));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[16]$_DFFE_PN0P__475  (.H(net525));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[17]$_DFFE_PN0P__476  (.H(net526));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[18]$_DFFE_PN0P__477  (.H(net527));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[19]$_DFFE_PN0P__478  (.H(net528));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[1]$_DFFE_PN0P__479  (.H(net529));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[20]$_DFFE_PN0P__480  (.H(net530));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[21]$_DFFE_PN0P__481  (.H(net531));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[22]$_DFFE_PN0P__482  (.H(net532));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[23]$_DFFE_PN0P__483  (.H(net533));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[24]$_DFFE_PN0P__484  (.H(net534));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[25]$_DFFE_PN0P__485  (.H(net535));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[26]$_DFFE_PN0P__486  (.H(net536));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[27]$_DFFE_PN0P__487  (.H(net537));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[28]$_DFFE_PN0P__488  (.H(net538));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[29]$_DFFE_PN0P__489  (.H(net539));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[2]$_DFFE_PN0P__490  (.H(net540));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[30]$_DFFE_PN0P__491  (.H(net541));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[31]$_DFFE_PN0P__492  (.H(net542));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[3]$_DFFE_PN0P__493  (.H(net543));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[4]$_DFFE_PN0P__494  (.H(net544));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[5]$_DFFE_PN0P__495  (.H(net545));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[6]$_DFFE_PN0P__496  (.H(net546));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[7]$_DFFE_PN0P__497  (.H(net547));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[8]$_DFFE_PN0P__498  (.H(net548));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_dscratch1_csr.rdata_q[9]$_DFFE_PN0P__499  (.H(net549));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[0]$_DFFE_PN0P__500  (.H(net550));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[1]$_DFFE_PN0P__501  (.H(net551));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[2]$_DFFE_PN0P__502  (.H(net552));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[3]$_DFFE_PN0P__503  (.H(net553));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[4]$_DFFE_PN0P__504  (.H(net554));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mcause_csr.rdata_q[5]$_DFFE_PN0P__505  (.H(net555));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[0]$_DFFE_PN0P__506  (.H(net556));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[10]$_DFFE_PN0P__507  (.H(net557));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[11]$_DFFE_PN0P__508  (.H(net558));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[12]$_DFFE_PN0P__509  (.H(net559));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[13]$_DFFE_PN0P__510  (.H(net560));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[14]$_DFFE_PN0P__511  (.H(net561));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[15]$_DFFE_PN0P__512  (.H(net562));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[16]$_DFFE_PN0P__513  (.H(net563));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[17]$_DFFE_PN0P__514  (.H(net564));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[18]$_DFFE_PN0P__515  (.H(net565));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[19]$_DFFE_PN0P__516  (.H(net566));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[1]$_DFFE_PN0P__517  (.H(net567));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[20]$_DFFE_PN0P__518  (.H(net568));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[21]$_DFFE_PN0P__519  (.H(net569));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[22]$_DFFE_PN0P__520  (.H(net570));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[23]$_DFFE_PN0P__521  (.H(net571));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[24]$_DFFE_PN0P__522  (.H(net572));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[25]$_DFFE_PN0P__523  (.H(net573));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[26]$_DFFE_PN0P__524  (.H(net574));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[27]$_DFFE_PN0P__525  (.H(net575));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[28]$_DFFE_PN0P__526  (.H(net576));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[29]$_DFFE_PN0P__527  (.H(net577));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[2]$_DFFE_PN0P__528  (.H(net578));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[30]$_DFFE_PN0P__529  (.H(net579));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[31]$_DFFE_PN0P__530  (.H(net580));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[3]$_DFFE_PN0P__531  (.H(net581));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[4]$_DFFE_PN0P__532  (.H(net582));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[5]$_DFFE_PN0P__533  (.H(net583));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[6]$_DFFE_PN0P__534  (.H(net584));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[7]$_DFFE_PN0P__535  (.H(net585));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[8]$_DFFE_PN0P__536  (.H(net586));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mepc_csr.rdata_q[9]$_DFFE_PN0P__537  (.H(net587));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[0]$_DFFE_PN0P__538  (.H(net588));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[10]$_DFFE_PN0P__539  (.H(net589));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[11]$_DFFE_PN0P__540  (.H(net590));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[12]$_DFFE_PN0P__541  (.H(net591));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[13]$_DFFE_PN0P__542  (.H(net592));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[14]$_DFFE_PN0P__543  (.H(net593));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[15]$_DFFE_PN0P__544  (.H(net594));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[16]$_DFFE_PN0P__545  (.H(net595));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[17]$_DFFE_PN0P__546  (.H(net596));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[1]$_DFFE_PN0P__547  (.H(net597));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[2]$_DFFE_PN0P__548  (.H(net598));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[3]$_DFFE_PN0P__549  (.H(net599));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[4]$_DFFE_PN0P__550  (.H(net600));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[5]$_DFFE_PN0P__551  (.H(net601));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[6]$_DFFE_PN0P__552  (.H(net602));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[7]$_DFFE_PN0P__553  (.H(net603));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[8]$_DFFE_PN0P__554  (.H(net604));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mie_csr.rdata_q[9]$_DFFE_PN0P__555  (.H(net605));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[0]$_DFFE_PN0P__556  (.H(net606));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[10]$_DFFE_PN0P__557  (.H(net607));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[11]$_DFFE_PN0P__558  (.H(net608));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[12]$_DFFE_PN0P__559  (.H(net609));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[13]$_DFFE_PN0P__560  (.H(net610));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[14]$_DFFE_PN0P__561  (.H(net611));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[15]$_DFFE_PN0P__562  (.H(net612));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[16]$_DFFE_PN0P__563  (.H(net613));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[17]$_DFFE_PN0P__564  (.H(net614));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[18]$_DFFE_PN0P__565  (.H(net615));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[19]$_DFFE_PN0P__566  (.H(net616));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[1]$_DFFE_PN0P__567  (.H(net617));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[20]$_DFFE_PN0P__568  (.H(net618));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[21]$_DFFE_PN0P__569  (.H(net619));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[22]$_DFFE_PN0P__570  (.H(net620));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[23]$_DFFE_PN0P__571  (.H(net621));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[24]$_DFFE_PN0P__572  (.H(net622));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[25]$_DFFE_PN0P__573  (.H(net623));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[26]$_DFFE_PN0P__574  (.H(net624));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[27]$_DFFE_PN0P__575  (.H(net625));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[28]$_DFFE_PN0P__576  (.H(net626));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[29]$_DFFE_PN0P__577  (.H(net627));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[2]$_DFFE_PN0P__578  (.H(net628));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[30]$_DFFE_PN0P__579  (.H(net629));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[31]$_DFFE_PN0P__580  (.H(net630));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[3]$_DFFE_PN0P__581  (.H(net631));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[4]$_DFFE_PN0P__582  (.H(net632));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[5]$_DFFE_PN0P__583  (.H(net633));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[6]$_DFFE_PN0P__584  (.H(net634));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[7]$_DFFE_PN0P__585  (.H(net635));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[8]$_DFFE_PN0P__586  (.H(net636));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mscratch_csr.rdata_q[9]$_DFFE_PN0P__587  (.H(net637));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[0]$_DFFE_PN0P__588  (.H(net638));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[1]$_DFFE_PN0P__589  (.H(net639));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[2]$_DFFE_PN0P__590  (.H(net640));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[3]$_DFFE_PN0P__591  (.H(net641));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[4]$_DFFE_PN0P__592  (.H(net642));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_cause_csr.rdata_q[5]$_DFFE_PN0P__593  (.H(net643));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rdata_q[0]$_DFFE_PN0P__594  (.H(net644));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rdata_q[1]$_DFFE_PN0P__595  (.H(net645));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_csr.rdata_q[2]$_DFFE_PN1P__596  (.H(net646));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[0]$_DFFE_PN0P__597  (.H(net647));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[10]$_DFFE_PN0P__598  (.H(net648));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[11]$_DFFE_PN0P__599  (.H(net649));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[12]$_DFFE_PN0P__600  (.H(net650));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[13]$_DFFE_PN0P__601  (.H(net651));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[14]$_DFFE_PN0P__602  (.H(net652));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[15]$_DFFE_PN0P__603  (.H(net653));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[16]$_DFFE_PN0P__604  (.H(net654));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[17]$_DFFE_PN0P__605  (.H(net655));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[18]$_DFFE_PN0P__606  (.H(net656));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[19]$_DFFE_PN0P__607  (.H(net657));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[1]$_DFFE_PN0P__608  (.H(net658));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[20]$_DFFE_PN0P__609  (.H(net659));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[21]$_DFFE_PN0P__610  (.H(net660));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[22]$_DFFE_PN0P__611  (.H(net661));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[23]$_DFFE_PN0P__612  (.H(net662));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[24]$_DFFE_PN0P__613  (.H(net663));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[25]$_DFFE_PN0P__614  (.H(net664));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[26]$_DFFE_PN0P__615  (.H(net665));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[27]$_DFFE_PN0P__616  (.H(net666));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[28]$_DFFE_PN0P__617  (.H(net667));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[29]$_DFFE_PN0P__618  (.H(net668));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[2]$_DFFE_PN0P__619  (.H(net669));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[30]$_DFFE_PN0P__620  (.H(net670));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[31]$_DFFE_PN0P__621  (.H(net671));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[3]$_DFFE_PN0P__622  (.H(net672));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[4]$_DFFE_PN0P__623  (.H(net673));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[5]$_DFFE_PN0P__624  (.H(net674));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[6]$_DFFE_PN0P__625  (.H(net675));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[7]$_DFFE_PN0P__626  (.H(net676));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[8]$_DFFE_PN0P__627  (.H(net677));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstack_epc_csr.rdata_q[9]$_DFFE_PN0P__628  (.H(net678));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[0]$_DFFE_PN0P__629  (.H(net679));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[1]$_DFFE_PN0P__630  (.H(net680));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[2]$_DFFE_PN0P__631  (.H(net681));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[3]$_DFFE_PN0P__632  (.H(net682));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[4]$_DFFE_PN1P__633  (.H(net683));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mstatus_csr.rdata_q[5]$_DFFE_PN0P__634  (.H(net684));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[0]$_DFFE_PN0P__635  (.H(net685));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[10]$_DFFE_PN0P__636  (.H(net686));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[11]$_DFFE_PN0P__637  (.H(net687));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[12]$_DFFE_PN0P__638  (.H(net688));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[13]$_DFFE_PN0P__639  (.H(net689));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[14]$_DFFE_PN0P__640  (.H(net690));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[15]$_DFFE_PN0P__641  (.H(net691));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[16]$_DFFE_PN0P__642  (.H(net692));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[17]$_DFFE_PN0P__643  (.H(net693));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[18]$_DFFE_PN0P__644  (.H(net694));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[19]$_DFFE_PN0P__645  (.H(net695));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[1]$_DFFE_PN0P__646  (.H(net696));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[20]$_DFFE_PN0P__647  (.H(net697));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[21]$_DFFE_PN0P__648  (.H(net698));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[22]$_DFFE_PN0P__649  (.H(net699));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[23]$_DFFE_PN0P__650  (.H(net700));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[24]$_DFFE_PN0P__651  (.H(net701));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[25]$_DFFE_PN0P__652  (.H(net702));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[26]$_DFFE_PN0P__653  (.H(net703));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[27]$_DFFE_PN0P__654  (.H(net704));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[28]$_DFFE_PN0P__655  (.H(net705));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[29]$_DFFE_PN0P__656  (.H(net706));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[2]$_DFFE_PN0P__657  (.H(net707));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[30]$_DFFE_PN0P__658  (.H(net708));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[31]$_DFFE_PN0P__659  (.H(net709));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[3]$_DFFE_PN0P__660  (.H(net710));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[4]$_DFFE_PN0P__661  (.H(net711));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[5]$_DFFE_PN0P__662  (.H(net712));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[6]$_DFFE_PN0P__663  (.H(net713));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[7]$_DFFE_PN0P__664  (.H(net714));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[8]$_DFFE_PN0P__665  (.H(net715));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtval_csr.rdata_q[9]$_DFFE_PN0P__666  (.H(net716));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[10]$_DFFE_PN0P__667  (.H(net717));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[11]$_DFFE_PN0P__668  (.H(net718));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[12]$_DFFE_PN0P__669  (.H(net719));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[13]$_DFFE_PN0P__670  (.H(net720));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[14]$_DFFE_PN0P__671  (.H(net721));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[15]$_DFFE_PN0P__672  (.H(net722));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[16]$_DFFE_PN0P__673  (.H(net723));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[17]$_DFFE_PN0P__674  (.H(net724));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[18]$_DFFE_PN0P__675  (.H(net725));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[19]$_DFFE_PN0P__676  (.H(net726));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[20]$_DFFE_PN0P__677  (.H(net727));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[21]$_DFFE_PN0P__678  (.H(net728));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[22]$_DFFE_PN0P__679  (.H(net729));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[23]$_DFFE_PN0P__680  (.H(net730));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[24]$_DFFE_PN0P__681  (.H(net731));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[25]$_DFFE_PN0P__682  (.H(net732));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[26]$_DFFE_PN0P__683  (.H(net733));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[27]$_DFFE_PN0P__684  (.H(net734));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[28]$_DFFE_PN0P__685  (.H(net735));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[29]$_DFFE_PN0P__686  (.H(net736));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[30]$_DFFE_PN0P__687  (.H(net737));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[31]$_DFFE_PN0P__688  (.H(net738));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[8]$_DFFE_PN0P__689  (.H(net739));
 TIEHIx1_ASAP7_75t_R \cs_registers_i.u_mtvec_csr.rdata_q[9]$_DFFE_PN0P__690  (.H(net740));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P__691  (.H(net741));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P__692  (.H(net742));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P__693  (.H(net743));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P__694  (.H(net744));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P__695  (.H(net745));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P__696  (.H(net746));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1__697  (.H(net747));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0__698  (.H(net748));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0__699  (.H(net749));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0__700  (.H(net750));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0__701  (.H(net751));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0__702  (.H(net752));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P__703  (.H(net753));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P__704  (.H(net754));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P__705  (.H(net755));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P__706  (.H(net756));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P__707  (.H(net757));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P__708  (.H(net758));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P__709  (.H(net759));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P__710  (.H(net760));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P__711  (.H(net761));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P__712  (.H(net762));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P__713  (.H(net763));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P__714  (.H(net764));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P__715  (.H(net765));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P__716  (.H(net766));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P__717  (.H(net767));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P__718  (.H(net768));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P__719  (.H(net769));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P__720  (.H(net770));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P__721  (.H(net771));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P__722  (.H(net772));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P__723  (.H(net773));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P__724  (.H(net774));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P__725  (.H(net775));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P__726  (.H(net776));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P__727  (.H(net777));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P__728  (.H(net778));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P__729  (.H(net779));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P__730  (.H(net780));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P__731  (.H(net781));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P__732  (.H(net782));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P__733  (.H(net783));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P__734  (.H(net784));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P__735  (.H(net785));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P__736  (.H(net786));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P__737  (.H(net787));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P__738  (.H(net788));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P__739  (.H(net789));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P__740  (.H(net790));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P__741  (.H(net791));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P__742  (.H(net792));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P__743  (.H(net793));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P__744  (.H(net794));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P__745  (.H(net795));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P__746  (.H(net796));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P__747  (.H(net797));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P__748  (.H(net798));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P__749  (.H(net799));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P__750  (.H(net800));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P__751  (.H(net801));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P__752  (.H(net802));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P__753  (.H(net803));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P__754  (.H(net804));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P__755  (.H(net805));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P__756  (.H(net806));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P__757  (.H(net807));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P__758  (.H(net808));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P__759  (.H(net809));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P__760  (.H(net810));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P__761  (.H(net811));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P__762  (.H(net812));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P__763  (.H(net813));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P__764  (.H(net814));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P__765  (.H(net815));
 TIEHIx1_ASAP7_75t_R \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P__766  (.H(net816));
 TIEHIx1_ASAP7_75t_R \fetch_enable_q$_DFFE_PN0P__767  (.H(net817));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[0]$_DFFE_PN0P__768  (.H(net818));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[100]$_DFFE_PN0P__769  (.H(net819));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[101]$_DFFE_PN0P__770  (.H(net820));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[102]$_DFFE_PN0P__771  (.H(net821));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[103]$_DFFE_PN0P__772  (.H(net822));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[104]$_DFFE_PN0P__773  (.H(net823));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[105]$_DFFE_PN0P__774  (.H(net824));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[106]$_DFFE_PN0P__775  (.H(net825));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[107]$_DFFE_PN0P__776  (.H(net826));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[108]$_DFFE_PN0P__777  (.H(net827));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[109]$_DFFE_PN0P__778  (.H(net828));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[10]$_DFFE_PN0P__779  (.H(net829));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[110]$_DFFE_PN0P__780  (.H(net830));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[111]$_DFFE_PN0P__781  (.H(net831));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[112]$_DFFE_PN0P__782  (.H(net832));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[113]$_DFFE_PN0P__783  (.H(net833));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[114]$_DFFE_PN0P__784  (.H(net834));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[115]$_DFFE_PN0P__785  (.H(net835));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[116]$_DFFE_PN0P__786  (.H(net836));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[117]$_DFFE_PN0P__787  (.H(net837));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[118]$_DFFE_PN0P__788  (.H(net838));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[119]$_DFFE_PN0P__789  (.H(net839));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[11]$_DFFE_PN0P__790  (.H(net840));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[120]$_DFFE_PN0P__791  (.H(net841));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[121]$_DFFE_PN0P__792  (.H(net842));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[122]$_DFFE_PN0P__793  (.H(net843));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[123]$_DFFE_PN0P__794  (.H(net844));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[124]$_DFFE_PN0P__795  (.H(net845));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[125]$_DFFE_PN0P__796  (.H(net846));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[126]$_DFFE_PN0P__797  (.H(net847));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[127]$_DFFE_PN0P__798  (.H(net848));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[128]$_DFFE_PN0P__799  (.H(net849));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[129]$_DFFE_PN0P__800  (.H(net850));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[12]$_DFFE_PN0P__801  (.H(net851));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[130]$_DFFE_PN0P__802  (.H(net852));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[131]$_DFFE_PN0P__803  (.H(net853));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[132]$_DFFE_PN0P__804  (.H(net854));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[133]$_DFFE_PN0P__805  (.H(net855));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[134]$_DFFE_PN0P__806  (.H(net856));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[135]$_DFFE_PN0P__807  (.H(net857));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[136]$_DFFE_PN0P__808  (.H(net858));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[137]$_DFFE_PN0P__809  (.H(net859));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[138]$_DFFE_PN0P__810  (.H(net860));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[139]$_DFFE_PN0P__811  (.H(net861));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[13]$_DFFE_PN0P__812  (.H(net862));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[140]$_DFFE_PN0P__813  (.H(net863));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[141]$_DFFE_PN0P__814  (.H(net864));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[142]$_DFFE_PN0P__815  (.H(net865));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[143]$_DFFE_PN0P__816  (.H(net866));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[144]$_DFFE_PN0P__817  (.H(net867));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[145]$_DFFE_PN0P__818  (.H(net868));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[146]$_DFFE_PN0P__819  (.H(net869));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[147]$_DFFE_PN0P__820  (.H(net870));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[148]$_DFFE_PN0P__821  (.H(net871));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[149]$_DFFE_PN0P__822  (.H(net872));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[14]$_DFFE_PN0P__823  (.H(net873));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[150]$_DFFE_PN0P__824  (.H(net874));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[151]$_DFFE_PN0P__825  (.H(net875));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[152]$_DFFE_PN0P__826  (.H(net876));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[153]$_DFFE_PN0P__827  (.H(net877));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[154]$_DFFE_PN0P__828  (.H(net878));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[155]$_DFFE_PN0P__829  (.H(net879));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[156]$_DFFE_PN0P__830  (.H(net880));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[157]$_DFFE_PN0P__831  (.H(net881));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[158]$_DFFE_PN0P__832  (.H(net882));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[159]$_DFFE_PN0P__833  (.H(net883));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[15]$_DFFE_PN0P__834  (.H(net884));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[160]$_DFFE_PN0P__835  (.H(net885));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[161]$_DFFE_PN0P__836  (.H(net886));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[162]$_DFFE_PN0P__837  (.H(net887));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[163]$_DFFE_PN0P__838  (.H(net888));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[164]$_DFFE_PN0P__839  (.H(net889));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[165]$_DFFE_PN0P__840  (.H(net890));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[166]$_DFFE_PN0P__841  (.H(net891));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[167]$_DFFE_PN0P__842  (.H(net892));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[168]$_DFFE_PN0P__843  (.H(net893));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[169]$_DFFE_PN0P__844  (.H(net894));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[16]$_DFFE_PN0P__845  (.H(net895));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[170]$_DFFE_PN0P__846  (.H(net896));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[171]$_DFFE_PN0P__847  (.H(net897));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[172]$_DFFE_PN0P__848  (.H(net898));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[173]$_DFFE_PN0P__849  (.H(net899));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[174]$_DFFE_PN0P__850  (.H(net900));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[175]$_DFFE_PN0P__851  (.H(net901));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[176]$_DFFE_PN0P__852  (.H(net902));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[177]$_DFFE_PN0P__853  (.H(net903));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[178]$_DFFE_PN0P__854  (.H(net904));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[179]$_DFFE_PN0P__855  (.H(net905));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[17]$_DFFE_PN0P__856  (.H(net906));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[180]$_DFFE_PN0P__857  (.H(net907));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[181]$_DFFE_PN0P__858  (.H(net908));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[182]$_DFFE_PN0P__859  (.H(net909));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[183]$_DFFE_PN0P__860  (.H(net910));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[184]$_DFFE_PN0P__861  (.H(net911));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[185]$_DFFE_PN0P__862  (.H(net912));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[186]$_DFFE_PN0P__863  (.H(net913));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[187]$_DFFE_PN0P__864  (.H(net914));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[188]$_DFFE_PN0P__865  (.H(net915));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[189]$_DFFE_PN0P__866  (.H(net916));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[18]$_DFFE_PN0P__867  (.H(net917));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[190]$_DFFE_PN0P__868  (.H(net918));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[191]$_DFFE_PN0P__869  (.H(net919));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[192]$_DFFE_PN0P__870  (.H(net920));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[193]$_DFFE_PN0P__871  (.H(net921));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[194]$_DFFE_PN0P__872  (.H(net922));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[195]$_DFFE_PN0P__873  (.H(net923));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[196]$_DFFE_PN0P__874  (.H(net924));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[197]$_DFFE_PN0P__875  (.H(net925));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[198]$_DFFE_PN0P__876  (.H(net926));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[199]$_DFFE_PN0P__877  (.H(net927));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[19]$_DFFE_PN0P__878  (.H(net928));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[1]$_DFFE_PN0P__879  (.H(net929));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[200]$_DFFE_PN0P__880  (.H(net930));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[201]$_DFFE_PN0P__881  (.H(net931));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[202]$_DFFE_PN0P__882  (.H(net932));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[203]$_DFFE_PN0P__883  (.H(net933));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[204]$_DFFE_PN0P__884  (.H(net934));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[205]$_DFFE_PN0P__885  (.H(net935));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[206]$_DFFE_PN0P__886  (.H(net936));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[207]$_DFFE_PN0P__887  (.H(net937));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[208]$_DFFE_PN0P__888  (.H(net938));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[209]$_DFFE_PN0P__889  (.H(net939));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[20]$_DFFE_PN0P__890  (.H(net940));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[210]$_DFFE_PN0P__891  (.H(net941));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[211]$_DFFE_PN0P__892  (.H(net942));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[212]$_DFFE_PN0P__893  (.H(net943));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[213]$_DFFE_PN0P__894  (.H(net944));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[214]$_DFFE_PN0P__895  (.H(net945));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[215]$_DFFE_PN0P__896  (.H(net946));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[216]$_DFFE_PN0P__897  (.H(net947));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[217]$_DFFE_PN0P__898  (.H(net948));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[218]$_DFFE_PN0P__899  (.H(net949));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[219]$_DFFE_PN0P__900  (.H(net950));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[21]$_DFFE_PN0P__901  (.H(net951));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[220]$_DFFE_PN0P__902  (.H(net952));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[221]$_DFFE_PN0P__903  (.H(net953));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[222]$_DFFE_PN0P__904  (.H(net954));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[223]$_DFFE_PN0P__905  (.H(net955));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[224]$_DFFE_PN0P__906  (.H(net956));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[225]$_DFFE_PN0P__907  (.H(net957));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[226]$_DFFE_PN0P__908  (.H(net958));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[227]$_DFFE_PN0P__909  (.H(net959));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[228]$_DFFE_PN0P__910  (.H(net960));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[229]$_DFFE_PN0P__911  (.H(net961));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[22]$_DFFE_PN0P__912  (.H(net962));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[230]$_DFFE_PN0P__913  (.H(net963));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[231]$_DFFE_PN0P__914  (.H(net964));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[232]$_DFFE_PN0P__915  (.H(net965));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[233]$_DFFE_PN0P__916  (.H(net966));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[234]$_DFFE_PN0P__917  (.H(net967));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[235]$_DFFE_PN0P__918  (.H(net968));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[236]$_DFFE_PN0P__919  (.H(net969));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[237]$_DFFE_PN0P__920  (.H(net970));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[238]$_DFFE_PN0P__921  (.H(net971));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[239]$_DFFE_PN0P__922  (.H(net972));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[23]$_DFFE_PN0P__923  (.H(net973));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[240]$_DFFE_PN0P__924  (.H(net974));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[241]$_DFFE_PN0P__925  (.H(net975));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[242]$_DFFE_PN0P__926  (.H(net976));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[243]$_DFFE_PN0P__927  (.H(net977));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[244]$_DFFE_PN0P__928  (.H(net978));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[245]$_DFFE_PN0P__929  (.H(net979));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[246]$_DFFE_PN0P__930  (.H(net980));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[247]$_DFFE_PN0P__931  (.H(net981));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[248]$_DFFE_PN0P__932  (.H(net982));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[249]$_DFFE_PN0P__933  (.H(net983));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[24]$_DFFE_PN0P__934  (.H(net984));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[250]$_DFFE_PN0P__935  (.H(net985));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[251]$_DFFE_PN0P__936  (.H(net986));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[252]$_DFFE_PN0P__937  (.H(net987));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[253]$_DFFE_PN0P__938  (.H(net988));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[254]$_DFFE_PN0P__939  (.H(net989));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[255]$_DFFE_PN0P__940  (.H(net990));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[256]$_DFFE_PN0P__941  (.H(net991));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[257]$_DFFE_PN0P__942  (.H(net992));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[258]$_DFFE_PN0P__943  (.H(net993));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[259]$_DFFE_PN0P__944  (.H(net994));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[25]$_DFFE_PN0P__945  (.H(net995));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[260]$_DFFE_PN0P__946  (.H(net996));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[261]$_DFFE_PN0P__947  (.H(net997));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[262]$_DFFE_PN0P__948  (.H(net998));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[263]$_DFFE_PN0P__949  (.H(net999));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[264]$_DFFE_PN0P__950  (.H(net1000));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[265]$_DFFE_PN0P__951  (.H(net1001));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[266]$_DFFE_PN0P__952  (.H(net1002));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[267]$_DFFE_PN0P__953  (.H(net1003));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[268]$_DFFE_PN0P__954  (.H(net1004));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[269]$_DFFE_PN0P__955  (.H(net1005));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[26]$_DFFE_PN0P__956  (.H(net1006));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[270]$_DFFE_PN0P__957  (.H(net1007));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[271]$_DFFE_PN0P__958  (.H(net1008));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[272]$_DFFE_PN0P__959  (.H(net1009));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[273]$_DFFE_PN0P__960  (.H(net1010));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[274]$_DFFE_PN0P__961  (.H(net1011));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[275]$_DFFE_PN0P__962  (.H(net1012));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[276]$_DFFE_PN0P__963  (.H(net1013));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[277]$_DFFE_PN0P__964  (.H(net1014));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[278]$_DFFE_PN0P__965  (.H(net1015));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[279]$_DFFE_PN0P__966  (.H(net1016));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[27]$_DFFE_PN0P__967  (.H(net1017));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[280]$_DFFE_PN0P__968  (.H(net1018));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[281]$_DFFE_PN0P__969  (.H(net1019));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[282]$_DFFE_PN0P__970  (.H(net1020));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[283]$_DFFE_PN0P__971  (.H(net1021));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[284]$_DFFE_PN0P__972  (.H(net1022));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[285]$_DFFE_PN0P__973  (.H(net1023));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[286]$_DFFE_PN0P__974  (.H(net1024));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[287]$_DFFE_PN0P__975  (.H(net1025));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[288]$_DFFE_PN0P__976  (.H(net1026));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[289]$_DFFE_PN0P__977  (.H(net1027));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[28]$_DFFE_PN0P__978  (.H(net1028));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[290]$_DFFE_PN0P__979  (.H(net1029));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[291]$_DFFE_PN0P__980  (.H(net1030));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[292]$_DFFE_PN0P__981  (.H(net1031));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[293]$_DFFE_PN0P__982  (.H(net1032));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[294]$_DFFE_PN0P__983  (.H(net1033));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[295]$_DFFE_PN0P__984  (.H(net1034));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[296]$_DFFE_PN0P__985  (.H(net1035));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[297]$_DFFE_PN0P__986  (.H(net1036));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[298]$_DFFE_PN0P__987  (.H(net1037));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[299]$_DFFE_PN0P__988  (.H(net1038));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[29]$_DFFE_PN0P__989  (.H(net1039));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[2]$_DFFE_PN0P__990  (.H(net1040));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[300]$_DFFE_PN0P__991  (.H(net1041));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[301]$_DFFE_PN0P__992  (.H(net1042));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[302]$_DFFE_PN0P__993  (.H(net1043));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[303]$_DFFE_PN0P__994  (.H(net1044));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[304]$_DFFE_PN0P__995  (.H(net1045));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[305]$_DFFE_PN0P__996  (.H(net1046));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[306]$_DFFE_PN0P__997  (.H(net1047));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[307]$_DFFE_PN0P__998  (.H(net1048));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[308]$_DFFE_PN0P__999  (.H(net1049));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[309]$_DFFE_PN0P__1000  (.H(net1050));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[30]$_DFFE_PN0P__1001  (.H(net1051));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[310]$_DFFE_PN0P__1002  (.H(net1052));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[311]$_DFFE_PN0P__1003  (.H(net1053));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[312]$_DFFE_PN0P__1004  (.H(net1054));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[313]$_DFFE_PN0P__1005  (.H(net1055));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[314]$_DFFE_PN0P__1006  (.H(net1056));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[315]$_DFFE_PN0P__1007  (.H(net1057));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[316]$_DFFE_PN0P__1008  (.H(net1058));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[317]$_DFFE_PN0P__1009  (.H(net1059));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[318]$_DFFE_PN0P__1010  (.H(net1060));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[319]$_DFFE_PN0P__1011  (.H(net1061));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[31]$_DFFE_PN0P__1012  (.H(net1062));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[320]$_DFFE_PN0P__1013  (.H(net1063));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[321]$_DFFE_PN0P__1014  (.H(net1064));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[322]$_DFFE_PN0P__1015  (.H(net1065));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[323]$_DFFE_PN0P__1016  (.H(net1066));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[324]$_DFFE_PN0P__1017  (.H(net1067));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[325]$_DFFE_PN0P__1018  (.H(net1068));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[326]$_DFFE_PN0P__1019  (.H(net1069));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[327]$_DFFE_PN0P__1020  (.H(net1070));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[328]$_DFFE_PN0P__1021  (.H(net1071));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[329]$_DFFE_PN0P__1022  (.H(net1072));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[32]$_DFFE_PN0P__1023  (.H(net1073));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[330]$_DFFE_PN0P__1024  (.H(net1074));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[331]$_DFFE_PN0P__1025  (.H(net1075));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[332]$_DFFE_PN0P__1026  (.H(net1076));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[333]$_DFFE_PN0P__1027  (.H(net1077));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[334]$_DFFE_PN0P__1028  (.H(net1078));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[335]$_DFFE_PN0P__1029  (.H(net1079));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[336]$_DFFE_PN0P__1030  (.H(net1080));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[337]$_DFFE_PN0P__1031  (.H(net1081));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[338]$_DFFE_PN0P__1032  (.H(net1082));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[339]$_DFFE_PN0P__1033  (.H(net1083));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[33]$_DFFE_PN0P__1034  (.H(net1084));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[340]$_DFFE_PN0P__1035  (.H(net1085));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[341]$_DFFE_PN0P__1036  (.H(net1086));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[342]$_DFFE_PN0P__1037  (.H(net1087));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[343]$_DFFE_PN0P__1038  (.H(net1088));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[344]$_DFFE_PN0P__1039  (.H(net1089));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[345]$_DFFE_PN0P__1040  (.H(net1090));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[346]$_DFFE_PN0P__1041  (.H(net1091));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[347]$_DFFE_PN0P__1042  (.H(net1092));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[348]$_DFFE_PN0P__1043  (.H(net1093));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[349]$_DFFE_PN0P__1044  (.H(net1094));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[34]$_DFFE_PN0P__1045  (.H(net1095));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[350]$_DFFE_PN0P__1046  (.H(net1096));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[351]$_DFFE_PN0P__1047  (.H(net1097));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[352]$_DFFE_PN0P__1048  (.H(net1098));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[353]$_DFFE_PN0P__1049  (.H(net1099));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[354]$_DFFE_PN0P__1050  (.H(net1100));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[355]$_DFFE_PN0P__1051  (.H(net1101));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[356]$_DFFE_PN0P__1052  (.H(net1102));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[357]$_DFFE_PN0P__1053  (.H(net1103));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[358]$_DFFE_PN0P__1054  (.H(net1104));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[359]$_DFFE_PN0P__1055  (.H(net1105));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[35]$_DFFE_PN0P__1056  (.H(net1106));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[360]$_DFFE_PN0P__1057  (.H(net1107));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[361]$_DFFE_PN0P__1058  (.H(net1108));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[362]$_DFFE_PN0P__1059  (.H(net1109));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[363]$_DFFE_PN0P__1060  (.H(net1110));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[364]$_DFFE_PN0P__1061  (.H(net1111));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[365]$_DFFE_PN0P__1062  (.H(net1112));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[366]$_DFFE_PN0P__1063  (.H(net1113));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[367]$_DFFE_PN0P__1064  (.H(net1114));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[368]$_DFFE_PN0P__1065  (.H(net1115));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[369]$_DFFE_PN0P__1066  (.H(net1116));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[36]$_DFFE_PN0P__1067  (.H(net1117));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[370]$_DFFE_PN0P__1068  (.H(net1118));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[371]$_DFFE_PN0P__1069  (.H(net1119));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[372]$_DFFE_PN0P__1070  (.H(net1120));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[373]$_DFFE_PN0P__1071  (.H(net1121));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[374]$_DFFE_PN0P__1072  (.H(net1122));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[375]$_DFFE_PN0P__1073  (.H(net1123));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[376]$_DFFE_PN0P__1074  (.H(net1124));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[377]$_DFFE_PN0P__1075  (.H(net1125));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[378]$_DFFE_PN0P__1076  (.H(net1126));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[379]$_DFFE_PN0P__1077  (.H(net1127));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[37]$_DFFE_PN0P__1078  (.H(net1128));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[380]$_DFFE_PN0P__1079  (.H(net1129));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[381]$_DFFE_PN0P__1080  (.H(net1130));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[382]$_DFFE_PN0P__1081  (.H(net1131));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[383]$_DFFE_PN0P__1082  (.H(net1132));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[384]$_DFFE_PN0P__1083  (.H(net1133));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[385]$_DFFE_PN0P__1084  (.H(net1134));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[386]$_DFFE_PN0P__1085  (.H(net1135));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[387]$_DFFE_PN0P__1086  (.H(net1136));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[388]$_DFFE_PN0P__1087  (.H(net1137));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[389]$_DFFE_PN0P__1088  (.H(net1138));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[38]$_DFFE_PN0P__1089  (.H(net1139));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[390]$_DFFE_PN0P__1090  (.H(net1140));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[391]$_DFFE_PN0P__1091  (.H(net1141));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[392]$_DFFE_PN0P__1092  (.H(net1142));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[393]$_DFFE_PN0P__1093  (.H(net1143));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[394]$_DFFE_PN0P__1094  (.H(net1144));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[395]$_DFFE_PN0P__1095  (.H(net1145));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[396]$_DFFE_PN0P__1096  (.H(net1146));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[397]$_DFFE_PN0P__1097  (.H(net1147));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[398]$_DFFE_PN0P__1098  (.H(net1148));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[399]$_DFFE_PN0P__1099  (.H(net1149));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[39]$_DFFE_PN0P__1100  (.H(net1150));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[3]$_DFFE_PN0P__1101  (.H(net1151));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[400]$_DFFE_PN0P__1102  (.H(net1152));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[401]$_DFFE_PN0P__1103  (.H(net1153));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[402]$_DFFE_PN0P__1104  (.H(net1154));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[403]$_DFFE_PN0P__1105  (.H(net1155));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[404]$_DFFE_PN0P__1106  (.H(net1156));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[405]$_DFFE_PN0P__1107  (.H(net1157));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[406]$_DFFE_PN0P__1108  (.H(net1158));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[407]$_DFFE_PN0P__1109  (.H(net1159));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[408]$_DFFE_PN0P__1110  (.H(net1160));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[409]$_DFFE_PN0P__1111  (.H(net1161));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[40]$_DFFE_PN0P__1112  (.H(net1162));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[410]$_DFFE_PN0P__1113  (.H(net1163));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[411]$_DFFE_PN0P__1114  (.H(net1164));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[412]$_DFFE_PN0P__1115  (.H(net1165));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[413]$_DFFE_PN0P__1116  (.H(net1166));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[414]$_DFFE_PN0P__1117  (.H(net1167));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[415]$_DFFE_PN0P__1118  (.H(net1168));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[416]$_DFFE_PN0P__1119  (.H(net1169));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[417]$_DFFE_PN0P__1120  (.H(net1170));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[418]$_DFFE_PN0P__1121  (.H(net1171));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[419]$_DFFE_PN0P__1122  (.H(net1172));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[41]$_DFFE_PN0P__1123  (.H(net1173));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[420]$_DFFE_PN0P__1124  (.H(net1174));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[421]$_DFFE_PN0P__1125  (.H(net1175));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[422]$_DFFE_PN0P__1126  (.H(net1176));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[423]$_DFFE_PN0P__1127  (.H(net1177));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[424]$_DFFE_PN0P__1128  (.H(net1178));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[425]$_DFFE_PN0P__1129  (.H(net1179));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[426]$_DFFE_PN0P__1130  (.H(net1180));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[427]$_DFFE_PN0P__1131  (.H(net1181));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[428]$_DFFE_PN0P__1132  (.H(net1182));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[429]$_DFFE_PN0P__1133  (.H(net1183));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[42]$_DFFE_PN0P__1134  (.H(net1184));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[430]$_DFFE_PN0P__1135  (.H(net1185));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[431]$_DFFE_PN0P__1136  (.H(net1186));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[432]$_DFFE_PN0P__1137  (.H(net1187));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[433]$_DFFE_PN0P__1138  (.H(net1188));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[434]$_DFFE_PN0P__1139  (.H(net1189));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[435]$_DFFE_PN0P__1140  (.H(net1190));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[436]$_DFFE_PN0P__1141  (.H(net1191));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[437]$_DFFE_PN0P__1142  (.H(net1192));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[438]$_DFFE_PN0P__1143  (.H(net1193));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[439]$_DFFE_PN0P__1144  (.H(net1194));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[43]$_DFFE_PN0P__1145  (.H(net1195));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[440]$_DFFE_PN0P__1146  (.H(net1196));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[441]$_DFFE_PN0P__1147  (.H(net1197));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[442]$_DFFE_PN0P__1148  (.H(net1198));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[443]$_DFFE_PN0P__1149  (.H(net1199));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[444]$_DFFE_PN0P__1150  (.H(net1200));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[445]$_DFFE_PN0P__1151  (.H(net1201));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[446]$_DFFE_PN0P__1152  (.H(net1202));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[447]$_DFFE_PN0P__1153  (.H(net1203));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[448]$_DFFE_PN0P__1154  (.H(net1204));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[449]$_DFFE_PN0P__1155  (.H(net1205));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[44]$_DFFE_PN0P__1156  (.H(net1206));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[450]$_DFFE_PN0P__1157  (.H(net1207));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[451]$_DFFE_PN0P__1158  (.H(net1208));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[452]$_DFFE_PN0P__1159  (.H(net1209));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[453]$_DFFE_PN0P__1160  (.H(net1210));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[454]$_DFFE_PN0P__1161  (.H(net1211));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[455]$_DFFE_PN0P__1162  (.H(net1212));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[456]$_DFFE_PN0P__1163  (.H(net1213));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[457]$_DFFE_PN0P__1164  (.H(net1214));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[458]$_DFFE_PN0P__1165  (.H(net1215));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[459]$_DFFE_PN0P__1166  (.H(net1216));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[45]$_DFFE_PN0P__1167  (.H(net1217));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[460]$_DFFE_PN0P__1168  (.H(net1218));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[461]$_DFFE_PN0P__1169  (.H(net1219));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[462]$_DFFE_PN0P__1170  (.H(net1220));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[463]$_DFFE_PN0P__1171  (.H(net1221));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[464]$_DFFE_PN0P__1172  (.H(net1222));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[465]$_DFFE_PN0P__1173  (.H(net1223));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[466]$_DFFE_PN0P__1174  (.H(net1224));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[467]$_DFFE_PN0P__1175  (.H(net1225));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[468]$_DFFE_PN0P__1176  (.H(net1226));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[469]$_DFFE_PN0P__1177  (.H(net1227));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[46]$_DFFE_PN0P__1178  (.H(net1228));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[470]$_DFFE_PN0P__1179  (.H(net1229));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[471]$_DFFE_PN0P__1180  (.H(net1230));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[472]$_DFFE_PN0P__1181  (.H(net1231));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[473]$_DFFE_PN0P__1182  (.H(net1232));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[474]$_DFFE_PN0P__1183  (.H(net1233));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[475]$_DFFE_PN0P__1184  (.H(net1234));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[476]$_DFFE_PN0P__1185  (.H(net1235));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[477]$_DFFE_PN0P__1186  (.H(net1236));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[478]$_DFFE_PN0P__1187  (.H(net1237));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[479]$_DFFE_PN0P__1188  (.H(net1238));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[47]$_DFFE_PN0P__1189  (.H(net1239));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[480]$_DFFE_PN0P__1190  (.H(net1240));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[481]$_DFFE_PN0P__1191  (.H(net1241));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[482]$_DFFE_PN0P__1192  (.H(net1242));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[483]$_DFFE_PN0P__1193  (.H(net1243));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[484]$_DFFE_PN0P__1194  (.H(net1244));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[485]$_DFFE_PN0P__1195  (.H(net1245));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[486]$_DFFE_PN0P__1196  (.H(net1246));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[487]$_DFFE_PN0P__1197  (.H(net1247));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[488]$_DFFE_PN0P__1198  (.H(net1248));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[489]$_DFFE_PN0P__1199  (.H(net1249));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[48]$_DFFE_PN0P__1200  (.H(net1250));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[490]$_DFFE_PN0P__1201  (.H(net1251));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[491]$_DFFE_PN0P__1202  (.H(net1252));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[492]$_DFFE_PN0P__1203  (.H(net1253));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[493]$_DFFE_PN0P__1204  (.H(net1254));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[494]$_DFFE_PN0P__1205  (.H(net1255));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[495]$_DFFE_PN0P__1206  (.H(net1256));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[496]$_DFFE_PN0P__1207  (.H(net1257));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[497]$_DFFE_PN0P__1208  (.H(net1258));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[498]$_DFFE_PN0P__1209  (.H(net1259));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[499]$_DFFE_PN0P__1210  (.H(net1260));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[49]$_DFFE_PN0P__1211  (.H(net1261));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[4]$_DFFE_PN0P__1212  (.H(net1262));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[500]$_DFFE_PN0P__1213  (.H(net1263));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[501]$_DFFE_PN0P__1214  (.H(net1264));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[502]$_DFFE_PN0P__1215  (.H(net1265));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[503]$_DFFE_PN0P__1216  (.H(net1266));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[504]$_DFFE_PN0P__1217  (.H(net1267));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[505]$_DFFE_PN0P__1218  (.H(net1268));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[506]$_DFFE_PN0P__1219  (.H(net1269));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[507]$_DFFE_PN0P__1220  (.H(net1270));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[508]$_DFFE_PN0P__1221  (.H(net1271));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[509]$_DFFE_PN0P__1222  (.H(net1272));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[50]$_DFFE_PN0P__1223  (.H(net1273));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[510]$_DFFE_PN0P__1224  (.H(net1274));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[511]$_DFFE_PN0P__1225  (.H(net1275));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[512]$_DFFE_PN0P__1226  (.H(net1276));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[513]$_DFFE_PN0P__1227  (.H(net1277));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[514]$_DFFE_PN0P__1228  (.H(net1278));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[515]$_DFFE_PN0P__1229  (.H(net1279));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[516]$_DFFE_PN0P__1230  (.H(net1280));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[517]$_DFFE_PN0P__1231  (.H(net1281));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[518]$_DFFE_PN0P__1232  (.H(net1282));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[519]$_DFFE_PN0P__1233  (.H(net1283));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[51]$_DFFE_PN0P__1234  (.H(net1284));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[520]$_DFFE_PN0P__1235  (.H(net1285));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[521]$_DFFE_PN0P__1236  (.H(net1286));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[522]$_DFFE_PN0P__1237  (.H(net1287));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[523]$_DFFE_PN0P__1238  (.H(net1288));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[524]$_DFFE_PN0P__1239  (.H(net1289));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[525]$_DFFE_PN0P__1240  (.H(net1290));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[526]$_DFFE_PN0P__1241  (.H(net1291));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[527]$_DFFE_PN0P__1242  (.H(net1292));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[528]$_DFFE_PN0P__1243  (.H(net1293));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[529]$_DFFE_PN0P__1244  (.H(net1294));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[52]$_DFFE_PN0P__1245  (.H(net1295));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[530]$_DFFE_PN0P__1246  (.H(net1296));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[531]$_DFFE_PN0P__1247  (.H(net1297));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[532]$_DFFE_PN0P__1248  (.H(net1298));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[533]$_DFFE_PN0P__1249  (.H(net1299));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[534]$_DFFE_PN0P__1250  (.H(net1300));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[535]$_DFFE_PN0P__1251  (.H(net1301));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[536]$_DFFE_PN0P__1252  (.H(net1302));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[537]$_DFFE_PN0P__1253  (.H(net1303));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[538]$_DFFE_PN0P__1254  (.H(net1304));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[539]$_DFFE_PN0P__1255  (.H(net1305));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[53]$_DFFE_PN0P__1256  (.H(net1306));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[540]$_DFFE_PN0P__1257  (.H(net1307));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[541]$_DFFE_PN0P__1258  (.H(net1308));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[542]$_DFFE_PN0P__1259  (.H(net1309));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[543]$_DFFE_PN0P__1260  (.H(net1310));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[544]$_DFFE_PN0P__1261  (.H(net1311));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[545]$_DFFE_PN0P__1262  (.H(net1312));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[546]$_DFFE_PN0P__1263  (.H(net1313));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[547]$_DFFE_PN0P__1264  (.H(net1314));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[548]$_DFFE_PN0P__1265  (.H(net1315));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[549]$_DFFE_PN0P__1266  (.H(net1316));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[54]$_DFFE_PN0P__1267  (.H(net1317));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[550]$_DFFE_PN0P__1268  (.H(net1318));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[551]$_DFFE_PN0P__1269  (.H(net1319));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[552]$_DFFE_PN0P__1270  (.H(net1320));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[553]$_DFFE_PN0P__1271  (.H(net1321));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[554]$_DFFE_PN0P__1272  (.H(net1322));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[555]$_DFFE_PN0P__1273  (.H(net1323));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[556]$_DFFE_PN0P__1274  (.H(net1324));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[557]$_DFFE_PN0P__1275  (.H(net1325));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[558]$_DFFE_PN0P__1276  (.H(net1326));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[559]$_DFFE_PN0P__1277  (.H(net1327));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[55]$_DFFE_PN0P__1278  (.H(net1328));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[560]$_DFFE_PN0P__1279  (.H(net1329));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[561]$_DFFE_PN0P__1280  (.H(net1330));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[562]$_DFFE_PN0P__1281  (.H(net1331));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[563]$_DFFE_PN0P__1282  (.H(net1332));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[564]$_DFFE_PN0P__1283  (.H(net1333));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[565]$_DFFE_PN0P__1284  (.H(net1334));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[566]$_DFFE_PN0P__1285  (.H(net1335));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[567]$_DFFE_PN0P__1286  (.H(net1336));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[568]$_DFFE_PN0P__1287  (.H(net1337));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[569]$_DFFE_PN0P__1288  (.H(net1338));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[56]$_DFFE_PN0P__1289  (.H(net1339));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[570]$_DFFE_PN0P__1290  (.H(net1340));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[571]$_DFFE_PN0P__1291  (.H(net1341));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[572]$_DFFE_PN0P__1292  (.H(net1342));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[573]$_DFFE_PN0P__1293  (.H(net1343));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[574]$_DFFE_PN0P__1294  (.H(net1344));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[575]$_DFFE_PN0P__1295  (.H(net1345));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[576]$_DFFE_PN0P__1296  (.H(net1346));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[577]$_DFFE_PN0P__1297  (.H(net1347));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[578]$_DFFE_PN0P__1298  (.H(net1348));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[579]$_DFFE_PN0P__1299  (.H(net1349));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[57]$_DFFE_PN0P__1300  (.H(net1350));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[580]$_DFFE_PN0P__1301  (.H(net1351));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[581]$_DFFE_PN0P__1302  (.H(net1352));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[582]$_DFFE_PN0P__1303  (.H(net1353));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[583]$_DFFE_PN0P__1304  (.H(net1354));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[584]$_DFFE_PN0P__1305  (.H(net1355));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[585]$_DFFE_PN0P__1306  (.H(net1356));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[586]$_DFFE_PN0P__1307  (.H(net1357));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[587]$_DFFE_PN0P__1308  (.H(net1358));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[588]$_DFFE_PN0P__1309  (.H(net1359));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[589]$_DFFE_PN0P__1310  (.H(net1360));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[58]$_DFFE_PN0P__1311  (.H(net1361));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[590]$_DFFE_PN0P__1312  (.H(net1362));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[591]$_DFFE_PN0P__1313  (.H(net1363));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[592]$_DFFE_PN0P__1314  (.H(net1364));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[593]$_DFFE_PN0P__1315  (.H(net1365));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[594]$_DFFE_PN0P__1316  (.H(net1366));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[595]$_DFFE_PN0P__1317  (.H(net1367));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[596]$_DFFE_PN0P__1318  (.H(net1368));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[597]$_DFFE_PN0P__1319  (.H(net1369));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[598]$_DFFE_PN0P__1320  (.H(net1370));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[599]$_DFFE_PN0P__1321  (.H(net1371));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[59]$_DFFE_PN0P__1322  (.H(net1372));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[5]$_DFFE_PN0P__1323  (.H(net1373));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[600]$_DFFE_PN0P__1324  (.H(net1374));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[601]$_DFFE_PN0P__1325  (.H(net1375));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[602]$_DFFE_PN0P__1326  (.H(net1376));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[603]$_DFFE_PN0P__1327  (.H(net1377));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[604]$_DFFE_PN0P__1328  (.H(net1378));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[605]$_DFFE_PN0P__1329  (.H(net1379));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[606]$_DFFE_PN0P__1330  (.H(net1380));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[607]$_DFFE_PN0P__1331  (.H(net1381));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[608]$_DFFE_PN0P__1332  (.H(net1382));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[609]$_DFFE_PN0P__1333  (.H(net1383));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[60]$_DFFE_PN0P__1334  (.H(net1384));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[610]$_DFFE_PN0P__1335  (.H(net1385));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[611]$_DFFE_PN0P__1336  (.H(net1386));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[612]$_DFFE_PN0P__1337  (.H(net1387));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[613]$_DFFE_PN0P__1338  (.H(net1388));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[614]$_DFFE_PN0P__1339  (.H(net1389));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[615]$_DFFE_PN0P__1340  (.H(net1390));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[616]$_DFFE_PN0P__1341  (.H(net1391));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[617]$_DFFE_PN0P__1342  (.H(net1392));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[618]$_DFFE_PN0P__1343  (.H(net1393));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[619]$_DFFE_PN0P__1344  (.H(net1394));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[61]$_DFFE_PN0P__1345  (.H(net1395));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[620]$_DFFE_PN0P__1346  (.H(net1396));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[621]$_DFFE_PN0P__1347  (.H(net1397));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[622]$_DFFE_PN0P__1348  (.H(net1398));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[623]$_DFFE_PN0P__1349  (.H(net1399));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[624]$_DFFE_PN0P__1350  (.H(net1400));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[625]$_DFFE_PN0P__1351  (.H(net1401));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[626]$_DFFE_PN0P__1352  (.H(net1402));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[627]$_DFFE_PN0P__1353  (.H(net1403));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[628]$_DFFE_PN0P__1354  (.H(net1404));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[629]$_DFFE_PN0P__1355  (.H(net1405));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[62]$_DFFE_PN0P__1356  (.H(net1406));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[630]$_DFFE_PN0P__1357  (.H(net1407));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[631]$_DFFE_PN0P__1358  (.H(net1408));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[632]$_DFFE_PN0P__1359  (.H(net1409));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[633]$_DFFE_PN0P__1360  (.H(net1410));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[634]$_DFFE_PN0P__1361  (.H(net1411));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[635]$_DFFE_PN0P__1362  (.H(net1412));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[636]$_DFFE_PN0P__1363  (.H(net1413));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[637]$_DFFE_PN0P__1364  (.H(net1414));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[638]$_DFFE_PN0P__1365  (.H(net1415));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[639]$_DFFE_PN0P__1366  (.H(net1416));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[63]$_DFFE_PN0P__1367  (.H(net1417));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[640]$_DFFE_PN0P__1368  (.H(net1418));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[641]$_DFFE_PN0P__1369  (.H(net1419));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[642]$_DFFE_PN0P__1370  (.H(net1420));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[643]$_DFFE_PN0P__1371  (.H(net1421));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[644]$_DFFE_PN0P__1372  (.H(net1422));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[645]$_DFFE_PN0P__1373  (.H(net1423));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[646]$_DFFE_PN0P__1374  (.H(net1424));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[647]$_DFFE_PN0P__1375  (.H(net1425));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[648]$_DFFE_PN0P__1376  (.H(net1426));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[649]$_DFFE_PN0P__1377  (.H(net1427));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[64]$_DFFE_PN0P__1378  (.H(net1428));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[650]$_DFFE_PN0P__1379  (.H(net1429));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[651]$_DFFE_PN0P__1380  (.H(net1430));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[652]$_DFFE_PN0P__1381  (.H(net1431));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[653]$_DFFE_PN0P__1382  (.H(net1432));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[654]$_DFFE_PN0P__1383  (.H(net1433));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[655]$_DFFE_PN0P__1384  (.H(net1434));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[656]$_DFFE_PN0P__1385  (.H(net1435));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[657]$_DFFE_PN0P__1386  (.H(net1436));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[658]$_DFFE_PN0P__1387  (.H(net1437));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[659]$_DFFE_PN0P__1388  (.H(net1438));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[65]$_DFFE_PN0P__1389  (.H(net1439));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[660]$_DFFE_PN0P__1390  (.H(net1440));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[661]$_DFFE_PN0P__1391  (.H(net1441));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[662]$_DFFE_PN0P__1392  (.H(net1442));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[663]$_DFFE_PN0P__1393  (.H(net1443));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[664]$_DFFE_PN0P__1394  (.H(net1444));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[665]$_DFFE_PN0P__1395  (.H(net1445));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[666]$_DFFE_PN0P__1396  (.H(net1446));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[667]$_DFFE_PN0P__1397  (.H(net1447));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[668]$_DFFE_PN0P__1398  (.H(net1448));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[669]$_DFFE_PN0P__1399  (.H(net1449));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[66]$_DFFE_PN0P__1400  (.H(net1450));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[670]$_DFFE_PN0P__1401  (.H(net1451));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[671]$_DFFE_PN0P__1402  (.H(net1452));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[672]$_DFFE_PN0P__1403  (.H(net1453));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[673]$_DFFE_PN0P__1404  (.H(net1454));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[674]$_DFFE_PN0P__1405  (.H(net1455));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[675]$_DFFE_PN0P__1406  (.H(net1456));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[676]$_DFFE_PN0P__1407  (.H(net1457));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[677]$_DFFE_PN0P__1408  (.H(net1458));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[678]$_DFFE_PN0P__1409  (.H(net1459));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[679]$_DFFE_PN0P__1410  (.H(net1460));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[67]$_DFFE_PN0P__1411  (.H(net1461));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[680]$_DFFE_PN0P__1412  (.H(net1462));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[681]$_DFFE_PN0P__1413  (.H(net1463));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[682]$_DFFE_PN0P__1414  (.H(net1464));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[683]$_DFFE_PN0P__1415  (.H(net1465));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[684]$_DFFE_PN0P__1416  (.H(net1466));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[685]$_DFFE_PN0P__1417  (.H(net1467));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[686]$_DFFE_PN0P__1418  (.H(net1468));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[687]$_DFFE_PN0P__1419  (.H(net1469));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[688]$_DFFE_PN0P__1420  (.H(net1470));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[689]$_DFFE_PN0P__1421  (.H(net1471));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[68]$_DFFE_PN0P__1422  (.H(net1472));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[690]$_DFFE_PN0P__1423  (.H(net1473));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[691]$_DFFE_PN0P__1424  (.H(net1474));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[692]$_DFFE_PN0P__1425  (.H(net1475));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[693]$_DFFE_PN0P__1426  (.H(net1476));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[694]$_DFFE_PN0P__1427  (.H(net1477));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[695]$_DFFE_PN0P__1428  (.H(net1478));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[696]$_DFFE_PN0P__1429  (.H(net1479));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[697]$_DFFE_PN0P__1430  (.H(net1480));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[698]$_DFFE_PN0P__1431  (.H(net1481));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[699]$_DFFE_PN0P__1432  (.H(net1482));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[69]$_DFFE_PN0P__1433  (.H(net1483));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[6]$_DFFE_PN0P__1434  (.H(net1484));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[700]$_DFFE_PN0P__1435  (.H(net1485));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[701]$_DFFE_PN0P__1436  (.H(net1486));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[702]$_DFFE_PN0P__1437  (.H(net1487));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[703]$_DFFE_PN0P__1438  (.H(net1488));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[704]$_DFFE_PN0P__1439  (.H(net1489));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[705]$_DFFE_PN0P__1440  (.H(net1490));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[706]$_DFFE_PN0P__1441  (.H(net1491));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[707]$_DFFE_PN0P__1442  (.H(net1492));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[708]$_DFFE_PN0P__1443  (.H(net1493));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[709]$_DFFE_PN0P__1444  (.H(net1494));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[70]$_DFFE_PN0P__1445  (.H(net1495));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[710]$_DFFE_PN0P__1446  (.H(net1496));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[711]$_DFFE_PN0P__1447  (.H(net1497));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[712]$_DFFE_PN0P__1448  (.H(net1498));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[713]$_DFFE_PN0P__1449  (.H(net1499));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[714]$_DFFE_PN0P__1450  (.H(net1500));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[715]$_DFFE_PN0P__1451  (.H(net1501));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[716]$_DFFE_PN0P__1452  (.H(net1502));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[717]$_DFFE_PN0P__1453  (.H(net1503));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[718]$_DFFE_PN0P__1454  (.H(net1504));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[719]$_DFFE_PN0P__1455  (.H(net1505));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[71]$_DFFE_PN0P__1456  (.H(net1506));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[720]$_DFFE_PN0P__1457  (.H(net1507));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[721]$_DFFE_PN0P__1458  (.H(net1508));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[722]$_DFFE_PN0P__1459  (.H(net1509));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[723]$_DFFE_PN0P__1460  (.H(net1510));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[724]$_DFFE_PN0P__1461  (.H(net1511));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[725]$_DFFE_PN0P__1462  (.H(net1512));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[726]$_DFFE_PN0P__1463  (.H(net1513));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[727]$_DFFE_PN0P__1464  (.H(net1514));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[728]$_DFFE_PN0P__1465  (.H(net1515));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[729]$_DFFE_PN0P__1466  (.H(net1516));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[72]$_DFFE_PN0P__1467  (.H(net1517));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[730]$_DFFE_PN0P__1468  (.H(net1518));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[731]$_DFFE_PN0P__1469  (.H(net1519));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[732]$_DFFE_PN0P__1470  (.H(net1520));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[733]$_DFFE_PN0P__1471  (.H(net1521));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[734]$_DFFE_PN0P__1472  (.H(net1522));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[735]$_DFFE_PN0P__1473  (.H(net1523));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[736]$_DFFE_PN0P__1474  (.H(net1524));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[737]$_DFFE_PN0P__1475  (.H(net1525));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[738]$_DFFE_PN0P__1476  (.H(net1526));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[739]$_DFFE_PN0P__1477  (.H(net1527));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[73]$_DFFE_PN0P__1478  (.H(net1528));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[740]$_DFFE_PN0P__1479  (.H(net1529));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[741]$_DFFE_PN0P__1480  (.H(net1530));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[742]$_DFFE_PN0P__1481  (.H(net1531));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[743]$_DFFE_PN0P__1482  (.H(net1532));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[744]$_DFFE_PN0P__1483  (.H(net1533));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[745]$_DFFE_PN0P__1484  (.H(net1534));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[746]$_DFFE_PN0P__1485  (.H(net1535));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[747]$_DFFE_PN0P__1486  (.H(net1536));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[748]$_DFFE_PN0P__1487  (.H(net1537));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[749]$_DFFE_PN0P__1488  (.H(net1538));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[74]$_DFFE_PN0P__1489  (.H(net1539));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[750]$_DFFE_PN0P__1490  (.H(net1540));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[751]$_DFFE_PN0P__1491  (.H(net1541));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[752]$_DFFE_PN0P__1492  (.H(net1542));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[753]$_DFFE_PN0P__1493  (.H(net1543));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[754]$_DFFE_PN0P__1494  (.H(net1544));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[755]$_DFFE_PN0P__1495  (.H(net1545));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[756]$_DFFE_PN0P__1496  (.H(net1546));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[757]$_DFFE_PN0P__1497  (.H(net1547));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[758]$_DFFE_PN0P__1498  (.H(net1548));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[759]$_DFFE_PN0P__1499  (.H(net1549));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[75]$_DFFE_PN0P__1500  (.H(net1550));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[760]$_DFFE_PN0P__1501  (.H(net1551));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[761]$_DFFE_PN0P__1502  (.H(net1552));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[762]$_DFFE_PN0P__1503  (.H(net1553));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[763]$_DFFE_PN0P__1504  (.H(net1554));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[764]$_DFFE_PN0P__1505  (.H(net1555));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[765]$_DFFE_PN0P__1506  (.H(net1556));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[766]$_DFFE_PN0P__1507  (.H(net1557));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[767]$_DFFE_PN0P__1508  (.H(net1558));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[768]$_DFFE_PN0P__1509  (.H(net1559));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[769]$_DFFE_PN0P__1510  (.H(net1560));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[76]$_DFFE_PN0P__1511  (.H(net1561));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[770]$_DFFE_PN0P__1512  (.H(net1562));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[771]$_DFFE_PN0P__1513  (.H(net1563));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[772]$_DFFE_PN0P__1514  (.H(net1564));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[773]$_DFFE_PN0P__1515  (.H(net1565));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[774]$_DFFE_PN0P__1516  (.H(net1566));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[775]$_DFFE_PN0P__1517  (.H(net1567));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[776]$_DFFE_PN0P__1518  (.H(net1568));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[777]$_DFFE_PN0P__1519  (.H(net1569));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[778]$_DFFE_PN0P__1520  (.H(net1570));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[779]$_DFFE_PN0P__1521  (.H(net1571));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[77]$_DFFE_PN0P__1522  (.H(net1572));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[780]$_DFFE_PN0P__1523  (.H(net1573));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[781]$_DFFE_PN0P__1524  (.H(net1574));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[782]$_DFFE_PN0P__1525  (.H(net1575));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[783]$_DFFE_PN0P__1526  (.H(net1576));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[784]$_DFFE_PN0P__1527  (.H(net1577));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[785]$_DFFE_PN0P__1528  (.H(net1578));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[786]$_DFFE_PN0P__1529  (.H(net1579));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[787]$_DFFE_PN0P__1530  (.H(net1580));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[788]$_DFFE_PN0P__1531  (.H(net1581));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[789]$_DFFE_PN0P__1532  (.H(net1582));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[78]$_DFFE_PN0P__1533  (.H(net1583));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[790]$_DFFE_PN0P__1534  (.H(net1584));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[791]$_DFFE_PN0P__1535  (.H(net1585));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[792]$_DFFE_PN0P__1536  (.H(net1586));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[793]$_DFFE_PN0P__1537  (.H(net1587));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[794]$_DFFE_PN0P__1538  (.H(net1588));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[795]$_DFFE_PN0P__1539  (.H(net1589));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[796]$_DFFE_PN0P__1540  (.H(net1590));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[797]$_DFFE_PN0P__1541  (.H(net1591));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[798]$_DFFE_PN0P__1542  (.H(net1592));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[799]$_DFFE_PN0P__1543  (.H(net1593));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[79]$_DFFE_PN0P__1544  (.H(net1594));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[7]$_DFFE_PN0P__1545  (.H(net1595));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[800]$_DFFE_PN0P__1546  (.H(net1596));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[801]$_DFFE_PN0P__1547  (.H(net1597));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[802]$_DFFE_PN0P__1548  (.H(net1598));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[803]$_DFFE_PN0P__1549  (.H(net1599));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[804]$_DFFE_PN0P__1550  (.H(net1600));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[805]$_DFFE_PN0P__1551  (.H(net1601));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[806]$_DFFE_PN0P__1552  (.H(net1602));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[807]$_DFFE_PN0P__1553  (.H(net1603));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[808]$_DFFE_PN0P__1554  (.H(net1604));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[809]$_DFFE_PN0P__1555  (.H(net1605));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[80]$_DFFE_PN0P__1556  (.H(net1606));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[810]$_DFFE_PN0P__1557  (.H(net1607));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[811]$_DFFE_PN0P__1558  (.H(net1608));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[812]$_DFFE_PN0P__1559  (.H(net1609));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[813]$_DFFE_PN0P__1560  (.H(net1610));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[814]$_DFFE_PN0P__1561  (.H(net1611));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[815]$_DFFE_PN0P__1562  (.H(net1612));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[816]$_DFFE_PN0P__1563  (.H(net1613));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[817]$_DFFE_PN0P__1564  (.H(net1614));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[818]$_DFFE_PN0P__1565  (.H(net1615));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[819]$_DFFE_PN0P__1566  (.H(net1616));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[81]$_DFFE_PN0P__1567  (.H(net1617));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[820]$_DFFE_PN0P__1568  (.H(net1618));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[821]$_DFFE_PN0P__1569  (.H(net1619));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[822]$_DFFE_PN0P__1570  (.H(net1620));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[823]$_DFFE_PN0P__1571  (.H(net1621));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[824]$_DFFE_PN0P__1572  (.H(net1622));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[825]$_DFFE_PN0P__1573  (.H(net1623));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[826]$_DFFE_PN0P__1574  (.H(net1624));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[827]$_DFFE_PN0P__1575  (.H(net1625));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[828]$_DFFE_PN0P__1576  (.H(net1626));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[829]$_DFFE_PN0P__1577  (.H(net1627));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[82]$_DFFE_PN0P__1578  (.H(net1628));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[830]$_DFFE_PN0P__1579  (.H(net1629));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[831]$_DFFE_PN0P__1580  (.H(net1630));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[832]$_DFFE_PN0P__1581  (.H(net1631));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[833]$_DFFE_PN0P__1582  (.H(net1632));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[834]$_DFFE_PN0P__1583  (.H(net1633));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[835]$_DFFE_PN0P__1584  (.H(net1634));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[836]$_DFFE_PN0P__1585  (.H(net1635));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[837]$_DFFE_PN0P__1586  (.H(net1636));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[838]$_DFFE_PN0P__1587  (.H(net1637));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[839]$_DFFE_PN0P__1588  (.H(net1638));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[83]$_DFFE_PN0P__1589  (.H(net1639));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[840]$_DFFE_PN0P__1590  (.H(net1640));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[841]$_DFFE_PN0P__1591  (.H(net1641));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[842]$_DFFE_PN0P__1592  (.H(net1642));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[843]$_DFFE_PN0P__1593  (.H(net1643));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[844]$_DFFE_PN0P__1594  (.H(net1644));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[845]$_DFFE_PN0P__1595  (.H(net1645));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[846]$_DFFE_PN0P__1596  (.H(net1646));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[847]$_DFFE_PN0P__1597  (.H(net1647));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[848]$_DFFE_PN0P__1598  (.H(net1648));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[849]$_DFFE_PN0P__1599  (.H(net1649));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[84]$_DFFE_PN0P__1600  (.H(net1650));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[850]$_DFFE_PN0P__1601  (.H(net1651));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[851]$_DFFE_PN0P__1602  (.H(net1652));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[852]$_DFFE_PN0P__1603  (.H(net1653));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[853]$_DFFE_PN0P__1604  (.H(net1654));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[854]$_DFFE_PN0P__1605  (.H(net1655));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[855]$_DFFE_PN0P__1606  (.H(net1656));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[856]$_DFFE_PN0P__1607  (.H(net1657));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[857]$_DFFE_PN0P__1608  (.H(net1658));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[858]$_DFFE_PN0P__1609  (.H(net1659));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[859]$_DFFE_PN0P__1610  (.H(net1660));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[85]$_DFFE_PN0P__1611  (.H(net1661));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[860]$_DFFE_PN0P__1612  (.H(net1662));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[861]$_DFFE_PN0P__1613  (.H(net1663));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[862]$_DFFE_PN0P__1614  (.H(net1664));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[863]$_DFFE_PN0P__1615  (.H(net1665));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[864]$_DFFE_PN0P__1616  (.H(net1666));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[865]$_DFFE_PN0P__1617  (.H(net1667));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[866]$_DFFE_PN0P__1618  (.H(net1668));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[867]$_DFFE_PN0P__1619  (.H(net1669));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[868]$_DFFE_PN0P__1620  (.H(net1670));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[869]$_DFFE_PN0P__1621  (.H(net1671));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[86]$_DFFE_PN0P__1622  (.H(net1672));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[870]$_DFFE_PN0P__1623  (.H(net1673));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[871]$_DFFE_PN0P__1624  (.H(net1674));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[872]$_DFFE_PN0P__1625  (.H(net1675));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[873]$_DFFE_PN0P__1626  (.H(net1676));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[874]$_DFFE_PN0P__1627  (.H(net1677));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[875]$_DFFE_PN0P__1628  (.H(net1678));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[876]$_DFFE_PN0P__1629  (.H(net1679));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[877]$_DFFE_PN0P__1630  (.H(net1680));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[878]$_DFFE_PN0P__1631  (.H(net1681));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[879]$_DFFE_PN0P__1632  (.H(net1682));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[87]$_DFFE_PN0P__1633  (.H(net1683));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[880]$_DFFE_PN0P__1634  (.H(net1684));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[881]$_DFFE_PN0P__1635  (.H(net1685));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[882]$_DFFE_PN0P__1636  (.H(net1686));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[883]$_DFFE_PN0P__1637  (.H(net1687));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[884]$_DFFE_PN0P__1638  (.H(net1688));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[885]$_DFFE_PN0P__1639  (.H(net1689));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[886]$_DFFE_PN0P__1640  (.H(net1690));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[887]$_DFFE_PN0P__1641  (.H(net1691));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[888]$_DFFE_PN0P__1642  (.H(net1692));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[889]$_DFFE_PN0P__1643  (.H(net1693));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[88]$_DFFE_PN0P__1644  (.H(net1694));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[890]$_DFFE_PN0P__1645  (.H(net1695));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[891]$_DFFE_PN0P__1646  (.H(net1696));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[892]$_DFFE_PN0P__1647  (.H(net1697));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[893]$_DFFE_PN0P__1648  (.H(net1698));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[894]$_DFFE_PN0P__1649  (.H(net1699));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[895]$_DFFE_PN0P__1650  (.H(net1700));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[896]$_DFFE_PN0P__1651  (.H(net1701));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[897]$_DFFE_PN0P__1652  (.H(net1702));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[898]$_DFFE_PN0P__1653  (.H(net1703));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[899]$_DFFE_PN0P__1654  (.H(net1704));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[89]$_DFFE_PN0P__1655  (.H(net1705));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[8]$_DFFE_PN0P__1656  (.H(net1706));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[900]$_DFFE_PN0P__1657  (.H(net1707));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[901]$_DFFE_PN0P__1658  (.H(net1708));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[902]$_DFFE_PN0P__1659  (.H(net1709));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[903]$_DFFE_PN0P__1660  (.H(net1710));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[904]$_DFFE_PN0P__1661  (.H(net1711));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[905]$_DFFE_PN0P__1662  (.H(net1712));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[906]$_DFFE_PN0P__1663  (.H(net1713));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[907]$_DFFE_PN0P__1664  (.H(net1714));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[908]$_DFFE_PN0P__1665  (.H(net1715));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[909]$_DFFE_PN0P__1666  (.H(net1716));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[90]$_DFFE_PN0P__1667  (.H(net1717));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[910]$_DFFE_PN0P__1668  (.H(net1718));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[911]$_DFFE_PN0P__1669  (.H(net1719));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[912]$_DFFE_PN0P__1670  (.H(net1720));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[913]$_DFFE_PN0P__1671  (.H(net1721));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[914]$_DFFE_PN0P__1672  (.H(net1722));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[915]$_DFFE_PN0P__1673  (.H(net1723));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[916]$_DFFE_PN0P__1674  (.H(net1724));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[917]$_DFFE_PN0P__1675  (.H(net1725));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[918]$_DFFE_PN0P__1676  (.H(net1726));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[919]$_DFFE_PN0P__1677  (.H(net1727));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[91]$_DFFE_PN0P__1678  (.H(net1728));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[920]$_DFFE_PN0P__1679  (.H(net1729));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[921]$_DFFE_PN0P__1680  (.H(net1730));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[922]$_DFFE_PN0P__1681  (.H(net1731));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[923]$_DFFE_PN0P__1682  (.H(net1732));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[924]$_DFFE_PN0P__1683  (.H(net1733));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[925]$_DFFE_PN0P__1684  (.H(net1734));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[926]$_DFFE_PN0P__1685  (.H(net1735));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[927]$_DFFE_PN0P__1686  (.H(net1736));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[928]$_DFFE_PN0P__1687  (.H(net1737));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[929]$_DFFE_PN0P__1688  (.H(net1738));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[92]$_DFFE_PN0P__1689  (.H(net1739));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[930]$_DFFE_PN0P__1690  (.H(net1740));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[931]$_DFFE_PN0P__1691  (.H(net1741));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[932]$_DFFE_PN0P__1692  (.H(net1742));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[933]$_DFFE_PN0P__1693  (.H(net1743));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[934]$_DFFE_PN0P__1694  (.H(net1744));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[935]$_DFFE_PN0P__1695  (.H(net1745));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[936]$_DFFE_PN0P__1696  (.H(net1746));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[937]$_DFFE_PN0P__1697  (.H(net1747));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[938]$_DFFE_PN0P__1698  (.H(net1748));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[939]$_DFFE_PN0P__1699  (.H(net1749));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[93]$_DFFE_PN0P__1700  (.H(net1750));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[940]$_DFFE_PN0P__1701  (.H(net1751));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[941]$_DFFE_PN0P__1702  (.H(net1752));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[942]$_DFFE_PN0P__1703  (.H(net1753));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[943]$_DFFE_PN0P__1704  (.H(net1754));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[944]$_DFFE_PN0P__1705  (.H(net1755));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[945]$_DFFE_PN0P__1706  (.H(net1756));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[946]$_DFFE_PN0P__1707  (.H(net1757));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[947]$_DFFE_PN0P__1708  (.H(net1758));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[948]$_DFFE_PN0P__1709  (.H(net1759));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[949]$_DFFE_PN0P__1710  (.H(net1760));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[94]$_DFFE_PN0P__1711  (.H(net1761));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[950]$_DFFE_PN0P__1712  (.H(net1762));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[951]$_DFFE_PN0P__1713  (.H(net1763));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[952]$_DFFE_PN0P__1714  (.H(net1764));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[953]$_DFFE_PN0P__1715  (.H(net1765));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[954]$_DFFE_PN0P__1716  (.H(net1766));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[955]$_DFFE_PN0P__1717  (.H(net1767));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[956]$_DFFE_PN0P__1718  (.H(net1768));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[957]$_DFFE_PN0P__1719  (.H(net1769));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[958]$_DFFE_PN0P__1720  (.H(net1770));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[959]$_DFFE_PN0P__1721  (.H(net1771));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[95]$_DFFE_PN0P__1722  (.H(net1772));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[960]$_DFFE_PN0P__1723  (.H(net1773));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[961]$_DFFE_PN0P__1724  (.H(net1774));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[962]$_DFFE_PN0P__1725  (.H(net1775));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[963]$_DFFE_PN0P__1726  (.H(net1776));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[964]$_DFFE_PN0P__1727  (.H(net1777));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[965]$_DFFE_PN0P__1728  (.H(net1778));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[966]$_DFFE_PN0P__1729  (.H(net1779));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[967]$_DFFE_PN0P__1730  (.H(net1780));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[968]$_DFFE_PN0P__1731  (.H(net1781));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[969]$_DFFE_PN0P__1732  (.H(net1782));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[96]$_DFFE_PN0P__1733  (.H(net1783));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[970]$_DFFE_PN0P__1734  (.H(net1784));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[971]$_DFFE_PN0P__1735  (.H(net1785));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[972]$_DFFE_PN0P__1736  (.H(net1786));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[973]$_DFFE_PN0P__1737  (.H(net1787));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[974]$_DFFE_PN0P__1738  (.H(net1788));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[975]$_DFFE_PN0P__1739  (.H(net1789));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[976]$_DFFE_PN0P__1740  (.H(net1790));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[977]$_DFFE_PN0P__1741  (.H(net1791));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[978]$_DFFE_PN0P__1742  (.H(net1792));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[979]$_DFFE_PN0P__1743  (.H(net1793));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[97]$_DFFE_PN0P__1744  (.H(net1794));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[980]$_DFFE_PN0P__1745  (.H(net1795));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[981]$_DFFE_PN0P__1746  (.H(net1796));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[982]$_DFFE_PN0P__1747  (.H(net1797));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[983]$_DFFE_PN0P__1748  (.H(net1798));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[984]$_DFFE_PN0P__1749  (.H(net1799));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[985]$_DFFE_PN0P__1750  (.H(net1800));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[986]$_DFFE_PN0P__1751  (.H(net1801));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[987]$_DFFE_PN0P__1752  (.H(net1802));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[988]$_DFFE_PN0P__1753  (.H(net1803));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[989]$_DFFE_PN0P__1754  (.H(net1804));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[98]$_DFFE_PN0P__1755  (.H(net1805));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[990]$_DFFE_PN0P__1756  (.H(net1806));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[991]$_DFFE_PN0P__1757  (.H(net1807));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[99]$_DFFE_PN0P__1758  (.H(net1808));
 TIEHIx1_ASAP7_75t_R \gen_regfile_ff.register_file_i.rf_reg_q[9]$_DFFE_PN0P__1759  (.H(net1809));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P__1760  (.H(net1810));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P__1761  (.H(net1811));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P__1762  (.H(net1812));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P__1763  (.H(net1813));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.debug_mode_q$_DFFE_PN0P__1764  (.H(net1814));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.exc_req_q$_DFF_PN0__1765  (.H(net1815));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0__1766  (.H(net1816));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.load_err_q$_DFF_PN0__1767  (.H(net1817));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.nmi_mode_q$_DFFE_PN0P__1768  (.H(net1818));
 TIEHIx1_ASAP7_75t_R \id_stage_i.controller_i.store_err_q$_DFF_PN0__1769  (.H(net1819));
 TIEHIx1_ASAP7_75t_R \id_stage_i.g_branch_set_flop.branch_set_q$_DFF_PN0__1770  (.H(net1820));
 TIEHIx1_ASAP7_75t_R \id_stage_i.id_fsm_q$_DFFE_PN0P__1771  (.H(net1821));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[0]$_DFFE_PN0P__1772  (.H(net1822));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[10]$_DFFE_PN0P__1773  (.H(net1823));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[11]$_DFFE_PN0P__1774  (.H(net1824));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[12]$_DFFE_PN0P__1775  (.H(net1825));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[13]$_DFFE_PN0P__1776  (.H(net1826));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[14]$_DFFE_PN0P__1777  (.H(net1827));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[15]$_DFFE_PN0P__1778  (.H(net1828));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[16]$_DFFE_PN0P__1779  (.H(net1829));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[17]$_DFFE_PN0P__1780  (.H(net1830));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[18]$_DFFE_PN0P__1781  (.H(net1831));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[19]$_DFFE_PN0P__1782  (.H(net1832));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[1]$_DFFE_PN0P__1783  (.H(net1833));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[20]$_DFFE_PN0P__1784  (.H(net1834));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[21]$_DFFE_PN0P__1785  (.H(net1835));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[22]$_DFFE_PN0P__1786  (.H(net1836));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[23]$_DFFE_PN0P__1787  (.H(net1837));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[24]$_DFFE_PN0P__1788  (.H(net1838));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[25]$_DFFE_PN0P__1789  (.H(net1839));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[26]$_DFFE_PN0P__1790  (.H(net1840));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[27]$_DFFE_PN0P__1791  (.H(net1841));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[28]$_DFFE_PN0P__1792  (.H(net1842));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[29]$_DFFE_PN0P__1793  (.H(net1843));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[2]$_DFFE_PN0P__1794  (.H(net1844));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[30]$_DFFE_PN0P__1795  (.H(net1845));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[31]$_DFFE_PN0P__1796  (.H(net1846));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[34]$_DFFE_PN0P__1797  (.H(net1847));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[35]$_DFFE_PN0P__1798  (.H(net1848));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[36]$_DFFE_PN0P__1799  (.H(net1849));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[37]$_DFFE_PN0P__1800  (.H(net1850));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[38]$_DFFE_PN0P__1801  (.H(net1851));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[39]$_DFFE_PN0P__1802  (.H(net1852));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[3]$_DFFE_PN0P__1803  (.H(net1853));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[40]$_DFFE_PN0P__1804  (.H(net1854));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[41]$_DFFE_PN0P__1805  (.H(net1855));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[42]$_DFFE_PN0P__1806  (.H(net1856));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[43]$_DFFE_PN0P__1807  (.H(net1857));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[44]$_DFFE_PN0P__1808  (.H(net1858));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[45]$_DFFE_PN0P__1809  (.H(net1859));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[46]$_DFFE_PN0P__1810  (.H(net1860));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[47]$_DFFE_PN0P__1811  (.H(net1861));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[48]$_DFFE_PN0P__1812  (.H(net1862));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[49]$_DFFE_PN0P__1813  (.H(net1863));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[4]$_DFFE_PN0P__1814  (.H(net1864));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[50]$_DFFE_PN0P__1815  (.H(net1865));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[51]$_DFFE_PN0P__1816  (.H(net1866));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[52]$_DFFE_PN0P__1817  (.H(net1867));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[53]$_DFFE_PN0P__1818  (.H(net1868));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[54]$_DFFE_PN0P__1819  (.H(net1869));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[55]$_DFFE_PN0P__1820  (.H(net1870));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[56]$_DFFE_PN0P__1821  (.H(net1871));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[57]$_DFFE_PN0P__1822  (.H(net1872));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[58]$_DFFE_PN0P__1823  (.H(net1873));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[59]$_DFFE_PN0P__1824  (.H(net1874));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[5]$_DFFE_PN0P__1825  (.H(net1875));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[60]$_DFFE_PN0P__1826  (.H(net1876));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[61]$_DFFE_PN0P__1827  (.H(net1877));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[62]$_DFFE_PN0P__1828  (.H(net1878));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[63]$_DFFE_PN0P__1829  (.H(net1879));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[64]$_DFFE_PN0P__1830  (.H(net1880));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[65]$_DFFE_PN0P__1831  (.H(net1881));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[66]$_DFFE_PN0P__1832  (.H(net1882));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[67]$_DFFE_PN0P__1833  (.H(net1883));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[6]$_DFFE_PN0P__1834  (.H(net1884));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[7]$_DFFE_PN0P__1835  (.H(net1885));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[8]$_DFFE_PN0P__1836  (.H(net1886));
 TIEHIx1_ASAP7_75t_R \id_stage_i.imd_val_q[9]$_DFFE_PN0P__1837  (.H(net1887));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0__1838  (.H(net1888));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0__1839  (.H(net1889));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0__1840  (.H(net1890));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0__1841  (.H(net1891));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0__1842  (.H(net1892));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0__1843  (.H(net1893));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0__1844  (.H(net1894));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0__1845  (.H(net1895));
 TIEHIx1_ASAP7_75t_R \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0__1846  (.H(net1896));
 TIEHIx1_ASAP7_75t_R \if_stage_i.instr_valid_id_q$_DFF_PN0__1847  (.H(net1897));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[0]$_DFFE_PN0P__1848  (.H(net1898));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[10]$_DFFE_PN0P__1849  (.H(net1899));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[11]$_DFFE_PN0P__1850  (.H(net1900));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[12]$_DFFE_PN0P__1851  (.H(net1901));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[13]$_DFFE_PN0P__1852  (.H(net1902));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[14]$_DFFE_PN0P__1853  (.H(net1903));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[15]$_DFFE_PN0P__1854  (.H(net1904));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[16]$_DFFE_PN0P__1855  (.H(net1905));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[17]$_DFFE_PN0P__1856  (.H(net1906));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[18]$_DFFE_PN0P__1857  (.H(net1907));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[19]$_DFFE_PN0P__1858  (.H(net1908));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[1]$_DFFE_PN0P__1859  (.H(net1909));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[20]$_DFFE_PN0P__1860  (.H(net1910));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[21]$_DFFE_PN0P__1861  (.H(net1911));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[22]$_DFFE_PN0P__1862  (.H(net1912));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[23]$_DFFE_PN0P__1863  (.H(net1913));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[24]$_DFFE_PN0P__1864  (.H(net1914));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[25]$_DFFE_PN0P__1865  (.H(net1915));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[26]$_DFFE_PN0P__1866  (.H(net1916));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[27]$_DFFE_PN0P__1867  (.H(net1917));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[28]$_DFFE_PN0P__1868  (.H(net1918));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[29]$_DFFE_PN0P__1869  (.H(net1919));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[2]$_DFFE_PN0P__1870  (.H(net1920));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[30]$_DFFE_PN0P__1871  (.H(net1921));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[31]$_DFFE_PN0P__1872  (.H(net1922));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[3]$_DFFE_PN0P__1873  (.H(net1923));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[4]$_DFFE_PN0P__1874  (.H(net1924));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[5]$_DFFE_PN0P__1875  (.H(net1925));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[6]$_DFFE_PN0P__1876  (.H(net1926));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[7]$_DFFE_PN0P__1877  (.H(net1927));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[8]$_DFFE_PN0P__1878  (.H(net1928));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.addr_last_q[9]$_DFFE_PN0P__1879  (.H(net1929));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P__1880  (.H(net1930));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.data_we_q$_DFFE_PN0P__1881  (.H(net1931));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P__1882  (.H(net1932));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P__1883  (.H(net1933));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P__1884  (.H(net1934));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P__1885  (.H(net1935));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.lsu_err_q$_DFFE_PN0P__1886  (.H(net1936));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P__1887  (.H(net1937));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P__1888  (.H(net1938));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[0]$_DFFE_PN0P__1889  (.H(net1939));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[10]$_DFFE_PN0P__1890  (.H(net1940));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[11]$_DFFE_PN0P__1891  (.H(net1941));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[12]$_DFFE_PN0P__1892  (.H(net1942));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[13]$_DFFE_PN0P__1893  (.H(net1943));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[14]$_DFFE_PN0P__1894  (.H(net1944));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[15]$_DFFE_PN0P__1895  (.H(net1945));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[16]$_DFFE_PN0P__1896  (.H(net1946));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[17]$_DFFE_PN0P__1897  (.H(net1947));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[18]$_DFFE_PN0P__1898  (.H(net1948));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[19]$_DFFE_PN0P__1899  (.H(net1949));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[1]$_DFFE_PN0P__1900  (.H(net1950));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[20]$_DFFE_PN0P__1901  (.H(net1951));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[21]$_DFFE_PN0P__1902  (.H(net1952));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[22]$_DFFE_PN0P__1903  (.H(net1953));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[23]$_DFFE_PN0P__1904  (.H(net1954));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[2]$_DFFE_PN0P__1905  (.H(net1955));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[3]$_DFFE_PN0P__1906  (.H(net1956));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[4]$_DFFE_PN0P__1907  (.H(net1957));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[5]$_DFFE_PN0P__1908  (.H(net1958));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[6]$_DFFE_PN0P__1909  (.H(net1959));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[7]$_DFFE_PN0P__1910  (.H(net1960));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[8]$_DFFE_PN0P__1911  (.H(net1961));
 TIEHIx1_ASAP7_75t_R \load_store_unit_i.rdata_q[9]$_DFFE_PN0P__1912  (.H(net1962));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk_i (.A(clk_i),
    .Y(clknet_0_clk_i));
 BUFx16f_ASAP7_75t_R clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_1_0__leaf_clk_i));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_0_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_1_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_2_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_3_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_4_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_5_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_6_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_7_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_8_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_9_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_10_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_11_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_12_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_13_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_14_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_15_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_16_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk_i_regs (.A(clknet_2_2__leaf_clk_i_regs),
    .Y(clknet_leaf_17_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_18_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_19_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_20_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_21_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_22_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_23_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_24_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_25_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_26_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_27_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_28_clk_i_regs (.A(clknet_2_3__leaf_clk_i_regs),
    .Y(clknet_leaf_28_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_29_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_29_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_30_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_30_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_31_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_31_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_32_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_32_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_33_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_33_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_34_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_34_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_35_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_35_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_36_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_36_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_37_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_37_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_38_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_38_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_39_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_39_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_40_clk_i_regs (.A(clknet_2_1__leaf_clk_i_regs),
    .Y(clknet_leaf_40_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_41_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_41_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_42_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_42_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_43_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_43_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_44_clk_i_regs (.A(clknet_2_0__leaf_clk_i_regs),
    .Y(clknet_leaf_44_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk_i_regs (.A(clk_i_regs),
    .Y(clknet_0_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_2_0__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Y(clknet_2_0__leaf_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_2_1__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Y(clknet_2_1__leaf_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_2_2__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Y(clknet_2_2__leaf_clk_i_regs));
 BUFx16f_ASAP7_75t_R clkbuf_2_3__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .Y(clknet_2_3__leaf_clk_i_regs));
 INVx8_ASAP7_75t_R clkload0 (.A(clknet_2_2__leaf_clk_i_regs));
 BUFx24_ASAP7_75t_R clkload1 (.A(clknet_2_3__leaf_clk_i_regs));
 BUFx8_ASAP7_75t_R clkload2 (.A(clknet_leaf_0_clk_i_regs));
 INVxp67_ASAP7_75t_R clkload3 (.A(clknet_leaf_1_clk_i_regs));
 INVxp67_ASAP7_75t_R clkload4 (.A(clknet_leaf_2_clk_i_regs));
 BUFx12_ASAP7_75t_R clkload5 (.A(clknet_leaf_4_clk_i_regs));
 BUFx8_ASAP7_75t_R clkload6 (.A(clknet_leaf_5_clk_i_regs));
 BUFx12_ASAP7_75t_R clkload7 (.A(clknet_leaf_6_clk_i_regs));
 CKINVDCx5p33_ASAP7_75t_R clkload8 (.A(clknet_leaf_7_clk_i_regs));
 INVxp67_ASAP7_75t_R clkload9 (.A(clknet_leaf_41_clk_i_regs));
 INVx5_ASAP7_75t_R clkload10 (.A(clknet_leaf_42_clk_i_regs));
 INVx3_ASAP7_75t_R clkload11 (.A(clknet_leaf_43_clk_i_regs));
 INVx4_ASAP7_75t_R clkload12 (.A(clknet_leaf_44_clk_i_regs));
 INVx5_ASAP7_75t_R clkload13 (.A(clknet_leaf_29_clk_i_regs));
 INVx4_ASAP7_75t_R clkload14 (.A(clknet_leaf_31_clk_i_regs));
 INVx3_ASAP7_75t_R clkload15 (.A(clknet_leaf_32_clk_i_regs));
 INVx3_ASAP7_75t_R clkload16 (.A(clknet_leaf_33_clk_i_regs));
 BUFx12_ASAP7_75t_R clkload17 (.A(clknet_leaf_34_clk_i_regs));
 BUFx8_ASAP7_75t_R clkload18 (.A(clknet_leaf_35_clk_i_regs));
 BUFx12_ASAP7_75t_R clkload19 (.A(clknet_leaf_37_clk_i_regs));
 CKINVDCx8_ASAP7_75t_R clkload20 (.A(clknet_leaf_38_clk_i_regs));
 CKINVDCx8_ASAP7_75t_R clkload21 (.A(clknet_leaf_39_clk_i_regs));
 INVx4_ASAP7_75t_R clkload22 (.A(clknet_leaf_40_clk_i_regs));
 CKINVDCx5p33_ASAP7_75t_R clkload23 (.A(clknet_leaf_8_clk_i_regs));
 BUFx12_ASAP7_75t_R clkload24 (.A(clknet_leaf_9_clk_i_regs));
 BUFx12_ASAP7_75t_R clkload25 (.A(clknet_leaf_10_clk_i_regs));
 INVxp67_ASAP7_75t_R clkload26 (.A(clknet_leaf_11_clk_i_regs));
 BUFx12_ASAP7_75t_R clkload27 (.A(clknet_leaf_12_clk_i_regs));
 BUFx8_ASAP7_75t_R clkload28 (.A(clknet_leaf_13_clk_i_regs));
 INVx11_ASAP7_75t_R clkload29 (.A(clknet_leaf_15_clk_i_regs));
 INVx3_ASAP7_75t_R clkload30 (.A(clknet_leaf_16_clk_i_regs));
 BUFx8_ASAP7_75t_R clkload31 (.A(clknet_leaf_17_clk_i_regs));
 CKINVDCx6p67_ASAP7_75t_R clkload32 (.A(clknet_leaf_19_clk_i_regs));
 CKINVDCx6p67_ASAP7_75t_R clkload33 (.A(clknet_leaf_20_clk_i_regs));
 INVx5_ASAP7_75t_R clkload34 (.A(clknet_leaf_21_clk_i_regs));
 INVxp67_ASAP7_75t_R clkload35 (.A(clknet_leaf_22_clk_i_regs));
 INVx5_ASAP7_75t_R clkload36 (.A(clknet_leaf_23_clk_i_regs));
 CKINVDCx12_ASAP7_75t_R clkload37 (.A(clknet_leaf_24_clk_i_regs));
 INVx13_ASAP7_75t_R clkload38 (.A(clknet_leaf_25_clk_i_regs));
 INVx5_ASAP7_75t_R clkload39 (.A(clknet_leaf_26_clk_i_regs));
 CKINVDCx6p67_ASAP7_75t_R clkload40 (.A(clknet_leaf_27_clk_i_regs));
 CKINVDCx5p33_ASAP7_75t_R clkload41 (.A(clknet_leaf_28_clk_i_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_1_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_2_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_3_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_4_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_5_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_6_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_7_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_8_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_9_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_11_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_14_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_15_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_18_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_19_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_21_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_23_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_24_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_25_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_26_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_27_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_28_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_28_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_29_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_29_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_30_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_30_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_31_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_31_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_32_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_32_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_33_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_33_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_34_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_34_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_35_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_35_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_36_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_36_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_37_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_37_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_38_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_38_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_39_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_39_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_40_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_40_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_41_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_41_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_42_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_42_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_43_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_43_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_44_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_44_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_45_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_45_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_46_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_46_clk));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_0_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_1_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_2_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_3_0_clk));
 CKINVDCx20_ASAP7_75t_R clkload42 (.A(clknet_2_0_0_clk));
 CKINVDCx12_ASAP7_75t_R clkload43 (.A(clknet_2_1_0_clk));
 CKINVDCx8_ASAP7_75t_R clkload44 (.A(clknet_leaf_37_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload45 (.A(clknet_leaf_38_clk));
 INVx5_ASAP7_75t_R clkload46 (.A(clknet_leaf_40_clk));
 INVx4_ASAP7_75t_R clkload47 (.A(clknet_leaf_41_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload48 (.A(clknet_leaf_42_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload49 (.A(clknet_leaf_43_clk));
 CKINVDCx8_ASAP7_75t_R clkload50 (.A(clknet_leaf_44_clk));
 INVxp67_ASAP7_75t_R clkload51 (.A(clknet_leaf_11_clk));
 INVx4_ASAP7_75t_R clkload52 (.A(clknet_leaf_28_clk));
 BUFx12_ASAP7_75t_R clkload53 (.A(clknet_leaf_29_clk));
 INVxp67_ASAP7_75t_R clkload54 (.A(clknet_leaf_30_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload55 (.A(clknet_leaf_31_clk));
 BUFx8_ASAP7_75t_R clkload56 (.A(clknet_leaf_32_clk));
 INVx3_ASAP7_75t_R clkload57 (.A(clknet_leaf_33_clk));
 BUFx12_ASAP7_75t_R clkload58 (.A(clknet_leaf_34_clk));
 INVx3_ASAP7_75t_R clkload59 (.A(clknet_leaf_35_clk));
 BUFx12_ASAP7_75t_R clkload60 (.A(clknet_leaf_36_clk));
 BUFx4f_ASAP7_75t_R clkload61 (.A(clknet_leaf_0_clk));
 INVxp67_ASAP7_75t_R clkload62 (.A(clknet_leaf_1_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload63 (.A(clknet_leaf_2_clk));
 BUFx4f_ASAP7_75t_R clkload64 (.A(clknet_leaf_4_clk));
 INVx3_ASAP7_75t_R clkload65 (.A(clknet_leaf_5_clk));
 BUFx8_ASAP7_75t_R clkload66 (.A(clknet_leaf_6_clk));
 INVxp67_ASAP7_75t_R clkload67 (.A(clknet_leaf_7_clk));
 BUFx5_ASAP7_75t_R clkload68 (.A(clknet_leaf_8_clk));
 INVx4_ASAP7_75t_R clkload69 (.A(clknet_leaf_9_clk));
 BUFx12_ASAP7_75t_R clkload70 (.A(clknet_leaf_13_clk));
 INVx5_ASAP7_75t_R clkload71 (.A(clknet_leaf_14_clk));
 INVx8_ASAP7_75t_R clkload72 (.A(clknet_leaf_45_clk));
 CKINVDCx11_ASAP7_75t_R clkload73 (.A(clknet_leaf_46_clk));
 INVx3_ASAP7_75t_R clkload74 (.A(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkload75 (.A(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkload76 (.A(clknet_leaf_15_clk));
 INVx5_ASAP7_75t_R clkload77 (.A(clknet_leaf_16_clk));
 INVx3_ASAP7_75t_R clkload78 (.A(clknet_leaf_17_clk));
 INVx3_ASAP7_75t_R clkload79 (.A(clknet_leaf_18_clk));
 BUFx8_ASAP7_75t_R clkload80 (.A(clknet_leaf_19_clk));
 BUFx12_ASAP7_75t_R clkload81 (.A(clknet_leaf_20_clk));
 BUFx8_ASAP7_75t_R clkload82 (.A(clknet_leaf_21_clk));
 BUFx8_ASAP7_75t_R clkload83 (.A(clknet_leaf_22_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload84 (.A(clknet_leaf_23_clk));
 BUFx8_ASAP7_75t_R clkload85 (.A(clknet_leaf_24_clk));
 INVx3_ASAP7_75t_R clkload86 (.A(clknet_leaf_25_clk));
 BUFx16f_ASAP7_75t_R delaybuf_0_core_clock (.A(delaynet_0_core_clock),
    .Y(delaynet_1_core_clock));
 BUFx16f_ASAP7_75t_R delaybuf_1_core_clock (.A(delaynet_1_core_clock),
    .Y(delaynet_2_core_clock));
 BUFx16f_ASAP7_75t_R delaybuf_2_core_clock (.A(delaynet_2_core_clock),
    .Y(clk_i_regs));
 BUFx3_ASAP7_75t_R rebuffer1 (.A(_18080_),
    .Y(net1963));
 BUFx2_ASAP7_75t_R rebuffer2 (.A(net1963),
    .Y(net1964));
 BUFx2_ASAP7_75t_R rebuffer3 (.A(net1964),
    .Y(net1965));
 BUFx2_ASAP7_75t_R rebuffer4 (.A(net1964),
    .Y(net1966));
 BUFx2_ASAP7_75t_R rebuffer5 (.A(net1966),
    .Y(net1967));
 BUFx2_ASAP7_75t_R rebuffer6 (.A(net1966),
    .Y(net1968));
 BUFx3_ASAP7_75t_R rebuffer7 (.A(_17962_),
    .Y(net1969));
 BUFx3_ASAP7_75t_R rebuffer8 (.A(net1969),
    .Y(net1970));
 BUFx2_ASAP7_75t_R rebuffer9 (.A(net1970),
    .Y(net1971));
 BUFx3_ASAP7_75t_R rebuffer10 (.A(net1971),
    .Y(net1972));
 BUFx3_ASAP7_75t_R rebuffer11 (.A(_02294_),
    .Y(net1973));
 BUFx3_ASAP7_75t_R rebuffer12 (.A(net1973),
    .Y(net1974));
 BUFx2_ASAP7_75t_R rebuffer13 (.A(net1974),
    .Y(net1975));
 BUFx3_ASAP7_75t_R rebuffer14 (.A(_00822_),
    .Y(net1976));
 BUFx2_ASAP7_75t_R rebuffer15 (.A(net1976),
    .Y(net1977));
 BUFx2_ASAP7_75t_R rebuffer16 (.A(net1977),
    .Y(net1978));
 BUFx2_ASAP7_75t_R rebuffer17 (.A(_00810_),
    .Y(net1979));
 BUFx2_ASAP7_75t_R rebuffer18 (.A(net1979),
    .Y(net1980));
 BUFx2_ASAP7_75t_R rebuffer19 (.A(_00805_),
    .Y(net1981));
 BUFx2_ASAP7_75t_R rebuffer20 (.A(net1981),
    .Y(net1982));
 BUFx3_ASAP7_75t_R rebuffer21 (.A(_00855_),
    .Y(net1983));
 BUFx2_ASAP7_75t_R rebuffer22 (.A(net1983),
    .Y(net1984));
 BUFx2_ASAP7_75t_R rebuffer23 (.A(net1984),
    .Y(net1985));
 BUFx2_ASAP7_75t_R rebuffer24 (.A(net1983),
    .Y(net1986));
 BUFx2_ASAP7_75t_R rebuffer25 (.A(net1986),
    .Y(net1987));
 BUFx2_ASAP7_75t_R rebuffer26 (.A(net1987),
    .Y(net1988));
 BUFx2_ASAP7_75t_R rebuffer27 (.A(_00813_),
    .Y(net1989));
 BUFx2_ASAP7_75t_R rebuffer28 (.A(_00406_),
    .Y(net1990));
 BUFx2_ASAP7_75t_R rebuffer29 (.A(_00793_),
    .Y(net1991));
 BUFx2_ASAP7_75t_R rebuffer30 (.A(net1991),
    .Y(net1992));
 BUFx2_ASAP7_75t_R rebuffer31 (.A(net1991),
    .Y(net1993));
 BUFx2_ASAP7_75t_R rebuffer32 (.A(net1993),
    .Y(net1994));
 BUFx2_ASAP7_75t_R rebuffer33 (.A(_02296_),
    .Y(net1995));
 BUFx2_ASAP7_75t_R rebuffer34 (.A(net1995),
    .Y(net1996));
 BUFx3_ASAP7_75t_R rebuffer35 (.A(_17914_),
    .Y(net1997));
 BUFx2_ASAP7_75t_R rebuffer36 (.A(net1997),
    .Y(net1998));
 BUFx2_ASAP7_75t_R rebuffer37 (.A(net1997),
    .Y(net1999));
 BUFx2_ASAP7_75t_R rebuffer38 (.A(_00401_),
    .Y(net2000));
 BUFx2_ASAP7_75t_R rebuffer39 (.A(net2000),
    .Y(net2001));
 BUFx2_ASAP7_75t_R rebuffer40 (.A(_18777_),
    .Y(net2002));
 BUFx2_ASAP7_75t_R clone41 (.A(_14921_),
    .Y(net2003));
 BUFx4_ASAP7_75t_R clone42 (.A(_13593_),
    .Y(net2004));
 BUFx4_ASAP7_75t_R clone43 (.A(_00401_),
    .Y(net2005));
 BUFx2_ASAP7_75t_R rebuffer44 (.A(_13559_),
    .Y(net2006));
 BUFx4_ASAP7_75t_R clone45 (.A(_14922_),
    .Y(net2007));
 BUFx2_ASAP7_75t_R rebuffer47 (.A(net2008),
    .Y(net2009));
 BUFx3_ASAP7_75t_R rebuffer48 (.A(_18114_),
    .Y(net2010));
 BUFx2_ASAP7_75t_R rebuffer49 (.A(net2010),
    .Y(net2011));
 BUFx2_ASAP7_75t_R rebuffer50 (.A(net2011),
    .Y(net2012));
 BUFx2_ASAP7_75t_R clone52 (.A(_00024_),
    .Y(net2014));
 BUFx2_ASAP7_75t_R rebuffer53 (.A(_00013_),
    .Y(net2015));
 BUFx2_ASAP7_75t_R rebuffer54 (.A(net2015),
    .Y(net2016));
 BUFx2_ASAP7_75t_R rebuffer55 (.A(net2015),
    .Y(net2017));
 BUFx2_ASAP7_75t_R rebuffer56 (.A(_01456_),
    .Y(net2018));
 BUFx2_ASAP7_75t_R rebuffer57 (.A(net2018),
    .Y(net2019));
 BUFx4_ASAP7_75t_R clone58 (.A(_13382_),
    .Y(net2020));
 BUFx16f_ASAP7_75t_R load_slew1 (.A(net59),
    .Y(net2021));
 BUFx3_ASAP7_75t_R rebuffer41 (.A(_00205_),
    .Y(net2022));
 AND2x4_ASAP7_75t_R clone44 (.A(_05168_),
    .B(_05309_),
    .Y(net2023));
 BUFx2_ASAP7_75t_R rebuffer45 (.A(_18143_),
    .Y(net2024));
 BUFx3_ASAP7_75t_R rebuffer51 (.A(net2024),
    .Y(net2025));
 BUFx3_ASAP7_75t_R rebuffer52 (.A(net2025),
    .Y(net2026));
 BUFx3_ASAP7_75t_R rebuffer58 (.A(net2026),
    .Y(net2027));
 BUFx2_ASAP7_75t_R rebuffer59 (.A(_00921_),
    .Y(net2028));
 BUFx2_ASAP7_75t_R rebuffer60 (.A(net2028),
    .Y(net2029));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662 ();
 DECAPx6_ASAP7_75t_R FILLER_0_684 ();
 FILLER_ASAP7_75t_R FILLER_0_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_828 ();
 FILLER_ASAP7_75t_R FILLER_0_842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_898 ();
 DECAPx1_ASAP7_75t_R FILLER_0_920 ();
 DECAPx4_ASAP7_75t_R FILLER_0_926 ();
 DECAPx4_ASAP7_75t_R FILLER_0_941 ();
 FILLER_ASAP7_75t_R FILLER_0_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_953 ();
 DECAPx10_ASAP7_75t_R FILLER_0_959 ();
 DECAPx10_ASAP7_75t_R FILLER_0_981 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1377 ();
 FILLER_ASAP7_75t_R FILLER_0_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1388 ();
 FILLER_ASAP7_75t_R FILLER_0_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_1_222 ();
 DECAPx10_ASAP7_75t_R FILLER_1_244 ();
 DECAPx10_ASAP7_75t_R FILLER_1_266 ();
 DECAPx10_ASAP7_75t_R FILLER_1_288 ();
 DECAPx10_ASAP7_75t_R FILLER_1_310 ();
 DECAPx10_ASAP7_75t_R FILLER_1_332 ();
 DECAPx10_ASAP7_75t_R FILLER_1_354 ();
 DECAPx10_ASAP7_75t_R FILLER_1_376 ();
 DECAPx10_ASAP7_75t_R FILLER_1_398 ();
 DECAPx10_ASAP7_75t_R FILLER_1_420 ();
 DECAPx10_ASAP7_75t_R FILLER_1_442 ();
 DECAPx10_ASAP7_75t_R FILLER_1_464 ();
 DECAPx10_ASAP7_75t_R FILLER_1_486 ();
 DECAPx10_ASAP7_75t_R FILLER_1_508 ();
 DECAPx10_ASAP7_75t_R FILLER_1_530 ();
 DECAPx10_ASAP7_75t_R FILLER_1_552 ();
 DECAPx10_ASAP7_75t_R FILLER_1_574 ();
 DECAPx10_ASAP7_75t_R FILLER_1_596 ();
 DECAPx10_ASAP7_75t_R FILLER_1_618 ();
 DECAPx10_ASAP7_75t_R FILLER_1_640 ();
 DECAPx10_ASAP7_75t_R FILLER_1_662 ();
 DECAPx10_ASAP7_75t_R FILLER_1_684 ();
 FILLER_ASAP7_75t_R FILLER_1_721 ();
 DECAPx4_ASAP7_75t_R FILLER_1_733 ();
 FILLER_ASAP7_75t_R FILLER_1_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_745 ();
 DECAPx10_ASAP7_75t_R FILLER_1_801 ();
 DECAPx10_ASAP7_75t_R FILLER_1_823 ();
 DECAPx10_ASAP7_75t_R FILLER_1_845 ();
 DECAPx10_ASAP7_75t_R FILLER_1_867 ();
 DECAPx10_ASAP7_75t_R FILLER_1_889 ();
 DECAPx4_ASAP7_75t_R FILLER_1_911 ();
 FILLER_ASAP7_75t_R FILLER_1_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_923 ();
 DECAPx10_ASAP7_75t_R FILLER_1_926 ();
 DECAPx10_ASAP7_75t_R FILLER_1_948 ();
 DECAPx10_ASAP7_75t_R FILLER_1_970 ();
 DECAPx10_ASAP7_75t_R FILLER_1_992 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_1_1388 ();
 FILLER_ASAP7_75t_R FILLER_1_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_2_222 ();
 DECAPx10_ASAP7_75t_R FILLER_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_2_266 ();
 DECAPx10_ASAP7_75t_R FILLER_2_288 ();
 DECAPx10_ASAP7_75t_R FILLER_2_310 ();
 DECAPx10_ASAP7_75t_R FILLER_2_332 ();
 DECAPx10_ASAP7_75t_R FILLER_2_354 ();
 DECAPx10_ASAP7_75t_R FILLER_2_376 ();
 DECAPx10_ASAP7_75t_R FILLER_2_398 ();
 DECAPx10_ASAP7_75t_R FILLER_2_420 ();
 DECAPx6_ASAP7_75t_R FILLER_2_442 ();
 DECAPx2_ASAP7_75t_R FILLER_2_456 ();
 DECAPx10_ASAP7_75t_R FILLER_2_464 ();
 DECAPx10_ASAP7_75t_R FILLER_2_486 ();
 DECAPx10_ASAP7_75t_R FILLER_2_508 ();
 DECAPx10_ASAP7_75t_R FILLER_2_530 ();
 DECAPx10_ASAP7_75t_R FILLER_2_552 ();
 DECAPx10_ASAP7_75t_R FILLER_2_574 ();
 DECAPx10_ASAP7_75t_R FILLER_2_596 ();
 DECAPx10_ASAP7_75t_R FILLER_2_618 ();
 DECAPx10_ASAP7_75t_R FILLER_2_640 ();
 DECAPx10_ASAP7_75t_R FILLER_2_662 ();
 DECAPx10_ASAP7_75t_R FILLER_2_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_706 ();
 DECAPx10_ASAP7_75t_R FILLER_2_712 ();
 DECAPx10_ASAP7_75t_R FILLER_2_734 ();
 DECAPx6_ASAP7_75t_R FILLER_2_756 ();
 DECAPx2_ASAP7_75t_R FILLER_2_770 ();
 DECAPx1_ASAP7_75t_R FILLER_2_781 ();
 DECAPx10_ASAP7_75t_R FILLER_2_790 ();
 DECAPx10_ASAP7_75t_R FILLER_2_812 ();
 DECAPx10_ASAP7_75t_R FILLER_2_834 ();
 DECAPx10_ASAP7_75t_R FILLER_2_856 ();
 DECAPx10_ASAP7_75t_R FILLER_2_878 ();
 DECAPx10_ASAP7_75t_R FILLER_2_900 ();
 DECAPx10_ASAP7_75t_R FILLER_2_922 ();
 DECAPx10_ASAP7_75t_R FILLER_2_944 ();
 DECAPx10_ASAP7_75t_R FILLER_2_966 ();
 DECAPx10_ASAP7_75t_R FILLER_2_988 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1362 ();
 FILLER_ASAP7_75t_R FILLER_2_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_2_1388 ();
 FILLER_ASAP7_75t_R FILLER_2_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_3_222 ();
 DECAPx10_ASAP7_75t_R FILLER_3_244 ();
 DECAPx10_ASAP7_75t_R FILLER_3_266 ();
 DECAPx10_ASAP7_75t_R FILLER_3_288 ();
 DECAPx10_ASAP7_75t_R FILLER_3_310 ();
 DECAPx10_ASAP7_75t_R FILLER_3_332 ();
 DECAPx10_ASAP7_75t_R FILLER_3_354 ();
 DECAPx10_ASAP7_75t_R FILLER_3_376 ();
 DECAPx10_ASAP7_75t_R FILLER_3_398 ();
 DECAPx10_ASAP7_75t_R FILLER_3_420 ();
 DECAPx10_ASAP7_75t_R FILLER_3_442 ();
 DECAPx10_ASAP7_75t_R FILLER_3_464 ();
 DECAPx10_ASAP7_75t_R FILLER_3_486 ();
 DECAPx10_ASAP7_75t_R FILLER_3_508 ();
 DECAPx10_ASAP7_75t_R FILLER_3_530 ();
 DECAPx10_ASAP7_75t_R FILLER_3_552 ();
 DECAPx10_ASAP7_75t_R FILLER_3_574 ();
 DECAPx10_ASAP7_75t_R FILLER_3_596 ();
 DECAPx10_ASAP7_75t_R FILLER_3_618 ();
 DECAPx10_ASAP7_75t_R FILLER_3_640 ();
 DECAPx10_ASAP7_75t_R FILLER_3_662 ();
 DECAPx10_ASAP7_75t_R FILLER_3_684 ();
 DECAPx10_ASAP7_75t_R FILLER_3_706 ();
 DECAPx10_ASAP7_75t_R FILLER_3_728 ();
 DECAPx10_ASAP7_75t_R FILLER_3_750 ();
 DECAPx10_ASAP7_75t_R FILLER_3_772 ();
 DECAPx10_ASAP7_75t_R FILLER_3_794 ();
 DECAPx10_ASAP7_75t_R FILLER_3_816 ();
 DECAPx10_ASAP7_75t_R FILLER_3_838 ();
 DECAPx10_ASAP7_75t_R FILLER_3_860 ();
 DECAPx10_ASAP7_75t_R FILLER_3_882 ();
 DECAPx6_ASAP7_75t_R FILLER_3_904 ();
 DECAPx2_ASAP7_75t_R FILLER_3_918 ();
 DECAPx10_ASAP7_75t_R FILLER_3_926 ();
 DECAPx10_ASAP7_75t_R FILLER_3_948 ();
 DECAPx10_ASAP7_75t_R FILLER_3_970 ();
 DECAPx10_ASAP7_75t_R FILLER_3_992 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1388 ();
 FILLER_ASAP7_75t_R FILLER_3_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_4_222 ();
 DECAPx10_ASAP7_75t_R FILLER_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_4_266 ();
 DECAPx10_ASAP7_75t_R FILLER_4_288 ();
 DECAPx10_ASAP7_75t_R FILLER_4_310 ();
 DECAPx10_ASAP7_75t_R FILLER_4_332 ();
 DECAPx10_ASAP7_75t_R FILLER_4_354 ();
 DECAPx10_ASAP7_75t_R FILLER_4_376 ();
 DECAPx10_ASAP7_75t_R FILLER_4_398 ();
 DECAPx10_ASAP7_75t_R FILLER_4_420 ();
 DECAPx6_ASAP7_75t_R FILLER_4_442 ();
 DECAPx2_ASAP7_75t_R FILLER_4_456 ();
 DECAPx10_ASAP7_75t_R FILLER_4_464 ();
 DECAPx10_ASAP7_75t_R FILLER_4_486 ();
 DECAPx10_ASAP7_75t_R FILLER_4_508 ();
 DECAPx10_ASAP7_75t_R FILLER_4_530 ();
 DECAPx10_ASAP7_75t_R FILLER_4_552 ();
 DECAPx10_ASAP7_75t_R FILLER_4_574 ();
 DECAPx10_ASAP7_75t_R FILLER_4_596 ();
 DECAPx10_ASAP7_75t_R FILLER_4_618 ();
 DECAPx10_ASAP7_75t_R FILLER_4_640 ();
 DECAPx10_ASAP7_75t_R FILLER_4_662 ();
 DECAPx10_ASAP7_75t_R FILLER_4_684 ();
 DECAPx10_ASAP7_75t_R FILLER_4_706 ();
 DECAPx10_ASAP7_75t_R FILLER_4_728 ();
 DECAPx10_ASAP7_75t_R FILLER_4_750 ();
 DECAPx10_ASAP7_75t_R FILLER_4_772 ();
 DECAPx10_ASAP7_75t_R FILLER_4_794 ();
 DECAPx10_ASAP7_75t_R FILLER_4_816 ();
 DECAPx10_ASAP7_75t_R FILLER_4_838 ();
 DECAPx10_ASAP7_75t_R FILLER_4_860 ();
 DECAPx10_ASAP7_75t_R FILLER_4_882 ();
 DECAPx10_ASAP7_75t_R FILLER_4_904 ();
 DECAPx10_ASAP7_75t_R FILLER_4_926 ();
 DECAPx10_ASAP7_75t_R FILLER_4_948 ();
 DECAPx10_ASAP7_75t_R FILLER_4_970 ();
 DECAPx10_ASAP7_75t_R FILLER_4_992 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1388 ();
 FILLER_ASAP7_75t_R FILLER_4_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx6_ASAP7_75t_R FILLER_5_46 ();
 FILLER_ASAP7_75t_R FILLER_5_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_62 ();
 DECAPx10_ASAP7_75t_R FILLER_5_74 ();
 DECAPx10_ASAP7_75t_R FILLER_5_96 ();
 DECAPx10_ASAP7_75t_R FILLER_5_118 ();
 DECAPx10_ASAP7_75t_R FILLER_5_140 ();
 DECAPx10_ASAP7_75t_R FILLER_5_162 ();
 DECAPx10_ASAP7_75t_R FILLER_5_184 ();
 DECAPx10_ASAP7_75t_R FILLER_5_206 ();
 DECAPx10_ASAP7_75t_R FILLER_5_228 ();
 DECAPx10_ASAP7_75t_R FILLER_5_250 ();
 DECAPx10_ASAP7_75t_R FILLER_5_272 ();
 DECAPx10_ASAP7_75t_R FILLER_5_294 ();
 DECAPx10_ASAP7_75t_R FILLER_5_316 ();
 DECAPx10_ASAP7_75t_R FILLER_5_338 ();
 DECAPx10_ASAP7_75t_R FILLER_5_360 ();
 DECAPx10_ASAP7_75t_R FILLER_5_382 ();
 DECAPx10_ASAP7_75t_R FILLER_5_404 ();
 DECAPx10_ASAP7_75t_R FILLER_5_426 ();
 DECAPx10_ASAP7_75t_R FILLER_5_448 ();
 DECAPx10_ASAP7_75t_R FILLER_5_470 ();
 DECAPx10_ASAP7_75t_R FILLER_5_492 ();
 DECAPx10_ASAP7_75t_R FILLER_5_514 ();
 DECAPx10_ASAP7_75t_R FILLER_5_536 ();
 DECAPx10_ASAP7_75t_R FILLER_5_558 ();
 DECAPx10_ASAP7_75t_R FILLER_5_580 ();
 DECAPx10_ASAP7_75t_R FILLER_5_602 ();
 DECAPx10_ASAP7_75t_R FILLER_5_624 ();
 DECAPx10_ASAP7_75t_R FILLER_5_646 ();
 DECAPx10_ASAP7_75t_R FILLER_5_668 ();
 DECAPx10_ASAP7_75t_R FILLER_5_690 ();
 DECAPx10_ASAP7_75t_R FILLER_5_712 ();
 DECAPx10_ASAP7_75t_R FILLER_5_734 ();
 DECAPx10_ASAP7_75t_R FILLER_5_756 ();
 DECAPx10_ASAP7_75t_R FILLER_5_778 ();
 DECAPx10_ASAP7_75t_R FILLER_5_800 ();
 DECAPx10_ASAP7_75t_R FILLER_5_822 ();
 DECAPx10_ASAP7_75t_R FILLER_5_844 ();
 DECAPx10_ASAP7_75t_R FILLER_5_866 ();
 DECAPx10_ASAP7_75t_R FILLER_5_888 ();
 DECAPx6_ASAP7_75t_R FILLER_5_910 ();
 DECAPx10_ASAP7_75t_R FILLER_5_926 ();
 DECAPx10_ASAP7_75t_R FILLER_5_948 ();
 DECAPx10_ASAP7_75t_R FILLER_5_970 ();
 DECAPx10_ASAP7_75t_R FILLER_5_992 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1388 ();
 FILLER_ASAP7_75t_R FILLER_5_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx2_ASAP7_75t_R FILLER_6_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_52 ();
 DECAPx10_ASAP7_75t_R FILLER_6_79 ();
 DECAPx10_ASAP7_75t_R FILLER_6_101 ();
 DECAPx10_ASAP7_75t_R FILLER_6_123 ();
 DECAPx10_ASAP7_75t_R FILLER_6_145 ();
 DECAPx10_ASAP7_75t_R FILLER_6_167 ();
 DECAPx10_ASAP7_75t_R FILLER_6_189 ();
 DECAPx10_ASAP7_75t_R FILLER_6_211 ();
 DECAPx10_ASAP7_75t_R FILLER_6_233 ();
 DECAPx10_ASAP7_75t_R FILLER_6_255 ();
 DECAPx10_ASAP7_75t_R FILLER_6_277 ();
 DECAPx10_ASAP7_75t_R FILLER_6_299 ();
 DECAPx10_ASAP7_75t_R FILLER_6_321 ();
 DECAPx10_ASAP7_75t_R FILLER_6_343 ();
 DECAPx10_ASAP7_75t_R FILLER_6_365 ();
 DECAPx10_ASAP7_75t_R FILLER_6_387 ();
 DECAPx10_ASAP7_75t_R FILLER_6_409 ();
 DECAPx10_ASAP7_75t_R FILLER_6_431 ();
 DECAPx2_ASAP7_75t_R FILLER_6_453 ();
 FILLER_ASAP7_75t_R FILLER_6_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_461 ();
 DECAPx10_ASAP7_75t_R FILLER_6_464 ();
 DECAPx10_ASAP7_75t_R FILLER_6_486 ();
 DECAPx10_ASAP7_75t_R FILLER_6_508 ();
 DECAPx10_ASAP7_75t_R FILLER_6_530 ();
 DECAPx10_ASAP7_75t_R FILLER_6_552 ();
 DECAPx10_ASAP7_75t_R FILLER_6_574 ();
 DECAPx10_ASAP7_75t_R FILLER_6_596 ();
 DECAPx10_ASAP7_75t_R FILLER_6_618 ();
 DECAPx10_ASAP7_75t_R FILLER_6_640 ();
 DECAPx10_ASAP7_75t_R FILLER_6_662 ();
 DECAPx10_ASAP7_75t_R FILLER_6_684 ();
 DECAPx10_ASAP7_75t_R FILLER_6_706 ();
 DECAPx10_ASAP7_75t_R FILLER_6_728 ();
 DECAPx10_ASAP7_75t_R FILLER_6_750 ();
 DECAPx10_ASAP7_75t_R FILLER_6_772 ();
 DECAPx10_ASAP7_75t_R FILLER_6_794 ();
 DECAPx10_ASAP7_75t_R FILLER_6_816 ();
 DECAPx10_ASAP7_75t_R FILLER_6_838 ();
 DECAPx10_ASAP7_75t_R FILLER_6_860 ();
 DECAPx10_ASAP7_75t_R FILLER_6_882 ();
 DECAPx10_ASAP7_75t_R FILLER_6_904 ();
 DECAPx10_ASAP7_75t_R FILLER_6_926 ();
 DECAPx10_ASAP7_75t_R FILLER_6_948 ();
 DECAPx10_ASAP7_75t_R FILLER_6_970 ();
 DECAPx10_ASAP7_75t_R FILLER_6_992 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_6_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_6_1388 ();
 FILLER_ASAP7_75t_R FILLER_6_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx6_ASAP7_75t_R FILLER_7_46 ();
 FILLER_ASAP7_75t_R FILLER_7_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_62 ();
 DECAPx10_ASAP7_75t_R FILLER_7_74 ();
 DECAPx10_ASAP7_75t_R FILLER_7_96 ();
 DECAPx10_ASAP7_75t_R FILLER_7_118 ();
 DECAPx10_ASAP7_75t_R FILLER_7_140 ();
 DECAPx10_ASAP7_75t_R FILLER_7_162 ();
 DECAPx10_ASAP7_75t_R FILLER_7_184 ();
 DECAPx10_ASAP7_75t_R FILLER_7_206 ();
 DECAPx10_ASAP7_75t_R FILLER_7_228 ();
 DECAPx10_ASAP7_75t_R FILLER_7_250 ();
 DECAPx10_ASAP7_75t_R FILLER_7_272 ();
 DECAPx10_ASAP7_75t_R FILLER_7_294 ();
 DECAPx10_ASAP7_75t_R FILLER_7_316 ();
 DECAPx10_ASAP7_75t_R FILLER_7_338 ();
 DECAPx10_ASAP7_75t_R FILLER_7_360 ();
 DECAPx10_ASAP7_75t_R FILLER_7_382 ();
 DECAPx10_ASAP7_75t_R FILLER_7_404 ();
 DECAPx10_ASAP7_75t_R FILLER_7_426 ();
 DECAPx10_ASAP7_75t_R FILLER_7_448 ();
 DECAPx10_ASAP7_75t_R FILLER_7_470 ();
 DECAPx10_ASAP7_75t_R FILLER_7_492 ();
 DECAPx10_ASAP7_75t_R FILLER_7_514 ();
 DECAPx10_ASAP7_75t_R FILLER_7_536 ();
 DECAPx10_ASAP7_75t_R FILLER_7_558 ();
 DECAPx10_ASAP7_75t_R FILLER_7_580 ();
 DECAPx10_ASAP7_75t_R FILLER_7_602 ();
 DECAPx10_ASAP7_75t_R FILLER_7_624 ();
 DECAPx10_ASAP7_75t_R FILLER_7_646 ();
 DECAPx10_ASAP7_75t_R FILLER_7_668 ();
 DECAPx10_ASAP7_75t_R FILLER_7_690 ();
 DECAPx10_ASAP7_75t_R FILLER_7_712 ();
 DECAPx10_ASAP7_75t_R FILLER_7_734 ();
 DECAPx10_ASAP7_75t_R FILLER_7_756 ();
 DECAPx10_ASAP7_75t_R FILLER_7_778 ();
 DECAPx10_ASAP7_75t_R FILLER_7_800 ();
 DECAPx10_ASAP7_75t_R FILLER_7_822 ();
 DECAPx10_ASAP7_75t_R FILLER_7_844 ();
 DECAPx10_ASAP7_75t_R FILLER_7_866 ();
 DECAPx10_ASAP7_75t_R FILLER_7_888 ();
 DECAPx6_ASAP7_75t_R FILLER_7_910 ();
 DECAPx10_ASAP7_75t_R FILLER_7_926 ();
 DECAPx10_ASAP7_75t_R FILLER_7_948 ();
 DECAPx10_ASAP7_75t_R FILLER_7_970 ();
 DECAPx10_ASAP7_75t_R FILLER_7_992 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_7_1388 ();
 FILLER_ASAP7_75t_R FILLER_7_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_8_222 ();
 DECAPx10_ASAP7_75t_R FILLER_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_8_266 ();
 DECAPx10_ASAP7_75t_R FILLER_8_288 ();
 DECAPx10_ASAP7_75t_R FILLER_8_310 ();
 DECAPx10_ASAP7_75t_R FILLER_8_332 ();
 DECAPx10_ASAP7_75t_R FILLER_8_354 ();
 DECAPx10_ASAP7_75t_R FILLER_8_376 ();
 DECAPx10_ASAP7_75t_R FILLER_8_398 ();
 DECAPx10_ASAP7_75t_R FILLER_8_420 ();
 DECAPx6_ASAP7_75t_R FILLER_8_442 ();
 DECAPx2_ASAP7_75t_R FILLER_8_456 ();
 DECAPx10_ASAP7_75t_R FILLER_8_464 ();
 DECAPx10_ASAP7_75t_R FILLER_8_486 ();
 DECAPx10_ASAP7_75t_R FILLER_8_508 ();
 DECAPx10_ASAP7_75t_R FILLER_8_530 ();
 DECAPx10_ASAP7_75t_R FILLER_8_552 ();
 DECAPx10_ASAP7_75t_R FILLER_8_574 ();
 DECAPx10_ASAP7_75t_R FILLER_8_596 ();
 DECAPx10_ASAP7_75t_R FILLER_8_618 ();
 DECAPx10_ASAP7_75t_R FILLER_8_640 ();
 DECAPx10_ASAP7_75t_R FILLER_8_662 ();
 DECAPx10_ASAP7_75t_R FILLER_8_684 ();
 DECAPx10_ASAP7_75t_R FILLER_8_706 ();
 DECAPx10_ASAP7_75t_R FILLER_8_728 ();
 DECAPx10_ASAP7_75t_R FILLER_8_750 ();
 DECAPx10_ASAP7_75t_R FILLER_8_772 ();
 DECAPx10_ASAP7_75t_R FILLER_8_794 ();
 DECAPx10_ASAP7_75t_R FILLER_8_816 ();
 DECAPx10_ASAP7_75t_R FILLER_8_838 ();
 DECAPx10_ASAP7_75t_R FILLER_8_860 ();
 DECAPx10_ASAP7_75t_R FILLER_8_882 ();
 DECAPx10_ASAP7_75t_R FILLER_8_904 ();
 DECAPx10_ASAP7_75t_R FILLER_8_926 ();
 DECAPx10_ASAP7_75t_R FILLER_8_948 ();
 DECAPx10_ASAP7_75t_R FILLER_8_970 ();
 DECAPx10_ASAP7_75t_R FILLER_8_992 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1388 ();
 FILLER_ASAP7_75t_R FILLER_8_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_9_222 ();
 DECAPx10_ASAP7_75t_R FILLER_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_9_266 ();
 DECAPx10_ASAP7_75t_R FILLER_9_288 ();
 DECAPx10_ASAP7_75t_R FILLER_9_310 ();
 DECAPx10_ASAP7_75t_R FILLER_9_332 ();
 DECAPx10_ASAP7_75t_R FILLER_9_354 ();
 DECAPx10_ASAP7_75t_R FILLER_9_376 ();
 DECAPx10_ASAP7_75t_R FILLER_9_398 ();
 DECAPx10_ASAP7_75t_R FILLER_9_420 ();
 DECAPx10_ASAP7_75t_R FILLER_9_442 ();
 DECAPx10_ASAP7_75t_R FILLER_9_464 ();
 DECAPx10_ASAP7_75t_R FILLER_9_486 ();
 DECAPx10_ASAP7_75t_R FILLER_9_508 ();
 DECAPx10_ASAP7_75t_R FILLER_9_530 ();
 DECAPx10_ASAP7_75t_R FILLER_9_552 ();
 DECAPx10_ASAP7_75t_R FILLER_9_574 ();
 DECAPx10_ASAP7_75t_R FILLER_9_596 ();
 DECAPx10_ASAP7_75t_R FILLER_9_618 ();
 DECAPx10_ASAP7_75t_R FILLER_9_640 ();
 DECAPx10_ASAP7_75t_R FILLER_9_662 ();
 DECAPx10_ASAP7_75t_R FILLER_9_684 ();
 DECAPx10_ASAP7_75t_R FILLER_9_706 ();
 DECAPx10_ASAP7_75t_R FILLER_9_728 ();
 DECAPx10_ASAP7_75t_R FILLER_9_750 ();
 DECAPx10_ASAP7_75t_R FILLER_9_772 ();
 DECAPx10_ASAP7_75t_R FILLER_9_794 ();
 DECAPx10_ASAP7_75t_R FILLER_9_816 ();
 DECAPx10_ASAP7_75t_R FILLER_9_838 ();
 DECAPx10_ASAP7_75t_R FILLER_9_860 ();
 DECAPx10_ASAP7_75t_R FILLER_9_882 ();
 DECAPx6_ASAP7_75t_R FILLER_9_904 ();
 DECAPx2_ASAP7_75t_R FILLER_9_918 ();
 DECAPx10_ASAP7_75t_R FILLER_9_926 ();
 DECAPx10_ASAP7_75t_R FILLER_9_948 ();
 DECAPx10_ASAP7_75t_R FILLER_9_970 ();
 DECAPx10_ASAP7_75t_R FILLER_9_992 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1388 ();
 FILLER_ASAP7_75t_R FILLER_9_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_10_200 ();
 DECAPx10_ASAP7_75t_R FILLER_10_222 ();
 DECAPx10_ASAP7_75t_R FILLER_10_244 ();
 DECAPx10_ASAP7_75t_R FILLER_10_266 ();
 DECAPx10_ASAP7_75t_R FILLER_10_288 ();
 DECAPx10_ASAP7_75t_R FILLER_10_310 ();
 DECAPx10_ASAP7_75t_R FILLER_10_332 ();
 DECAPx10_ASAP7_75t_R FILLER_10_354 ();
 DECAPx10_ASAP7_75t_R FILLER_10_376 ();
 DECAPx10_ASAP7_75t_R FILLER_10_398 ();
 DECAPx10_ASAP7_75t_R FILLER_10_420 ();
 DECAPx6_ASAP7_75t_R FILLER_10_442 ();
 DECAPx2_ASAP7_75t_R FILLER_10_456 ();
 DECAPx10_ASAP7_75t_R FILLER_10_464 ();
 DECAPx10_ASAP7_75t_R FILLER_10_486 ();
 DECAPx10_ASAP7_75t_R FILLER_10_508 ();
 DECAPx10_ASAP7_75t_R FILLER_10_530 ();
 DECAPx10_ASAP7_75t_R FILLER_10_552 ();
 DECAPx10_ASAP7_75t_R FILLER_10_574 ();
 DECAPx10_ASAP7_75t_R FILLER_10_596 ();
 DECAPx10_ASAP7_75t_R FILLER_10_618 ();
 DECAPx10_ASAP7_75t_R FILLER_10_640 ();
 DECAPx10_ASAP7_75t_R FILLER_10_662 ();
 DECAPx10_ASAP7_75t_R FILLER_10_684 ();
 DECAPx10_ASAP7_75t_R FILLER_10_706 ();
 DECAPx10_ASAP7_75t_R FILLER_10_728 ();
 DECAPx10_ASAP7_75t_R FILLER_10_750 ();
 DECAPx10_ASAP7_75t_R FILLER_10_772 ();
 DECAPx10_ASAP7_75t_R FILLER_10_794 ();
 DECAPx10_ASAP7_75t_R FILLER_10_816 ();
 DECAPx10_ASAP7_75t_R FILLER_10_838 ();
 DECAPx10_ASAP7_75t_R FILLER_10_860 ();
 DECAPx10_ASAP7_75t_R FILLER_10_882 ();
 DECAPx10_ASAP7_75t_R FILLER_10_904 ();
 DECAPx10_ASAP7_75t_R FILLER_10_926 ();
 DECAPx10_ASAP7_75t_R FILLER_10_948 ();
 DECAPx10_ASAP7_75t_R FILLER_10_970 ();
 DECAPx10_ASAP7_75t_R FILLER_10_992 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1388 ();
 FILLER_ASAP7_75t_R FILLER_10_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_11_112 ();
 DECAPx10_ASAP7_75t_R FILLER_11_134 ();
 DECAPx10_ASAP7_75t_R FILLER_11_156 ();
 DECAPx10_ASAP7_75t_R FILLER_11_178 ();
 DECAPx10_ASAP7_75t_R FILLER_11_200 ();
 DECAPx10_ASAP7_75t_R FILLER_11_222 ();
 DECAPx10_ASAP7_75t_R FILLER_11_244 ();
 DECAPx10_ASAP7_75t_R FILLER_11_266 ();
 DECAPx10_ASAP7_75t_R FILLER_11_288 ();
 DECAPx10_ASAP7_75t_R FILLER_11_310 ();
 DECAPx10_ASAP7_75t_R FILLER_11_332 ();
 DECAPx10_ASAP7_75t_R FILLER_11_354 ();
 DECAPx10_ASAP7_75t_R FILLER_11_376 ();
 DECAPx10_ASAP7_75t_R FILLER_11_398 ();
 DECAPx10_ASAP7_75t_R FILLER_11_420 ();
 DECAPx10_ASAP7_75t_R FILLER_11_442 ();
 DECAPx10_ASAP7_75t_R FILLER_11_464 ();
 DECAPx10_ASAP7_75t_R FILLER_11_486 ();
 DECAPx10_ASAP7_75t_R FILLER_11_508 ();
 DECAPx10_ASAP7_75t_R FILLER_11_530 ();
 DECAPx10_ASAP7_75t_R FILLER_11_552 ();
 DECAPx10_ASAP7_75t_R FILLER_11_574 ();
 DECAPx10_ASAP7_75t_R FILLER_11_596 ();
 DECAPx10_ASAP7_75t_R FILLER_11_618 ();
 DECAPx10_ASAP7_75t_R FILLER_11_640 ();
 DECAPx10_ASAP7_75t_R FILLER_11_662 ();
 DECAPx10_ASAP7_75t_R FILLER_11_684 ();
 DECAPx10_ASAP7_75t_R FILLER_11_706 ();
 DECAPx10_ASAP7_75t_R FILLER_11_728 ();
 DECAPx10_ASAP7_75t_R FILLER_11_750 ();
 DECAPx10_ASAP7_75t_R FILLER_11_772 ();
 DECAPx10_ASAP7_75t_R FILLER_11_794 ();
 DECAPx10_ASAP7_75t_R FILLER_11_816 ();
 DECAPx10_ASAP7_75t_R FILLER_11_838 ();
 DECAPx10_ASAP7_75t_R FILLER_11_860 ();
 DECAPx10_ASAP7_75t_R FILLER_11_882 ();
 DECAPx6_ASAP7_75t_R FILLER_11_904 ();
 DECAPx2_ASAP7_75t_R FILLER_11_918 ();
 DECAPx10_ASAP7_75t_R FILLER_11_926 ();
 DECAPx10_ASAP7_75t_R FILLER_11_948 ();
 DECAPx10_ASAP7_75t_R FILLER_11_970 ();
 DECAPx10_ASAP7_75t_R FILLER_11_992 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_11_1388 ();
 FILLER_ASAP7_75t_R FILLER_11_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_12_112 ();
 DECAPx10_ASAP7_75t_R FILLER_12_134 ();
 DECAPx10_ASAP7_75t_R FILLER_12_156 ();
 DECAPx10_ASAP7_75t_R FILLER_12_178 ();
 DECAPx10_ASAP7_75t_R FILLER_12_200 ();
 DECAPx10_ASAP7_75t_R FILLER_12_222 ();
 DECAPx10_ASAP7_75t_R FILLER_12_244 ();
 DECAPx10_ASAP7_75t_R FILLER_12_266 ();
 DECAPx10_ASAP7_75t_R FILLER_12_288 ();
 DECAPx10_ASAP7_75t_R FILLER_12_310 ();
 DECAPx10_ASAP7_75t_R FILLER_12_332 ();
 DECAPx10_ASAP7_75t_R FILLER_12_354 ();
 DECAPx10_ASAP7_75t_R FILLER_12_376 ();
 DECAPx10_ASAP7_75t_R FILLER_12_398 ();
 DECAPx10_ASAP7_75t_R FILLER_12_420 ();
 DECAPx6_ASAP7_75t_R FILLER_12_442 ();
 DECAPx2_ASAP7_75t_R FILLER_12_456 ();
 DECAPx10_ASAP7_75t_R FILLER_12_464 ();
 DECAPx10_ASAP7_75t_R FILLER_12_486 ();
 DECAPx10_ASAP7_75t_R FILLER_12_508 ();
 DECAPx10_ASAP7_75t_R FILLER_12_530 ();
 DECAPx10_ASAP7_75t_R FILLER_12_552 ();
 DECAPx10_ASAP7_75t_R FILLER_12_574 ();
 DECAPx10_ASAP7_75t_R FILLER_12_596 ();
 DECAPx10_ASAP7_75t_R FILLER_12_618 ();
 DECAPx10_ASAP7_75t_R FILLER_12_640 ();
 DECAPx10_ASAP7_75t_R FILLER_12_662 ();
 DECAPx10_ASAP7_75t_R FILLER_12_684 ();
 DECAPx10_ASAP7_75t_R FILLER_12_706 ();
 DECAPx10_ASAP7_75t_R FILLER_12_728 ();
 DECAPx10_ASAP7_75t_R FILLER_12_750 ();
 DECAPx10_ASAP7_75t_R FILLER_12_772 ();
 DECAPx10_ASAP7_75t_R FILLER_12_794 ();
 DECAPx10_ASAP7_75t_R FILLER_12_816 ();
 DECAPx6_ASAP7_75t_R FILLER_12_838 ();
 FILLER_ASAP7_75t_R FILLER_12_852 ();
 DECAPx10_ASAP7_75t_R FILLER_12_857 ();
 DECAPx10_ASAP7_75t_R FILLER_12_879 ();
 DECAPx10_ASAP7_75t_R FILLER_12_901 ();
 DECAPx10_ASAP7_75t_R FILLER_12_923 ();
 DECAPx10_ASAP7_75t_R FILLER_12_945 ();
 DECAPx10_ASAP7_75t_R FILLER_12_967 ();
 DECAPx10_ASAP7_75t_R FILLER_12_989 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_12_1388 ();
 FILLER_ASAP7_75t_R FILLER_12_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_13_112 ();
 DECAPx10_ASAP7_75t_R FILLER_13_134 ();
 DECAPx10_ASAP7_75t_R FILLER_13_156 ();
 DECAPx10_ASAP7_75t_R FILLER_13_178 ();
 DECAPx10_ASAP7_75t_R FILLER_13_200 ();
 DECAPx10_ASAP7_75t_R FILLER_13_222 ();
 DECAPx10_ASAP7_75t_R FILLER_13_244 ();
 DECAPx10_ASAP7_75t_R FILLER_13_266 ();
 DECAPx10_ASAP7_75t_R FILLER_13_288 ();
 DECAPx10_ASAP7_75t_R FILLER_13_310 ();
 DECAPx10_ASAP7_75t_R FILLER_13_332 ();
 DECAPx10_ASAP7_75t_R FILLER_13_354 ();
 DECAPx10_ASAP7_75t_R FILLER_13_376 ();
 DECAPx10_ASAP7_75t_R FILLER_13_398 ();
 DECAPx10_ASAP7_75t_R FILLER_13_420 ();
 DECAPx10_ASAP7_75t_R FILLER_13_442 ();
 DECAPx10_ASAP7_75t_R FILLER_13_464 ();
 DECAPx10_ASAP7_75t_R FILLER_13_486 ();
 DECAPx10_ASAP7_75t_R FILLER_13_508 ();
 DECAPx10_ASAP7_75t_R FILLER_13_530 ();
 DECAPx10_ASAP7_75t_R FILLER_13_552 ();
 DECAPx10_ASAP7_75t_R FILLER_13_574 ();
 DECAPx10_ASAP7_75t_R FILLER_13_596 ();
 DECAPx10_ASAP7_75t_R FILLER_13_618 ();
 DECAPx10_ASAP7_75t_R FILLER_13_640 ();
 DECAPx10_ASAP7_75t_R FILLER_13_662 ();
 DECAPx10_ASAP7_75t_R FILLER_13_684 ();
 DECAPx10_ASAP7_75t_R FILLER_13_706 ();
 DECAPx2_ASAP7_75t_R FILLER_13_728 ();
 FILLER_ASAP7_75t_R FILLER_13_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_736 ();
 DECAPx10_ASAP7_75t_R FILLER_13_740 ();
 FILLER_ASAP7_75t_R FILLER_13_762 ();
 DECAPx1_ASAP7_75t_R FILLER_13_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_786 ();
 FILLER_ASAP7_75t_R FILLER_13_797 ();
 DECAPx6_ASAP7_75t_R FILLER_13_819 ();
 FILLER_ASAP7_75t_R FILLER_13_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_835 ();
 FILLER_ASAP7_75t_R FILLER_13_842 ();
 FILLER_ASAP7_75t_R FILLER_13_850 ();
 DECAPx1_ASAP7_75t_R FILLER_13_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_880 ();
 FILLER_ASAP7_75t_R FILLER_13_887 ();
 DECAPx10_ASAP7_75t_R FILLER_13_895 ();
 DECAPx2_ASAP7_75t_R FILLER_13_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_923 ();
 DECAPx10_ASAP7_75t_R FILLER_13_926 ();
 DECAPx10_ASAP7_75t_R FILLER_13_948 ();
 DECAPx10_ASAP7_75t_R FILLER_13_970 ();
 DECAPx10_ASAP7_75t_R FILLER_13_992 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_13_1388 ();
 FILLER_ASAP7_75t_R FILLER_13_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_14_68 ();
 DECAPx10_ASAP7_75t_R FILLER_14_90 ();
 DECAPx10_ASAP7_75t_R FILLER_14_112 ();
 DECAPx10_ASAP7_75t_R FILLER_14_134 ();
 DECAPx10_ASAP7_75t_R FILLER_14_156 ();
 DECAPx10_ASAP7_75t_R FILLER_14_178 ();
 DECAPx10_ASAP7_75t_R FILLER_14_200 ();
 DECAPx10_ASAP7_75t_R FILLER_14_222 ();
 DECAPx10_ASAP7_75t_R FILLER_14_244 ();
 DECAPx10_ASAP7_75t_R FILLER_14_266 ();
 DECAPx10_ASAP7_75t_R FILLER_14_288 ();
 DECAPx10_ASAP7_75t_R FILLER_14_310 ();
 DECAPx10_ASAP7_75t_R FILLER_14_332 ();
 DECAPx10_ASAP7_75t_R FILLER_14_354 ();
 DECAPx10_ASAP7_75t_R FILLER_14_376 ();
 DECAPx10_ASAP7_75t_R FILLER_14_398 ();
 DECAPx10_ASAP7_75t_R FILLER_14_420 ();
 DECAPx6_ASAP7_75t_R FILLER_14_442 ();
 DECAPx2_ASAP7_75t_R FILLER_14_456 ();
 DECAPx10_ASAP7_75t_R FILLER_14_464 ();
 DECAPx10_ASAP7_75t_R FILLER_14_486 ();
 DECAPx10_ASAP7_75t_R FILLER_14_508 ();
 DECAPx10_ASAP7_75t_R FILLER_14_530 ();
 DECAPx10_ASAP7_75t_R FILLER_14_552 ();
 DECAPx10_ASAP7_75t_R FILLER_14_574 ();
 DECAPx10_ASAP7_75t_R FILLER_14_596 ();
 DECAPx10_ASAP7_75t_R FILLER_14_618 ();
 DECAPx10_ASAP7_75t_R FILLER_14_640 ();
 DECAPx10_ASAP7_75t_R FILLER_14_662 ();
 DECAPx4_ASAP7_75t_R FILLER_14_684 ();
 FILLER_ASAP7_75t_R FILLER_14_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_696 ();
 DECAPx10_ASAP7_75t_R FILLER_14_707 ();
 DECAPx1_ASAP7_75t_R FILLER_14_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_733 ();
 FILLER_ASAP7_75t_R FILLER_14_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_748 ();
 FILLER_ASAP7_75t_R FILLER_14_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_754 ();
 FILLER_ASAP7_75t_R FILLER_14_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_797 ();
 DECAPx1_ASAP7_75t_R FILLER_14_824 ();
 FILLER_ASAP7_75t_R FILLER_14_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_876 ();
 FILLER_ASAP7_75t_R FILLER_14_891 ();
 DECAPx2_ASAP7_75t_R FILLER_14_913 ();
 FILLER_ASAP7_75t_R FILLER_14_925 ();
 DECAPx10_ASAP7_75t_R FILLER_14_930 ();
 DECAPx10_ASAP7_75t_R FILLER_14_952 ();
 DECAPx10_ASAP7_75t_R FILLER_14_974 ();
 DECAPx10_ASAP7_75t_R FILLER_14_996 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_14_1370 ();
 FILLER_ASAP7_75t_R FILLER_14_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_14_1388 ();
 FILLER_ASAP7_75t_R FILLER_14_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_15_68 ();
 DECAPx10_ASAP7_75t_R FILLER_15_90 ();
 DECAPx10_ASAP7_75t_R FILLER_15_112 ();
 DECAPx10_ASAP7_75t_R FILLER_15_134 ();
 DECAPx10_ASAP7_75t_R FILLER_15_156 ();
 DECAPx10_ASAP7_75t_R FILLER_15_178 ();
 DECAPx10_ASAP7_75t_R FILLER_15_200 ();
 DECAPx10_ASAP7_75t_R FILLER_15_222 ();
 DECAPx10_ASAP7_75t_R FILLER_15_244 ();
 DECAPx10_ASAP7_75t_R FILLER_15_266 ();
 DECAPx10_ASAP7_75t_R FILLER_15_288 ();
 DECAPx10_ASAP7_75t_R FILLER_15_310 ();
 DECAPx10_ASAP7_75t_R FILLER_15_332 ();
 DECAPx10_ASAP7_75t_R FILLER_15_354 ();
 DECAPx10_ASAP7_75t_R FILLER_15_376 ();
 DECAPx10_ASAP7_75t_R FILLER_15_398 ();
 DECAPx10_ASAP7_75t_R FILLER_15_420 ();
 DECAPx10_ASAP7_75t_R FILLER_15_442 ();
 DECAPx10_ASAP7_75t_R FILLER_15_464 ();
 DECAPx10_ASAP7_75t_R FILLER_15_486 ();
 DECAPx10_ASAP7_75t_R FILLER_15_508 ();
 DECAPx10_ASAP7_75t_R FILLER_15_530 ();
 DECAPx10_ASAP7_75t_R FILLER_15_552 ();
 DECAPx10_ASAP7_75t_R FILLER_15_574 ();
 DECAPx10_ASAP7_75t_R FILLER_15_596 ();
 DECAPx10_ASAP7_75t_R FILLER_15_618 ();
 DECAPx10_ASAP7_75t_R FILLER_15_640 ();
 DECAPx10_ASAP7_75t_R FILLER_15_662 ();
 DECAPx6_ASAP7_75t_R FILLER_15_684 ();
 FILLER_ASAP7_75t_R FILLER_15_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_700 ();
 DECAPx6_ASAP7_75t_R FILLER_15_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_753 ();
 FILLER_ASAP7_75t_R FILLER_15_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_766 ();
 DECAPx1_ASAP7_75t_R FILLER_15_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_794 ();
 DECAPx1_ASAP7_75t_R FILLER_15_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_811 ();
 DECAPx1_ASAP7_75t_R FILLER_15_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_836 ();
 DECAPx2_ASAP7_75t_R FILLER_15_843 ();
 DECAPx2_ASAP7_75t_R FILLER_15_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_858 ();
 DECAPx2_ASAP7_75t_R FILLER_15_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_880 ();
 FILLER_ASAP7_75t_R FILLER_15_887 ();
 DECAPx1_ASAP7_75t_R FILLER_15_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_902 ();
 DECAPx1_ASAP7_75t_R FILLER_15_909 ();
 DECAPx1_ASAP7_75t_R FILLER_15_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_923 ();
 DECAPx10_ASAP7_75t_R FILLER_15_940 ();
 DECAPx10_ASAP7_75t_R FILLER_15_962 ();
 DECAPx10_ASAP7_75t_R FILLER_15_984 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1358 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1380 ();
 FILLER_ASAP7_75t_R FILLER_15_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_16_68 ();
 DECAPx10_ASAP7_75t_R FILLER_16_90 ();
 DECAPx10_ASAP7_75t_R FILLER_16_112 ();
 DECAPx10_ASAP7_75t_R FILLER_16_134 ();
 DECAPx10_ASAP7_75t_R FILLER_16_156 ();
 DECAPx10_ASAP7_75t_R FILLER_16_178 ();
 DECAPx10_ASAP7_75t_R FILLER_16_200 ();
 DECAPx10_ASAP7_75t_R FILLER_16_222 ();
 DECAPx10_ASAP7_75t_R FILLER_16_244 ();
 DECAPx10_ASAP7_75t_R FILLER_16_266 ();
 DECAPx10_ASAP7_75t_R FILLER_16_288 ();
 DECAPx10_ASAP7_75t_R FILLER_16_310 ();
 DECAPx10_ASAP7_75t_R FILLER_16_332 ();
 DECAPx10_ASAP7_75t_R FILLER_16_354 ();
 DECAPx10_ASAP7_75t_R FILLER_16_376 ();
 DECAPx10_ASAP7_75t_R FILLER_16_398 ();
 DECAPx10_ASAP7_75t_R FILLER_16_420 ();
 DECAPx6_ASAP7_75t_R FILLER_16_442 ();
 DECAPx2_ASAP7_75t_R FILLER_16_456 ();
 DECAPx10_ASAP7_75t_R FILLER_16_464 ();
 DECAPx10_ASAP7_75t_R FILLER_16_486 ();
 DECAPx10_ASAP7_75t_R FILLER_16_508 ();
 DECAPx10_ASAP7_75t_R FILLER_16_530 ();
 DECAPx10_ASAP7_75t_R FILLER_16_552 ();
 DECAPx10_ASAP7_75t_R FILLER_16_574 ();
 DECAPx10_ASAP7_75t_R FILLER_16_596 ();
 DECAPx10_ASAP7_75t_R FILLER_16_618 ();
 DECAPx10_ASAP7_75t_R FILLER_16_640 ();
 DECAPx10_ASAP7_75t_R FILLER_16_662 ();
 DECAPx6_ASAP7_75t_R FILLER_16_684 ();
 DECAPx1_ASAP7_75t_R FILLER_16_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_702 ();
 DECAPx1_ASAP7_75t_R FILLER_16_713 ();
 FILLER_ASAP7_75t_R FILLER_16_738 ();
 DECAPx2_ASAP7_75t_R FILLER_16_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_758 ();
 DECAPx6_ASAP7_75t_R FILLER_16_769 ();
 FILLER_ASAP7_75t_R FILLER_16_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_785 ();
 DECAPx10_ASAP7_75t_R FILLER_16_789 ();
 DECAPx2_ASAP7_75t_R FILLER_16_811 ();
 DECAPx2_ASAP7_75t_R FILLER_16_840 ();
 DECAPx4_ASAP7_75t_R FILLER_16_849 ();
 FILLER_ASAP7_75t_R FILLER_16_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_861 ();
 DECAPx4_ASAP7_75t_R FILLER_16_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_886 ();
 DECAPx2_ASAP7_75t_R FILLER_16_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_896 ();
 DECAPx1_ASAP7_75t_R FILLER_16_914 ();
 FILLER_ASAP7_75t_R FILLER_16_924 ();
 DECAPx10_ASAP7_75t_R FILLER_16_946 ();
 DECAPx10_ASAP7_75t_R FILLER_16_968 ();
 DECAPx10_ASAP7_75t_R FILLER_16_990 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_16_1388 ();
 FILLER_ASAP7_75t_R FILLER_16_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_17_68 ();
 DECAPx10_ASAP7_75t_R FILLER_17_90 ();
 DECAPx10_ASAP7_75t_R FILLER_17_112 ();
 DECAPx10_ASAP7_75t_R FILLER_17_134 ();
 DECAPx10_ASAP7_75t_R FILLER_17_156 ();
 DECAPx10_ASAP7_75t_R FILLER_17_178 ();
 DECAPx10_ASAP7_75t_R FILLER_17_200 ();
 DECAPx10_ASAP7_75t_R FILLER_17_222 ();
 DECAPx10_ASAP7_75t_R FILLER_17_244 ();
 DECAPx10_ASAP7_75t_R FILLER_17_266 ();
 DECAPx10_ASAP7_75t_R FILLER_17_288 ();
 DECAPx10_ASAP7_75t_R FILLER_17_310 ();
 DECAPx10_ASAP7_75t_R FILLER_17_332 ();
 DECAPx10_ASAP7_75t_R FILLER_17_354 ();
 DECAPx10_ASAP7_75t_R FILLER_17_376 ();
 DECAPx10_ASAP7_75t_R FILLER_17_398 ();
 DECAPx10_ASAP7_75t_R FILLER_17_420 ();
 DECAPx10_ASAP7_75t_R FILLER_17_442 ();
 DECAPx10_ASAP7_75t_R FILLER_17_464 ();
 DECAPx10_ASAP7_75t_R FILLER_17_486 ();
 DECAPx10_ASAP7_75t_R FILLER_17_508 ();
 DECAPx10_ASAP7_75t_R FILLER_17_530 ();
 DECAPx10_ASAP7_75t_R FILLER_17_552 ();
 DECAPx10_ASAP7_75t_R FILLER_17_574 ();
 DECAPx10_ASAP7_75t_R FILLER_17_596 ();
 DECAPx10_ASAP7_75t_R FILLER_17_618 ();
 DECAPx10_ASAP7_75t_R FILLER_17_640 ();
 DECAPx10_ASAP7_75t_R FILLER_17_662 ();
 DECAPx2_ASAP7_75t_R FILLER_17_684 ();
 FILLER_ASAP7_75t_R FILLER_17_690 ();
 DECAPx6_ASAP7_75t_R FILLER_17_702 ();
 DECAPx10_ASAP7_75t_R FILLER_17_728 ();
 DECAPx10_ASAP7_75t_R FILLER_17_750 ();
 DECAPx4_ASAP7_75t_R FILLER_17_772 ();
 FILLER_ASAP7_75t_R FILLER_17_782 ();
 DECAPx1_ASAP7_75t_R FILLER_17_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_800 ();
 DECAPx2_ASAP7_75t_R FILLER_17_820 ();
 DECAPx2_ASAP7_75t_R FILLER_17_829 ();
 DECAPx1_ASAP7_75t_R FILLER_17_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_842 ();
 DECAPx4_ASAP7_75t_R FILLER_17_860 ();
 DECAPx1_ASAP7_75t_R FILLER_17_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_877 ();
 DECAPx10_ASAP7_75t_R FILLER_17_881 ();
 FILLER_ASAP7_75t_R FILLER_17_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_908 ();
 DECAPx4_ASAP7_75t_R FILLER_17_912 ();
 FILLER_ASAP7_75t_R FILLER_17_922 ();
 DECAPx10_ASAP7_75t_R FILLER_17_932 ();
 DECAPx2_ASAP7_75t_R FILLER_17_954 ();
 FILLER_ASAP7_75t_R FILLER_17_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_962 ();
 DECAPx10_ASAP7_75t_R FILLER_17_968 ();
 DECAPx10_ASAP7_75t_R FILLER_17_990 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1386 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_18_90 ();
 DECAPx10_ASAP7_75t_R FILLER_18_112 ();
 DECAPx10_ASAP7_75t_R FILLER_18_134 ();
 DECAPx10_ASAP7_75t_R FILLER_18_156 ();
 DECAPx10_ASAP7_75t_R FILLER_18_178 ();
 DECAPx10_ASAP7_75t_R FILLER_18_200 ();
 DECAPx10_ASAP7_75t_R FILLER_18_222 ();
 DECAPx10_ASAP7_75t_R FILLER_18_244 ();
 DECAPx10_ASAP7_75t_R FILLER_18_266 ();
 DECAPx10_ASAP7_75t_R FILLER_18_288 ();
 DECAPx10_ASAP7_75t_R FILLER_18_310 ();
 DECAPx10_ASAP7_75t_R FILLER_18_332 ();
 DECAPx10_ASAP7_75t_R FILLER_18_354 ();
 DECAPx10_ASAP7_75t_R FILLER_18_376 ();
 DECAPx10_ASAP7_75t_R FILLER_18_398 ();
 DECAPx10_ASAP7_75t_R FILLER_18_420 ();
 DECAPx6_ASAP7_75t_R FILLER_18_442 ();
 DECAPx2_ASAP7_75t_R FILLER_18_456 ();
 DECAPx10_ASAP7_75t_R FILLER_18_464 ();
 DECAPx10_ASAP7_75t_R FILLER_18_486 ();
 DECAPx10_ASAP7_75t_R FILLER_18_508 ();
 DECAPx10_ASAP7_75t_R FILLER_18_530 ();
 DECAPx10_ASAP7_75t_R FILLER_18_552 ();
 DECAPx10_ASAP7_75t_R FILLER_18_574 ();
 DECAPx10_ASAP7_75t_R FILLER_18_596 ();
 DECAPx10_ASAP7_75t_R FILLER_18_618 ();
 DECAPx10_ASAP7_75t_R FILLER_18_640 ();
 DECAPx10_ASAP7_75t_R FILLER_18_662 ();
 DECAPx6_ASAP7_75t_R FILLER_18_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_698 ();
 DECAPx2_ASAP7_75t_R FILLER_18_709 ();
 DECAPx6_ASAP7_75t_R FILLER_18_732 ();
 FILLER_ASAP7_75t_R FILLER_18_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_748 ();
 FILLER_ASAP7_75t_R FILLER_18_773 ();
 DECAPx2_ASAP7_75t_R FILLER_18_795 ();
 FILLER_ASAP7_75t_R FILLER_18_801 ();
 DECAPx2_ASAP7_75t_R FILLER_18_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_857 ();
 DECAPx4_ASAP7_75t_R FILLER_18_867 ();
 FILLER_ASAP7_75t_R FILLER_18_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_879 ();
 DECAPx6_ASAP7_75t_R FILLER_18_894 ();
 DECAPx1_ASAP7_75t_R FILLER_18_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_964 ();
 DECAPx10_ASAP7_75t_R FILLER_18_977 ();
 DECAPx10_ASAP7_75t_R FILLER_18_999 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1351 ();
 DECAPx4_ASAP7_75t_R FILLER_18_1373 ();
 FILLER_ASAP7_75t_R FILLER_18_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1388 ();
 FILLER_ASAP7_75t_R FILLER_18_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_19_68 ();
 DECAPx10_ASAP7_75t_R FILLER_19_90 ();
 DECAPx10_ASAP7_75t_R FILLER_19_112 ();
 DECAPx10_ASAP7_75t_R FILLER_19_134 ();
 DECAPx10_ASAP7_75t_R FILLER_19_156 ();
 DECAPx10_ASAP7_75t_R FILLER_19_178 ();
 DECAPx10_ASAP7_75t_R FILLER_19_200 ();
 DECAPx10_ASAP7_75t_R FILLER_19_222 ();
 DECAPx10_ASAP7_75t_R FILLER_19_244 ();
 DECAPx10_ASAP7_75t_R FILLER_19_266 ();
 DECAPx10_ASAP7_75t_R FILLER_19_288 ();
 DECAPx10_ASAP7_75t_R FILLER_19_310 ();
 DECAPx10_ASAP7_75t_R FILLER_19_332 ();
 DECAPx10_ASAP7_75t_R FILLER_19_354 ();
 DECAPx10_ASAP7_75t_R FILLER_19_376 ();
 DECAPx10_ASAP7_75t_R FILLER_19_398 ();
 DECAPx10_ASAP7_75t_R FILLER_19_420 ();
 DECAPx10_ASAP7_75t_R FILLER_19_442 ();
 DECAPx10_ASAP7_75t_R FILLER_19_464 ();
 DECAPx10_ASAP7_75t_R FILLER_19_486 ();
 DECAPx10_ASAP7_75t_R FILLER_19_508 ();
 DECAPx10_ASAP7_75t_R FILLER_19_530 ();
 DECAPx10_ASAP7_75t_R FILLER_19_552 ();
 DECAPx10_ASAP7_75t_R FILLER_19_574 ();
 DECAPx10_ASAP7_75t_R FILLER_19_596 ();
 DECAPx10_ASAP7_75t_R FILLER_19_618 ();
 DECAPx10_ASAP7_75t_R FILLER_19_640 ();
 DECAPx10_ASAP7_75t_R FILLER_19_662 ();
 FILLER_ASAP7_75t_R FILLER_19_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_686 ();
 FILLER_ASAP7_75t_R FILLER_19_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_716 ();
 DECAPx4_ASAP7_75t_R FILLER_19_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_805 ();
 DECAPx2_ASAP7_75t_R FILLER_19_818 ();
 DECAPx2_ASAP7_75t_R FILLER_19_836 ();
 FILLER_ASAP7_75t_R FILLER_19_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_888 ();
 FILLER_ASAP7_75t_R FILLER_19_898 ();
 DECAPx1_ASAP7_75t_R FILLER_19_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_913 ();
 FILLER_ASAP7_75t_R FILLER_19_936 ();
 DECAPx10_ASAP7_75t_R FILLER_19_980 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1354 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1398 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_20_90 ();
 DECAPx10_ASAP7_75t_R FILLER_20_112 ();
 DECAPx10_ASAP7_75t_R FILLER_20_134 ();
 DECAPx10_ASAP7_75t_R FILLER_20_156 ();
 DECAPx10_ASAP7_75t_R FILLER_20_178 ();
 DECAPx10_ASAP7_75t_R FILLER_20_200 ();
 DECAPx10_ASAP7_75t_R FILLER_20_222 ();
 DECAPx10_ASAP7_75t_R FILLER_20_244 ();
 DECAPx10_ASAP7_75t_R FILLER_20_266 ();
 DECAPx10_ASAP7_75t_R FILLER_20_288 ();
 DECAPx10_ASAP7_75t_R FILLER_20_310 ();
 DECAPx10_ASAP7_75t_R FILLER_20_332 ();
 DECAPx10_ASAP7_75t_R FILLER_20_354 ();
 DECAPx10_ASAP7_75t_R FILLER_20_376 ();
 DECAPx10_ASAP7_75t_R FILLER_20_398 ();
 DECAPx10_ASAP7_75t_R FILLER_20_420 ();
 DECAPx6_ASAP7_75t_R FILLER_20_442 ();
 DECAPx2_ASAP7_75t_R FILLER_20_456 ();
 DECAPx10_ASAP7_75t_R FILLER_20_464 ();
 DECAPx10_ASAP7_75t_R FILLER_20_486 ();
 DECAPx10_ASAP7_75t_R FILLER_20_508 ();
 DECAPx10_ASAP7_75t_R FILLER_20_530 ();
 DECAPx10_ASAP7_75t_R FILLER_20_552 ();
 DECAPx10_ASAP7_75t_R FILLER_20_574 ();
 DECAPx10_ASAP7_75t_R FILLER_20_596 ();
 DECAPx10_ASAP7_75t_R FILLER_20_618 ();
 DECAPx10_ASAP7_75t_R FILLER_20_640 ();
 DECAPx1_ASAP7_75t_R FILLER_20_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_666 ();
 DECAPx6_ASAP7_75t_R FILLER_20_677 ();
 FILLER_ASAP7_75t_R FILLER_20_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_693 ();
 FILLER_ASAP7_75t_R FILLER_20_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_706 ();
 DECAPx2_ASAP7_75t_R FILLER_20_724 ();
 FILLER_ASAP7_75t_R FILLER_20_730 ();
 DECAPx2_ASAP7_75t_R FILLER_20_746 ();
 FILLER_ASAP7_75t_R FILLER_20_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_754 ();
 DECAPx1_ASAP7_75t_R FILLER_20_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_771 ();
 DECAPx2_ASAP7_75t_R FILLER_20_775 ();
 FILLER_ASAP7_75t_R FILLER_20_781 ();
 DECAPx1_ASAP7_75t_R FILLER_20_786 ();
 DECAPx1_ASAP7_75t_R FILLER_20_793 ();
 FILLER_ASAP7_75t_R FILLER_20_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_802 ();
 DECAPx6_ASAP7_75t_R FILLER_20_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_820 ();
 DECAPx1_ASAP7_75t_R FILLER_20_831 ();
 DECAPx10_ASAP7_75t_R FILLER_20_841 ();
 DECAPx2_ASAP7_75t_R FILLER_20_863 ();
 DECAPx1_ASAP7_75t_R FILLER_20_889 ();
 DECAPx1_ASAP7_75t_R FILLER_20_921 ();
 DECAPx2_ASAP7_75t_R FILLER_20_931 ();
 FILLER_ASAP7_75t_R FILLER_20_937 ();
 DECAPx6_ASAP7_75t_R FILLER_20_953 ();
 FILLER_ASAP7_75t_R FILLER_20_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_969 ();
 DECAPx10_ASAP7_75t_R FILLER_20_982 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1378 ();
 FILLER_ASAP7_75t_R FILLER_20_1384 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1388 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1392 ();
 DECAPx10_ASAP7_75t_R FILLER_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_21_90 ();
 DECAPx10_ASAP7_75t_R FILLER_21_112 ();
 DECAPx10_ASAP7_75t_R FILLER_21_134 ();
 DECAPx10_ASAP7_75t_R FILLER_21_156 ();
 DECAPx10_ASAP7_75t_R FILLER_21_178 ();
 DECAPx10_ASAP7_75t_R FILLER_21_200 ();
 DECAPx10_ASAP7_75t_R FILLER_21_222 ();
 DECAPx10_ASAP7_75t_R FILLER_21_244 ();
 DECAPx10_ASAP7_75t_R FILLER_21_266 ();
 DECAPx10_ASAP7_75t_R FILLER_21_288 ();
 DECAPx10_ASAP7_75t_R FILLER_21_310 ();
 DECAPx10_ASAP7_75t_R FILLER_21_332 ();
 DECAPx10_ASAP7_75t_R FILLER_21_354 ();
 DECAPx10_ASAP7_75t_R FILLER_21_376 ();
 DECAPx10_ASAP7_75t_R FILLER_21_398 ();
 DECAPx10_ASAP7_75t_R FILLER_21_420 ();
 DECAPx10_ASAP7_75t_R FILLER_21_442 ();
 DECAPx10_ASAP7_75t_R FILLER_21_464 ();
 DECAPx10_ASAP7_75t_R FILLER_21_486 ();
 DECAPx10_ASAP7_75t_R FILLER_21_508 ();
 DECAPx10_ASAP7_75t_R FILLER_21_530 ();
 DECAPx10_ASAP7_75t_R FILLER_21_552 ();
 DECAPx10_ASAP7_75t_R FILLER_21_574 ();
 DECAPx10_ASAP7_75t_R FILLER_21_596 ();
 DECAPx10_ASAP7_75t_R FILLER_21_618 ();
 DECAPx10_ASAP7_75t_R FILLER_21_640 ();
 DECAPx1_ASAP7_75t_R FILLER_21_662 ();
 DECAPx1_ASAP7_75t_R FILLER_21_676 ();
 DECAPx6_ASAP7_75t_R FILLER_21_692 ();
 FILLER_ASAP7_75t_R FILLER_21_706 ();
 DECAPx1_ASAP7_75t_R FILLER_21_714 ();
 DECAPx4_ASAP7_75t_R FILLER_21_721 ();
 FILLER_ASAP7_75t_R FILLER_21_731 ();
 FILLER_ASAP7_75t_R FILLER_21_739 ();
 DECAPx1_ASAP7_75t_R FILLER_21_755 ();
 DECAPx2_ASAP7_75t_R FILLER_21_765 ();
 DECAPx2_ASAP7_75t_R FILLER_21_774 ();
 FILLER_ASAP7_75t_R FILLER_21_780 ();
 DECAPx1_ASAP7_75t_R FILLER_21_788 ();
 DECAPx1_ASAP7_75t_R FILLER_21_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_830 ();
 DECAPx6_ASAP7_75t_R FILLER_21_848 ();
 DECAPx1_ASAP7_75t_R FILLER_21_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_886 ();
 DECAPx4_ASAP7_75t_R FILLER_21_890 ();
 FILLER_ASAP7_75t_R FILLER_21_900 ();
 DECAPx2_ASAP7_75t_R FILLER_21_908 ();
 FILLER_ASAP7_75t_R FILLER_21_914 ();
 DECAPx1_ASAP7_75t_R FILLER_21_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_923 ();
 DECAPx10_ASAP7_75t_R FILLER_21_926 ();
 DECAPx4_ASAP7_75t_R FILLER_21_948 ();
 FILLER_ASAP7_75t_R FILLER_21_958 ();
 DECAPx1_ASAP7_75t_R FILLER_21_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_978 ();
 DECAPx10_ASAP7_75t_R FILLER_21_991 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1365 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1387 ();
 DECAPx1_ASAP7_75t_R FILLER_21_1401 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_22_112 ();
 DECAPx10_ASAP7_75t_R FILLER_22_134 ();
 DECAPx10_ASAP7_75t_R FILLER_22_156 ();
 DECAPx10_ASAP7_75t_R FILLER_22_178 ();
 DECAPx10_ASAP7_75t_R FILLER_22_200 ();
 DECAPx10_ASAP7_75t_R FILLER_22_222 ();
 DECAPx10_ASAP7_75t_R FILLER_22_244 ();
 DECAPx10_ASAP7_75t_R FILLER_22_266 ();
 DECAPx10_ASAP7_75t_R FILLER_22_288 ();
 DECAPx10_ASAP7_75t_R FILLER_22_310 ();
 DECAPx10_ASAP7_75t_R FILLER_22_332 ();
 DECAPx10_ASAP7_75t_R FILLER_22_354 ();
 DECAPx10_ASAP7_75t_R FILLER_22_376 ();
 DECAPx10_ASAP7_75t_R FILLER_22_398 ();
 DECAPx10_ASAP7_75t_R FILLER_22_420 ();
 DECAPx6_ASAP7_75t_R FILLER_22_442 ();
 DECAPx2_ASAP7_75t_R FILLER_22_456 ();
 DECAPx10_ASAP7_75t_R FILLER_22_464 ();
 DECAPx10_ASAP7_75t_R FILLER_22_486 ();
 DECAPx10_ASAP7_75t_R FILLER_22_508 ();
 DECAPx10_ASAP7_75t_R FILLER_22_530 ();
 DECAPx10_ASAP7_75t_R FILLER_22_552 ();
 DECAPx10_ASAP7_75t_R FILLER_22_574 ();
 DECAPx10_ASAP7_75t_R FILLER_22_596 ();
 DECAPx10_ASAP7_75t_R FILLER_22_618 ();
 DECAPx4_ASAP7_75t_R FILLER_22_640 ();
 FILLER_ASAP7_75t_R FILLER_22_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_652 ();
 DECAPx4_ASAP7_75t_R FILLER_22_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_675 ();
 DECAPx2_ASAP7_75t_R FILLER_22_690 ();
 FILLER_ASAP7_75t_R FILLER_22_696 ();
 DECAPx1_ASAP7_75t_R FILLER_22_704 ();
 DECAPx2_ASAP7_75t_R FILLER_22_714 ();
 FILLER_ASAP7_75t_R FILLER_22_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_722 ();
 DECAPx4_ASAP7_75t_R FILLER_22_741 ();
 FILLER_ASAP7_75t_R FILLER_22_754 ();
 FILLER_ASAP7_75t_R FILLER_22_768 ();
 DECAPx6_ASAP7_75t_R FILLER_22_798 ();
 FILLER_ASAP7_75t_R FILLER_22_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_824 ();
 DECAPx1_ASAP7_75t_R FILLER_22_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_867 ();
 DECAPx2_ASAP7_75t_R FILLER_22_878 ();
 DECAPx1_ASAP7_75t_R FILLER_22_898 ();
 DECAPx1_ASAP7_75t_R FILLER_22_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_923 ();
 DECAPx1_ASAP7_75t_R FILLER_22_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_942 ();
 DECAPx4_ASAP7_75t_R FILLER_22_971 ();
 FILLER_ASAP7_75t_R FILLER_22_981 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_22_1388 ();
 FILLER_ASAP7_75t_R FILLER_22_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_23_68 ();
 DECAPx10_ASAP7_75t_R FILLER_23_90 ();
 DECAPx10_ASAP7_75t_R FILLER_23_112 ();
 DECAPx10_ASAP7_75t_R FILLER_23_134 ();
 DECAPx10_ASAP7_75t_R FILLER_23_156 ();
 DECAPx10_ASAP7_75t_R FILLER_23_178 ();
 DECAPx10_ASAP7_75t_R FILLER_23_200 ();
 DECAPx10_ASAP7_75t_R FILLER_23_222 ();
 DECAPx10_ASAP7_75t_R FILLER_23_244 ();
 DECAPx10_ASAP7_75t_R FILLER_23_266 ();
 DECAPx10_ASAP7_75t_R FILLER_23_288 ();
 DECAPx10_ASAP7_75t_R FILLER_23_310 ();
 DECAPx10_ASAP7_75t_R FILLER_23_332 ();
 DECAPx10_ASAP7_75t_R FILLER_23_354 ();
 DECAPx10_ASAP7_75t_R FILLER_23_376 ();
 DECAPx10_ASAP7_75t_R FILLER_23_398 ();
 DECAPx10_ASAP7_75t_R FILLER_23_420 ();
 DECAPx10_ASAP7_75t_R FILLER_23_442 ();
 DECAPx10_ASAP7_75t_R FILLER_23_464 ();
 DECAPx10_ASAP7_75t_R FILLER_23_486 ();
 DECAPx10_ASAP7_75t_R FILLER_23_508 ();
 DECAPx10_ASAP7_75t_R FILLER_23_530 ();
 DECAPx10_ASAP7_75t_R FILLER_23_552 ();
 DECAPx10_ASAP7_75t_R FILLER_23_574 ();
 DECAPx10_ASAP7_75t_R FILLER_23_596 ();
 DECAPx10_ASAP7_75t_R FILLER_23_618 ();
 DECAPx4_ASAP7_75t_R FILLER_23_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_650 ();
 DECAPx4_ASAP7_75t_R FILLER_23_665 ();
 FILLER_ASAP7_75t_R FILLER_23_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_700 ();
 DECAPx1_ASAP7_75t_R FILLER_23_707 ();
 DECAPx1_ASAP7_75t_R FILLER_23_749 ();
 DECAPx10_ASAP7_75t_R FILLER_23_770 ();
 FILLER_ASAP7_75t_R FILLER_23_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_794 ();
 DECAPx1_ASAP7_75t_R FILLER_23_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_802 ();
 DECAPx10_ASAP7_75t_R FILLER_23_809 ();
 DECAPx1_ASAP7_75t_R FILLER_23_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_835 ();
 FILLER_ASAP7_75t_R FILLER_23_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_855 ();
 DECAPx1_ASAP7_75t_R FILLER_23_876 ();
 FILLER_ASAP7_75t_R FILLER_23_900 ();
 FILLER_ASAP7_75t_R FILLER_23_922 ();
 DECAPx2_ASAP7_75t_R FILLER_23_943 ();
 FILLER_ASAP7_75t_R FILLER_23_949 ();
 FILLER_ASAP7_75t_R FILLER_23_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_961 ();
 DECAPx10_ASAP7_75t_R FILLER_23_998 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1350 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1372 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx10_ASAP7_75t_R FILLER_24_112 ();
 DECAPx10_ASAP7_75t_R FILLER_24_134 ();
 DECAPx10_ASAP7_75t_R FILLER_24_156 ();
 DECAPx10_ASAP7_75t_R FILLER_24_178 ();
 DECAPx10_ASAP7_75t_R FILLER_24_200 ();
 DECAPx10_ASAP7_75t_R FILLER_24_222 ();
 DECAPx10_ASAP7_75t_R FILLER_24_244 ();
 DECAPx10_ASAP7_75t_R FILLER_24_266 ();
 DECAPx10_ASAP7_75t_R FILLER_24_288 ();
 DECAPx10_ASAP7_75t_R FILLER_24_310 ();
 DECAPx10_ASAP7_75t_R FILLER_24_332 ();
 DECAPx10_ASAP7_75t_R FILLER_24_354 ();
 DECAPx10_ASAP7_75t_R FILLER_24_376 ();
 DECAPx10_ASAP7_75t_R FILLER_24_398 ();
 DECAPx10_ASAP7_75t_R FILLER_24_420 ();
 DECAPx6_ASAP7_75t_R FILLER_24_442 ();
 DECAPx2_ASAP7_75t_R FILLER_24_456 ();
 DECAPx10_ASAP7_75t_R FILLER_24_464 ();
 DECAPx10_ASAP7_75t_R FILLER_24_486 ();
 DECAPx10_ASAP7_75t_R FILLER_24_508 ();
 DECAPx10_ASAP7_75t_R FILLER_24_530 ();
 DECAPx10_ASAP7_75t_R FILLER_24_552 ();
 DECAPx10_ASAP7_75t_R FILLER_24_574 ();
 DECAPx10_ASAP7_75t_R FILLER_24_596 ();
 DECAPx10_ASAP7_75t_R FILLER_24_618 ();
 DECAPx4_ASAP7_75t_R FILLER_24_640 ();
 FILLER_ASAP7_75t_R FILLER_24_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_661 ();
 DECAPx1_ASAP7_75t_R FILLER_24_665 ();
 DECAPx4_ASAP7_75t_R FILLER_24_683 ();
 DECAPx4_ASAP7_75t_R FILLER_24_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_723 ();
 FILLER_ASAP7_75t_R FILLER_24_730 ();
 DECAPx1_ASAP7_75t_R FILLER_24_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_748 ();
 DECAPx2_ASAP7_75t_R FILLER_24_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_758 ();
 DECAPx6_ASAP7_75t_R FILLER_24_796 ();
 DECAPx1_ASAP7_75t_R FILLER_24_810 ();
 DECAPx10_ASAP7_75t_R FILLER_24_831 ();
 FILLER_ASAP7_75t_R FILLER_24_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_855 ();
 DECAPx6_ASAP7_75t_R FILLER_24_859 ();
 DECAPx4_ASAP7_75t_R FILLER_24_882 ();
 FILLER_ASAP7_75t_R FILLER_24_892 ();
 DECAPx2_ASAP7_75t_R FILLER_24_906 ();
 FILLER_ASAP7_75t_R FILLER_24_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_914 ();
 DECAPx1_ASAP7_75t_R FILLER_24_921 ();
 DECAPx4_ASAP7_75t_R FILLER_24_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_958 ();
 DECAPx10_ASAP7_75t_R FILLER_24_974 ();
 DECAPx10_ASAP7_75t_R FILLER_24_996 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_24_1370 ();
 FILLER_ASAP7_75t_R FILLER_24_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_24_1388 ();
 FILLER_ASAP7_75t_R FILLER_24_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_25_90 ();
 DECAPx10_ASAP7_75t_R FILLER_25_112 ();
 DECAPx10_ASAP7_75t_R FILLER_25_134 ();
 DECAPx10_ASAP7_75t_R FILLER_25_156 ();
 DECAPx10_ASAP7_75t_R FILLER_25_178 ();
 DECAPx10_ASAP7_75t_R FILLER_25_200 ();
 DECAPx10_ASAP7_75t_R FILLER_25_222 ();
 DECAPx10_ASAP7_75t_R FILLER_25_244 ();
 DECAPx10_ASAP7_75t_R FILLER_25_266 ();
 DECAPx10_ASAP7_75t_R FILLER_25_288 ();
 DECAPx10_ASAP7_75t_R FILLER_25_310 ();
 DECAPx10_ASAP7_75t_R FILLER_25_332 ();
 DECAPx10_ASAP7_75t_R FILLER_25_354 ();
 DECAPx6_ASAP7_75t_R FILLER_25_376 ();
 DECAPx10_ASAP7_75t_R FILLER_25_393 ();
 DECAPx10_ASAP7_75t_R FILLER_25_415 ();
 DECAPx10_ASAP7_75t_R FILLER_25_437 ();
 DECAPx10_ASAP7_75t_R FILLER_25_459 ();
 DECAPx10_ASAP7_75t_R FILLER_25_481 ();
 DECAPx10_ASAP7_75t_R FILLER_25_503 ();
 DECAPx10_ASAP7_75t_R FILLER_25_525 ();
 DECAPx10_ASAP7_75t_R FILLER_25_547 ();
 DECAPx10_ASAP7_75t_R FILLER_25_569 ();
 DECAPx10_ASAP7_75t_R FILLER_25_591 ();
 DECAPx6_ASAP7_75t_R FILLER_25_613 ();
 FILLER_ASAP7_75t_R FILLER_25_627 ();
 DECAPx6_ASAP7_75t_R FILLER_25_635 ();
 FILLER_ASAP7_75t_R FILLER_25_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_661 ();
 DECAPx10_ASAP7_75t_R FILLER_25_688 ();
 DECAPx4_ASAP7_75t_R FILLER_25_710 ();
 FILLER_ASAP7_75t_R FILLER_25_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_722 ();
 DECAPx4_ASAP7_75t_R FILLER_25_743 ();
 FILLER_ASAP7_75t_R FILLER_25_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_755 ();
 DECAPx4_ASAP7_75t_R FILLER_25_762 ();
 DECAPx2_ASAP7_75t_R FILLER_25_775 ();
 FILLER_ASAP7_75t_R FILLER_25_781 ();
 FILLER_ASAP7_75t_R FILLER_25_789 ();
 FILLER_ASAP7_75t_R FILLER_25_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_825 ();
 DECAPx2_ASAP7_75t_R FILLER_25_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_835 ();
 DECAPx4_ASAP7_75t_R FILLER_25_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_849 ();
 DECAPx1_ASAP7_75t_R FILLER_25_853 ();
 DECAPx10_ASAP7_75t_R FILLER_25_860 ();
 DECAPx2_ASAP7_75t_R FILLER_25_882 ();
 FILLER_ASAP7_75t_R FILLER_25_888 ();
 DECAPx2_ASAP7_75t_R FILLER_25_904 ();
 DECAPx1_ASAP7_75t_R FILLER_25_913 ();
 DECAPx1_ASAP7_75t_R FILLER_25_920 ();
 DECAPx6_ASAP7_75t_R FILLER_25_929 ();
 DECAPx4_ASAP7_75t_R FILLER_25_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_967 ();
 DECAPx4_ASAP7_75t_R FILLER_25_971 ();
 FILLER_ASAP7_75t_R FILLER_25_981 ();
 DECAPx10_ASAP7_75t_R FILLER_25_995 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1369 ();
 DECAPx6_ASAP7_75t_R FILLER_25_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 DECAPx10_ASAP7_75t_R FILLER_26_112 ();
 DECAPx10_ASAP7_75t_R FILLER_26_134 ();
 DECAPx10_ASAP7_75t_R FILLER_26_156 ();
 DECAPx10_ASAP7_75t_R FILLER_26_178 ();
 DECAPx10_ASAP7_75t_R FILLER_26_200 ();
 DECAPx10_ASAP7_75t_R FILLER_26_222 ();
 DECAPx4_ASAP7_75t_R FILLER_26_244 ();
 FILLER_ASAP7_75t_R FILLER_26_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_285 ();
 FILLER_ASAP7_75t_R FILLER_26_318 ();
 DECAPx2_ASAP7_75t_R FILLER_26_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_352 ();
 DECAPx6_ASAP7_75t_R FILLER_26_357 ();
 DECAPx1_ASAP7_75t_R FILLER_26_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_375 ();
 DECAPx10_ASAP7_75t_R FILLER_26_402 ();
 DECAPx10_ASAP7_75t_R FILLER_26_424 ();
 DECAPx6_ASAP7_75t_R FILLER_26_446 ();
 FILLER_ASAP7_75t_R FILLER_26_460 ();
 DECAPx10_ASAP7_75t_R FILLER_26_464 ();
 DECAPx10_ASAP7_75t_R FILLER_26_486 ();
 DECAPx10_ASAP7_75t_R FILLER_26_508 ();
 DECAPx10_ASAP7_75t_R FILLER_26_530 ();
 DECAPx10_ASAP7_75t_R FILLER_26_552 ();
 DECAPx10_ASAP7_75t_R FILLER_26_574 ();
 DECAPx10_ASAP7_75t_R FILLER_26_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_618 ();
 DECAPx1_ASAP7_75t_R FILLER_26_639 ();
 DECAPx4_ASAP7_75t_R FILLER_26_657 ();
 FILLER_ASAP7_75t_R FILLER_26_667 ();
 DECAPx6_ASAP7_75t_R FILLER_26_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_692 ();
 DECAPx4_ASAP7_75t_R FILLER_26_705 ();
 FILLER_ASAP7_75t_R FILLER_26_715 ();
 DECAPx2_ASAP7_75t_R FILLER_26_723 ();
 FILLER_ASAP7_75t_R FILLER_26_729 ();
 FILLER_ASAP7_75t_R FILLER_26_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_748 ();
 DECAPx2_ASAP7_75t_R FILLER_26_772 ();
 FILLER_ASAP7_75t_R FILLER_26_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_780 ();
 DECAPx2_ASAP7_75t_R FILLER_26_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_807 ();
 DECAPx2_ASAP7_75t_R FILLER_26_825 ();
 FILLER_ASAP7_75t_R FILLER_26_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_847 ();
 FILLER_ASAP7_75t_R FILLER_26_868 ();
 DECAPx4_ASAP7_75t_R FILLER_26_904 ();
 FILLER_ASAP7_75t_R FILLER_26_914 ();
 DECAPx4_ASAP7_75t_R FILLER_26_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_940 ();
 DECAPx10_ASAP7_75t_R FILLER_26_995 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1347 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1369 ();
 FILLER_ASAP7_75t_R FILLER_26_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1388 ();
 FILLER_ASAP7_75t_R FILLER_26_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_27_90 ();
 DECAPx10_ASAP7_75t_R FILLER_27_112 ();
 DECAPx10_ASAP7_75t_R FILLER_27_134 ();
 DECAPx10_ASAP7_75t_R FILLER_27_156 ();
 DECAPx10_ASAP7_75t_R FILLER_27_178 ();
 DECAPx10_ASAP7_75t_R FILLER_27_200 ();
 DECAPx10_ASAP7_75t_R FILLER_27_222 ();
 DECAPx6_ASAP7_75t_R FILLER_27_244 ();
 DECAPx2_ASAP7_75t_R FILLER_27_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_264 ();
 FILLER_ASAP7_75t_R FILLER_27_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_299 ();
 DECAPx1_ASAP7_75t_R FILLER_27_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_330 ();
 FILLER_ASAP7_75t_R FILLER_27_390 ();
 DECAPx2_ASAP7_75t_R FILLER_27_424 ();
 DECAPx10_ASAP7_75t_R FILLER_27_433 ();
 DECAPx10_ASAP7_75t_R FILLER_27_455 ();
 DECAPx10_ASAP7_75t_R FILLER_27_477 ();
 DECAPx10_ASAP7_75t_R FILLER_27_499 ();
 DECAPx10_ASAP7_75t_R FILLER_27_521 ();
 DECAPx10_ASAP7_75t_R FILLER_27_543 ();
 DECAPx10_ASAP7_75t_R FILLER_27_565 ();
 DECAPx10_ASAP7_75t_R FILLER_27_587 ();
 DECAPx6_ASAP7_75t_R FILLER_27_609 ();
 FILLER_ASAP7_75t_R FILLER_27_623 ();
 DECAPx1_ASAP7_75t_R FILLER_27_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_688 ();
 FILLER_ASAP7_75t_R FILLER_27_715 ();
 DECAPx2_ASAP7_75t_R FILLER_27_729 ();
 FILLER_ASAP7_75t_R FILLER_27_735 ();
 DECAPx6_ASAP7_75t_R FILLER_27_740 ();
 DECAPx1_ASAP7_75t_R FILLER_27_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_758 ();
 DECAPx10_ASAP7_75t_R FILLER_27_765 ();
 DECAPx2_ASAP7_75t_R FILLER_27_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_793 ();
 DECAPx1_ASAP7_75t_R FILLER_27_797 ();
 DECAPx6_ASAP7_75t_R FILLER_27_804 ();
 DECAPx2_ASAP7_75t_R FILLER_27_821 ();
 FILLER_ASAP7_75t_R FILLER_27_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_857 ();
 DECAPx1_ASAP7_75t_R FILLER_27_881 ();
 FILLER_ASAP7_75t_R FILLER_27_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_890 ();
 FILLER_ASAP7_75t_R FILLER_27_897 ();
 FILLER_ASAP7_75t_R FILLER_27_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_923 ();
 FILLER_ASAP7_75t_R FILLER_27_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_933 ();
 DECAPx6_ASAP7_75t_R FILLER_27_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_966 ();
 DECAPx1_ASAP7_75t_R FILLER_27_970 ();
 DECAPx10_ASAP7_75t_R FILLER_27_989 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1363 ();
 DECAPx6_ASAP7_75t_R FILLER_27_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_28_68 ();
 DECAPx10_ASAP7_75t_R FILLER_28_90 ();
 DECAPx10_ASAP7_75t_R FILLER_28_112 ();
 DECAPx10_ASAP7_75t_R FILLER_28_134 ();
 DECAPx10_ASAP7_75t_R FILLER_28_156 ();
 DECAPx10_ASAP7_75t_R FILLER_28_178 ();
 DECAPx10_ASAP7_75t_R FILLER_28_200 ();
 DECAPx10_ASAP7_75t_R FILLER_28_222 ();
 DECAPx10_ASAP7_75t_R FILLER_28_244 ();
 FILLER_ASAP7_75t_R FILLER_28_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_319 ();
 FILLER_ASAP7_75t_R FILLER_28_339 ();
 DECAPx1_ASAP7_75t_R FILLER_28_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_373 ();
 FILLER_ASAP7_75t_R FILLER_28_393 ();
 FILLER_ASAP7_75t_R FILLER_28_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_403 ();
 DECAPx6_ASAP7_75t_R FILLER_28_445 ();
 FILLER_ASAP7_75t_R FILLER_28_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_461 ();
 DECAPx10_ASAP7_75t_R FILLER_28_464 ();
 DECAPx10_ASAP7_75t_R FILLER_28_486 ();
 DECAPx10_ASAP7_75t_R FILLER_28_508 ();
 DECAPx10_ASAP7_75t_R FILLER_28_530 ();
 DECAPx10_ASAP7_75t_R FILLER_28_552 ();
 DECAPx10_ASAP7_75t_R FILLER_28_574 ();
 DECAPx10_ASAP7_75t_R FILLER_28_596 ();
 DECAPx4_ASAP7_75t_R FILLER_28_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_628 ();
 DECAPx2_ASAP7_75t_R FILLER_28_639 ();
 FILLER_ASAP7_75t_R FILLER_28_645 ();
 DECAPx2_ASAP7_75t_R FILLER_28_653 ();
 DECAPx4_ASAP7_75t_R FILLER_28_662 ();
 FILLER_ASAP7_75t_R FILLER_28_731 ();
 DECAPx2_ASAP7_75t_R FILLER_28_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_759 ();
 DECAPx6_ASAP7_75t_R FILLER_28_763 ();
 DECAPx1_ASAP7_75t_R FILLER_28_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_781 ();
 DECAPx4_ASAP7_75t_R FILLER_28_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_836 ();
 FILLER_ASAP7_75t_R FILLER_28_843 ();
 DECAPx2_ASAP7_75t_R FILLER_28_867 ();
 FILLER_ASAP7_75t_R FILLER_28_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_875 ();
 DECAPx1_ASAP7_75t_R FILLER_28_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_883 ();
 DECAPx2_ASAP7_75t_R FILLER_28_887 ();
 FILLER_ASAP7_75t_R FILLER_28_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_920 ();
 DECAPx4_ASAP7_75t_R FILLER_28_952 ();
 FILLER_ASAP7_75t_R FILLER_28_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_964 ();
 DECAPx10_ASAP7_75t_R FILLER_28_982 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1378 ();
 FILLER_ASAP7_75t_R FILLER_28_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_28_1388 ();
 FILLER_ASAP7_75t_R FILLER_28_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_29_68 ();
 DECAPx10_ASAP7_75t_R FILLER_29_90 ();
 DECAPx10_ASAP7_75t_R FILLER_29_112 ();
 DECAPx10_ASAP7_75t_R FILLER_29_134 ();
 DECAPx10_ASAP7_75t_R FILLER_29_156 ();
 DECAPx10_ASAP7_75t_R FILLER_29_178 ();
 DECAPx10_ASAP7_75t_R FILLER_29_200 ();
 DECAPx10_ASAP7_75t_R FILLER_29_222 ();
 DECAPx10_ASAP7_75t_R FILLER_29_244 ();
 DECAPx4_ASAP7_75t_R FILLER_29_266 ();
 DECAPx4_ASAP7_75t_R FILLER_29_279 ();
 DECAPx10_ASAP7_75t_R FILLER_29_292 ();
 DECAPx10_ASAP7_75t_R FILLER_29_314 ();
 DECAPx10_ASAP7_75t_R FILLER_29_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_358 ();
 DECAPx1_ASAP7_75t_R FILLER_29_385 ();
 DECAPx6_ASAP7_75t_R FILLER_29_427 ();
 DECAPx1_ASAP7_75t_R FILLER_29_441 ();
 DECAPx10_ASAP7_75t_R FILLER_29_454 ();
 DECAPx10_ASAP7_75t_R FILLER_29_476 ();
 DECAPx10_ASAP7_75t_R FILLER_29_498 ();
 DECAPx10_ASAP7_75t_R FILLER_29_520 ();
 DECAPx10_ASAP7_75t_R FILLER_29_542 ();
 DECAPx10_ASAP7_75t_R FILLER_29_564 ();
 DECAPx10_ASAP7_75t_R FILLER_29_586 ();
 DECAPx10_ASAP7_75t_R FILLER_29_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_650 ();
 DECAPx1_ASAP7_75t_R FILLER_29_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_682 ();
 FILLER_ASAP7_75t_R FILLER_29_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_688 ();
 FILLER_ASAP7_75t_R FILLER_29_704 ();
 DECAPx1_ASAP7_75t_R FILLER_29_712 ();
 DECAPx2_ASAP7_75t_R FILLER_29_719 ();
 FILLER_ASAP7_75t_R FILLER_29_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_727 ();
 FILLER_ASAP7_75t_R FILLER_29_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_733 ();
 FILLER_ASAP7_75t_R FILLER_29_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_770 ();
 DECAPx2_ASAP7_75t_R FILLER_29_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_787 ();
 FILLER_ASAP7_75t_R FILLER_29_794 ();
 DECAPx6_ASAP7_75t_R FILLER_29_841 ();
 DECAPx6_ASAP7_75t_R FILLER_29_900 ();
 DECAPx1_ASAP7_75t_R FILLER_29_914 ();
 DECAPx4_ASAP7_75t_R FILLER_29_940 ();
 FILLER_ASAP7_75t_R FILLER_29_950 ();
 DECAPx4_ASAP7_75t_R FILLER_29_958 ();
 FILLER_ASAP7_75t_R FILLER_29_968 ();
 DECAPx10_ASAP7_75t_R FILLER_29_985 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1359 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1381 ();
 FILLER_ASAP7_75t_R FILLER_29_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_30_68 ();
 DECAPx10_ASAP7_75t_R FILLER_30_90 ();
 DECAPx10_ASAP7_75t_R FILLER_30_112 ();
 DECAPx10_ASAP7_75t_R FILLER_30_134 ();
 DECAPx10_ASAP7_75t_R FILLER_30_156 ();
 DECAPx10_ASAP7_75t_R FILLER_30_178 ();
 DECAPx10_ASAP7_75t_R FILLER_30_200 ();
 DECAPx4_ASAP7_75t_R FILLER_30_222 ();
 FILLER_ASAP7_75t_R FILLER_30_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_234 ();
 DECAPx6_ASAP7_75t_R FILLER_30_267 ();
 FILLER_ASAP7_75t_R FILLER_30_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_283 ();
 DECAPx1_ASAP7_75t_R FILLER_30_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_328 ();
 DECAPx1_ASAP7_75t_R FILLER_30_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_359 ();
 FILLER_ASAP7_75t_R FILLER_30_372 ();
 DECAPx1_ASAP7_75t_R FILLER_30_377 ();
 DECAPx4_ASAP7_75t_R FILLER_30_385 ();
 FILLER_ASAP7_75t_R FILLER_30_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_397 ();
 DECAPx2_ASAP7_75t_R FILLER_30_404 ();
 DECAPx10_ASAP7_75t_R FILLER_30_464 ();
 DECAPx10_ASAP7_75t_R FILLER_30_486 ();
 DECAPx10_ASAP7_75t_R FILLER_30_508 ();
 DECAPx10_ASAP7_75t_R FILLER_30_530 ();
 DECAPx10_ASAP7_75t_R FILLER_30_552 ();
 DECAPx10_ASAP7_75t_R FILLER_30_574 ();
 DECAPx10_ASAP7_75t_R FILLER_30_596 ();
 DECAPx10_ASAP7_75t_R FILLER_30_618 ();
 DECAPx6_ASAP7_75t_R FILLER_30_640 ();
 DECAPx2_ASAP7_75t_R FILLER_30_654 ();
 DECAPx2_ASAP7_75t_R FILLER_30_663 ();
 DECAPx10_ASAP7_75t_R FILLER_30_672 ();
 DECAPx6_ASAP7_75t_R FILLER_30_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_708 ();
 DECAPx6_ASAP7_75t_R FILLER_30_712 ();
 FILLER_ASAP7_75t_R FILLER_30_726 ();
 DECAPx2_ASAP7_75t_R FILLER_30_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_769 ();
 FILLER_ASAP7_75t_R FILLER_30_773 ();
 DECAPx2_ASAP7_75t_R FILLER_30_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_804 ();
 FILLER_ASAP7_75t_R FILLER_30_835 ();
 DECAPx2_ASAP7_75t_R FILLER_30_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_872 ();
 FILLER_ASAP7_75t_R FILLER_30_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_889 ();
 DECAPx6_ASAP7_75t_R FILLER_30_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_924 ();
 DECAPx4_ASAP7_75t_R FILLER_30_928 ();
 FILLER_ASAP7_75t_R FILLER_30_938 ();
 DECAPx1_ASAP7_75t_R FILLER_30_943 ();
 DECAPx10_ASAP7_75t_R FILLER_30_989 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1388 ();
 FILLER_ASAP7_75t_R FILLER_30_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_31_68 ();
 DECAPx10_ASAP7_75t_R FILLER_31_90 ();
 DECAPx10_ASAP7_75t_R FILLER_31_112 ();
 DECAPx10_ASAP7_75t_R FILLER_31_134 ();
 DECAPx10_ASAP7_75t_R FILLER_31_156 ();
 DECAPx10_ASAP7_75t_R FILLER_31_178 ();
 DECAPx10_ASAP7_75t_R FILLER_31_200 ();
 DECAPx2_ASAP7_75t_R FILLER_31_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_254 ();
 FILLER_ASAP7_75t_R FILLER_31_299 ();
 FILLER_ASAP7_75t_R FILLER_31_330 ();
 DECAPx4_ASAP7_75t_R FILLER_31_351 ();
 FILLER_ASAP7_75t_R FILLER_31_361 ();
 DECAPx2_ASAP7_75t_R FILLER_31_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_375 ();
 DECAPx6_ASAP7_75t_R FILLER_31_379 ();
 DECAPx2_ASAP7_75t_R FILLER_31_393 ();
 DECAPx1_ASAP7_75t_R FILLER_31_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_409 ();
 FILLER_ASAP7_75t_R FILLER_31_413 ();
 DECAPx2_ASAP7_75t_R FILLER_31_424 ();
 FILLER_ASAP7_75t_R FILLER_31_433 ();
 FILLER_ASAP7_75t_R FILLER_31_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_440 ();
 DECAPx2_ASAP7_75t_R FILLER_31_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_456 ();
 DECAPx10_ASAP7_75t_R FILLER_31_463 ();
 DECAPx10_ASAP7_75t_R FILLER_31_485 ();
 DECAPx10_ASAP7_75t_R FILLER_31_507 ();
 DECAPx10_ASAP7_75t_R FILLER_31_529 ();
 DECAPx10_ASAP7_75t_R FILLER_31_551 ();
 DECAPx10_ASAP7_75t_R FILLER_31_573 ();
 DECAPx10_ASAP7_75t_R FILLER_31_595 ();
 DECAPx4_ASAP7_75t_R FILLER_31_617 ();
 FILLER_ASAP7_75t_R FILLER_31_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_629 ();
 DECAPx4_ASAP7_75t_R FILLER_31_642 ();
 DECAPx6_ASAP7_75t_R FILLER_31_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_684 ();
 DECAPx6_ASAP7_75t_R FILLER_31_699 ();
 DECAPx1_ASAP7_75t_R FILLER_31_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_717 ();
 DECAPx6_ASAP7_75t_R FILLER_31_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_752 ();
 DECAPx4_ASAP7_75t_R FILLER_31_756 ();
 DECAPx1_ASAP7_75t_R FILLER_31_769 ();
 DECAPx4_ASAP7_75t_R FILLER_31_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_800 ();
 DECAPx2_ASAP7_75t_R FILLER_31_807 ();
 FILLER_ASAP7_75t_R FILLER_31_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_815 ();
 DECAPx10_ASAP7_75t_R FILLER_31_819 ();
 DECAPx4_ASAP7_75t_R FILLER_31_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_851 ();
 FILLER_ASAP7_75t_R FILLER_31_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_857 ();
 DECAPx4_ASAP7_75t_R FILLER_31_864 ();
 DECAPx4_ASAP7_75t_R FILLER_31_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_898 ();
 DECAPx2_ASAP7_75t_R FILLER_31_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_923 ();
 DECAPx2_ASAP7_75t_R FILLER_31_926 ();
 FILLER_ASAP7_75t_R FILLER_31_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_934 ();
 DECAPx4_ASAP7_75t_R FILLER_31_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_948 ();
 FILLER_ASAP7_75t_R FILLER_31_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_954 ();
 DECAPx1_ASAP7_75t_R FILLER_31_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_976 ();
 DECAPx10_ASAP7_75t_R FILLER_31_989 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1363 ();
 DECAPx6_ASAP7_75t_R FILLER_31_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_32_68 ();
 DECAPx10_ASAP7_75t_R FILLER_32_90 ();
 DECAPx10_ASAP7_75t_R FILLER_32_112 ();
 DECAPx10_ASAP7_75t_R FILLER_32_134 ();
 DECAPx10_ASAP7_75t_R FILLER_32_156 ();
 DECAPx10_ASAP7_75t_R FILLER_32_178 ();
 DECAPx10_ASAP7_75t_R FILLER_32_200 ();
 DECAPx6_ASAP7_75t_R FILLER_32_222 ();
 FILLER_ASAP7_75t_R FILLER_32_236 ();
 FILLER_ASAP7_75t_R FILLER_32_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_249 ();
 FILLER_ASAP7_75t_R FILLER_32_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_255 ();
 DECAPx2_ASAP7_75t_R FILLER_32_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_269 ();
 DECAPx2_ASAP7_75t_R FILLER_32_285 ();
 FILLER_ASAP7_75t_R FILLER_32_291 ();
 DECAPx1_ASAP7_75t_R FILLER_32_306 ();
 FILLER_ASAP7_75t_R FILLER_32_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_318 ();
 DECAPx2_ASAP7_75t_R FILLER_32_325 ();
 DECAPx2_ASAP7_75t_R FILLER_32_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_343 ();
 DECAPx4_ASAP7_75t_R FILLER_32_350 ();
 FILLER_ASAP7_75t_R FILLER_32_360 ();
 DECAPx2_ASAP7_75t_R FILLER_32_391 ();
 DECAPx10_ASAP7_75t_R FILLER_32_403 ();
 DECAPx6_ASAP7_75t_R FILLER_32_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_439 ();
 DECAPx2_ASAP7_75t_R FILLER_32_448 ();
 FILLER_ASAP7_75t_R FILLER_32_454 ();
 FILLER_ASAP7_75t_R FILLER_32_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_492 ();
 DECAPx10_ASAP7_75t_R FILLER_32_515 ();
 DECAPx10_ASAP7_75t_R FILLER_32_537 ();
 DECAPx10_ASAP7_75t_R FILLER_32_559 ();
 DECAPx10_ASAP7_75t_R FILLER_32_581 ();
 DECAPx6_ASAP7_75t_R FILLER_32_603 ();
 DECAPx1_ASAP7_75t_R FILLER_32_617 ();
 FILLER_ASAP7_75t_R FILLER_32_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_643 ();
 DECAPx1_ASAP7_75t_R FILLER_32_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_654 ();
 DECAPx1_ASAP7_75t_R FILLER_32_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_702 ();
 FILLER_ASAP7_75t_R FILLER_32_720 ();
 FILLER_ASAP7_75t_R FILLER_32_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_727 ();
 FILLER_ASAP7_75t_R FILLER_32_737 ();
 DECAPx6_ASAP7_75t_R FILLER_32_742 ();
 DECAPx2_ASAP7_75t_R FILLER_32_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_762 ();
 DECAPx4_ASAP7_75t_R FILLER_32_776 ();
 DECAPx2_ASAP7_75t_R FILLER_32_792 ();
 FILLER_ASAP7_75t_R FILLER_32_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_800 ();
 DECAPx4_ASAP7_75t_R FILLER_32_811 ();
 FILLER_ASAP7_75t_R FILLER_32_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_823 ();
 DECAPx2_ASAP7_75t_R FILLER_32_866 ();
 FILLER_ASAP7_75t_R FILLER_32_872 ();
 DECAPx2_ASAP7_75t_R FILLER_32_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_886 ();
 FILLER_ASAP7_75t_R FILLER_32_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_906 ();
 DECAPx2_ASAP7_75t_R FILLER_32_949 ();
 DECAPx2_ASAP7_75t_R FILLER_32_958 ();
 FILLER_ASAP7_75t_R FILLER_32_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_966 ();
 DECAPx2_ASAP7_75t_R FILLER_32_970 ();
 DECAPx10_ASAP7_75t_R FILLER_32_979 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1388 ();
 FILLER_ASAP7_75t_R FILLER_32_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_33_68 ();
 DECAPx10_ASAP7_75t_R FILLER_33_90 ();
 DECAPx10_ASAP7_75t_R FILLER_33_112 ();
 DECAPx10_ASAP7_75t_R FILLER_33_134 ();
 DECAPx10_ASAP7_75t_R FILLER_33_156 ();
 DECAPx10_ASAP7_75t_R FILLER_33_178 ();
 DECAPx10_ASAP7_75t_R FILLER_33_200 ();
 DECAPx10_ASAP7_75t_R FILLER_33_222 ();
 FILLER_ASAP7_75t_R FILLER_33_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_246 ();
 DECAPx10_ASAP7_75t_R FILLER_33_273 ();
 DECAPx4_ASAP7_75t_R FILLER_33_301 ();
 FILLER_ASAP7_75t_R FILLER_33_311 ();
 DECAPx2_ASAP7_75t_R FILLER_33_371 ();
 FILLER_ASAP7_75t_R FILLER_33_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_379 ();
 FILLER_ASAP7_75t_R FILLER_33_409 ();
 DECAPx2_ASAP7_75t_R FILLER_33_437 ();
 FILLER_ASAP7_75t_R FILLER_33_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_471 ();
 FILLER_ASAP7_75t_R FILLER_33_475 ();
 DECAPx10_ASAP7_75t_R FILLER_33_481 ();
 DECAPx10_ASAP7_75t_R FILLER_33_503 ();
 DECAPx10_ASAP7_75t_R FILLER_33_525 ();
 DECAPx10_ASAP7_75t_R FILLER_33_547 ();
 DECAPx10_ASAP7_75t_R FILLER_33_569 ();
 DECAPx10_ASAP7_75t_R FILLER_33_591 ();
 FILLER_ASAP7_75t_R FILLER_33_613 ();
 DECAPx4_ASAP7_75t_R FILLER_33_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_640 ();
 DECAPx10_ASAP7_75t_R FILLER_33_653 ();
 FILLER_ASAP7_75t_R FILLER_33_675 ();
 FILLER_ASAP7_75t_R FILLER_33_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_685 ();
 FILLER_ASAP7_75t_R FILLER_33_689 ();
 DECAPx1_ASAP7_75t_R FILLER_33_747 ();
 FILLER_ASAP7_75t_R FILLER_33_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_759 ();
 DECAPx6_ASAP7_75t_R FILLER_33_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_777 ();
 DECAPx2_ASAP7_75t_R FILLER_33_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_826 ();
 FILLER_ASAP7_75t_R FILLER_33_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_849 ();
 DECAPx6_ASAP7_75t_R FILLER_33_867 ();
 DECAPx1_ASAP7_75t_R FILLER_33_881 ();
 DECAPx6_ASAP7_75t_R FILLER_33_888 ();
 FILLER_ASAP7_75t_R FILLER_33_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_904 ();
 DECAPx1_ASAP7_75t_R FILLER_33_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_923 ();
 DECAPx2_ASAP7_75t_R FILLER_33_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_939 ();
 DECAPx6_ASAP7_75t_R FILLER_33_957 ();
 DECAPx1_ASAP7_75t_R FILLER_33_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_975 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1377 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_34_68 ();
 DECAPx10_ASAP7_75t_R FILLER_34_90 ();
 DECAPx10_ASAP7_75t_R FILLER_34_112 ();
 DECAPx10_ASAP7_75t_R FILLER_34_134 ();
 DECAPx10_ASAP7_75t_R FILLER_34_156 ();
 DECAPx10_ASAP7_75t_R FILLER_34_178 ();
 DECAPx6_ASAP7_75t_R FILLER_34_200 ();
 DECAPx2_ASAP7_75t_R FILLER_34_214 ();
 DECAPx2_ASAP7_75t_R FILLER_34_252 ();
 DECAPx4_ASAP7_75t_R FILLER_34_277 ();
 FILLER_ASAP7_75t_R FILLER_34_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_289 ();
 DECAPx4_ASAP7_75t_R FILLER_34_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_326 ();
 DECAPx1_ASAP7_75t_R FILLER_34_330 ();
 DECAPx2_ASAP7_75t_R FILLER_34_337 ();
 FILLER_ASAP7_75t_R FILLER_34_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_352 ();
 DECAPx4_ASAP7_75t_R FILLER_34_382 ();
 FILLER_ASAP7_75t_R FILLER_34_392 ();
 FILLER_ASAP7_75t_R FILLER_34_400 ();
 FILLER_ASAP7_75t_R FILLER_34_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_461 ();
 DECAPx1_ASAP7_75t_R FILLER_34_464 ();
 DECAPx10_ASAP7_75t_R FILLER_34_494 ();
 DECAPx10_ASAP7_75t_R FILLER_34_516 ();
 DECAPx10_ASAP7_75t_R FILLER_34_538 ();
 DECAPx10_ASAP7_75t_R FILLER_34_560 ();
 DECAPx10_ASAP7_75t_R FILLER_34_582 ();
 DECAPx2_ASAP7_75t_R FILLER_34_604 ();
 FILLER_ASAP7_75t_R FILLER_34_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_627 ();
 FILLER_ASAP7_75t_R FILLER_34_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_644 ();
 DECAPx6_ASAP7_75t_R FILLER_34_673 ();
 DECAPx2_ASAP7_75t_R FILLER_34_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_693 ();
 DECAPx1_ASAP7_75t_R FILLER_34_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_701 ();
 DECAPx4_ASAP7_75t_R FILLER_34_720 ();
 FILLER_ASAP7_75t_R FILLER_34_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_732 ();
 DECAPx4_ASAP7_75t_R FILLER_34_739 ();
 FILLER_ASAP7_75t_R FILLER_34_749 ();
 DECAPx4_ASAP7_75t_R FILLER_34_774 ();
 FILLER_ASAP7_75t_R FILLER_34_784 ();
 DECAPx2_ASAP7_75t_R FILLER_34_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_813 ();
 DECAPx1_ASAP7_75t_R FILLER_34_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_853 ();
 DECAPx1_ASAP7_75t_R FILLER_34_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_861 ();
 DECAPx4_ASAP7_75t_R FILLER_34_865 ();
 DECAPx1_ASAP7_75t_R FILLER_34_884 ();
 DECAPx1_ASAP7_75t_R FILLER_34_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_904 ();
 DECAPx4_ASAP7_75t_R FILLER_34_908 ();
 FILLER_ASAP7_75t_R FILLER_34_918 ();
 FILLER_ASAP7_75t_R FILLER_34_951 ();
 DECAPx2_ASAP7_75t_R FILLER_34_959 ();
 FILLER_ASAP7_75t_R FILLER_34_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_967 ();
 FILLER_ASAP7_75t_R FILLER_34_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_979 ();
 DECAPx10_ASAP7_75t_R FILLER_34_989 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_34_1388 ();
 FILLER_ASAP7_75t_R FILLER_34_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_35_68 ();
 DECAPx10_ASAP7_75t_R FILLER_35_90 ();
 DECAPx10_ASAP7_75t_R FILLER_35_112 ();
 DECAPx10_ASAP7_75t_R FILLER_35_134 ();
 DECAPx10_ASAP7_75t_R FILLER_35_156 ();
 DECAPx10_ASAP7_75t_R FILLER_35_178 ();
 DECAPx10_ASAP7_75t_R FILLER_35_200 ();
 DECAPx4_ASAP7_75t_R FILLER_35_222 ();
 FILLER_ASAP7_75t_R FILLER_35_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_234 ();
 FILLER_ASAP7_75t_R FILLER_35_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_240 ();
 DECAPx4_ASAP7_75t_R FILLER_35_250 ();
 FILLER_ASAP7_75t_R FILLER_35_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_266 ();
 DECAPx6_ASAP7_75t_R FILLER_35_273 ();
 DECAPx1_ASAP7_75t_R FILLER_35_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_291 ();
 FILLER_ASAP7_75t_R FILLER_35_298 ();
 DECAPx6_ASAP7_75t_R FILLER_35_342 ();
 FILLER_ASAP7_75t_R FILLER_35_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_358 ();
 FILLER_ASAP7_75t_R FILLER_35_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_364 ();
 DECAPx1_ASAP7_75t_R FILLER_35_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_395 ();
 DECAPx2_ASAP7_75t_R FILLER_35_399 ();
 FILLER_ASAP7_75t_R FILLER_35_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_407 ();
 FILLER_ASAP7_75t_R FILLER_35_426 ();
 DECAPx10_ASAP7_75t_R FILLER_35_450 ();
 DECAPx4_ASAP7_75t_R FILLER_35_472 ();
 DECAPx10_ASAP7_75t_R FILLER_35_511 ();
 DECAPx10_ASAP7_75t_R FILLER_35_533 ();
 DECAPx10_ASAP7_75t_R FILLER_35_555 ();
 DECAPx10_ASAP7_75t_R FILLER_35_577 ();
 DECAPx6_ASAP7_75t_R FILLER_35_599 ();
 DECAPx6_ASAP7_75t_R FILLER_35_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_641 ();
 DECAPx1_ASAP7_75t_R FILLER_35_648 ();
 DECAPx2_ASAP7_75t_R FILLER_35_655 ();
 FILLER_ASAP7_75t_R FILLER_35_661 ();
 FILLER_ASAP7_75t_R FILLER_35_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_672 ();
 FILLER_ASAP7_75t_R FILLER_35_676 ();
 FILLER_ASAP7_75t_R FILLER_35_681 ();
 DECAPx1_ASAP7_75t_R FILLER_35_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_690 ();
 DECAPx6_ASAP7_75t_R FILLER_35_694 ();
 DECAPx10_ASAP7_75t_R FILLER_35_714 ();
 DECAPx1_ASAP7_75t_R FILLER_35_736 ();
 DECAPx1_ASAP7_75t_R FILLER_35_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_747 ();
 FILLER_ASAP7_75t_R FILLER_35_762 ();
 DECAPx6_ASAP7_75t_R FILLER_35_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_804 ();
 DECAPx4_ASAP7_75t_R FILLER_35_822 ();
 DECAPx1_ASAP7_75t_R FILLER_35_835 ();
 DECAPx4_ASAP7_75t_R FILLER_35_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_861 ();
 DECAPx10_ASAP7_75t_R FILLER_35_871 ();
 DECAPx4_ASAP7_75t_R FILLER_35_893 ();
 DECAPx4_ASAP7_75t_R FILLER_35_912 ();
 FILLER_ASAP7_75t_R FILLER_35_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_940 ();
 DECAPx2_ASAP7_75t_R FILLER_35_944 ();
 FILLER_ASAP7_75t_R FILLER_35_950 ();
 DECAPx10_ASAP7_75t_R FILLER_35_989 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1363 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_36_68 ();
 DECAPx10_ASAP7_75t_R FILLER_36_90 ();
 DECAPx10_ASAP7_75t_R FILLER_36_112 ();
 DECAPx10_ASAP7_75t_R FILLER_36_134 ();
 DECAPx10_ASAP7_75t_R FILLER_36_156 ();
 DECAPx10_ASAP7_75t_R FILLER_36_178 ();
 DECAPx4_ASAP7_75t_R FILLER_36_200 ();
 FILLER_ASAP7_75t_R FILLER_36_210 ();
 DECAPx1_ASAP7_75t_R FILLER_36_244 ();
 DECAPx1_ASAP7_75t_R FILLER_36_274 ();
 FILLER_ASAP7_75t_R FILLER_36_310 ();
 DECAPx6_ASAP7_75t_R FILLER_36_341 ();
 FILLER_ASAP7_75t_R FILLER_36_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_370 ();
 FILLER_ASAP7_75t_R FILLER_36_374 ();
 DECAPx6_ASAP7_75t_R FILLER_36_408 ();
 DECAPx1_ASAP7_75t_R FILLER_36_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_429 ();
 DECAPx2_ASAP7_75t_R FILLER_36_464 ();
 FILLER_ASAP7_75t_R FILLER_36_470 ();
 FILLER_ASAP7_75t_R FILLER_36_484 ();
 FILLER_ASAP7_75t_R FILLER_36_498 ();
 DECAPx10_ASAP7_75t_R FILLER_36_526 ();
 DECAPx10_ASAP7_75t_R FILLER_36_548 ();
 DECAPx10_ASAP7_75t_R FILLER_36_570 ();
 DECAPx10_ASAP7_75t_R FILLER_36_592 ();
 DECAPx2_ASAP7_75t_R FILLER_36_614 ();
 FILLER_ASAP7_75t_R FILLER_36_620 ();
 DECAPx6_ASAP7_75t_R FILLER_36_639 ();
 DECAPx2_ASAP7_75t_R FILLER_36_653 ();
 DECAPx2_ASAP7_75t_R FILLER_36_676 ();
 FILLER_ASAP7_75t_R FILLER_36_682 ();
 DECAPx6_ASAP7_75t_R FILLER_36_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_715 ();
 DECAPx6_ASAP7_75t_R FILLER_36_719 ();
 FILLER_ASAP7_75t_R FILLER_36_733 ();
 DECAPx2_ASAP7_75t_R FILLER_36_758 ();
 DECAPx2_ASAP7_75t_R FILLER_36_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_773 ();
 DECAPx2_ASAP7_75t_R FILLER_36_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_783 ();
 DECAPx2_ASAP7_75t_R FILLER_36_798 ();
 DECAPx1_ASAP7_75t_R FILLER_36_818 ();
 DECAPx4_ASAP7_75t_R FILLER_36_828 ();
 DECAPx4_ASAP7_75t_R FILLER_36_847 ();
 FILLER_ASAP7_75t_R FILLER_36_857 ();
 FILLER_ASAP7_75t_R FILLER_36_915 ();
 FILLER_ASAP7_75t_R FILLER_36_920 ();
 DECAPx6_ASAP7_75t_R FILLER_36_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_939 ();
 DECAPx10_ASAP7_75t_R FILLER_36_943 ();
 DECAPx10_ASAP7_75t_R FILLER_36_988 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1362 ();
 FILLER_ASAP7_75t_R FILLER_36_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1388 ();
 FILLER_ASAP7_75t_R FILLER_36_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_37_24 ();
 DECAPx10_ASAP7_75t_R FILLER_37_46 ();
 DECAPx10_ASAP7_75t_R FILLER_37_68 ();
 DECAPx10_ASAP7_75t_R FILLER_37_90 ();
 DECAPx10_ASAP7_75t_R FILLER_37_112 ();
 DECAPx10_ASAP7_75t_R FILLER_37_134 ();
 DECAPx10_ASAP7_75t_R FILLER_37_156 ();
 DECAPx10_ASAP7_75t_R FILLER_37_178 ();
 DECAPx10_ASAP7_75t_R FILLER_37_200 ();
 DECAPx1_ASAP7_75t_R FILLER_37_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_230 ();
 DECAPx2_ASAP7_75t_R FILLER_37_264 ();
 FILLER_ASAP7_75t_R FILLER_37_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_281 ();
 FILLER_ASAP7_75t_R FILLER_37_285 ();
 DECAPx4_ASAP7_75t_R FILLER_37_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_306 ();
 FILLER_ASAP7_75t_R FILLER_37_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_328 ();
 DECAPx4_ASAP7_75t_R FILLER_37_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_378 ();
 DECAPx2_ASAP7_75t_R FILLER_37_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_388 ();
 DECAPx2_ASAP7_75t_R FILLER_37_395 ();
 FILLER_ASAP7_75t_R FILLER_37_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_403 ();
 DECAPx6_ASAP7_75t_R FILLER_37_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_424 ();
 DECAPx2_ASAP7_75t_R FILLER_37_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_470 ();
 DECAPx2_ASAP7_75t_R FILLER_37_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_480 ();
 DECAPx1_ASAP7_75t_R FILLER_37_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_488 ();
 FILLER_ASAP7_75t_R FILLER_37_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_499 ();
 DECAPx2_ASAP7_75t_R FILLER_37_503 ();
 DECAPx10_ASAP7_75t_R FILLER_37_535 ();
 DECAPx10_ASAP7_75t_R FILLER_37_557 ();
 DECAPx10_ASAP7_75t_R FILLER_37_579 ();
 DECAPx6_ASAP7_75t_R FILLER_37_601 ();
 DECAPx4_ASAP7_75t_R FILLER_37_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_631 ();
 DECAPx2_ASAP7_75t_R FILLER_37_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_661 ();
 DECAPx1_ASAP7_75t_R FILLER_37_665 ();
 FILLER_ASAP7_75t_R FILLER_37_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_680 ();
 FILLER_ASAP7_75t_R FILLER_37_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_686 ();
 DECAPx2_ASAP7_75t_R FILLER_37_701 ();
 FILLER_ASAP7_75t_R FILLER_37_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_709 ();
 FILLER_ASAP7_75t_R FILLER_37_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_751 ();
 FILLER_ASAP7_75t_R FILLER_37_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_768 ();
 DECAPx6_ASAP7_75t_R FILLER_37_772 ();
 DECAPx2_ASAP7_75t_R FILLER_37_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_795 ();
 DECAPx6_ASAP7_75t_R FILLER_37_799 ();
 FILLER_ASAP7_75t_R FILLER_37_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_815 ();
 DECAPx1_ASAP7_75t_R FILLER_37_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_823 ();
 DECAPx1_ASAP7_75t_R FILLER_37_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_847 ();
 FILLER_ASAP7_75t_R FILLER_37_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_913 ();
 DECAPx1_ASAP7_75t_R FILLER_37_935 ();
 DECAPx6_ASAP7_75t_R FILLER_37_962 ();
 FILLER_ASAP7_75t_R FILLER_37_976 ();
 DECAPx10_ASAP7_75t_R FILLER_37_981 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1377 ();
 DECAPx2_ASAP7_75t_R FILLER_37_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_38_24 ();
 DECAPx10_ASAP7_75t_R FILLER_38_46 ();
 DECAPx10_ASAP7_75t_R FILLER_38_68 ();
 DECAPx10_ASAP7_75t_R FILLER_38_90 ();
 DECAPx10_ASAP7_75t_R FILLER_38_112 ();
 DECAPx10_ASAP7_75t_R FILLER_38_134 ();
 DECAPx10_ASAP7_75t_R FILLER_38_156 ();
 DECAPx10_ASAP7_75t_R FILLER_38_178 ();
 DECAPx1_ASAP7_75t_R FILLER_38_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_230 ();
 DECAPx6_ASAP7_75t_R FILLER_38_243 ();
 DECAPx1_ASAP7_75t_R FILLER_38_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_261 ();
 DECAPx1_ASAP7_75t_R FILLER_38_326 ();
 DECAPx1_ASAP7_75t_R FILLER_38_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_343 ();
 FILLER_ASAP7_75t_R FILLER_38_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_349 ();
 DECAPx10_ASAP7_75t_R FILLER_38_362 ();
 DECAPx4_ASAP7_75t_R FILLER_38_384 ();
 DECAPx4_ASAP7_75t_R FILLER_38_452 ();
 DECAPx4_ASAP7_75t_R FILLER_38_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_474 ();
 DECAPx10_ASAP7_75t_R FILLER_38_478 ();
 FILLER_ASAP7_75t_R FILLER_38_500 ();
 DECAPx1_ASAP7_75t_R FILLER_38_508 ();
 DECAPx10_ASAP7_75t_R FILLER_38_527 ();
 DECAPx10_ASAP7_75t_R FILLER_38_549 ();
 DECAPx10_ASAP7_75t_R FILLER_38_571 ();
 DECAPx10_ASAP7_75t_R FILLER_38_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_639 ();
 FILLER_ASAP7_75t_R FILLER_38_666 ();
 FILLER_ASAP7_75t_R FILLER_38_696 ();
 DECAPx1_ASAP7_75t_R FILLER_38_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_731 ();
 DECAPx4_ASAP7_75t_R FILLER_38_735 ();
 FILLER_ASAP7_75t_R FILLER_38_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_747 ();
 DECAPx6_ASAP7_75t_R FILLER_38_751 ();
 DECAPx1_ASAP7_75t_R FILLER_38_765 ();
 DECAPx10_ASAP7_75t_R FILLER_38_797 ();
 DECAPx6_ASAP7_75t_R FILLER_38_819 ();
 FILLER_ASAP7_75t_R FILLER_38_833 ();
 FILLER_ASAP7_75t_R FILLER_38_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_879 ();
 DECAPx2_ASAP7_75t_R FILLER_38_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_891 ();
 DECAPx4_ASAP7_75t_R FILLER_38_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_978 ();
 DECAPx10_ASAP7_75t_R FILLER_38_982 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1378 ();
 FILLER_ASAP7_75t_R FILLER_38_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1388 ();
 FILLER_ASAP7_75t_R FILLER_38_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_39_24 ();
 DECAPx10_ASAP7_75t_R FILLER_39_46 ();
 DECAPx10_ASAP7_75t_R FILLER_39_68 ();
 DECAPx10_ASAP7_75t_R FILLER_39_90 ();
 DECAPx10_ASAP7_75t_R FILLER_39_112 ();
 DECAPx10_ASAP7_75t_R FILLER_39_134 ();
 DECAPx10_ASAP7_75t_R FILLER_39_156 ();
 DECAPx10_ASAP7_75t_R FILLER_39_178 ();
 DECAPx6_ASAP7_75t_R FILLER_39_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_221 ();
 DECAPx2_ASAP7_75t_R FILLER_39_225 ();
 DECAPx6_ASAP7_75t_R FILLER_39_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_290 ();
 DECAPx6_ASAP7_75t_R FILLER_39_294 ();
 DECAPx2_ASAP7_75t_R FILLER_39_308 ();
 DECAPx10_ASAP7_75t_R FILLER_39_317 ();
 DECAPx4_ASAP7_75t_R FILLER_39_339 ();
 FILLER_ASAP7_75t_R FILLER_39_349 ();
 DECAPx6_ASAP7_75t_R FILLER_39_360 ();
 FILLER_ASAP7_75t_R FILLER_39_374 ();
 DECAPx2_ASAP7_75t_R FILLER_39_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_388 ();
 DECAPx2_ASAP7_75t_R FILLER_39_392 ();
 FILLER_ASAP7_75t_R FILLER_39_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_400 ();
 DECAPx1_ASAP7_75t_R FILLER_39_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_411 ();
 DECAPx2_ASAP7_75t_R FILLER_39_415 ();
 FILLER_ASAP7_75t_R FILLER_39_421 ();
 DECAPx2_ASAP7_75t_R FILLER_39_429 ();
 FILLER_ASAP7_75t_R FILLER_39_438 ();
 FILLER_ASAP7_75t_R FILLER_39_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_448 ();
 DECAPx1_ASAP7_75t_R FILLER_39_487 ();
 DECAPx4_ASAP7_75t_R FILLER_39_494 ();
 FILLER_ASAP7_75t_R FILLER_39_513 ();
 DECAPx4_ASAP7_75t_R FILLER_39_518 ();
 FILLER_ASAP7_75t_R FILLER_39_528 ();
 DECAPx10_ASAP7_75t_R FILLER_39_536 ();
 DECAPx10_ASAP7_75t_R FILLER_39_558 ();
 DECAPx10_ASAP7_75t_R FILLER_39_580 ();
 DECAPx4_ASAP7_75t_R FILLER_39_602 ();
 DECAPx4_ASAP7_75t_R FILLER_39_626 ();
 DECAPx2_ASAP7_75t_R FILLER_39_639 ();
 FILLER_ASAP7_75t_R FILLER_39_645 ();
 DECAPx4_ASAP7_75t_R FILLER_39_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_688 ();
 DECAPx2_ASAP7_75t_R FILLER_39_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_698 ();
 DECAPx2_ASAP7_75t_R FILLER_39_702 ();
 FILLER_ASAP7_75t_R FILLER_39_708 ();
 DECAPx2_ASAP7_75t_R FILLER_39_713 ();
 FILLER_ASAP7_75t_R FILLER_39_719 ();
 DECAPx1_ASAP7_75t_R FILLER_39_738 ();
 FILLER_ASAP7_75t_R FILLER_39_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_750 ();
 DECAPx2_ASAP7_75t_R FILLER_39_754 ();
 FILLER_ASAP7_75t_R FILLER_39_760 ();
 DECAPx2_ASAP7_75t_R FILLER_39_768 ();
 FILLER_ASAP7_75t_R FILLER_39_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_776 ();
 DECAPx2_ASAP7_75t_R FILLER_39_800 ();
 DECAPx10_ASAP7_75t_R FILLER_39_835 ();
 DECAPx10_ASAP7_75t_R FILLER_39_857 ();
 DECAPx10_ASAP7_75t_R FILLER_39_879 ();
 DECAPx6_ASAP7_75t_R FILLER_39_901 ();
 DECAPx2_ASAP7_75t_R FILLER_39_918 ();
 DECAPx6_ASAP7_75t_R FILLER_39_926 ();
 FILLER_ASAP7_75t_R FILLER_39_940 ();
 DECAPx2_ASAP7_75t_R FILLER_39_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_972 ();
 DECAPx10_ASAP7_75t_R FILLER_39_990 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1386 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx10_ASAP7_75t_R FILLER_40_24 ();
 DECAPx10_ASAP7_75t_R FILLER_40_46 ();
 DECAPx10_ASAP7_75t_R FILLER_40_68 ();
 DECAPx10_ASAP7_75t_R FILLER_40_90 ();
 DECAPx10_ASAP7_75t_R FILLER_40_112 ();
 DECAPx10_ASAP7_75t_R FILLER_40_134 ();
 DECAPx10_ASAP7_75t_R FILLER_40_156 ();
 DECAPx10_ASAP7_75t_R FILLER_40_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_230 ();
 DECAPx2_ASAP7_75t_R FILLER_40_264 ();
 FILLER_ASAP7_75t_R FILLER_40_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_272 ();
 DECAPx2_ASAP7_75t_R FILLER_40_276 ();
 DECAPx4_ASAP7_75t_R FILLER_40_285 ();
 FILLER_ASAP7_75t_R FILLER_40_295 ();
 FILLER_ASAP7_75t_R FILLER_40_323 ();
 DECAPx1_ASAP7_75t_R FILLER_40_337 ();
 FILLER_ASAP7_75t_R FILLER_40_367 ();
 DECAPx4_ASAP7_75t_R FILLER_40_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_411 ();
 DECAPx1_ASAP7_75t_R FILLER_40_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_422 ();
 DECAPx2_ASAP7_75t_R FILLER_40_426 ();
 FILLER_ASAP7_75t_R FILLER_40_432 ();
 FILLER_ASAP7_75t_R FILLER_40_460 ();
 DECAPx2_ASAP7_75t_R FILLER_40_467 ();
 DECAPx2_ASAP7_75t_R FILLER_40_499 ();
 FILLER_ASAP7_75t_R FILLER_40_505 ();
 DECAPx4_ASAP7_75t_R FILLER_40_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_523 ();
 DECAPx10_ASAP7_75t_R FILLER_40_556 ();
 DECAPx10_ASAP7_75t_R FILLER_40_578 ();
 DECAPx10_ASAP7_75t_R FILLER_40_600 ();
 DECAPx2_ASAP7_75t_R FILLER_40_625 ();
 FILLER_ASAP7_75t_R FILLER_40_631 ();
 DECAPx6_ASAP7_75t_R FILLER_40_639 ();
 DECAPx2_ASAP7_75t_R FILLER_40_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_659 ();
 FILLER_ASAP7_75t_R FILLER_40_663 ();
 DECAPx2_ASAP7_75t_R FILLER_40_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_674 ();
 DECAPx2_ASAP7_75t_R FILLER_40_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_722 ();
 DECAPx2_ASAP7_75t_R FILLER_40_726 ();
 DECAPx2_ASAP7_75t_R FILLER_40_780 ();
 FILLER_ASAP7_75t_R FILLER_40_786 ();
 FILLER_ASAP7_75t_R FILLER_40_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_820 ();
 DECAPx6_ASAP7_75t_R FILLER_40_852 ();
 FILLER_ASAP7_75t_R FILLER_40_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_868 ();
 FILLER_ASAP7_75t_R FILLER_40_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_889 ();
 DECAPx2_ASAP7_75t_R FILLER_40_899 ();
 FILLER_ASAP7_75t_R FILLER_40_905 ();
 DECAPx2_ASAP7_75t_R FILLER_40_925 ();
 DECAPx1_ASAP7_75t_R FILLER_40_940 ();
 DECAPx6_ASAP7_75t_R FILLER_40_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_967 ();
 DECAPx10_ASAP7_75t_R FILLER_40_985 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1388 ();
 FILLER_ASAP7_75t_R FILLER_40_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_24 ();
 DECAPx10_ASAP7_75t_R FILLER_41_46 ();
 DECAPx10_ASAP7_75t_R FILLER_41_68 ();
 DECAPx10_ASAP7_75t_R FILLER_41_90 ();
 DECAPx10_ASAP7_75t_R FILLER_41_112 ();
 DECAPx10_ASAP7_75t_R FILLER_41_134 ();
 DECAPx10_ASAP7_75t_R FILLER_41_156 ();
 DECAPx2_ASAP7_75t_R FILLER_41_178 ();
 FILLER_ASAP7_75t_R FILLER_41_184 ();
 DECAPx4_ASAP7_75t_R FILLER_41_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_222 ();
 DECAPx4_ASAP7_75t_R FILLER_41_255 ();
 FILLER_ASAP7_75t_R FILLER_41_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_306 ();
 DECAPx1_ASAP7_75t_R FILLER_41_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_349 ();
 DECAPx1_ASAP7_75t_R FILLER_41_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_366 ();
 DECAPx1_ASAP7_75t_R FILLER_41_399 ();
 FILLER_ASAP7_75t_R FILLER_41_435 ();
 DECAPx2_ASAP7_75t_R FILLER_41_443 ();
 DECAPx6_ASAP7_75t_R FILLER_41_475 ();
 FILLER_ASAP7_75t_R FILLER_41_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_491 ();
 FILLER_ASAP7_75t_R FILLER_41_518 ();
 DECAPx10_ASAP7_75t_R FILLER_41_555 ();
 DECAPx6_ASAP7_75t_R FILLER_41_577 ();
 DECAPx1_ASAP7_75t_R FILLER_41_591 ();
 DECAPx4_ASAP7_75t_R FILLER_41_605 ();
 DECAPx2_ASAP7_75t_R FILLER_41_624 ();
 FILLER_ASAP7_75t_R FILLER_41_630 ();
 DECAPx4_ASAP7_75t_R FILLER_41_647 ();
 FILLER_ASAP7_75t_R FILLER_41_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_662 ();
 DECAPx4_ASAP7_75t_R FILLER_41_675 ();
 FILLER_ASAP7_75t_R FILLER_41_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_702 ();
 DECAPx4_ASAP7_75t_R FILLER_41_726 ();
 FILLER_ASAP7_75t_R FILLER_41_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_741 ();
 DECAPx6_ASAP7_75t_R FILLER_41_748 ();
 DECAPx2_ASAP7_75t_R FILLER_41_762 ();
 DECAPx1_ASAP7_75t_R FILLER_41_785 ();
 FILLER_ASAP7_75t_R FILLER_41_834 ();
 DECAPx4_ASAP7_75t_R FILLER_41_845 ();
 FILLER_ASAP7_75t_R FILLER_41_855 ();
 DECAPx2_ASAP7_75t_R FILLER_41_872 ();
 DECAPx6_ASAP7_75t_R FILLER_41_890 ();
 FILLER_ASAP7_75t_R FILLER_41_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_923 ();
 FILLER_ASAP7_75t_R FILLER_41_926 ();
 DECAPx1_ASAP7_75t_R FILLER_41_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_939 ();
 DECAPx6_ASAP7_75t_R FILLER_41_947 ();
 DECAPx2_ASAP7_75t_R FILLER_41_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_967 ();
 DECAPx10_ASAP7_75t_R FILLER_41_982 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1356 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx10_ASAP7_75t_R FILLER_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_42_68 ();
 DECAPx10_ASAP7_75t_R FILLER_42_90 ();
 DECAPx10_ASAP7_75t_R FILLER_42_112 ();
 DECAPx10_ASAP7_75t_R FILLER_42_134 ();
 DECAPx6_ASAP7_75t_R FILLER_42_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_170 ();
 FILLER_ASAP7_75t_R FILLER_42_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_199 ();
 DECAPx1_ASAP7_75t_R FILLER_42_203 ();
 DECAPx10_ASAP7_75t_R FILLER_42_213 ();
 FILLER_ASAP7_75t_R FILLER_42_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_241 ();
 DECAPx2_ASAP7_75t_R FILLER_42_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_277 ();
 DECAPx2_ASAP7_75t_R FILLER_42_281 ();
 DECAPx10_ASAP7_75t_R FILLER_42_293 ();
 DECAPx2_ASAP7_75t_R FILLER_42_315 ();
 DECAPx2_ASAP7_75t_R FILLER_42_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_333 ();
 DECAPx6_ASAP7_75t_R FILLER_42_337 ();
 FILLER_ASAP7_75t_R FILLER_42_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_353 ();
 DECAPx1_ASAP7_75t_R FILLER_42_380 ();
 DECAPx4_ASAP7_75t_R FILLER_42_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_426 ();
 FILLER_ASAP7_75t_R FILLER_42_433 ();
 DECAPx4_ASAP7_75t_R FILLER_42_443 ();
 FILLER_ASAP7_75t_R FILLER_42_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_461 ();
 DECAPx1_ASAP7_75t_R FILLER_42_472 ();
 DECAPx2_ASAP7_75t_R FILLER_42_482 ();
 FILLER_ASAP7_75t_R FILLER_42_491 ();
 DECAPx1_ASAP7_75t_R FILLER_42_503 ();
 DECAPx1_ASAP7_75t_R FILLER_42_513 ();
 DECAPx2_ASAP7_75t_R FILLER_42_520 ();
 FILLER_ASAP7_75t_R FILLER_42_529 ();
 DECAPx1_ASAP7_75t_R FILLER_42_537 ();
 DECAPx4_ASAP7_75t_R FILLER_42_544 ();
 FILLER_ASAP7_75t_R FILLER_42_554 ();
 FILLER_ASAP7_75t_R FILLER_42_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_564 ();
 DECAPx6_ASAP7_75t_R FILLER_42_568 ();
 DECAPx2_ASAP7_75t_R FILLER_42_582 ();
 DECAPx1_ASAP7_75t_R FILLER_42_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_608 ();
 DECAPx6_ASAP7_75t_R FILLER_42_649 ();
 DECAPx2_ASAP7_75t_R FILLER_42_683 ();
 FILLER_ASAP7_75t_R FILLER_42_689 ();
 DECAPx6_ASAP7_75t_R FILLER_42_697 ();
 FILLER_ASAP7_75t_R FILLER_42_711 ();
 DECAPx1_ASAP7_75t_R FILLER_42_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_723 ();
 DECAPx2_ASAP7_75t_R FILLER_42_738 ();
 DECAPx2_ASAP7_75t_R FILLER_42_761 ();
 FILLER_ASAP7_75t_R FILLER_42_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_769 ();
 DECAPx6_ASAP7_75t_R FILLER_42_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_799 ();
 DECAPx2_ASAP7_75t_R FILLER_42_816 ();
 FILLER_ASAP7_75t_R FILLER_42_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_876 ();
 DECAPx1_ASAP7_75t_R FILLER_42_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_908 ();
 DECAPx1_ASAP7_75t_R FILLER_42_942 ();
 DECAPx10_ASAP7_75t_R FILLER_42_978 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1352 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1374 ();
 FILLER_ASAP7_75t_R FILLER_42_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_42_1388 ();
 FILLER_ASAP7_75t_R FILLER_42_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx10_ASAP7_75t_R FILLER_43_24 ();
 DECAPx10_ASAP7_75t_R FILLER_43_46 ();
 DECAPx10_ASAP7_75t_R FILLER_43_68 ();
 DECAPx10_ASAP7_75t_R FILLER_43_90 ();
 DECAPx10_ASAP7_75t_R FILLER_43_112 ();
 DECAPx2_ASAP7_75t_R FILLER_43_134 ();
 FILLER_ASAP7_75t_R FILLER_43_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_142 ();
 FILLER_ASAP7_75t_R FILLER_43_169 ();
 DECAPx2_ASAP7_75t_R FILLER_43_177 ();
 FILLER_ASAP7_75t_R FILLER_43_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_185 ();
 DECAPx1_ASAP7_75t_R FILLER_43_189 ();
 DECAPx2_ASAP7_75t_R FILLER_43_199 ();
 DECAPx4_ASAP7_75t_R FILLER_43_231 ();
 FILLER_ASAP7_75t_R FILLER_43_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_243 ();
 FILLER_ASAP7_75t_R FILLER_43_250 ();
 DECAPx1_ASAP7_75t_R FILLER_43_290 ();
 DECAPx6_ASAP7_75t_R FILLER_43_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_334 ();
 DECAPx2_ASAP7_75t_R FILLER_43_348 ();
 FILLER_ASAP7_75t_R FILLER_43_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_356 ();
 DECAPx2_ASAP7_75t_R FILLER_43_363 ();
 FILLER_ASAP7_75t_R FILLER_43_372 ();
 DECAPx2_ASAP7_75t_R FILLER_43_380 ();
 FILLER_ASAP7_75t_R FILLER_43_386 ();
 DECAPx2_ASAP7_75t_R FILLER_43_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_407 ();
 DECAPx2_ASAP7_75t_R FILLER_43_419 ();
 DECAPx1_ASAP7_75t_R FILLER_43_451 ();
 FILLER_ASAP7_75t_R FILLER_43_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_463 ();
 DECAPx4_ASAP7_75t_R FILLER_43_467 ();
 DECAPx4_ASAP7_75t_R FILLER_43_483 ();
 FILLER_ASAP7_75t_R FILLER_43_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_495 ();
 DECAPx6_ASAP7_75t_R FILLER_43_499 ();
 DECAPx1_ASAP7_75t_R FILLER_43_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_517 ();
 DECAPx10_ASAP7_75t_R FILLER_43_524 ();
 DECAPx1_ASAP7_75t_R FILLER_43_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_576 ();
 DECAPx10_ASAP7_75t_R FILLER_43_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_613 ();
 DECAPx2_ASAP7_75t_R FILLER_43_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_642 ();
 DECAPx2_ASAP7_75t_R FILLER_43_649 ();
 DECAPx2_ASAP7_75t_R FILLER_43_658 ();
 DECAPx4_ASAP7_75t_R FILLER_43_667 ();
 FILLER_ASAP7_75t_R FILLER_43_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_679 ();
 FILLER_ASAP7_75t_R FILLER_43_690 ();
 DECAPx6_ASAP7_75t_R FILLER_43_702 ();
 FILLER_ASAP7_75t_R FILLER_43_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_718 ();
 DECAPx2_ASAP7_75t_R FILLER_43_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_742 ();
 DECAPx2_ASAP7_75t_R FILLER_43_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_763 ();
 FILLER_ASAP7_75t_R FILLER_43_770 ();
 DECAPx2_ASAP7_75t_R FILLER_43_786 ();
 FILLER_ASAP7_75t_R FILLER_43_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_794 ();
 DECAPx2_ASAP7_75t_R FILLER_43_801 ();
 FILLER_ASAP7_75t_R FILLER_43_807 ();
 DECAPx10_ASAP7_75t_R FILLER_43_819 ();
 DECAPx2_ASAP7_75t_R FILLER_43_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_847 ();
 FILLER_ASAP7_75t_R FILLER_43_904 ();
 DECAPx2_ASAP7_75t_R FILLER_43_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_934 ();
 DECAPx1_ASAP7_75t_R FILLER_43_947 ();
 DECAPx1_ASAP7_75t_R FILLER_43_959 ();
 DECAPx10_ASAP7_75t_R FILLER_43_979 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1397 ();
 FILLER_ASAP7_75t_R FILLER_43_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_44_24 ();
 DECAPx10_ASAP7_75t_R FILLER_44_46 ();
 DECAPx10_ASAP7_75t_R FILLER_44_68 ();
 DECAPx10_ASAP7_75t_R FILLER_44_90 ();
 DECAPx10_ASAP7_75t_R FILLER_44_112 ();
 DECAPx6_ASAP7_75t_R FILLER_44_134 ();
 FILLER_ASAP7_75t_R FILLER_44_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_150 ();
 FILLER_ASAP7_75t_R FILLER_44_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_199 ();
 DECAPx10_ASAP7_75t_R FILLER_44_236 ();
 DECAPx2_ASAP7_75t_R FILLER_44_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_264 ();
 DECAPx4_ASAP7_75t_R FILLER_44_271 ();
 FILLER_ASAP7_75t_R FILLER_44_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_283 ();
 DECAPx4_ASAP7_75t_R FILLER_44_293 ();
 FILLER_ASAP7_75t_R FILLER_44_303 ();
 DECAPx4_ASAP7_75t_R FILLER_44_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_331 ();
 DECAPx2_ASAP7_75t_R FILLER_44_358 ();
 FILLER_ASAP7_75t_R FILLER_44_364 ();
 DECAPx10_ASAP7_75t_R FILLER_44_373 ();
 DECAPx6_ASAP7_75t_R FILLER_44_395 ();
 DECAPx1_ASAP7_75t_R FILLER_44_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_413 ();
 DECAPx2_ASAP7_75t_R FILLER_44_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_427 ();
 DECAPx1_ASAP7_75t_R FILLER_44_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_438 ();
 FILLER_ASAP7_75t_R FILLER_44_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_448 ();
 DECAPx2_ASAP7_75t_R FILLER_44_456 ();
 DECAPx6_ASAP7_75t_R FILLER_44_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_508 ();
 FILLER_ASAP7_75t_R FILLER_44_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_543 ();
 FILLER_ASAP7_75t_R FILLER_44_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_560 ();
 DECAPx10_ASAP7_75t_R FILLER_44_577 ();
 DECAPx4_ASAP7_75t_R FILLER_44_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_609 ();
 DECAPx6_ASAP7_75t_R FILLER_44_628 ();
 DECAPx10_ASAP7_75t_R FILLER_44_670 ();
 FILLER_ASAP7_75t_R FILLER_44_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_694 ();
 FILLER_ASAP7_75t_R FILLER_44_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_711 ();
 DECAPx2_ASAP7_75t_R FILLER_44_715 ();
 FILLER_ASAP7_75t_R FILLER_44_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_723 ();
 DECAPx4_ASAP7_75t_R FILLER_44_741 ();
 FILLER_ASAP7_75t_R FILLER_44_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_759 ();
 DECAPx10_ASAP7_75t_R FILLER_44_792 ();
 DECAPx10_ASAP7_75t_R FILLER_44_814 ();
 DECAPx6_ASAP7_75t_R FILLER_44_836 ();
 DECAPx1_ASAP7_75t_R FILLER_44_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_873 ();
 FILLER_ASAP7_75t_R FILLER_44_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_883 ();
 DECAPx1_ASAP7_75t_R FILLER_44_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_894 ();
 DECAPx10_ASAP7_75t_R FILLER_44_902 ();
 DECAPx10_ASAP7_75t_R FILLER_44_924 ();
 DECAPx2_ASAP7_75t_R FILLER_44_946 ();
 FILLER_ASAP7_75t_R FILLER_44_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_954 ();
 DECAPx4_ASAP7_75t_R FILLER_44_958 ();
 DECAPx10_ASAP7_75t_R FILLER_44_976 ();
 DECAPx10_ASAP7_75t_R FILLER_44_998 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1372 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1388 ();
 FILLER_ASAP7_75t_R FILLER_44_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_45_24 ();
 DECAPx10_ASAP7_75t_R FILLER_45_46 ();
 DECAPx10_ASAP7_75t_R FILLER_45_68 ();
 DECAPx10_ASAP7_75t_R FILLER_45_90 ();
 DECAPx4_ASAP7_75t_R FILLER_45_112 ();
 FILLER_ASAP7_75t_R FILLER_45_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_124 ();
 FILLER_ASAP7_75t_R FILLER_45_220 ();
 FILLER_ASAP7_75t_R FILLER_45_225 ();
 DECAPx1_ASAP7_75t_R FILLER_45_253 ();
 DECAPx10_ASAP7_75t_R FILLER_45_260 ();
 DECAPx10_ASAP7_75t_R FILLER_45_282 ();
 DECAPx1_ASAP7_75t_R FILLER_45_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_308 ();
 DECAPx10_ASAP7_75t_R FILLER_45_316 ();
 DECAPx2_ASAP7_75t_R FILLER_45_338 ();
 FILLER_ASAP7_75t_R FILLER_45_344 ();
 DECAPx4_ASAP7_75t_R FILLER_45_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_359 ();
 DECAPx4_ASAP7_75t_R FILLER_45_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_448 ();
 DECAPx2_ASAP7_75t_R FILLER_45_478 ();
 DECAPx1_ASAP7_75t_R FILLER_45_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_495 ();
 FILLER_ASAP7_75t_R FILLER_45_522 ();
 DECAPx2_ASAP7_75t_R FILLER_45_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_562 ();
 DECAPx4_ASAP7_75t_R FILLER_45_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_583 ();
 DECAPx4_ASAP7_75t_R FILLER_45_598 ();
 FILLER_ASAP7_75t_R FILLER_45_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_630 ();
 DECAPx2_ASAP7_75t_R FILLER_45_637 ();
 DECAPx2_ASAP7_75t_R FILLER_45_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_663 ();
 DECAPx2_ASAP7_75t_R FILLER_45_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_696 ();
 FILLER_ASAP7_75t_R FILLER_45_720 ();
 DECAPx4_ASAP7_75t_R FILLER_45_739 ();
 FILLER_ASAP7_75t_R FILLER_45_749 ();
 DECAPx6_ASAP7_75t_R FILLER_45_760 ();
 DECAPx4_ASAP7_75t_R FILLER_45_788 ();
 FILLER_ASAP7_75t_R FILLER_45_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_800 ();
 DECAPx2_ASAP7_75t_R FILLER_45_816 ();
 FILLER_ASAP7_75t_R FILLER_45_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_861 ();
 DECAPx6_ASAP7_75t_R FILLER_45_869 ();
 DECAPx10_ASAP7_75t_R FILLER_45_889 ();
 DECAPx4_ASAP7_75t_R FILLER_45_911 ();
 FILLER_ASAP7_75t_R FILLER_45_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_923 ();
 DECAPx1_ASAP7_75t_R FILLER_45_941 ();
 FILLER_ASAP7_75t_R FILLER_45_952 ();
 FILLER_ASAP7_75t_R FILLER_45_980 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_46_24 ();
 DECAPx10_ASAP7_75t_R FILLER_46_46 ();
 DECAPx10_ASAP7_75t_R FILLER_46_68 ();
 DECAPx10_ASAP7_75t_R FILLER_46_90 ();
 DECAPx6_ASAP7_75t_R FILLER_46_112 ();
 DECAPx2_ASAP7_75t_R FILLER_46_126 ();
 DECAPx10_ASAP7_75t_R FILLER_46_148 ();
 FILLER_ASAP7_75t_R FILLER_46_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_172 ();
 DECAPx6_ASAP7_75t_R FILLER_46_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_190 ();
 DECAPx10_ASAP7_75t_R FILLER_46_200 ();
 DECAPx2_ASAP7_75t_R FILLER_46_222 ();
 FILLER_ASAP7_75t_R FILLER_46_228 ();
 FILLER_ASAP7_75t_R FILLER_46_237 ();
 DECAPx10_ASAP7_75t_R FILLER_46_268 ();
 DECAPx2_ASAP7_75t_R FILLER_46_290 ();
 FILLER_ASAP7_75t_R FILLER_46_296 ();
 DECAPx10_ASAP7_75t_R FILLER_46_330 ();
 DECAPx6_ASAP7_75t_R FILLER_46_352 ();
 FILLER_ASAP7_75t_R FILLER_46_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_368 ();
 FILLER_ASAP7_75t_R FILLER_46_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_377 ();
 DECAPx1_ASAP7_75t_R FILLER_46_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_385 ();
 FILLER_ASAP7_75t_R FILLER_46_399 ();
 DECAPx4_ASAP7_75t_R FILLER_46_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_414 ();
 DECAPx2_ASAP7_75t_R FILLER_46_421 ();
 DECAPx6_ASAP7_75t_R FILLER_46_430 ();
 DECAPx2_ASAP7_75t_R FILLER_46_444 ();
 DECAPx2_ASAP7_75t_R FILLER_46_456 ();
 FILLER_ASAP7_75t_R FILLER_46_464 ();
 DECAPx2_ASAP7_75t_R FILLER_46_473 ();
 DECAPx2_ASAP7_75t_R FILLER_46_482 ();
 DECAPx1_ASAP7_75t_R FILLER_46_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_498 ();
 DECAPx1_ASAP7_75t_R FILLER_46_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_519 ();
 FILLER_ASAP7_75t_R FILLER_46_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_531 ();
 FILLER_ASAP7_75t_R FILLER_46_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_546 ();
 DECAPx10_ASAP7_75t_R FILLER_46_559 ();
 DECAPx2_ASAP7_75t_R FILLER_46_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_587 ();
 DECAPx1_ASAP7_75t_R FILLER_46_610 ();
 FILLER_ASAP7_75t_R FILLER_46_620 ();
 DECAPx1_ASAP7_75t_R FILLER_46_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_652 ();
 FILLER_ASAP7_75t_R FILLER_46_679 ();
 DECAPx1_ASAP7_75t_R FILLER_46_698 ();
 DECAPx6_ASAP7_75t_R FILLER_46_719 ();
 DECAPx2_ASAP7_75t_R FILLER_46_733 ();
 DECAPx10_ASAP7_75t_R FILLER_46_753 ();
 DECAPx2_ASAP7_75t_R FILLER_46_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_800 ();
 DECAPx10_ASAP7_75t_R FILLER_46_867 ();
 DECAPx1_ASAP7_75t_R FILLER_46_889 ();
 DECAPx2_ASAP7_75t_R FILLER_46_903 ();
 FILLER_ASAP7_75t_R FILLER_46_927 ();
 FILLER_ASAP7_75t_R FILLER_46_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_993 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1388 ();
 FILLER_ASAP7_75t_R FILLER_46_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx10_ASAP7_75t_R FILLER_47_24 ();
 DECAPx10_ASAP7_75t_R FILLER_47_46 ();
 DECAPx10_ASAP7_75t_R FILLER_47_68 ();
 DECAPx10_ASAP7_75t_R FILLER_47_90 ();
 DECAPx10_ASAP7_75t_R FILLER_47_112 ();
 DECAPx6_ASAP7_75t_R FILLER_47_134 ();
 DECAPx2_ASAP7_75t_R FILLER_47_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_154 ();
 DECAPx10_ASAP7_75t_R FILLER_47_181 ();
 DECAPx4_ASAP7_75t_R FILLER_47_203 ();
 FILLER_ASAP7_75t_R FILLER_47_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_215 ();
 DECAPx1_ASAP7_75t_R FILLER_47_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_227 ();
 FILLER_ASAP7_75t_R FILLER_47_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_233 ();
 DECAPx10_ASAP7_75t_R FILLER_47_240 ();
 DECAPx1_ASAP7_75t_R FILLER_47_262 ();
 DECAPx2_ASAP7_75t_R FILLER_47_279 ();
 FILLER_ASAP7_75t_R FILLER_47_285 ();
 DECAPx6_ASAP7_75t_R FILLER_47_293 ();
 DECAPx1_ASAP7_75t_R FILLER_47_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_311 ();
 DECAPx10_ASAP7_75t_R FILLER_47_315 ();
 DECAPx2_ASAP7_75t_R FILLER_47_337 ();
 FILLER_ASAP7_75t_R FILLER_47_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_345 ();
 DECAPx2_ASAP7_75t_R FILLER_47_352 ();
 FILLER_ASAP7_75t_R FILLER_47_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_360 ();
 DECAPx10_ASAP7_75t_R FILLER_47_367 ();
 FILLER_ASAP7_75t_R FILLER_47_389 ();
 DECAPx6_ASAP7_75t_R FILLER_47_407 ();
 DECAPx1_ASAP7_75t_R FILLER_47_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_451 ();
 DECAPx4_ASAP7_75t_R FILLER_47_455 ();
 DECAPx2_ASAP7_75t_R FILLER_47_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_497 ();
 DECAPx6_ASAP7_75t_R FILLER_47_501 ();
 DECAPx1_ASAP7_75t_R FILLER_47_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_519 ();
 DECAPx1_ASAP7_75t_R FILLER_47_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_558 ();
 DECAPx1_ASAP7_75t_R FILLER_47_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_573 ();
 DECAPx10_ASAP7_75t_R FILLER_47_577 ();
 DECAPx6_ASAP7_75t_R FILLER_47_599 ();
 FILLER_ASAP7_75t_R FILLER_47_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_634 ();
 DECAPx2_ASAP7_75t_R FILLER_47_644 ();
 FILLER_ASAP7_75t_R FILLER_47_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_652 ();
 DECAPx1_ASAP7_75t_R FILLER_47_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_675 ();
 FILLER_ASAP7_75t_R FILLER_47_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_681 ();
 DECAPx6_ASAP7_75t_R FILLER_47_699 ();
 FILLER_ASAP7_75t_R FILLER_47_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_715 ();
 DECAPx6_ASAP7_75t_R FILLER_47_725 ();
 FILLER_ASAP7_75t_R FILLER_47_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_741 ();
 DECAPx10_ASAP7_75t_R FILLER_47_757 ();
 DECAPx1_ASAP7_75t_R FILLER_47_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_783 ();
 DECAPx1_ASAP7_75t_R FILLER_47_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_808 ();
 DECAPx1_ASAP7_75t_R FILLER_47_823 ();
 DECAPx10_ASAP7_75t_R FILLER_47_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_869 ();
 DECAPx2_ASAP7_75t_R FILLER_47_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_884 ();
 DECAPx6_ASAP7_75t_R FILLER_47_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_923 ();
 DECAPx4_ASAP7_75t_R FILLER_47_926 ();
 DECAPx1_ASAP7_75t_R FILLER_47_948 ();
 FILLER_ASAP7_75t_R FILLER_47_967 ();
 DECAPx2_ASAP7_75t_R FILLER_47_972 ();
 FILLER_ASAP7_75t_R FILLER_47_978 ();
 FILLER_ASAP7_75t_R FILLER_47_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_985 ();
 FILLER_ASAP7_75t_R FILLER_47_994 ();
 DECAPx1_ASAP7_75t_R FILLER_47_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1351 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1373 ();
 DECAPx4_ASAP7_75t_R FILLER_47_1395 ();
 DECAPx10_ASAP7_75t_R FILLER_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_48_68 ();
 DECAPx10_ASAP7_75t_R FILLER_48_90 ();
 DECAPx2_ASAP7_75t_R FILLER_48_112 ();
 DECAPx4_ASAP7_75t_R FILLER_48_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_168 ();
 FILLER_ASAP7_75t_R FILLER_48_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_174 ();
 FILLER_ASAP7_75t_R FILLER_48_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_203 ();
 DECAPx2_ASAP7_75t_R FILLER_48_207 ();
 DECAPx10_ASAP7_75t_R FILLER_48_239 ();
 DECAPx1_ASAP7_75t_R FILLER_48_261 ();
 DECAPx6_ASAP7_75t_R FILLER_48_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_287 ();
 DECAPx10_ASAP7_75t_R FILLER_48_296 ();
 DECAPx4_ASAP7_75t_R FILLER_48_318 ();
 DECAPx2_ASAP7_75t_R FILLER_48_334 ();
 FILLER_ASAP7_75t_R FILLER_48_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_342 ();
 DECAPx1_ASAP7_75t_R FILLER_48_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_355 ();
 DECAPx2_ASAP7_75t_R FILLER_48_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_388 ();
 FILLER_ASAP7_75t_R FILLER_48_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_417 ();
 DECAPx1_ASAP7_75t_R FILLER_48_421 ();
 DECAPx1_ASAP7_75t_R FILLER_48_432 ();
 FILLER_ASAP7_75t_R FILLER_48_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_466 ();
 DECAPx1_ASAP7_75t_R FILLER_48_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_477 ();
 DECAPx6_ASAP7_75t_R FILLER_48_514 ();
 DECAPx1_ASAP7_75t_R FILLER_48_528 ();
 DECAPx10_ASAP7_75t_R FILLER_48_588 ();
 DECAPx6_ASAP7_75t_R FILLER_48_610 ();
 FILLER_ASAP7_75t_R FILLER_48_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_626 ();
 DECAPx2_ASAP7_75t_R FILLER_48_630 ();
 DECAPx1_ASAP7_75t_R FILLER_48_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_668 ();
 DECAPx6_ASAP7_75t_R FILLER_48_672 ();
 DECAPx1_ASAP7_75t_R FILLER_48_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_693 ();
 DECAPx6_ASAP7_75t_R FILLER_48_702 ();
 FILLER_ASAP7_75t_R FILLER_48_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_733 ();
 FILLER_ASAP7_75t_R FILLER_48_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_763 ();
 DECAPx10_ASAP7_75t_R FILLER_48_778 ();
 DECAPx1_ASAP7_75t_R FILLER_48_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_804 ();
 DECAPx6_ASAP7_75t_R FILLER_48_811 ();
 DECAPx1_ASAP7_75t_R FILLER_48_825 ();
 FILLER_ASAP7_75t_R FILLER_48_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_843 ();
 DECAPx2_ASAP7_75t_R FILLER_48_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_878 ();
 DECAPx2_ASAP7_75t_R FILLER_48_887 ();
 FILLER_ASAP7_75t_R FILLER_48_893 ();
 DECAPx6_ASAP7_75t_R FILLER_48_903 ();
 FILLER_ASAP7_75t_R FILLER_48_917 ();
 DECAPx2_ASAP7_75t_R FILLER_48_929 ();
 FILLER_ASAP7_75t_R FILLER_48_935 ();
 DECAPx4_ASAP7_75t_R FILLER_48_940 ();
 FILLER_ASAP7_75t_R FILLER_48_950 ();
 DECAPx10_ASAP7_75t_R FILLER_48_958 ();
 DECAPx10_ASAP7_75t_R FILLER_48_980 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1049 ();
 FILLER_ASAP7_75t_R FILLER_48_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1382 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1388 ();
 FILLER_ASAP7_75t_R FILLER_48_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_49_68 ();
 DECAPx6_ASAP7_75t_R FILLER_49_90 ();
 DECAPx1_ASAP7_75t_R FILLER_49_107 ();
 FILLER_ASAP7_75t_R FILLER_49_144 ();
 DECAPx1_ASAP7_75t_R FILLER_49_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_221 ();
 FILLER_ASAP7_75t_R FILLER_49_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_262 ();
 DECAPx10_ASAP7_75t_R FILLER_49_269 ();
 DECAPx2_ASAP7_75t_R FILLER_49_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_297 ();
 DECAPx2_ASAP7_75t_R FILLER_49_304 ();
 FILLER_ASAP7_75t_R FILLER_49_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_327 ();
 DECAPx10_ASAP7_75t_R FILLER_49_334 ();
 FILLER_ASAP7_75t_R FILLER_49_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_358 ();
 FILLER_ASAP7_75t_R FILLER_49_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_375 ();
 DECAPx2_ASAP7_75t_R FILLER_49_389 ();
 FILLER_ASAP7_75t_R FILLER_49_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_436 ();
 DECAPx2_ASAP7_75t_R FILLER_49_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_482 ();
 DECAPx10_ASAP7_75t_R FILLER_49_489 ();
 DECAPx4_ASAP7_75t_R FILLER_49_511 ();
 FILLER_ASAP7_75t_R FILLER_49_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_538 ();
 FILLER_ASAP7_75t_R FILLER_49_542 ();
 DECAPx2_ASAP7_75t_R FILLER_49_570 ();
 FILLER_ASAP7_75t_R FILLER_49_576 ();
 DECAPx1_ASAP7_75t_R FILLER_49_586 ();
 DECAPx6_ASAP7_75t_R FILLER_49_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_616 ();
 DECAPx4_ASAP7_75t_R FILLER_49_626 ();
 FILLER_ASAP7_75t_R FILLER_49_636 ();
 DECAPx2_ASAP7_75t_R FILLER_49_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_664 ();
 FILLER_ASAP7_75t_R FILLER_49_682 ();
 FILLER_ASAP7_75t_R FILLER_49_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_689 ();
 DECAPx2_ASAP7_75t_R FILLER_49_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_731 ();
 DECAPx6_ASAP7_75t_R FILLER_49_744 ();
 DECAPx1_ASAP7_75t_R FILLER_49_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_762 ();
 FILLER_ASAP7_75t_R FILLER_49_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_777 ();
 DECAPx4_ASAP7_75t_R FILLER_49_787 ();
 DECAPx1_ASAP7_75t_R FILLER_49_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_807 ();
 DECAPx10_ASAP7_75t_R FILLER_49_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_842 ();
 DECAPx4_ASAP7_75t_R FILLER_49_849 ();
 FILLER_ASAP7_75t_R FILLER_49_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_878 ();
 DECAPx1_ASAP7_75t_R FILLER_49_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_897 ();
 DECAPx1_ASAP7_75t_R FILLER_49_906 ();
 DECAPx1_ASAP7_75t_R FILLER_49_920 ();
 DECAPx2_ASAP7_75t_R FILLER_49_952 ();
 FILLER_ASAP7_75t_R FILLER_49_958 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1015 ();
 FILLER_ASAP7_75t_R FILLER_49_1025 ();
 FILLER_ASAP7_75t_R FILLER_49_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1130 ();
 FILLER_ASAP7_75t_R FILLER_49_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1388 ();
 FILLER_ASAP7_75t_R FILLER_49_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_50_68 ();
 DECAPx2_ASAP7_75t_R FILLER_50_116 ();
 FILLER_ASAP7_75t_R FILLER_50_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_138 ();
 DECAPx1_ASAP7_75t_R FILLER_50_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_155 ();
 DECAPx1_ASAP7_75t_R FILLER_50_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_166 ();
 DECAPx6_ASAP7_75t_R FILLER_50_170 ();
 FILLER_ASAP7_75t_R FILLER_50_200 ();
 DECAPx2_ASAP7_75t_R FILLER_50_228 ();
 FILLER_ASAP7_75t_R FILLER_50_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_244 ();
 DECAPx10_ASAP7_75t_R FILLER_50_248 ();
 DECAPx10_ASAP7_75t_R FILLER_50_270 ();
 DECAPx10_ASAP7_75t_R FILLER_50_292 ();
 DECAPx10_ASAP7_75t_R FILLER_50_314 ();
 DECAPx10_ASAP7_75t_R FILLER_50_336 ();
 FILLER_ASAP7_75t_R FILLER_50_358 ();
 FILLER_ASAP7_75t_R FILLER_50_366 ();
 DECAPx2_ASAP7_75t_R FILLER_50_394 ();
 FILLER_ASAP7_75t_R FILLER_50_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_402 ();
 DECAPx10_ASAP7_75t_R FILLER_50_409 ();
 DECAPx2_ASAP7_75t_R FILLER_50_431 ();
 FILLER_ASAP7_75t_R FILLER_50_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_439 ();
 DECAPx4_ASAP7_75t_R FILLER_50_443 ();
 FILLER_ASAP7_75t_R FILLER_50_453 ();
 DECAPx4_ASAP7_75t_R FILLER_50_473 ();
 FILLER_ASAP7_75t_R FILLER_50_483 ();
 FILLER_ASAP7_75t_R FILLER_50_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_513 ();
 DECAPx2_ASAP7_75t_R FILLER_50_552 ();
 DECAPx2_ASAP7_75t_R FILLER_50_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_573 ();
 FILLER_ASAP7_75t_R FILLER_50_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_612 ();
 DECAPx6_ASAP7_75t_R FILLER_50_633 ();
 DECAPx2_ASAP7_75t_R FILLER_50_647 ();
 DECAPx10_ASAP7_75t_R FILLER_50_681 ();
 FILLER_ASAP7_75t_R FILLER_50_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_705 ();
 DECAPx6_ASAP7_75t_R FILLER_50_709 ();
 DECAPx6_ASAP7_75t_R FILLER_50_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_757 ();
 DECAPx2_ASAP7_75t_R FILLER_50_782 ();
 FILLER_ASAP7_75t_R FILLER_50_788 ();
 DECAPx1_ASAP7_75t_R FILLER_50_803 ();
 DECAPx6_ASAP7_75t_R FILLER_50_821 ();
 DECAPx2_ASAP7_75t_R FILLER_50_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_841 ();
 DECAPx4_ASAP7_75t_R FILLER_50_860 ();
 FILLER_ASAP7_75t_R FILLER_50_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_878 ();
 DECAPx1_ASAP7_75t_R FILLER_50_891 ();
 DECAPx6_ASAP7_75t_R FILLER_50_921 ();
 DECAPx2_ASAP7_75t_R FILLER_50_935 ();
 DECAPx1_ASAP7_75t_R FILLER_50_944 ();
 DECAPx1_ASAP7_75t_R FILLER_50_982 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1023 ();
 FILLER_ASAP7_75t_R FILLER_50_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1076 ();
 FILLER_ASAP7_75t_R FILLER_50_1082 ();
 FILLER_ASAP7_75t_R FILLER_50_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1361 ();
 FILLER_ASAP7_75t_R FILLER_50_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1388 ();
 FILLER_ASAP7_75t_R FILLER_50_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_51_24 ();
 DECAPx6_ASAP7_75t_R FILLER_51_46 ();
 DECAPx1_ASAP7_75t_R FILLER_51_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_116 ();
 DECAPx4_ASAP7_75t_R FILLER_51_120 ();
 FILLER_ASAP7_75t_R FILLER_51_130 ();
 DECAPx10_ASAP7_75t_R FILLER_51_175 ();
 DECAPx2_ASAP7_75t_R FILLER_51_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_203 ();
 DECAPx10_ASAP7_75t_R FILLER_51_220 ();
 DECAPx10_ASAP7_75t_R FILLER_51_242 ();
 FILLER_ASAP7_75t_R FILLER_51_264 ();
 DECAPx10_ASAP7_75t_R FILLER_51_272 ();
 DECAPx6_ASAP7_75t_R FILLER_51_294 ();
 DECAPx2_ASAP7_75t_R FILLER_51_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_314 ();
 DECAPx10_ASAP7_75t_R FILLER_51_321 ();
 FILLER_ASAP7_75t_R FILLER_51_343 ();
 FILLER_ASAP7_75t_R FILLER_51_351 ();
 DECAPx1_ASAP7_75t_R FILLER_51_393 ();
 FILLER_ASAP7_75t_R FILLER_51_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_412 ();
 DECAPx10_ASAP7_75t_R FILLER_51_416 ();
 DECAPx10_ASAP7_75t_R FILLER_51_438 ();
 DECAPx10_ASAP7_75t_R FILLER_51_460 ();
 FILLER_ASAP7_75t_R FILLER_51_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_498 ();
 DECAPx6_ASAP7_75t_R FILLER_51_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_539 ();
 DECAPx2_ASAP7_75t_R FILLER_51_543 ();
 FILLER_ASAP7_75t_R FILLER_51_549 ();
 DECAPx2_ASAP7_75t_R FILLER_51_557 ();
 FILLER_ASAP7_75t_R FILLER_51_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_565 ();
 DECAPx10_ASAP7_75t_R FILLER_51_569 ();
 DECAPx6_ASAP7_75t_R FILLER_51_603 ();
 DECAPx2_ASAP7_75t_R FILLER_51_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_638 ();
 DECAPx6_ASAP7_75t_R FILLER_51_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_662 ();
 DECAPx4_ASAP7_75t_R FILLER_51_666 ();
 FILLER_ASAP7_75t_R FILLER_51_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_678 ();
 DECAPx4_ASAP7_75t_R FILLER_51_682 ();
 FILLER_ASAP7_75t_R FILLER_51_706 ();
 FILLER_ASAP7_75t_R FILLER_51_711 ();
 DECAPx10_ASAP7_75t_R FILLER_51_725 ();
 FILLER_ASAP7_75t_R FILLER_51_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_768 ();
 DECAPx2_ASAP7_75t_R FILLER_51_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_794 ();
 FILLER_ASAP7_75t_R FILLER_51_816 ();
 FILLER_ASAP7_75t_R FILLER_51_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_842 ();
 FILLER_ASAP7_75t_R FILLER_51_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_857 ();
 DECAPx10_ASAP7_75t_R FILLER_51_868 ();
 FILLER_ASAP7_75t_R FILLER_51_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_892 ();
 DECAPx2_ASAP7_75t_R FILLER_51_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_909 ();
 DECAPx4_ASAP7_75t_R FILLER_51_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_926 ();
 DECAPx2_ASAP7_75t_R FILLER_51_966 ();
 FILLER_ASAP7_75t_R FILLER_51_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_974 ();
 DECAPx6_ASAP7_75t_R FILLER_51_978 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1358 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1380 ();
 FILLER_ASAP7_75t_R FILLER_51_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_52_2 ();
 DECAPx10_ASAP7_75t_R FILLER_52_24 ();
 DECAPx10_ASAP7_75t_R FILLER_52_46 ();
 DECAPx6_ASAP7_75t_R FILLER_52_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_82 ();
 DECAPx1_ASAP7_75t_R FILLER_52_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_90 ();
 DECAPx1_ASAP7_75t_R FILLER_52_103 ();
 DECAPx2_ASAP7_75t_R FILLER_52_133 ();
 FILLER_ASAP7_75t_R FILLER_52_165 ();
 DECAPx2_ASAP7_75t_R FILLER_52_193 ();
 FILLER_ASAP7_75t_R FILLER_52_199 ();
 DECAPx10_ASAP7_75t_R FILLER_52_207 ();
 DECAPx1_ASAP7_75t_R FILLER_52_229 ();
 FILLER_ASAP7_75t_R FILLER_52_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_249 ();
 DECAPx4_ASAP7_75t_R FILLER_52_256 ();
 FILLER_ASAP7_75t_R FILLER_52_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_268 ();
 DECAPx4_ASAP7_75t_R FILLER_52_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_287 ();
 DECAPx6_ASAP7_75t_R FILLER_52_302 ();
 DECAPx1_ASAP7_75t_R FILLER_52_316 ();
 DECAPx4_ASAP7_75t_R FILLER_52_328 ();
 FILLER_ASAP7_75t_R FILLER_52_338 ();
 DECAPx2_ASAP7_75t_R FILLER_52_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_354 ();
 DECAPx1_ASAP7_75t_R FILLER_52_381 ();
 DECAPx2_ASAP7_75t_R FILLER_52_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_397 ();
 DECAPx2_ASAP7_75t_R FILLER_52_456 ();
 DECAPx2_ASAP7_75t_R FILLER_52_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_513 ();
 DECAPx6_ASAP7_75t_R FILLER_52_517 ();
 FILLER_ASAP7_75t_R FILLER_52_531 ();
 DECAPx2_ASAP7_75t_R FILLER_52_539 ();
 DECAPx2_ASAP7_75t_R FILLER_52_577 ();
 DECAPx4_ASAP7_75t_R FILLER_52_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_637 ();
 DECAPx2_ASAP7_75t_R FILLER_52_655 ();
 FILLER_ASAP7_75t_R FILLER_52_675 ();
 FILLER_ASAP7_75t_R FILLER_52_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_691 ();
 FILLER_ASAP7_75t_R FILLER_52_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_708 ();
 DECAPx2_ASAP7_75t_R FILLER_52_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_729 ();
 DECAPx1_ASAP7_75t_R FILLER_52_739 ();
 DECAPx2_ASAP7_75t_R FILLER_52_755 ();
 FILLER_ASAP7_75t_R FILLER_52_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_763 ();
 DECAPx1_ASAP7_75t_R FILLER_52_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_796 ();
 DECAPx10_ASAP7_75t_R FILLER_52_809 ();
 DECAPx2_ASAP7_75t_R FILLER_52_831 ();
 DECAPx2_ASAP7_75t_R FILLER_52_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_883 ();
 DECAPx4_ASAP7_75t_R FILLER_52_890 ();
 DECAPx6_ASAP7_75t_R FILLER_52_908 ();
 FILLER_ASAP7_75t_R FILLER_52_922 ();
 DECAPx1_ASAP7_75t_R FILLER_52_936 ();
 DECAPx1_ASAP7_75t_R FILLER_52_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_957 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1013 ();
 FILLER_ASAP7_75t_R FILLER_52_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1046 ();
 FILLER_ASAP7_75t_R FILLER_52_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1104 ();
 FILLER_ASAP7_75t_R FILLER_52_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1370 ();
 FILLER_ASAP7_75t_R FILLER_52_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1388 ();
 FILLER_ASAP7_75t_R FILLER_52_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_53_2 ();
 DECAPx1_ASAP7_75t_R FILLER_53_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_28 ();
 FILLER_ASAP7_75t_R FILLER_53_59 ();
 DECAPx1_ASAP7_75t_R FILLER_53_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_68 ();
 DECAPx1_ASAP7_75t_R FILLER_53_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_103 ();
 DECAPx6_ASAP7_75t_R FILLER_53_107 ();
 DECAPx2_ASAP7_75t_R FILLER_53_194 ();
 DECAPx6_ASAP7_75t_R FILLER_53_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_228 ();
 DECAPx10_ASAP7_75t_R FILLER_53_265 ();
 DECAPx1_ASAP7_75t_R FILLER_53_287 ();
 DECAPx10_ASAP7_75t_R FILLER_53_297 ();
 DECAPx6_ASAP7_75t_R FILLER_53_319 ();
 FILLER_ASAP7_75t_R FILLER_53_333 ();
 DECAPx6_ASAP7_75t_R FILLER_53_341 ();
 DECAPx2_ASAP7_75t_R FILLER_53_355 ();
 DECAPx6_ASAP7_75t_R FILLER_53_367 ();
 FILLER_ASAP7_75t_R FILLER_53_381 ();
 DECAPx1_ASAP7_75t_R FILLER_53_434 ();
 FILLER_ASAP7_75t_R FILLER_53_525 ();
 DECAPx2_ASAP7_75t_R FILLER_53_553 ();
 FILLER_ASAP7_75t_R FILLER_53_559 ();
 FILLER_ASAP7_75t_R FILLER_53_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_597 ();
 DECAPx6_ASAP7_75t_R FILLER_53_601 ();
 FILLER_ASAP7_75t_R FILLER_53_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_626 ();
 DECAPx1_ASAP7_75t_R FILLER_53_644 ();
 DECAPx6_ASAP7_75t_R FILLER_53_676 ();
 DECAPx1_ASAP7_75t_R FILLER_53_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_694 ();
 DECAPx1_ASAP7_75t_R FILLER_53_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_711 ();
 DECAPx4_ASAP7_75t_R FILLER_53_715 ();
 DECAPx1_ASAP7_75t_R FILLER_53_754 ();
 FILLER_ASAP7_75t_R FILLER_53_779 ();
 FILLER_ASAP7_75t_R FILLER_53_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_795 ();
 DECAPx6_ASAP7_75t_R FILLER_53_802 ();
 FILLER_ASAP7_75t_R FILLER_53_816 ();
 DECAPx10_ASAP7_75t_R FILLER_53_826 ();
 DECAPx4_ASAP7_75t_R FILLER_53_848 ();
 FILLER_ASAP7_75t_R FILLER_53_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_860 ();
 DECAPx6_ASAP7_75t_R FILLER_53_867 ();
 FILLER_ASAP7_75t_R FILLER_53_900 ();
 DECAPx1_ASAP7_75t_R FILLER_53_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_912 ();
 DECAPx1_ASAP7_75t_R FILLER_53_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_923 ();
 DECAPx1_ASAP7_75t_R FILLER_53_939 ();
 DECAPx6_ASAP7_75t_R FILLER_53_993 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1022 ();
 FILLER_ASAP7_75t_R FILLER_53_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1101 ();
 FILLER_ASAP7_75t_R FILLER_53_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1109 ();
 FILLER_ASAP7_75t_R FILLER_53_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1119 ();
 FILLER_ASAP7_75t_R FILLER_53_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1386 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_54_2 ();
 FILLER_ASAP7_75t_R FILLER_54_24 ();
 DECAPx4_ASAP7_75t_R FILLER_54_96 ();
 FILLER_ASAP7_75t_R FILLER_54_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_108 ();
 FILLER_ASAP7_75t_R FILLER_54_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_126 ();
 DECAPx2_ASAP7_75t_R FILLER_54_145 ();
 FILLER_ASAP7_75t_R FILLER_54_151 ();
 DECAPx2_ASAP7_75t_R FILLER_54_156 ();
 FILLER_ASAP7_75t_R FILLER_54_162 ();
 DECAPx4_ASAP7_75t_R FILLER_54_186 ();
 DECAPx1_ASAP7_75t_R FILLER_54_216 ();
 DECAPx1_ASAP7_75t_R FILLER_54_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_230 ();
 FILLER_ASAP7_75t_R FILLER_54_237 ();
 DECAPx1_ASAP7_75t_R FILLER_54_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_249 ();
 DECAPx10_ASAP7_75t_R FILLER_54_258 ();
 DECAPx10_ASAP7_75t_R FILLER_54_280 ();
 FILLER_ASAP7_75t_R FILLER_54_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_304 ();
 DECAPx4_ASAP7_75t_R FILLER_54_325 ();
 FILLER_ASAP7_75t_R FILLER_54_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_337 ();
 DECAPx6_ASAP7_75t_R FILLER_54_344 ();
 DECAPx1_ASAP7_75t_R FILLER_54_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_362 ();
 FILLER_ASAP7_75t_R FILLER_54_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_401 ();
 DECAPx2_ASAP7_75t_R FILLER_54_410 ();
 FILLER_ASAP7_75t_R FILLER_54_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_439 ();
 DECAPx6_ASAP7_75t_R FILLER_54_446 ();
 FILLER_ASAP7_75t_R FILLER_54_460 ();
 DECAPx2_ASAP7_75t_R FILLER_54_464 ();
 FILLER_ASAP7_75t_R FILLER_54_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_472 ();
 FILLER_ASAP7_75t_R FILLER_54_489 ();
 DECAPx6_ASAP7_75t_R FILLER_54_494 ();
 FILLER_ASAP7_75t_R FILLER_54_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_516 ();
 DECAPx1_ASAP7_75t_R FILLER_54_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_540 ();
 DECAPx6_ASAP7_75t_R FILLER_54_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_558 ();
 DECAPx6_ASAP7_75t_R FILLER_54_567 ();
 FILLER_ASAP7_75t_R FILLER_54_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_583 ();
 DECAPx1_ASAP7_75t_R FILLER_54_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_591 ();
 DECAPx2_ASAP7_75t_R FILLER_54_601 ();
 DECAPx10_ASAP7_75t_R FILLER_54_627 ();
 DECAPx4_ASAP7_75t_R FILLER_54_649 ();
 DECAPx4_ASAP7_75t_R FILLER_54_662 ();
 FILLER_ASAP7_75t_R FILLER_54_672 ();
 DECAPx2_ASAP7_75t_R FILLER_54_677 ();
 DECAPx1_ASAP7_75t_R FILLER_54_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_707 ();
 DECAPx10_ASAP7_75t_R FILLER_54_714 ();
 DECAPx2_ASAP7_75t_R FILLER_54_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_742 ();
 DECAPx1_ASAP7_75t_R FILLER_54_767 ();
 DECAPx6_ASAP7_75t_R FILLER_54_789 ();
 DECAPx1_ASAP7_75t_R FILLER_54_803 ();
 DECAPx2_ASAP7_75t_R FILLER_54_813 ();
 FILLER_ASAP7_75t_R FILLER_54_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_821 ();
 DECAPx4_ASAP7_75t_R FILLER_54_832 ();
 DECAPx4_ASAP7_75t_R FILLER_54_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_858 ();
 DECAPx1_ASAP7_75t_R FILLER_54_875 ();
 DECAPx2_ASAP7_75t_R FILLER_54_885 ();
 FILLER_ASAP7_75t_R FILLER_54_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_893 ();
 DECAPx2_ASAP7_75t_R FILLER_54_900 ();
 DECAPx10_ASAP7_75t_R FILLER_54_928 ();
 FILLER_ASAP7_75t_R FILLER_54_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_961 ();
 DECAPx1_ASAP7_75t_R FILLER_54_972 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1019 ();
 FILLER_ASAP7_75t_R FILLER_54_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1073 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1100 ();
 FILLER_ASAP7_75t_R FILLER_54_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1388 ();
 FILLER_ASAP7_75t_R FILLER_54_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_55_2 ();
 DECAPx6_ASAP7_75t_R FILLER_55_24 ();
 DECAPx2_ASAP7_75t_R FILLER_55_38 ();
 FILLER_ASAP7_75t_R FILLER_55_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_49 ();
 DECAPx6_ASAP7_75t_R FILLER_55_56 ();
 FILLER_ASAP7_75t_R FILLER_55_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_72 ();
 FILLER_ASAP7_75t_R FILLER_55_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_84 ();
 DECAPx10_ASAP7_75t_R FILLER_55_88 ();
 DECAPx10_ASAP7_75t_R FILLER_55_110 ();
 DECAPx2_ASAP7_75t_R FILLER_55_132 ();
 FILLER_ASAP7_75t_R FILLER_55_138 ();
 FILLER_ASAP7_75t_R FILLER_55_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_149 ();
 DECAPx10_ASAP7_75t_R FILLER_55_156 ();
 DECAPx10_ASAP7_75t_R FILLER_55_178 ();
 DECAPx1_ASAP7_75t_R FILLER_55_214 ();
 DECAPx2_ASAP7_75t_R FILLER_55_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_238 ();
 DECAPx6_ASAP7_75t_R FILLER_55_251 ();
 FILLER_ASAP7_75t_R FILLER_55_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_275 ();
 DECAPx1_ASAP7_75t_R FILLER_55_288 ();
 DECAPx6_ASAP7_75t_R FILLER_55_298 ();
 DECAPx2_ASAP7_75t_R FILLER_55_326 ();
 FILLER_ASAP7_75t_R FILLER_55_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_334 ();
 DECAPx2_ASAP7_75t_R FILLER_55_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_348 ();
 DECAPx4_ASAP7_75t_R FILLER_55_352 ();
 FILLER_ASAP7_75t_R FILLER_55_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_364 ();
 DECAPx10_ASAP7_75t_R FILLER_55_381 ();
 DECAPx6_ASAP7_75t_R FILLER_55_403 ();
 FILLER_ASAP7_75t_R FILLER_55_417 ();
 FILLER_ASAP7_75t_R FILLER_55_431 ();
 DECAPx6_ASAP7_75t_R FILLER_55_449 ();
 DECAPx4_ASAP7_75t_R FILLER_55_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_480 ();
 DECAPx2_ASAP7_75t_R FILLER_55_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_513 ();
 DECAPx10_ASAP7_75t_R FILLER_55_517 ();
 DECAPx2_ASAP7_75t_R FILLER_55_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_545 ();
 DECAPx2_ASAP7_75t_R FILLER_55_572 ();
 FILLER_ASAP7_75t_R FILLER_55_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_580 ();
 DECAPx2_ASAP7_75t_R FILLER_55_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_616 ();
 FILLER_ASAP7_75t_R FILLER_55_623 ();
 DECAPx1_ASAP7_75t_R FILLER_55_628 ();
 DECAPx6_ASAP7_75t_R FILLER_55_635 ();
 FILLER_ASAP7_75t_R FILLER_55_649 ();
 DECAPx1_ASAP7_75t_R FILLER_55_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_658 ();
 DECAPx4_ASAP7_75t_R FILLER_55_662 ();
 FILLER_ASAP7_75t_R FILLER_55_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_699 ();
 FILLER_ASAP7_75t_R FILLER_55_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_731 ();
 DECAPx2_ASAP7_75t_R FILLER_55_738 ();
 FILLER_ASAP7_75t_R FILLER_55_744 ();
 DECAPx10_ASAP7_75t_R FILLER_55_766 ();
 DECAPx6_ASAP7_75t_R FILLER_55_788 ();
 DECAPx1_ASAP7_75t_R FILLER_55_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_806 ();
 DECAPx1_ASAP7_75t_R FILLER_55_819 ();
 FILLER_ASAP7_75t_R FILLER_55_844 ();
 DECAPx1_ASAP7_75t_R FILLER_55_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_853 ();
 DECAPx2_ASAP7_75t_R FILLER_55_868 ();
 FILLER_ASAP7_75t_R FILLER_55_874 ();
 FILLER_ASAP7_75t_R FILLER_55_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_888 ();
 FILLER_ASAP7_75t_R FILLER_55_901 ();
 DECAPx2_ASAP7_75t_R FILLER_55_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_915 ();
 FILLER_ASAP7_75t_R FILLER_55_922 ();
 DECAPx2_ASAP7_75t_R FILLER_55_936 ();
 FILLER_ASAP7_75t_R FILLER_55_942 ();
 DECAPx1_ASAP7_75t_R FILLER_55_986 ();
 DECAPx1_ASAP7_75t_R FILLER_55_993 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1007 ();
 FILLER_ASAP7_75t_R FILLER_55_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_55_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1124 ();
 FILLER_ASAP7_75t_R FILLER_55_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1359 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1381 ();
 FILLER_ASAP7_75t_R FILLER_55_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_56_2 ();
 DECAPx2_ASAP7_75t_R FILLER_56_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_30 ();
 DECAPx10_ASAP7_75t_R FILLER_56_40 ();
 DECAPx2_ASAP7_75t_R FILLER_56_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_68 ();
 DECAPx10_ASAP7_75t_R FILLER_56_72 ();
 FILLER_ASAP7_75t_R FILLER_56_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_110 ();
 DECAPx6_ASAP7_75t_R FILLER_56_119 ();
 FILLER_ASAP7_75t_R FILLER_56_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_135 ();
 DECAPx2_ASAP7_75t_R FILLER_56_162 ();
 DECAPx4_ASAP7_75t_R FILLER_56_174 ();
 FILLER_ASAP7_75t_R FILLER_56_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_192 ();
 DECAPx2_ASAP7_75t_R FILLER_56_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_211 ();
 DECAPx4_ASAP7_75t_R FILLER_56_218 ();
 DECAPx2_ASAP7_75t_R FILLER_56_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_241 ();
 DECAPx2_ASAP7_75t_R FILLER_56_248 ();
 FILLER_ASAP7_75t_R FILLER_56_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_256 ();
 DECAPx4_ASAP7_75t_R FILLER_56_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_315 ();
 DECAPx4_ASAP7_75t_R FILLER_56_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_333 ();
 DECAPx2_ASAP7_75t_R FILLER_56_360 ();
 DECAPx6_ASAP7_75t_R FILLER_56_369 ();
 DECAPx1_ASAP7_75t_R FILLER_56_383 ();
 DECAPx10_ASAP7_75t_R FILLER_56_413 ();
 DECAPx4_ASAP7_75t_R FILLER_56_435 ();
 DECAPx1_ASAP7_75t_R FILLER_56_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_461 ();
 DECAPx4_ASAP7_75t_R FILLER_56_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_500 ();
 DECAPx1_ASAP7_75t_R FILLER_56_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_531 ();
 DECAPx4_ASAP7_75t_R FILLER_56_535 ();
 FILLER_ASAP7_75t_R FILLER_56_545 ();
 DECAPx2_ASAP7_75t_R FILLER_56_554 ();
 FILLER_ASAP7_75t_R FILLER_56_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_588 ();
 DECAPx10_ASAP7_75t_R FILLER_56_595 ();
 DECAPx2_ASAP7_75t_R FILLER_56_617 ();
 FILLER_ASAP7_75t_R FILLER_56_623 ();
 FILLER_ASAP7_75t_R FILLER_56_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_641 ();
 FILLER_ASAP7_75t_R FILLER_56_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_657 ();
 DECAPx6_ASAP7_75t_R FILLER_56_675 ();
 FILLER_ASAP7_75t_R FILLER_56_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_691 ();
 DECAPx4_ASAP7_75t_R FILLER_56_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_732 ();
 DECAPx2_ASAP7_75t_R FILLER_56_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_750 ();
 DECAPx6_ASAP7_75t_R FILLER_56_758 ();
 FILLER_ASAP7_75t_R FILLER_56_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_797 ();
 FILLER_ASAP7_75t_R FILLER_56_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_806 ();
 DECAPx1_ASAP7_75t_R FILLER_56_821 ();
 FILLER_ASAP7_75t_R FILLER_56_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_841 ();
 FILLER_ASAP7_75t_R FILLER_56_872 ();
 DECAPx2_ASAP7_75t_R FILLER_56_900 ();
 FILLER_ASAP7_75t_R FILLER_56_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_908 ();
 FILLER_ASAP7_75t_R FILLER_56_916 ();
 DECAPx6_ASAP7_75t_R FILLER_56_944 ();
 DECAPx2_ASAP7_75t_R FILLER_56_961 ();
 FILLER_ASAP7_75t_R FILLER_56_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_969 ();
 DECAPx2_ASAP7_75t_R FILLER_56_978 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1000 ();
 FILLER_ASAP7_75t_R FILLER_56_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1023 ();
 FILLER_ASAP7_75t_R FILLER_56_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1049 ();
 FILLER_ASAP7_75t_R FILLER_56_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1077 ();
 FILLER_ASAP7_75t_R FILLER_56_1089 ();
 FILLER_ASAP7_75t_R FILLER_56_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1125 ();
 FILLER_ASAP7_75t_R FILLER_56_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1142 ();
 FILLER_ASAP7_75t_R FILLER_56_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1382 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1388 ();
 FILLER_ASAP7_75t_R FILLER_56_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_57_2 ();
 FILLER_ASAP7_75t_R FILLER_57_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_53 ();
 FILLER_ASAP7_75t_R FILLER_57_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_85 ();
 DECAPx1_ASAP7_75t_R FILLER_57_112 ();
 FILLER_ASAP7_75t_R FILLER_57_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_127 ();
 DECAPx2_ASAP7_75t_R FILLER_57_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_185 ();
 DECAPx1_ASAP7_75t_R FILLER_57_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_215 ();
 FILLER_ASAP7_75t_R FILLER_57_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_246 ();
 DECAPx4_ASAP7_75t_R FILLER_57_261 ();
 FILLER_ASAP7_75t_R FILLER_57_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_305 ();
 FILLER_ASAP7_75t_R FILLER_57_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_334 ();
 DECAPx1_ASAP7_75t_R FILLER_57_341 ();
 DECAPx6_ASAP7_75t_R FILLER_57_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_391 ();
 DECAPx4_ASAP7_75t_R FILLER_57_408 ();
 FILLER_ASAP7_75t_R FILLER_57_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_420 ();
 DECAPx6_ASAP7_75t_R FILLER_57_433 ();
 DECAPx4_ASAP7_75t_R FILLER_57_453 ();
 FILLER_ASAP7_75t_R FILLER_57_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_465 ();
 FILLER_ASAP7_75t_R FILLER_57_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_474 ();
 FILLER_ASAP7_75t_R FILLER_57_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_480 ();
 DECAPx2_ASAP7_75t_R FILLER_57_487 ();
 FILLER_ASAP7_75t_R FILLER_57_493 ();
 FILLER_ASAP7_75t_R FILLER_57_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_511 ();
 DECAPx1_ASAP7_75t_R FILLER_57_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_558 ();
 DECAPx1_ASAP7_75t_R FILLER_57_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_589 ();
 FILLER_ASAP7_75t_R FILLER_57_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_598 ();
 FILLER_ASAP7_75t_R FILLER_57_602 ();
 DECAPx2_ASAP7_75t_R FILLER_57_612 ();
 FILLER_ASAP7_75t_R FILLER_57_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_673 ();
 DECAPx6_ASAP7_75t_R FILLER_57_683 ();
 DECAPx1_ASAP7_75t_R FILLER_57_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_701 ();
 DECAPx1_ASAP7_75t_R FILLER_57_705 ();
 FILLER_ASAP7_75t_R FILLER_57_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_744 ();
 DECAPx2_ASAP7_75t_R FILLER_57_763 ();
 FILLER_ASAP7_75t_R FILLER_57_769 ();
 DECAPx1_ASAP7_75t_R FILLER_57_783 ();
 DECAPx6_ASAP7_75t_R FILLER_57_807 ();
 DECAPx1_ASAP7_75t_R FILLER_57_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_825 ();
 FILLER_ASAP7_75t_R FILLER_57_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_831 ();
 DECAPx4_ASAP7_75t_R FILLER_57_847 ();
 FILLER_ASAP7_75t_R FILLER_57_857 ();
 DECAPx4_ASAP7_75t_R FILLER_57_871 ();
 DECAPx2_ASAP7_75t_R FILLER_57_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_897 ();
 DECAPx6_ASAP7_75t_R FILLER_57_910 ();
 DECAPx1_ASAP7_75t_R FILLER_57_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_930 ();
 DECAPx6_ASAP7_75t_R FILLER_57_950 ();
 DECAPx6_ASAP7_75t_R FILLER_57_976 ();
 DECAPx2_ASAP7_75t_R FILLER_57_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_57_1037 ();
 FILLER_ASAP7_75t_R FILLER_57_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_57_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1072 ();
 FILLER_ASAP7_75t_R FILLER_57_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_58_2 ();
 DECAPx1_ASAP7_75t_R FILLER_58_24 ();
 DECAPx2_ASAP7_75t_R FILLER_58_37 ();
 FILLER_ASAP7_75t_R FILLER_58_84 ();
 FILLER_ASAP7_75t_R FILLER_58_98 ();
 DECAPx1_ASAP7_75t_R FILLER_58_103 ();
 DECAPx2_ASAP7_75t_R FILLER_58_149 ();
 FILLER_ASAP7_75t_R FILLER_58_155 ();
 DECAPx1_ASAP7_75t_R FILLER_58_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_179 ();
 FILLER_ASAP7_75t_R FILLER_58_194 ();
 FILLER_ASAP7_75t_R FILLER_58_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_214 ();
 DECAPx6_ASAP7_75t_R FILLER_58_228 ();
 DECAPx1_ASAP7_75t_R FILLER_58_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_252 ();
 DECAPx10_ASAP7_75t_R FILLER_58_265 ();
 DECAPx2_ASAP7_75t_R FILLER_58_287 ();
 FILLER_ASAP7_75t_R FILLER_58_293 ();
 DECAPx4_ASAP7_75t_R FILLER_58_301 ();
 DECAPx1_ASAP7_75t_R FILLER_58_347 ();
 DECAPx4_ASAP7_75t_R FILLER_58_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_383 ();
 DECAPx6_ASAP7_75t_R FILLER_58_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_404 ();
 DECAPx6_ASAP7_75t_R FILLER_58_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_461 ();
 DECAPx6_ASAP7_75t_R FILLER_58_464 ();
 DECAPx1_ASAP7_75t_R FILLER_58_478 ();
 DECAPx6_ASAP7_75t_R FILLER_58_488 ();
 FILLER_ASAP7_75t_R FILLER_58_502 ();
 DECAPx2_ASAP7_75t_R FILLER_58_510 ();
 FILLER_ASAP7_75t_R FILLER_58_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_528 ();
 DECAPx2_ASAP7_75t_R FILLER_58_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_542 ();
 DECAPx1_ASAP7_75t_R FILLER_58_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_550 ();
 FILLER_ASAP7_75t_R FILLER_58_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_559 ();
 DECAPx4_ASAP7_75t_R FILLER_58_563 ();
 FILLER_ASAP7_75t_R FILLER_58_573 ();
 DECAPx2_ASAP7_75t_R FILLER_58_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_617 ();
 DECAPx10_ASAP7_75t_R FILLER_58_632 ();
 DECAPx2_ASAP7_75t_R FILLER_58_668 ();
 FILLER_ASAP7_75t_R FILLER_58_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_676 ();
 FILLER_ASAP7_75t_R FILLER_58_686 ();
 DECAPx6_ASAP7_75t_R FILLER_58_702 ();
 DECAPx1_ASAP7_75t_R FILLER_58_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_720 ();
 FILLER_ASAP7_75t_R FILLER_58_739 ();
 FILLER_ASAP7_75t_R FILLER_58_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_764 ();
 DECAPx1_ASAP7_75t_R FILLER_58_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_794 ();
 DECAPx1_ASAP7_75t_R FILLER_58_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_805 ();
 FILLER_ASAP7_75t_R FILLER_58_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_820 ();
 DECAPx4_ASAP7_75t_R FILLER_58_827 ();
 DECAPx2_ASAP7_75t_R FILLER_58_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_846 ();
 DECAPx4_ASAP7_75t_R FILLER_58_850 ();
 FILLER_ASAP7_75t_R FILLER_58_860 ();
 FILLER_ASAP7_75t_R FILLER_58_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_870 ();
 DECAPx1_ASAP7_75t_R FILLER_58_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_878 ();
 DECAPx10_ASAP7_75t_R FILLER_58_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_919 ();
 DECAPx4_ASAP7_75t_R FILLER_58_929 ();
 DECAPx1_ASAP7_75t_R FILLER_58_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_959 ();
 FILLER_ASAP7_75t_R FILLER_58_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_994 ();
 DECAPx4_ASAP7_75t_R FILLER_58_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1027 ();
 FILLER_ASAP7_75t_R FILLER_58_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1099 ();
 FILLER_ASAP7_75t_R FILLER_58_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1123 ();
 FILLER_ASAP7_75t_R FILLER_58_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1158 ();
 FILLER_ASAP7_75t_R FILLER_58_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1370 ();
 FILLER_ASAP7_75t_R FILLER_58_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1388 ();
 FILLER_ASAP7_75t_R FILLER_58_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_59_2 ();
 FILLER_ASAP7_75t_R FILLER_59_16 ();
 DECAPx1_ASAP7_75t_R FILLER_59_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_51 ();
 FILLER_ASAP7_75t_R FILLER_59_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_60 ();
 DECAPx4_ASAP7_75t_R FILLER_59_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_80 ();
 FILLER_ASAP7_75t_R FILLER_59_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_97 ();
 DECAPx2_ASAP7_75t_R FILLER_59_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_110 ();
 DECAPx10_ASAP7_75t_R FILLER_59_123 ();
 DECAPx6_ASAP7_75t_R FILLER_59_145 ();
 DECAPx1_ASAP7_75t_R FILLER_59_159 ();
 DECAPx4_ASAP7_75t_R FILLER_59_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_210 ();
 DECAPx10_ASAP7_75t_R FILLER_59_217 ();
 DECAPx2_ASAP7_75t_R FILLER_59_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_245 ();
 DECAPx6_ASAP7_75t_R FILLER_59_254 ();
 DECAPx2_ASAP7_75t_R FILLER_59_268 ();
 DECAPx10_ASAP7_75t_R FILLER_59_284 ();
 DECAPx2_ASAP7_75t_R FILLER_59_306 ();
 FILLER_ASAP7_75t_R FILLER_59_312 ();
 DECAPx6_ASAP7_75t_R FILLER_59_320 ();
 DECAPx10_ASAP7_75t_R FILLER_59_340 ();
 DECAPx6_ASAP7_75t_R FILLER_59_362 ();
 DECAPx2_ASAP7_75t_R FILLER_59_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_382 ();
 DECAPx10_ASAP7_75t_R FILLER_59_391 ();
 DECAPx6_ASAP7_75t_R FILLER_59_413 ();
 FILLER_ASAP7_75t_R FILLER_59_427 ();
 DECAPx2_ASAP7_75t_R FILLER_59_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_441 ();
 DECAPx10_ASAP7_75t_R FILLER_59_456 ();
 DECAPx10_ASAP7_75t_R FILLER_59_504 ();
 FILLER_ASAP7_75t_R FILLER_59_526 ();
 DECAPx4_ASAP7_75t_R FILLER_59_554 ();
 DECAPx6_ASAP7_75t_R FILLER_59_570 ();
 DECAPx1_ASAP7_75t_R FILLER_59_584 ();
 DECAPx2_ASAP7_75t_R FILLER_59_606 ();
 DECAPx1_ASAP7_75t_R FILLER_59_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_619 ();
 DECAPx1_ASAP7_75t_R FILLER_59_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_630 ();
 DECAPx2_ASAP7_75t_R FILLER_59_634 ();
 DECAPx4_ASAP7_75t_R FILLER_59_652 ();
 FILLER_ASAP7_75t_R FILLER_59_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_664 ();
 FILLER_ASAP7_75t_R FILLER_59_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_701 ();
 DECAPx1_ASAP7_75t_R FILLER_59_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_729 ();
 DECAPx6_ASAP7_75t_R FILLER_59_736 ();
 FILLER_ASAP7_75t_R FILLER_59_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_752 ();
 DECAPx10_ASAP7_75t_R FILLER_59_759 ();
 DECAPx4_ASAP7_75t_R FILLER_59_781 ();
 FILLER_ASAP7_75t_R FILLER_59_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_808 ();
 DECAPx2_ASAP7_75t_R FILLER_59_812 ();
 FILLER_ASAP7_75t_R FILLER_59_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_842 ();
 DECAPx1_ASAP7_75t_R FILLER_59_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_864 ();
 DECAPx6_ASAP7_75t_R FILLER_59_871 ();
 DECAPx2_ASAP7_75t_R FILLER_59_907 ();
 FILLER_ASAP7_75t_R FILLER_59_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_923 ();
 DECAPx6_ASAP7_75t_R FILLER_59_932 ();
 DECAPx2_ASAP7_75t_R FILLER_59_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_952 ();
 FILLER_ASAP7_75t_R FILLER_59_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_981 ();
 DECAPx2_ASAP7_75t_R FILLER_59_998 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1020 ();
 FILLER_ASAP7_75t_R FILLER_59_1027 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1035 ();
 FILLER_ASAP7_75t_R FILLER_59_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1059 ();
 FILLER_ASAP7_75t_R FILLER_59_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1141 ();
 FILLER_ASAP7_75t_R FILLER_59_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1368 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1390 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_60_2 ();
 DECAPx2_ASAP7_75t_R FILLER_60_24 ();
 FILLER_ASAP7_75t_R FILLER_60_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_32 ();
 DECAPx10_ASAP7_75t_R FILLER_60_39 ();
 DECAPx10_ASAP7_75t_R FILLER_60_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_109 ();
 FILLER_ASAP7_75t_R FILLER_60_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_169 ();
 DECAPx10_ASAP7_75t_R FILLER_60_182 ();
 FILLER_ASAP7_75t_R FILLER_60_204 ();
 DECAPx4_ASAP7_75t_R FILLER_60_212 ();
 FILLER_ASAP7_75t_R FILLER_60_222 ();
 DECAPx6_ASAP7_75t_R FILLER_60_238 ();
 FILLER_ASAP7_75t_R FILLER_60_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_254 ();
 DECAPx4_ASAP7_75t_R FILLER_60_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_295 ();
 DECAPx6_ASAP7_75t_R FILLER_60_306 ();
 DECAPx2_ASAP7_75t_R FILLER_60_320 ();
 DECAPx6_ASAP7_75t_R FILLER_60_332 ();
 DECAPx1_ASAP7_75t_R FILLER_60_346 ();
 DECAPx6_ASAP7_75t_R FILLER_60_362 ();
 DECAPx2_ASAP7_75t_R FILLER_60_376 ();
 DECAPx6_ASAP7_75t_R FILLER_60_388 ();
 DECAPx1_ASAP7_75t_R FILLER_60_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_406 ();
 DECAPx2_ASAP7_75t_R FILLER_60_419 ();
 DECAPx4_ASAP7_75t_R FILLER_60_431 ();
 FILLER_ASAP7_75t_R FILLER_60_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_443 ();
 DECAPx1_ASAP7_75t_R FILLER_60_450 ();
 FILLER_ASAP7_75t_R FILLER_60_460 ();
 DECAPx2_ASAP7_75t_R FILLER_60_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_495 ();
 DECAPx2_ASAP7_75t_R FILLER_60_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_528 ();
 DECAPx10_ASAP7_75t_R FILLER_60_535 ();
 DECAPx2_ASAP7_75t_R FILLER_60_557 ();
 DECAPx2_ASAP7_75t_R FILLER_60_589 ();
 FILLER_ASAP7_75t_R FILLER_60_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_624 ();
 FILLER_ASAP7_75t_R FILLER_60_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_633 ();
 DECAPx10_ASAP7_75t_R FILLER_60_648 ();
 DECAPx6_ASAP7_75t_R FILLER_60_676 ();
 FILLER_ASAP7_75t_R FILLER_60_690 ();
 DECAPx1_ASAP7_75t_R FILLER_60_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_708 ();
 FILLER_ASAP7_75t_R FILLER_60_715 ();
 DECAPx10_ASAP7_75t_R FILLER_60_723 ();
 DECAPx2_ASAP7_75t_R FILLER_60_745 ();
 DECAPx10_ASAP7_75t_R FILLER_60_757 ();
 DECAPx1_ASAP7_75t_R FILLER_60_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_789 ();
 DECAPx4_ASAP7_75t_R FILLER_60_810 ();
 FILLER_ASAP7_75t_R FILLER_60_820 ();
 DECAPx2_ASAP7_75t_R FILLER_60_825 ();
 DECAPx2_ASAP7_75t_R FILLER_60_840 ();
 FILLER_ASAP7_75t_R FILLER_60_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_848 ();
 DECAPx4_ASAP7_75t_R FILLER_60_852 ();
 FILLER_ASAP7_75t_R FILLER_60_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_864 ();
 DECAPx10_ASAP7_75t_R FILLER_60_871 ();
 DECAPx2_ASAP7_75t_R FILLER_60_893 ();
 DECAPx10_ASAP7_75t_R FILLER_60_925 ();
 DECAPx2_ASAP7_75t_R FILLER_60_947 ();
 FILLER_ASAP7_75t_R FILLER_60_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_955 ();
 DECAPx2_ASAP7_75t_R FILLER_60_959 ();
 FILLER_ASAP7_75t_R FILLER_60_965 ();
 DECAPx1_ASAP7_75t_R FILLER_60_970 ();
 DECAPx2_ASAP7_75t_R FILLER_60_977 ();
 FILLER_ASAP7_75t_R FILLER_60_983 ();
 DECAPx6_ASAP7_75t_R FILLER_60_991 ();
 FILLER_ASAP7_75t_R FILLER_60_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1063 ();
 FILLER_ASAP7_75t_R FILLER_60_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1071 ();
 FILLER_ASAP7_75t_R FILLER_60_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1082 ();
 FILLER_ASAP7_75t_R FILLER_60_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1388 ();
 FILLER_ASAP7_75t_R FILLER_60_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_61_2 ();
 FILLER_ASAP7_75t_R FILLER_61_24 ();
 DECAPx1_ASAP7_75t_R FILLER_61_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_67 ();
 DECAPx4_ASAP7_75t_R FILLER_61_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_84 ();
 FILLER_ASAP7_75t_R FILLER_61_91 ();
 FILLER_ASAP7_75t_R FILLER_61_96 ();
 DECAPx4_ASAP7_75t_R FILLER_61_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_111 ();
 DECAPx1_ASAP7_75t_R FILLER_61_126 ();
 DECAPx1_ASAP7_75t_R FILLER_61_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_160 ();
 FILLER_ASAP7_75t_R FILLER_61_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_171 ();
 DECAPx1_ASAP7_75t_R FILLER_61_184 ();
 FILLER_ASAP7_75t_R FILLER_61_194 ();
 DECAPx1_ASAP7_75t_R FILLER_61_203 ();
 DECAPx4_ASAP7_75t_R FILLER_61_213 ();
 FILLER_ASAP7_75t_R FILLER_61_237 ();
 DECAPx2_ASAP7_75t_R FILLER_61_249 ();
 FILLER_ASAP7_75t_R FILLER_61_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_257 ();
 DECAPx2_ASAP7_75t_R FILLER_61_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_296 ();
 DECAPx4_ASAP7_75t_R FILLER_61_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_335 ();
 DECAPx2_ASAP7_75t_R FILLER_61_342 ();
 FILLER_ASAP7_75t_R FILLER_61_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_350 ();
 DECAPx2_ASAP7_75t_R FILLER_61_373 ();
 FILLER_ASAP7_75t_R FILLER_61_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_381 ();
 DECAPx2_ASAP7_75t_R FILLER_61_388 ();
 FILLER_ASAP7_75t_R FILLER_61_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_418 ();
 DECAPx6_ASAP7_75t_R FILLER_61_425 ();
 DECAPx1_ASAP7_75t_R FILLER_61_439 ();
 DECAPx10_ASAP7_75t_R FILLER_61_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_473 ();
 DECAPx2_ASAP7_75t_R FILLER_61_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_487 ();
 DECAPx6_ASAP7_75t_R FILLER_61_491 ();
 FILLER_ASAP7_75t_R FILLER_61_505 ();
 DECAPx2_ASAP7_75t_R FILLER_61_542 ();
 FILLER_ASAP7_75t_R FILLER_61_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_576 ();
 FILLER_ASAP7_75t_R FILLER_61_580 ();
 DECAPx4_ASAP7_75t_R FILLER_61_586 ();
 DECAPx2_ASAP7_75t_R FILLER_61_608 ();
 FILLER_ASAP7_75t_R FILLER_61_614 ();
 DECAPx4_ASAP7_75t_R FILLER_61_639 ();
 FILLER_ASAP7_75t_R FILLER_61_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_658 ();
 DECAPx6_ASAP7_75t_R FILLER_61_685 ();
 FILLER_ASAP7_75t_R FILLER_61_699 ();
 DECAPx2_ASAP7_75t_R FILLER_61_704 ();
 DECAPx6_ASAP7_75t_R FILLER_61_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_740 ();
 FILLER_ASAP7_75t_R FILLER_61_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_761 ();
 DECAPx1_ASAP7_75t_R FILLER_61_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_778 ();
 FILLER_ASAP7_75t_R FILLER_61_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_795 ();
 FILLER_ASAP7_75t_R FILLER_61_811 ();
 DECAPx4_ASAP7_75t_R FILLER_61_825 ();
 FILLER_ASAP7_75t_R FILLER_61_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_840 ();
 DECAPx2_ASAP7_75t_R FILLER_61_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_865 ();
 DECAPx1_ASAP7_75t_R FILLER_61_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_876 ();
 FILLER_ASAP7_75t_R FILLER_61_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_899 ();
 FILLER_ASAP7_75t_R FILLER_61_912 ();
 DECAPx2_ASAP7_75t_R FILLER_61_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_923 ();
 DECAPx6_ASAP7_75t_R FILLER_61_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_940 ();
 DECAPx6_ASAP7_75t_R FILLER_61_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_987 ();
 DECAPx2_ASAP7_75t_R FILLER_61_995 ();
 FILLER_ASAP7_75t_R FILLER_61_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1083 ();
 FILLER_ASAP7_75t_R FILLER_61_1108 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1128 ();
 FILLER_ASAP7_75t_R FILLER_61_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1352 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1374 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1396 ();
 FILLER_ASAP7_75t_R FILLER_61_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_62_2 ();
 DECAPx4_ASAP7_75t_R FILLER_62_24 ();
 DECAPx4_ASAP7_75t_R FILLER_62_104 ();
 DECAPx1_ASAP7_75t_R FILLER_62_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_124 ();
 FILLER_ASAP7_75t_R FILLER_62_128 ();
 FILLER_ASAP7_75t_R FILLER_62_143 ();
 DECAPx2_ASAP7_75t_R FILLER_62_148 ();
 FILLER_ASAP7_75t_R FILLER_62_174 ();
 DECAPx2_ASAP7_75t_R FILLER_62_218 ();
 FILLER_ASAP7_75t_R FILLER_62_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_226 ();
 DECAPx4_ASAP7_75t_R FILLER_62_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_261 ();
 DECAPx2_ASAP7_75t_R FILLER_62_290 ();
 FILLER_ASAP7_75t_R FILLER_62_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_298 ();
 DECAPx6_ASAP7_75t_R FILLER_62_307 ();
 DECAPx2_ASAP7_75t_R FILLER_62_321 ();
 DECAPx10_ASAP7_75t_R FILLER_62_333 ();
 DECAPx10_ASAP7_75t_R FILLER_62_355 ();
 DECAPx1_ASAP7_75t_R FILLER_62_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_381 ();
 DECAPx2_ASAP7_75t_R FILLER_62_388 ();
 FILLER_ASAP7_75t_R FILLER_62_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_396 ();
 DECAPx4_ASAP7_75t_R FILLER_62_419 ();
 DECAPx6_ASAP7_75t_R FILLER_62_445 ();
 FILLER_ASAP7_75t_R FILLER_62_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_461 ();
 DECAPx4_ASAP7_75t_R FILLER_62_464 ();
 DECAPx1_ASAP7_75t_R FILLER_62_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_529 ();
 DECAPx2_ASAP7_75t_R FILLER_62_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_565 ();
 DECAPx6_ASAP7_75t_R FILLER_62_572 ();
 DECAPx2_ASAP7_75t_R FILLER_62_586 ();
 DECAPx2_ASAP7_75t_R FILLER_62_618 ();
 DECAPx2_ASAP7_75t_R FILLER_62_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_655 ();
 DECAPx1_ASAP7_75t_R FILLER_62_679 ();
 FILLER_ASAP7_75t_R FILLER_62_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_702 ();
 DECAPx1_ASAP7_75t_R FILLER_62_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_734 ();
 DECAPx2_ASAP7_75t_R FILLER_62_741 ();
 FILLER_ASAP7_75t_R FILLER_62_764 ();
 FILLER_ASAP7_75t_R FILLER_62_789 ();
 DECAPx6_ASAP7_75t_R FILLER_62_794 ();
 DECAPx1_ASAP7_75t_R FILLER_62_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_828 ();
 FILLER_ASAP7_75t_R FILLER_62_843 ();
 DECAPx4_ASAP7_75t_R FILLER_62_848 ();
 DECAPx2_ASAP7_75t_R FILLER_62_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_885 ();
 DECAPx1_ASAP7_75t_R FILLER_62_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_900 ();
 DECAPx1_ASAP7_75t_R FILLER_62_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_961 ();
 DECAPx4_ASAP7_75t_R FILLER_62_976 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1016 ();
 FILLER_ASAP7_75t_R FILLER_62_1026 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1036 ();
 FILLER_ASAP7_75t_R FILLER_62_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1093 ();
 FILLER_ASAP7_75t_R FILLER_62_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1115 ();
 FILLER_ASAP7_75t_R FILLER_62_1129 ();
 FILLER_ASAP7_75t_R FILLER_62_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1372 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1388 ();
 FILLER_ASAP7_75t_R FILLER_62_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_63_2 ();
 FILLER_ASAP7_75t_R FILLER_63_78 ();
 DECAPx10_ASAP7_75t_R FILLER_63_86 ();
 DECAPx10_ASAP7_75t_R FILLER_63_108 ();
 DECAPx10_ASAP7_75t_R FILLER_63_130 ();
 DECAPx2_ASAP7_75t_R FILLER_63_152 ();
 FILLER_ASAP7_75t_R FILLER_63_158 ();
 DECAPx2_ASAP7_75t_R FILLER_63_174 ();
 FILLER_ASAP7_75t_R FILLER_63_180 ();
 FILLER_ASAP7_75t_R FILLER_63_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_198 ();
 DECAPx2_ASAP7_75t_R FILLER_63_205 ();
 FILLER_ASAP7_75t_R FILLER_63_211 ();
 FILLER_ASAP7_75t_R FILLER_63_219 ();
 DECAPx6_ASAP7_75t_R FILLER_63_227 ();
 DECAPx1_ASAP7_75t_R FILLER_63_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_258 ();
 DECAPx10_ASAP7_75t_R FILLER_63_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_287 ();
 FILLER_ASAP7_75t_R FILLER_63_302 ();
 DECAPx6_ASAP7_75t_R FILLER_63_311 ();
 DECAPx1_ASAP7_75t_R FILLER_63_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_329 ();
 DECAPx2_ASAP7_75t_R FILLER_63_344 ();
 DECAPx10_ASAP7_75t_R FILLER_63_362 ();
 DECAPx2_ASAP7_75t_R FILLER_63_384 ();
 DECAPx10_ASAP7_75t_R FILLER_63_414 ();
 DECAPx2_ASAP7_75t_R FILLER_63_436 ();
 FILLER_ASAP7_75t_R FILLER_63_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_451 ();
 DECAPx4_ASAP7_75t_R FILLER_63_464 ();
 FILLER_ASAP7_75t_R FILLER_63_474 ();
 DECAPx2_ASAP7_75t_R FILLER_63_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_488 ();
 FILLER_ASAP7_75t_R FILLER_63_511 ();
 DECAPx2_ASAP7_75t_R FILLER_63_522 ();
 FILLER_ASAP7_75t_R FILLER_63_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_530 ();
 DECAPx4_ASAP7_75t_R FILLER_63_557 ();
 FILLER_ASAP7_75t_R FILLER_63_567 ();
 DECAPx2_ASAP7_75t_R FILLER_63_601 ();
 DECAPx6_ASAP7_75t_R FILLER_63_618 ();
 FILLER_ASAP7_75t_R FILLER_63_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_634 ();
 FILLER_ASAP7_75t_R FILLER_63_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_663 ();
 DECAPx4_ASAP7_75t_R FILLER_63_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_677 ();
 DECAPx2_ASAP7_75t_R FILLER_63_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_710 ();
 FILLER_ASAP7_75t_R FILLER_63_717 ();
 DECAPx1_ASAP7_75t_R FILLER_63_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_749 ();
 DECAPx4_ASAP7_75t_R FILLER_63_753 ();
 FILLER_ASAP7_75t_R FILLER_63_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_765 ();
 DECAPx2_ASAP7_75t_R FILLER_63_780 ();
 DECAPx2_ASAP7_75t_R FILLER_63_795 ();
 FILLER_ASAP7_75t_R FILLER_63_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_803 ();
 DECAPx2_ASAP7_75t_R FILLER_63_807 ();
 DECAPx10_ASAP7_75t_R FILLER_63_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_838 ();
 FILLER_ASAP7_75t_R FILLER_63_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_850 ();
 FILLER_ASAP7_75t_R FILLER_63_874 ();
 DECAPx4_ASAP7_75t_R FILLER_63_896 ();
 DECAPx1_ASAP7_75t_R FILLER_63_932 ();
 DECAPx2_ASAP7_75t_R FILLER_63_962 ();
 DECAPx6_ASAP7_75t_R FILLER_63_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_985 ();
 DECAPx2_ASAP7_75t_R FILLER_63_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_63_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1101 ();
 FILLER_ASAP7_75t_R FILLER_63_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1368 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1390 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_64_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_72 ();
 DECAPx1_ASAP7_75t_R FILLER_64_105 ();
 DECAPx2_ASAP7_75t_R FILLER_64_138 ();
 DECAPx4_ASAP7_75t_R FILLER_64_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_167 ();
 DECAPx10_ASAP7_75t_R FILLER_64_176 ();
 DECAPx6_ASAP7_75t_R FILLER_64_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_212 ();
 DECAPx10_ASAP7_75t_R FILLER_64_219 ();
 DECAPx2_ASAP7_75t_R FILLER_64_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_247 ();
 FILLER_ASAP7_75t_R FILLER_64_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_266 ();
 DECAPx2_ASAP7_75t_R FILLER_64_281 ();
 FILLER_ASAP7_75t_R FILLER_64_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_289 ();
 DECAPx2_ASAP7_75t_R FILLER_64_306 ();
 DECAPx10_ASAP7_75t_R FILLER_64_320 ();
 DECAPx2_ASAP7_75t_R FILLER_64_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_356 ();
 DECAPx10_ASAP7_75t_R FILLER_64_365 ();
 DECAPx6_ASAP7_75t_R FILLER_64_387 ();
 DECAPx2_ASAP7_75t_R FILLER_64_401 ();
 DECAPx1_ASAP7_75t_R FILLER_64_413 ();
 DECAPx10_ASAP7_75t_R FILLER_64_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_461 ();
 DECAPx1_ASAP7_75t_R FILLER_64_464 ();
 DECAPx4_ASAP7_75t_R FILLER_64_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_488 ();
 DECAPx6_ASAP7_75t_R FILLER_64_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_539 ();
 DECAPx2_ASAP7_75t_R FILLER_64_549 ();
 FILLER_ASAP7_75t_R FILLER_64_555 ();
 DECAPx1_ASAP7_75t_R FILLER_64_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_571 ();
 DECAPx10_ASAP7_75t_R FILLER_64_594 ();
 DECAPx6_ASAP7_75t_R FILLER_64_616 ();
 DECAPx1_ASAP7_75t_R FILLER_64_630 ();
 FILLER_ASAP7_75t_R FILLER_64_651 ();
 DECAPx2_ASAP7_75t_R FILLER_64_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_671 ();
 DECAPx2_ASAP7_75t_R FILLER_64_681 ();
 FILLER_ASAP7_75t_R FILLER_64_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_689 ();
 DECAPx1_ASAP7_75t_R FILLER_64_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_700 ();
 DECAPx2_ASAP7_75t_R FILLER_64_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_741 ();
 DECAPx10_ASAP7_75t_R FILLER_64_745 ();
 DECAPx6_ASAP7_75t_R FILLER_64_767 ();
 DECAPx1_ASAP7_75t_R FILLER_64_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_785 ();
 DECAPx1_ASAP7_75t_R FILLER_64_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_793 ();
 DECAPx2_ASAP7_75t_R FILLER_64_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_812 ();
 DECAPx1_ASAP7_75t_R FILLER_64_827 ();
 DECAPx10_ASAP7_75t_R FILLER_64_843 ();
 DECAPx4_ASAP7_75t_R FILLER_64_865 ();
 FILLER_ASAP7_75t_R FILLER_64_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_877 ();
 FILLER_ASAP7_75t_R FILLER_64_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_893 ();
 FILLER_ASAP7_75t_R FILLER_64_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_914 ();
 DECAPx1_ASAP7_75t_R FILLER_64_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_922 ();
 DECAPx2_ASAP7_75t_R FILLER_64_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_935 ();
 DECAPx2_ASAP7_75t_R FILLER_64_944 ();
 DECAPx10_ASAP7_75t_R FILLER_64_985 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1007 ();
 FILLER_ASAP7_75t_R FILLER_64_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1061 ();
 FILLER_ASAP7_75t_R FILLER_64_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1143 ();
 FILLER_ASAP7_75t_R FILLER_64_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1388 ();
 FILLER_ASAP7_75t_R FILLER_64_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_65_2 ();
 DECAPx1_ASAP7_75t_R FILLER_65_24 ();
 DECAPx2_ASAP7_75t_R FILLER_65_31 ();
 DECAPx2_ASAP7_75t_R FILLER_65_40 ();
 FILLER_ASAP7_75t_R FILLER_65_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_48 ();
 DECAPx4_ASAP7_75t_R FILLER_65_58 ();
 FILLER_ASAP7_75t_R FILLER_65_68 ();
 FILLER_ASAP7_75t_R FILLER_65_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_75 ();
 DECAPx1_ASAP7_75t_R FILLER_65_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_127 ();
 DECAPx1_ASAP7_75t_R FILLER_65_154 ();
 DECAPx10_ASAP7_75t_R FILLER_65_184 ();
 DECAPx6_ASAP7_75t_R FILLER_65_226 ();
 FILLER_ASAP7_75t_R FILLER_65_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_242 ();
 DECAPx4_ASAP7_75t_R FILLER_65_255 ();
 FILLER_ASAP7_75t_R FILLER_65_265 ();
 DECAPx2_ASAP7_75t_R FILLER_65_281 ();
 FILLER_ASAP7_75t_R FILLER_65_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_302 ();
 DECAPx1_ASAP7_75t_R FILLER_65_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_313 ();
 DECAPx2_ASAP7_75t_R FILLER_65_324 ();
 FILLER_ASAP7_75t_R FILLER_65_330 ();
 DECAPx6_ASAP7_75t_R FILLER_65_340 ();
 DECAPx4_ASAP7_75t_R FILLER_65_360 ();
 DECAPx4_ASAP7_75t_R FILLER_65_376 ();
 FILLER_ASAP7_75t_R FILLER_65_386 ();
 FILLER_ASAP7_75t_R FILLER_65_400 ();
 DECAPx6_ASAP7_75t_R FILLER_65_418 ();
 FILLER_ASAP7_75t_R FILLER_65_432 ();
 DECAPx10_ASAP7_75t_R FILLER_65_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_470 ();
 FILLER_ASAP7_75t_R FILLER_65_485 ();
 FILLER_ASAP7_75t_R FILLER_65_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_527 ();
 DECAPx2_ASAP7_75t_R FILLER_65_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_541 ();
 FILLER_ASAP7_75t_R FILLER_65_545 ();
 DECAPx2_ASAP7_75t_R FILLER_65_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_563 ();
 DECAPx4_ASAP7_75t_R FILLER_65_570 ();
 FILLER_ASAP7_75t_R FILLER_65_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_582 ();
 DECAPx1_ASAP7_75t_R FILLER_65_603 ();
 FILLER_ASAP7_75t_R FILLER_65_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_635 ();
 DECAPx2_ASAP7_75t_R FILLER_65_642 ();
 FILLER_ASAP7_75t_R FILLER_65_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_650 ();
 DECAPx10_ASAP7_75t_R FILLER_65_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_702 ();
 DECAPx10_ASAP7_75t_R FILLER_65_706 ();
 DECAPx6_ASAP7_75t_R FILLER_65_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_756 ();
 DECAPx1_ASAP7_75t_R FILLER_65_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_776 ();
 FILLER_ASAP7_75t_R FILLER_65_780 ();
 DECAPx2_ASAP7_75t_R FILLER_65_791 ();
 FILLER_ASAP7_75t_R FILLER_65_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_799 ();
 DECAPx6_ASAP7_75t_R FILLER_65_812 ();
 FILLER_ASAP7_75t_R FILLER_65_826 ();
 DECAPx6_ASAP7_75t_R FILLER_65_849 ();
 DECAPx1_ASAP7_75t_R FILLER_65_894 ();
 DECAPx1_ASAP7_75t_R FILLER_65_912 ();
 DECAPx1_ASAP7_75t_R FILLER_65_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_938 ();
 DECAPx1_ASAP7_75t_R FILLER_65_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_949 ();
 DECAPx10_ASAP7_75t_R FILLER_65_960 ();
 FILLER_ASAP7_75t_R FILLER_65_982 ();
 DECAPx10_ASAP7_75t_R FILLER_65_997 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1092 ();
 FILLER_ASAP7_75t_R FILLER_65_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1121 ();
 FILLER_ASAP7_75t_R FILLER_65_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1147 ();
 FILLER_ASAP7_75t_R FILLER_65_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1386 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1404 ();
 FILLER_ASAP7_75t_R FILLER_66_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_40 ();
 DECAPx2_ASAP7_75t_R FILLER_66_70 ();
 DECAPx1_ASAP7_75t_R FILLER_66_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_86 ();
 DECAPx2_ASAP7_75t_R FILLER_66_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_96 ();
 DECAPx2_ASAP7_75t_R FILLER_66_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_112 ();
 DECAPx6_ASAP7_75t_R FILLER_66_122 ();
 DECAPx2_ASAP7_75t_R FILLER_66_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_146 ();
 DECAPx2_ASAP7_75t_R FILLER_66_154 ();
 FILLER_ASAP7_75t_R FILLER_66_160 ();
 FILLER_ASAP7_75t_R FILLER_66_190 ();
 FILLER_ASAP7_75t_R FILLER_66_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_228 ();
 DECAPx10_ASAP7_75t_R FILLER_66_259 ();
 DECAPx10_ASAP7_75t_R FILLER_66_281 ();
 DECAPx10_ASAP7_75t_R FILLER_66_303 ();
 DECAPx2_ASAP7_75t_R FILLER_66_325 ();
 FILLER_ASAP7_75t_R FILLER_66_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_333 ();
 DECAPx4_ASAP7_75t_R FILLER_66_340 ();
 FILLER_ASAP7_75t_R FILLER_66_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_352 ();
 DECAPx4_ASAP7_75t_R FILLER_66_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_371 ();
 FILLER_ASAP7_75t_R FILLER_66_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_382 ();
 DECAPx10_ASAP7_75t_R FILLER_66_389 ();
 DECAPx1_ASAP7_75t_R FILLER_66_411 ();
 DECAPx2_ASAP7_75t_R FILLER_66_421 ();
 DECAPx10_ASAP7_75t_R FILLER_66_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_461 ();
 DECAPx2_ASAP7_75t_R FILLER_66_476 ();
 FILLER_ASAP7_75t_R FILLER_66_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_484 ();
 DECAPx6_ASAP7_75t_R FILLER_66_491 ();
 DECAPx1_ASAP7_75t_R FILLER_66_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_509 ();
 DECAPx4_ASAP7_75t_R FILLER_66_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_526 ();
 DECAPx1_ASAP7_75t_R FILLER_66_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_616 ();
 FILLER_ASAP7_75t_R FILLER_66_623 ();
 FILLER_ASAP7_75t_R FILLER_66_628 ();
 DECAPx2_ASAP7_75t_R FILLER_66_638 ();
 FILLER_ASAP7_75t_R FILLER_66_644 ();
 DECAPx2_ASAP7_75t_R FILLER_66_649 ();
 DECAPx2_ASAP7_75t_R FILLER_66_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_664 ();
 FILLER_ASAP7_75t_R FILLER_66_682 ();
 DECAPx6_ASAP7_75t_R FILLER_66_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_717 ();
 DECAPx1_ASAP7_75t_R FILLER_66_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_725 ();
 DECAPx2_ASAP7_75t_R FILLER_66_729 ();
 FILLER_ASAP7_75t_R FILLER_66_735 ();
 FILLER_ASAP7_75t_R FILLER_66_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_759 ();
 DECAPx2_ASAP7_75t_R FILLER_66_769 ();
 FILLER_ASAP7_75t_R FILLER_66_775 ();
 FILLER_ASAP7_75t_R FILLER_66_780 ();
 FILLER_ASAP7_75t_R FILLER_66_794 ();
 DECAPx1_ASAP7_75t_R FILLER_66_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_814 ();
 FILLER_ASAP7_75t_R FILLER_66_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_837 ();
 FILLER_ASAP7_75t_R FILLER_66_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_871 ();
 DECAPx10_ASAP7_75t_R FILLER_66_878 ();
 DECAPx10_ASAP7_75t_R FILLER_66_900 ();
 DECAPx2_ASAP7_75t_R FILLER_66_922 ();
 FILLER_ASAP7_75t_R FILLER_66_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_938 ();
 DECAPx10_ASAP7_75t_R FILLER_66_945 ();
 DECAPx4_ASAP7_75t_R FILLER_66_987 ();
 FILLER_ASAP7_75t_R FILLER_66_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_999 ();
 FILLER_ASAP7_75t_R FILLER_66_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1018 ();
 FILLER_ASAP7_75t_R FILLER_66_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1076 ();
 FILLER_ASAP7_75t_R FILLER_66_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1159 ();
 FILLER_ASAP7_75t_R FILLER_66_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1388 ();
 FILLER_ASAP7_75t_R FILLER_66_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_67_2 ();
 FILLER_ASAP7_75t_R FILLER_67_44 ();
 DECAPx4_ASAP7_75t_R FILLER_67_84 ();
 DECAPx1_ASAP7_75t_R FILLER_67_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_130 ();
 DECAPx1_ASAP7_75t_R FILLER_67_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_167 ();
 DECAPx1_ASAP7_75t_R FILLER_67_174 ();
 DECAPx1_ASAP7_75t_R FILLER_67_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_232 ();
 DECAPx6_ASAP7_75t_R FILLER_67_239 ();
 DECAPx1_ASAP7_75t_R FILLER_67_253 ();
 DECAPx6_ASAP7_75t_R FILLER_67_263 ();
 DECAPx2_ASAP7_75t_R FILLER_67_277 ();
 DECAPx10_ASAP7_75t_R FILLER_67_297 ();
 DECAPx4_ASAP7_75t_R FILLER_67_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_329 ();
 DECAPx1_ASAP7_75t_R FILLER_67_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_369 ();
 DECAPx4_ASAP7_75t_R FILLER_67_382 ();
 DECAPx10_ASAP7_75t_R FILLER_67_398 ();
 FILLER_ASAP7_75t_R FILLER_67_420 ();
 DECAPx6_ASAP7_75t_R FILLER_67_428 ();
 DECAPx2_ASAP7_75t_R FILLER_67_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_448 ();
 FILLER_ASAP7_75t_R FILLER_67_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_469 ();
 FILLER_ASAP7_75t_R FILLER_67_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_478 ();
 DECAPx2_ASAP7_75t_R FILLER_67_485 ();
 FILLER_ASAP7_75t_R FILLER_67_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_493 ();
 DECAPx4_ASAP7_75t_R FILLER_67_514 ();
 FILLER_ASAP7_75t_R FILLER_67_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_526 ();
 DECAPx2_ASAP7_75t_R FILLER_67_539 ();
 FILLER_ASAP7_75t_R FILLER_67_545 ();
 DECAPx4_ASAP7_75t_R FILLER_67_555 ();
 FILLER_ASAP7_75t_R FILLER_67_565 ();
 DECAPx2_ASAP7_75t_R FILLER_67_626 ();
 FILLER_ASAP7_75t_R FILLER_67_632 ();
 DECAPx4_ASAP7_75t_R FILLER_67_637 ();
 FILLER_ASAP7_75t_R FILLER_67_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_663 ();
 DECAPx1_ASAP7_75t_R FILLER_67_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_705 ();
 DECAPx1_ASAP7_75t_R FILLER_67_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_722 ();
 DECAPx2_ASAP7_75t_R FILLER_67_737 ();
 FILLER_ASAP7_75t_R FILLER_67_743 ();
 DECAPx1_ASAP7_75t_R FILLER_67_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_764 ();
 FILLER_ASAP7_75t_R FILLER_67_794 ();
 DECAPx6_ASAP7_75t_R FILLER_67_805 ();
 FILLER_ASAP7_75t_R FILLER_67_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_821 ();
 DECAPx6_ASAP7_75t_R FILLER_67_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_850 ();
 FILLER_ASAP7_75t_R FILLER_67_866 ();
 DECAPx2_ASAP7_75t_R FILLER_67_888 ();
 DECAPx2_ASAP7_75t_R FILLER_67_918 ();
 DECAPx4_ASAP7_75t_R FILLER_67_926 ();
 FILLER_ASAP7_75t_R FILLER_67_936 ();
 DECAPx1_ASAP7_75t_R FILLER_67_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_964 ();
 DECAPx1_ASAP7_75t_R FILLER_67_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_979 ();
 DECAPx1_ASAP7_75t_R FILLER_67_990 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1025 ();
 FILLER_ASAP7_75t_R FILLER_67_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1121 ();
 FILLER_ASAP7_75t_R FILLER_67_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1129 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1138 ();
 FILLER_ASAP7_75t_R FILLER_67_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1154 ();
 FILLER_ASAP7_75t_R FILLER_67_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1397 ();
 FILLER_ASAP7_75t_R FILLER_67_1403 ();
 DECAPx4_ASAP7_75t_R FILLER_68_2 ();
 FILLER_ASAP7_75t_R FILLER_68_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_14 ();
 FILLER_ASAP7_75t_R FILLER_68_18 ();
 FILLER_ASAP7_75t_R FILLER_68_34 ();
 DECAPx1_ASAP7_75t_R FILLER_68_42 ();
 FILLER_ASAP7_75t_R FILLER_68_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_54 ();
 DECAPx2_ASAP7_75t_R FILLER_68_58 ();
 FILLER_ASAP7_75t_R FILLER_68_70 ();
 DECAPx2_ASAP7_75t_R FILLER_68_75 ();
 FILLER_ASAP7_75t_R FILLER_68_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_86 ();
 DECAPx6_ASAP7_75t_R FILLER_68_90 ();
 DECAPx1_ASAP7_75t_R FILLER_68_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_108 ();
 DECAPx2_ASAP7_75t_R FILLER_68_112 ();
 FILLER_ASAP7_75t_R FILLER_68_118 ();
 FILLER_ASAP7_75t_R FILLER_68_126 ();
 DECAPx4_ASAP7_75t_R FILLER_68_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_144 ();
 DECAPx10_ASAP7_75t_R FILLER_68_148 ();
 DECAPx6_ASAP7_75t_R FILLER_68_170 ();
 DECAPx2_ASAP7_75t_R FILLER_68_184 ();
 DECAPx2_ASAP7_75t_R FILLER_68_204 ();
 FILLER_ASAP7_75t_R FILLER_68_210 ();
 DECAPx4_ASAP7_75t_R FILLER_68_218 ();
 FILLER_ASAP7_75t_R FILLER_68_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_230 ();
 DECAPx6_ASAP7_75t_R FILLER_68_239 ();
 DECAPx4_ASAP7_75t_R FILLER_68_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_271 ();
 DECAPx6_ASAP7_75t_R FILLER_68_286 ();
 DECAPx2_ASAP7_75t_R FILLER_68_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_306 ();
 DECAPx6_ASAP7_75t_R FILLER_68_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_345 ();
 FILLER_ASAP7_75t_R FILLER_68_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_354 ();
 DECAPx1_ASAP7_75t_R FILLER_68_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_371 ();
 FILLER_ASAP7_75t_R FILLER_68_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_382 ();
 DECAPx2_ASAP7_75t_R FILLER_68_414 ();
 FILLER_ASAP7_75t_R FILLER_68_420 ();
 DECAPx4_ASAP7_75t_R FILLER_68_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_446 ();
 DECAPx1_ASAP7_75t_R FILLER_68_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_461 ();
 DECAPx1_ASAP7_75t_R FILLER_68_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_476 ();
 DECAPx1_ASAP7_75t_R FILLER_68_519 ();
 DECAPx10_ASAP7_75t_R FILLER_68_529 ();
 DECAPx4_ASAP7_75t_R FILLER_68_551 ();
 FILLER_ASAP7_75t_R FILLER_68_561 ();
 DECAPx1_ASAP7_75t_R FILLER_68_589 ();
 FILLER_ASAP7_75t_R FILLER_68_605 ();
 DECAPx2_ASAP7_75t_R FILLER_68_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_651 ();
 DECAPx1_ASAP7_75t_R FILLER_68_661 ();
 DECAPx2_ASAP7_75t_R FILLER_68_679 ();
 FILLER_ASAP7_75t_R FILLER_68_685 ();
 DECAPx1_ASAP7_75t_R FILLER_68_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_700 ();
 FILLER_ASAP7_75t_R FILLER_68_721 ();
 FILLER_ASAP7_75t_R FILLER_68_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_739 ();
 DECAPx4_ASAP7_75t_R FILLER_68_749 ();
 FILLER_ASAP7_75t_R FILLER_68_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_761 ();
 DECAPx10_ASAP7_75t_R FILLER_68_776 ();
 DECAPx4_ASAP7_75t_R FILLER_68_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_840 ();
 DECAPx6_ASAP7_75t_R FILLER_68_848 ();
 DECAPx2_ASAP7_75t_R FILLER_68_870 ();
 FILLER_ASAP7_75t_R FILLER_68_876 ();
 FILLER_ASAP7_75t_R FILLER_68_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_894 ();
 DECAPx2_ASAP7_75t_R FILLER_68_917 ();
 FILLER_ASAP7_75t_R FILLER_68_923 ();
 DECAPx1_ASAP7_75t_R FILLER_68_941 ();
 FILLER_ASAP7_75t_R FILLER_68_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_953 ();
 DECAPx2_ASAP7_75t_R FILLER_68_962 ();
 DECAPx1_ASAP7_75t_R FILLER_68_981 ();
 DECAPx1_ASAP7_75t_R FILLER_68_991 ();
 FILLER_ASAP7_75t_R FILLER_68_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1022 ();
 FILLER_ASAP7_75t_R FILLER_68_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1079 ();
 FILLER_ASAP7_75t_R FILLER_68_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1098 ();
 FILLER_ASAP7_75t_R FILLER_68_1104 ();
 FILLER_ASAP7_75t_R FILLER_68_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1141 ();
 FILLER_ASAP7_75t_R FILLER_68_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1370 ();
 FILLER_ASAP7_75t_R FILLER_68_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1388 ();
 FILLER_ASAP7_75t_R FILLER_68_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_69_2 ();
 DECAPx2_ASAP7_75t_R FILLER_69_24 ();
 FILLER_ASAP7_75t_R FILLER_69_30 ();
 DECAPx4_ASAP7_75t_R FILLER_69_35 ();
 DECAPx6_ASAP7_75t_R FILLER_69_48 ();
 DECAPx1_ASAP7_75t_R FILLER_69_68 ();
 DECAPx6_ASAP7_75t_R FILLER_69_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_112 ();
 DECAPx2_ASAP7_75t_R FILLER_69_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_145 ();
 DECAPx10_ASAP7_75t_R FILLER_69_172 ();
 FILLER_ASAP7_75t_R FILLER_69_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_196 ();
 DECAPx10_ASAP7_75t_R FILLER_69_203 ();
 DECAPx6_ASAP7_75t_R FILLER_69_225 ();
 DECAPx1_ASAP7_75t_R FILLER_69_245 ();
 DECAPx10_ASAP7_75t_R FILLER_69_269 ();
 DECAPx6_ASAP7_75t_R FILLER_69_291 ();
 DECAPx1_ASAP7_75t_R FILLER_69_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_309 ();
 DECAPx10_ASAP7_75t_R FILLER_69_326 ();
 DECAPx10_ASAP7_75t_R FILLER_69_348 ();
 DECAPx1_ASAP7_75t_R FILLER_69_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_374 ();
 DECAPx6_ASAP7_75t_R FILLER_69_381 ();
 DECAPx2_ASAP7_75t_R FILLER_69_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_401 ();
 DECAPx6_ASAP7_75t_R FILLER_69_416 ();
 DECAPx1_ASAP7_75t_R FILLER_69_430 ();
 DECAPx1_ASAP7_75t_R FILLER_69_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_444 ();
 DECAPx2_ASAP7_75t_R FILLER_69_466 ();
 FILLER_ASAP7_75t_R FILLER_69_472 ();
 DECAPx2_ASAP7_75t_R FILLER_69_488 ();
 DECAPx4_ASAP7_75t_R FILLER_69_514 ();
 FILLER_ASAP7_75t_R FILLER_69_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_526 ();
 DECAPx1_ASAP7_75t_R FILLER_69_539 ();
 FILLER_ASAP7_75t_R FILLER_69_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_561 ();
 FILLER_ASAP7_75t_R FILLER_69_575 ();
 DECAPx1_ASAP7_75t_R FILLER_69_606 ();
 FILLER_ASAP7_75t_R FILLER_69_628 ();
 DECAPx10_ASAP7_75t_R FILLER_69_656 ();
 DECAPx4_ASAP7_75t_R FILLER_69_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_688 ();
 DECAPx2_ASAP7_75t_R FILLER_69_695 ();
 FILLER_ASAP7_75t_R FILLER_69_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_703 ();
 FILLER_ASAP7_75t_R FILLER_69_718 ();
 FILLER_ASAP7_75t_R FILLER_69_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_740 ();
 DECAPx4_ASAP7_75t_R FILLER_69_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_754 ();
 DECAPx2_ASAP7_75t_R FILLER_69_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_776 ();
 DECAPx2_ASAP7_75t_R FILLER_69_780 ();
 FILLER_ASAP7_75t_R FILLER_69_786 ();
 DECAPx1_ASAP7_75t_R FILLER_69_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_798 ();
 DECAPx10_ASAP7_75t_R FILLER_69_806 ();
 DECAPx4_ASAP7_75t_R FILLER_69_828 ();
 FILLER_ASAP7_75t_R FILLER_69_838 ();
 DECAPx4_ASAP7_75t_R FILLER_69_867 ();
 FILLER_ASAP7_75t_R FILLER_69_877 ();
 DECAPx1_ASAP7_75t_R FILLER_69_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_892 ();
 DECAPx4_ASAP7_75t_R FILLER_69_899 ();
 FILLER_ASAP7_75t_R FILLER_69_909 ();
 DECAPx1_ASAP7_75t_R FILLER_69_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_930 ();
 DECAPx2_ASAP7_75t_R FILLER_69_939 ();
 FILLER_ASAP7_75t_R FILLER_69_945 ();
 DECAPx2_ASAP7_75t_R FILLER_69_961 ();
 DECAPx2_ASAP7_75t_R FILLER_69_973 ();
 FILLER_ASAP7_75t_R FILLER_69_979 ();
 DECAPx6_ASAP7_75t_R FILLER_69_991 ();
 FILLER_ASAP7_75t_R FILLER_69_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1022 ();
 FILLER_ASAP7_75t_R FILLER_69_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1060 ();
 FILLER_ASAP7_75t_R FILLER_69_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1124 ();
 FILLER_ASAP7_75t_R FILLER_69_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1397 ();
 FILLER_ASAP7_75t_R FILLER_69_1403 ();
 DECAPx4_ASAP7_75t_R FILLER_70_2 ();
 FILLER_ASAP7_75t_R FILLER_70_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_18 ();
 DECAPx1_ASAP7_75t_R FILLER_70_29 ();
 FILLER_ASAP7_75t_R FILLER_70_62 ();
 FILLER_ASAP7_75t_R FILLER_70_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_110 ();
 DECAPx1_ASAP7_75t_R FILLER_70_123 ();
 FILLER_ASAP7_75t_R FILLER_70_139 ();
 FILLER_ASAP7_75t_R FILLER_70_147 ();
 DECAPx2_ASAP7_75t_R FILLER_70_182 ();
 DECAPx2_ASAP7_75t_R FILLER_70_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_214 ();
 DECAPx2_ASAP7_75t_R FILLER_70_221 ();
 FILLER_ASAP7_75t_R FILLER_70_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_236 ();
 DECAPx6_ASAP7_75t_R FILLER_70_257 ();
 FILLER_ASAP7_75t_R FILLER_70_271 ();
 FILLER_ASAP7_75t_R FILLER_70_307 ();
 DECAPx6_ASAP7_75t_R FILLER_70_317 ();
 FILLER_ASAP7_75t_R FILLER_70_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_333 ();
 DECAPx10_ASAP7_75t_R FILLER_70_342 ();
 DECAPx10_ASAP7_75t_R FILLER_70_364 ();
 DECAPx10_ASAP7_75t_R FILLER_70_386 ();
 DECAPx6_ASAP7_75t_R FILLER_70_408 ();
 FILLER_ASAP7_75t_R FILLER_70_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_424 ();
 DECAPx6_ASAP7_75t_R FILLER_70_445 ();
 FILLER_ASAP7_75t_R FILLER_70_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_461 ();
 DECAPx10_ASAP7_75t_R FILLER_70_464 ();
 DECAPx10_ASAP7_75t_R FILLER_70_486 ();
 DECAPx6_ASAP7_75t_R FILLER_70_508 ();
 DECAPx2_ASAP7_75t_R FILLER_70_522 ();
 FILLER_ASAP7_75t_R FILLER_70_548 ();
 DECAPx10_ASAP7_75t_R FILLER_70_566 ();
 DECAPx2_ASAP7_75t_R FILLER_70_588 ();
 DECAPx4_ASAP7_75t_R FILLER_70_597 ();
 FILLER_ASAP7_75t_R FILLER_70_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_643 ();
 DECAPx6_ASAP7_75t_R FILLER_70_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_661 ();
 DECAPx2_ASAP7_75t_R FILLER_70_665 ();
 DECAPx1_ASAP7_75t_R FILLER_70_674 ();
 DECAPx10_ASAP7_75t_R FILLER_70_692 ();
 DECAPx4_ASAP7_75t_R FILLER_70_714 ();
 FILLER_ASAP7_75t_R FILLER_70_724 ();
 DECAPx1_ASAP7_75t_R FILLER_70_738 ();
 FILLER_ASAP7_75t_R FILLER_70_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_747 ();
 DECAPx1_ASAP7_75t_R FILLER_70_800 ();
 DECAPx1_ASAP7_75t_R FILLER_70_827 ();
 DECAPx4_ASAP7_75t_R FILLER_70_843 ();
 FILLER_ASAP7_75t_R FILLER_70_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_855 ();
 FILLER_ASAP7_75t_R FILLER_70_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_868 ();
 DECAPx4_ASAP7_75t_R FILLER_70_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_899 ();
 DECAPx4_ASAP7_75t_R FILLER_70_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_918 ();
 FILLER_ASAP7_75t_R FILLER_70_932 ();
 DECAPx4_ASAP7_75t_R FILLER_70_950 ();
 FILLER_ASAP7_75t_R FILLER_70_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_962 ();
 DECAPx1_ASAP7_75t_R FILLER_70_969 ();
 DECAPx10_ASAP7_75t_R FILLER_70_996 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1057 ();
 FILLER_ASAP7_75t_R FILLER_70_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1121 ();
 FILLER_ASAP7_75t_R FILLER_70_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1129 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1187 ();
 FILLER_ASAP7_75t_R FILLER_70_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1352 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1374 ();
 FILLER_ASAP7_75t_R FILLER_70_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1388 ();
 FILLER_ASAP7_75t_R FILLER_70_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_71_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_52 ();
 DECAPx2_ASAP7_75t_R FILLER_71_152 ();
 FILLER_ASAP7_75t_R FILLER_71_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_160 ();
 FILLER_ASAP7_75t_R FILLER_71_164 ();
 FILLER_ASAP7_75t_R FILLER_71_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_181 ();
 FILLER_ASAP7_75t_R FILLER_71_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_215 ();
 DECAPx4_ASAP7_75t_R FILLER_71_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_260 ();
 DECAPx4_ASAP7_75t_R FILLER_71_271 ();
 FILLER_ASAP7_75t_R FILLER_71_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_283 ();
 DECAPx10_ASAP7_75t_R FILLER_71_290 ();
 DECAPx2_ASAP7_75t_R FILLER_71_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_318 ();
 DECAPx2_ASAP7_75t_R FILLER_71_327 ();
 DECAPx2_ASAP7_75t_R FILLER_71_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_365 ();
 DECAPx10_ASAP7_75t_R FILLER_71_379 ();
 DECAPx10_ASAP7_75t_R FILLER_71_401 ();
 DECAPx2_ASAP7_75t_R FILLER_71_423 ();
 FILLER_ASAP7_75t_R FILLER_71_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_431 ();
 DECAPx6_ASAP7_75t_R FILLER_71_438 ();
 DECAPx6_ASAP7_75t_R FILLER_71_466 ();
 DECAPx1_ASAP7_75t_R FILLER_71_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_484 ();
 DECAPx10_ASAP7_75t_R FILLER_71_497 ();
 DECAPx10_ASAP7_75t_R FILLER_71_519 ();
 DECAPx2_ASAP7_75t_R FILLER_71_541 ();
 FILLER_ASAP7_75t_R FILLER_71_547 ();
 DECAPx4_ASAP7_75t_R FILLER_71_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_571 ();
 DECAPx2_ASAP7_75t_R FILLER_71_578 ();
 FILLER_ASAP7_75t_R FILLER_71_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_586 ();
 DECAPx10_ASAP7_75t_R FILLER_71_590 ();
 DECAPx4_ASAP7_75t_R FILLER_71_612 ();
 FILLER_ASAP7_75t_R FILLER_71_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_624 ();
 DECAPx6_ASAP7_75t_R FILLER_71_635 ();
 FILLER_ASAP7_75t_R FILLER_71_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_651 ();
 DECAPx2_ASAP7_75t_R FILLER_71_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_661 ();
 FILLER_ASAP7_75t_R FILLER_71_674 ();
 DECAPx4_ASAP7_75t_R FILLER_71_696 ();
 FILLER_ASAP7_75t_R FILLER_71_706 ();
 DECAPx2_ASAP7_75t_R FILLER_71_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_727 ();
 FILLER_ASAP7_75t_R FILLER_71_742 ();
 FILLER_ASAP7_75t_R FILLER_71_753 ();
 DECAPx4_ASAP7_75t_R FILLER_71_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_777 ();
 DECAPx2_ASAP7_75t_R FILLER_71_795 ();
 FILLER_ASAP7_75t_R FILLER_71_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_803 ();
 DECAPx4_ASAP7_75t_R FILLER_71_811 ();
 FILLER_ASAP7_75t_R FILLER_71_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_849 ();
 DECAPx6_ASAP7_75t_R FILLER_71_880 ();
 DECAPx2_ASAP7_75t_R FILLER_71_894 ();
 FILLER_ASAP7_75t_R FILLER_71_922 ();
 DECAPx2_ASAP7_75t_R FILLER_71_934 ();
 FILLER_ASAP7_75t_R FILLER_71_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_969 ();
 FILLER_ASAP7_75t_R FILLER_71_983 ();
 DECAPx6_ASAP7_75t_R FILLER_71_992 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1040 ();
 FILLER_ASAP7_75t_R FILLER_71_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1077 ();
 FILLER_ASAP7_75t_R FILLER_71_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1159 ();
 FILLER_ASAP7_75t_R FILLER_71_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1368 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1390 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_72_2 ();
 FILLER_ASAP7_75t_R FILLER_72_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_14 ();
 DECAPx2_ASAP7_75t_R FILLER_72_41 ();
 DECAPx2_ASAP7_75t_R FILLER_72_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_56 ();
 DECAPx1_ASAP7_75t_R FILLER_72_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_67 ();
 DECAPx2_ASAP7_75t_R FILLER_72_101 ();
 DECAPx1_ASAP7_75t_R FILLER_72_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_117 ();
 DECAPx10_ASAP7_75t_R FILLER_72_121 ();
 DECAPx10_ASAP7_75t_R FILLER_72_143 ();
 DECAPx1_ASAP7_75t_R FILLER_72_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_169 ();
 DECAPx2_ASAP7_75t_R FILLER_72_173 ();
 DECAPx2_ASAP7_75t_R FILLER_72_185 ();
 FILLER_ASAP7_75t_R FILLER_72_191 ();
 DECAPx1_ASAP7_75t_R FILLER_72_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_209 ();
 DECAPx6_ASAP7_75t_R FILLER_72_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_230 ();
 DECAPx10_ASAP7_75t_R FILLER_72_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_267 ();
 DECAPx10_ASAP7_75t_R FILLER_72_275 ();
 DECAPx10_ASAP7_75t_R FILLER_72_297 ();
 FILLER_ASAP7_75t_R FILLER_72_319 ();
 DECAPx10_ASAP7_75t_R FILLER_72_330 ();
 DECAPx2_ASAP7_75t_R FILLER_72_352 ();
 FILLER_ASAP7_75t_R FILLER_72_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_360 ();
 DECAPx1_ASAP7_75t_R FILLER_72_374 ();
 FILLER_ASAP7_75t_R FILLER_72_405 ();
 DECAPx1_ASAP7_75t_R FILLER_72_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_419 ();
 FILLER_ASAP7_75t_R FILLER_72_430 ();
 DECAPx4_ASAP7_75t_R FILLER_72_440 ();
 DECAPx2_ASAP7_75t_R FILLER_72_472 ();
 FILLER_ASAP7_75t_R FILLER_72_478 ();
 DECAPx10_ASAP7_75t_R FILLER_72_494 ();
 DECAPx2_ASAP7_75t_R FILLER_72_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_522 ();
 DECAPx10_ASAP7_75t_R FILLER_72_533 ();
 DECAPx4_ASAP7_75t_R FILLER_72_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_565 ();
 DECAPx2_ASAP7_75t_R FILLER_72_607 ();
 DECAPx10_ASAP7_75t_R FILLER_72_619 ();
 FILLER_ASAP7_75t_R FILLER_72_641 ();
 DECAPx1_ASAP7_75t_R FILLER_72_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_672 ();
 DECAPx1_ASAP7_75t_R FILLER_72_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_700 ();
 FILLER_ASAP7_75t_R FILLER_72_715 ();
 FILLER_ASAP7_75t_R FILLER_72_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_754 ();
 DECAPx10_ASAP7_75t_R FILLER_72_758 ();
 DECAPx1_ASAP7_75t_R FILLER_72_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_784 ();
 DECAPx6_ASAP7_75t_R FILLER_72_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_806 ();
 DECAPx1_ASAP7_75t_R FILLER_72_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_837 ();
 DECAPx2_ASAP7_75t_R FILLER_72_841 ();
 DECAPx4_ASAP7_75t_R FILLER_72_852 ();
 FILLER_ASAP7_75t_R FILLER_72_862 ();
 DECAPx1_ASAP7_75t_R FILLER_72_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_876 ();
 DECAPx2_ASAP7_75t_R FILLER_72_889 ();
 FILLER_ASAP7_75t_R FILLER_72_895 ();
 DECAPx10_ASAP7_75t_R FILLER_72_915 ();
 DECAPx6_ASAP7_75t_R FILLER_72_937 ();
 DECAPx1_ASAP7_75t_R FILLER_72_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_955 ();
 DECAPx10_ASAP7_75t_R FILLER_72_963 ();
 DECAPx6_ASAP7_75t_R FILLER_72_985 ();
 DECAPx2_ASAP7_75t_R FILLER_72_999 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1023 ();
 FILLER_ASAP7_75t_R FILLER_72_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1046 ();
 FILLER_ASAP7_75t_R FILLER_72_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1086 ();
 FILLER_ASAP7_75t_R FILLER_72_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1113 ();
 FILLER_ASAP7_75t_R FILLER_72_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1362 ();
 FILLER_ASAP7_75t_R FILLER_72_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1388 ();
 FILLER_ASAP7_75t_R FILLER_72_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_73_2 ();
 DECAPx1_ASAP7_75t_R FILLER_73_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_27 ();
 FILLER_ASAP7_75t_R FILLER_73_37 ();
 DECAPx1_ASAP7_75t_R FILLER_73_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_52 ();
 DECAPx10_ASAP7_75t_R FILLER_73_59 ();
 DECAPx6_ASAP7_75t_R FILLER_73_107 ();
 FILLER_ASAP7_75t_R FILLER_73_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_123 ();
 DECAPx2_ASAP7_75t_R FILLER_73_130 ();
 FILLER_ASAP7_75t_R FILLER_73_139 ();
 FILLER_ASAP7_75t_R FILLER_73_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_149 ();
 DECAPx1_ASAP7_75t_R FILLER_73_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_161 ();
 DECAPx6_ASAP7_75t_R FILLER_73_165 ();
 FILLER_ASAP7_75t_R FILLER_73_179 ();
 DECAPx10_ASAP7_75t_R FILLER_73_189 ();
 DECAPx2_ASAP7_75t_R FILLER_73_211 ();
 FILLER_ASAP7_75t_R FILLER_73_217 ();
 DECAPx6_ASAP7_75t_R FILLER_73_233 ();
 DECAPx1_ASAP7_75t_R FILLER_73_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_251 ();
 DECAPx1_ASAP7_75t_R FILLER_73_258 ();
 DECAPx10_ASAP7_75t_R FILLER_73_294 ();
 DECAPx1_ASAP7_75t_R FILLER_73_316 ();
 DECAPx10_ASAP7_75t_R FILLER_73_326 ();
 FILLER_ASAP7_75t_R FILLER_73_348 ();
 DECAPx10_ASAP7_75t_R FILLER_73_356 ();
 DECAPx10_ASAP7_75t_R FILLER_73_378 ();
 DECAPx1_ASAP7_75t_R FILLER_73_400 ();
 DECAPx10_ASAP7_75t_R FILLER_73_412 ();
 DECAPx6_ASAP7_75t_R FILLER_73_434 ();
 FILLER_ASAP7_75t_R FILLER_73_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_450 ();
 DECAPx4_ASAP7_75t_R FILLER_73_457 ();
 FILLER_ASAP7_75t_R FILLER_73_467 ();
 DECAPx2_ASAP7_75t_R FILLER_73_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_487 ();
 DECAPx1_ASAP7_75t_R FILLER_73_497 ();
 FILLER_ASAP7_75t_R FILLER_73_517 ();
 DECAPx1_ASAP7_75t_R FILLER_73_537 ();
 FILLER_ASAP7_75t_R FILLER_73_547 ();
 DECAPx2_ASAP7_75t_R FILLER_73_555 ();
 FILLER_ASAP7_75t_R FILLER_73_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_605 ();
 DECAPx4_ASAP7_75t_R FILLER_73_670 ();
 FILLER_ASAP7_75t_R FILLER_73_680 ();
 FILLER_ASAP7_75t_R FILLER_73_691 ();
 FILLER_ASAP7_75t_R FILLER_73_696 ();
 DECAPx2_ASAP7_75t_R FILLER_73_722 ();
 FILLER_ASAP7_75t_R FILLER_73_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_730 ();
 DECAPx10_ASAP7_75t_R FILLER_73_740 ();
 DECAPx2_ASAP7_75t_R FILLER_73_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_768 ();
 DECAPx10_ASAP7_75t_R FILLER_73_779 ();
 FILLER_ASAP7_75t_R FILLER_73_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_803 ();
 FILLER_ASAP7_75t_R FILLER_73_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_827 ();
 FILLER_ASAP7_75t_R FILLER_73_842 ();
 DECAPx1_ASAP7_75t_R FILLER_73_858 ();
 FILLER_ASAP7_75t_R FILLER_73_868 ();
 DECAPx1_ASAP7_75t_R FILLER_73_884 ();
 DECAPx6_ASAP7_75t_R FILLER_73_899 ();
 DECAPx1_ASAP7_75t_R FILLER_73_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_926 ();
 DECAPx10_ASAP7_75t_R FILLER_73_943 ();
 FILLER_ASAP7_75t_R FILLER_73_975 ();
 DECAPx6_ASAP7_75t_R FILLER_73_985 ();
 FILLER_ASAP7_75t_R FILLER_73_999 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1058 ();
 FILLER_ASAP7_75t_R FILLER_73_1064 ();
 FILLER_ASAP7_75t_R FILLER_73_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1100 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1160 ();
 FILLER_ASAP7_75t_R FILLER_73_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1168 ();
 FILLER_ASAP7_75t_R FILLER_73_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1357 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1379 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1401 ();
 DECAPx6_ASAP7_75t_R FILLER_74_2 ();
 DECAPx1_ASAP7_75t_R FILLER_74_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_20 ();
 DECAPx4_ASAP7_75t_R FILLER_74_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_37 ();
 FILLER_ASAP7_75t_R FILLER_74_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_79 ();
 DECAPx1_ASAP7_75t_R FILLER_74_92 ();
 DECAPx2_ASAP7_75t_R FILLER_74_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_105 ();
 DECAPx2_ASAP7_75t_R FILLER_74_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_184 ();
 DECAPx1_ASAP7_75t_R FILLER_74_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_199 ();
 DECAPx6_ASAP7_75t_R FILLER_74_206 ();
 DECAPx1_ASAP7_75t_R FILLER_74_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_246 ();
 DECAPx2_ASAP7_75t_R FILLER_74_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_275 ();
 DECAPx1_ASAP7_75t_R FILLER_74_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_295 ();
 DECAPx4_ASAP7_75t_R FILLER_74_329 ();
 DECAPx6_ASAP7_75t_R FILLER_74_361 ();
 DECAPx2_ASAP7_75t_R FILLER_74_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_381 ();
 DECAPx4_ASAP7_75t_R FILLER_74_396 ();
 DECAPx2_ASAP7_75t_R FILLER_74_415 ();
 FILLER_ASAP7_75t_R FILLER_74_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_423 ();
 DECAPx6_ASAP7_75t_R FILLER_74_438 ();
 DECAPx1_ASAP7_75t_R FILLER_74_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_470 ();
 DECAPx2_ASAP7_75t_R FILLER_74_477 ();
 FILLER_ASAP7_75t_R FILLER_74_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_485 ();
 DECAPx10_ASAP7_75t_R FILLER_74_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_518 ();
 DECAPx1_ASAP7_75t_R FILLER_74_535 ();
 FILLER_ASAP7_75t_R FILLER_74_549 ();
 DECAPx2_ASAP7_75t_R FILLER_74_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_567 ();
 DECAPx2_ASAP7_75t_R FILLER_74_575 ();
 FILLER_ASAP7_75t_R FILLER_74_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_583 ();
 DECAPx6_ASAP7_75t_R FILLER_74_587 ();
 DECAPx2_ASAP7_75t_R FILLER_74_636 ();
 FILLER_ASAP7_75t_R FILLER_74_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_644 ();
 DECAPx6_ASAP7_75t_R FILLER_74_662 ();
 DECAPx1_ASAP7_75t_R FILLER_74_676 ();
 DECAPx1_ASAP7_75t_R FILLER_74_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_699 ();
 DECAPx10_ASAP7_75t_R FILLER_74_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_736 ();
 DECAPx6_ASAP7_75t_R FILLER_74_740 ();
 DECAPx2_ASAP7_75t_R FILLER_74_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_780 ();
 FILLER_ASAP7_75t_R FILLER_74_787 ();
 DECAPx10_ASAP7_75t_R FILLER_74_828 ();
 DECAPx4_ASAP7_75t_R FILLER_74_850 ();
 DECAPx6_ASAP7_75t_R FILLER_74_866 ();
 FILLER_ASAP7_75t_R FILLER_74_880 ();
 DECAPx1_ASAP7_75t_R FILLER_74_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_892 ();
 FILLER_ASAP7_75t_R FILLER_74_910 ();
 DECAPx2_ASAP7_75t_R FILLER_74_918 ();
 DECAPx2_ASAP7_75t_R FILLER_74_954 ();
 FILLER_ASAP7_75t_R FILLER_74_972 ();
 DECAPx2_ASAP7_75t_R FILLER_74_981 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1128 ();
 FILLER_ASAP7_75t_R FILLER_74_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1175 ();
 FILLER_ASAP7_75t_R FILLER_74_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1388 ();
 FILLER_ASAP7_75t_R FILLER_74_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_75_37 ();
 FILLER_ASAP7_75t_R FILLER_75_51 ();
 FILLER_ASAP7_75t_R FILLER_75_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_58 ();
 DECAPx6_ASAP7_75t_R FILLER_75_88 ();
 DECAPx10_ASAP7_75t_R FILLER_75_128 ();
 DECAPx2_ASAP7_75t_R FILLER_75_150 ();
 DECAPx6_ASAP7_75t_R FILLER_75_162 ();
 FILLER_ASAP7_75t_R FILLER_75_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_178 ();
 DECAPx1_ASAP7_75t_R FILLER_75_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_225 ();
 DECAPx10_ASAP7_75t_R FILLER_75_232 ();
 DECAPx1_ASAP7_75t_R FILLER_75_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_258 ();
 DECAPx4_ASAP7_75t_R FILLER_75_265 ();
 FILLER_ASAP7_75t_R FILLER_75_275 ();
 DECAPx10_ASAP7_75t_R FILLER_75_291 ();
 FILLER_ASAP7_75t_R FILLER_75_313 ();
 DECAPx10_ASAP7_75t_R FILLER_75_321 ();
 DECAPx10_ASAP7_75t_R FILLER_75_343 ();
 DECAPx6_ASAP7_75t_R FILLER_75_365 ();
 FILLER_ASAP7_75t_R FILLER_75_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_381 ();
 DECAPx10_ASAP7_75t_R FILLER_75_388 ();
 DECAPx6_ASAP7_75t_R FILLER_75_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_424 ();
 DECAPx10_ASAP7_75t_R FILLER_75_439 ();
 DECAPx4_ASAP7_75t_R FILLER_75_475 ();
 FILLER_ASAP7_75t_R FILLER_75_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_487 ();
 DECAPx10_ASAP7_75t_R FILLER_75_500 ();
 DECAPx4_ASAP7_75t_R FILLER_75_522 ();
 FILLER_ASAP7_75t_R FILLER_75_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_534 ();
 DECAPx10_ASAP7_75t_R FILLER_75_547 ();
 DECAPx1_ASAP7_75t_R FILLER_75_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_573 ();
 DECAPx4_ASAP7_75t_R FILLER_75_580 ();
 DECAPx4_ASAP7_75t_R FILLER_75_593 ();
 FILLER_ASAP7_75t_R FILLER_75_603 ();
 DECAPx4_ASAP7_75t_R FILLER_75_611 ();
 DECAPx2_ASAP7_75t_R FILLER_75_624 ();
 FILLER_ASAP7_75t_R FILLER_75_630 ();
 DECAPx10_ASAP7_75t_R FILLER_75_638 ();
 DECAPx10_ASAP7_75t_R FILLER_75_660 ();
 DECAPx6_ASAP7_75t_R FILLER_75_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_696 ();
 DECAPx10_ASAP7_75t_R FILLER_75_705 ();
 DECAPx10_ASAP7_75t_R FILLER_75_727 ();
 DECAPx2_ASAP7_75t_R FILLER_75_749 ();
 FILLER_ASAP7_75t_R FILLER_75_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_757 ();
 FILLER_ASAP7_75t_R FILLER_75_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_766 ();
 DECAPx1_ASAP7_75t_R FILLER_75_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_778 ();
 DECAPx6_ASAP7_75t_R FILLER_75_797 ();
 DECAPx6_ASAP7_75t_R FILLER_75_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_831 ();
 DECAPx4_ASAP7_75t_R FILLER_75_839 ();
 FILLER_ASAP7_75t_R FILLER_75_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_851 ();
 DECAPx1_ASAP7_75t_R FILLER_75_862 ();
 DECAPx1_ASAP7_75t_R FILLER_75_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_876 ();
 FILLER_ASAP7_75t_R FILLER_75_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_892 ();
 DECAPx1_ASAP7_75t_R FILLER_75_899 ();
 DECAPx1_ASAP7_75t_R FILLER_75_909 ();
 FILLER_ASAP7_75t_R FILLER_75_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_923 ();
 FILLER_ASAP7_75t_R FILLER_75_926 ();
 DECAPx1_ASAP7_75t_R FILLER_75_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_938 ();
 DECAPx1_ASAP7_75t_R FILLER_75_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_946 ();
 DECAPx6_ASAP7_75t_R FILLER_75_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_975 ();
 DECAPx4_ASAP7_75t_R FILLER_75_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_999 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1028 ();
 FILLER_ASAP7_75t_R FILLER_75_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1077 ();
 FILLER_ASAP7_75t_R FILLER_75_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1386 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_76_34 ();
 DECAPx6_ASAP7_75t_R FILLER_76_50 ();
 FILLER_ASAP7_75t_R FILLER_76_64 ();
 DECAPx1_ASAP7_75t_R FILLER_76_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_106 ();
 DECAPx2_ASAP7_75t_R FILLER_76_145 ();
 FILLER_ASAP7_75t_R FILLER_76_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_160 ();
 FILLER_ASAP7_75t_R FILLER_76_167 ();
 DECAPx4_ASAP7_75t_R FILLER_76_176 ();
 FILLER_ASAP7_75t_R FILLER_76_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_188 ();
 DECAPx6_ASAP7_75t_R FILLER_76_223 ();
 DECAPx1_ASAP7_75t_R FILLER_76_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_241 ();
 DECAPx10_ASAP7_75t_R FILLER_76_248 ();
 DECAPx2_ASAP7_75t_R FILLER_76_270 ();
 FILLER_ASAP7_75t_R FILLER_76_276 ();
 DECAPx4_ASAP7_75t_R FILLER_76_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_296 ();
 FILLER_ASAP7_75t_R FILLER_76_304 ();
 DECAPx1_ASAP7_75t_R FILLER_76_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_316 ();
 DECAPx1_ASAP7_75t_R FILLER_76_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_327 ();
 DECAPx4_ASAP7_75t_R FILLER_76_334 ();
 FILLER_ASAP7_75t_R FILLER_76_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_346 ();
 DECAPx10_ASAP7_75t_R FILLER_76_353 ();
 DECAPx10_ASAP7_75t_R FILLER_76_375 ();
 DECAPx1_ASAP7_75t_R FILLER_76_397 ();
 DECAPx2_ASAP7_75t_R FILLER_76_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_415 ();
 DECAPx6_ASAP7_75t_R FILLER_76_426 ();
 FILLER_ASAP7_75t_R FILLER_76_440 ();
 DECAPx4_ASAP7_75t_R FILLER_76_450 ();
 FILLER_ASAP7_75t_R FILLER_76_460 ();
 DECAPx4_ASAP7_75t_R FILLER_76_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_488 ();
 DECAPx10_ASAP7_75t_R FILLER_76_501 ();
 DECAPx2_ASAP7_75t_R FILLER_76_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_529 ();
 DECAPx4_ASAP7_75t_R FILLER_76_542 ();
 DECAPx4_ASAP7_75t_R FILLER_76_558 ();
 DECAPx2_ASAP7_75t_R FILLER_76_601 ();
 FILLER_ASAP7_75t_R FILLER_76_607 ();
 DECAPx6_ASAP7_75t_R FILLER_76_612 ();
 DECAPx1_ASAP7_75t_R FILLER_76_626 ();
 DECAPx4_ASAP7_75t_R FILLER_76_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_666 ();
 DECAPx10_ASAP7_75t_R FILLER_76_670 ();
 FILLER_ASAP7_75t_R FILLER_76_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_694 ();
 DECAPx4_ASAP7_75t_R FILLER_76_703 ();
 FILLER_ASAP7_75t_R FILLER_76_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_715 ();
 FILLER_ASAP7_75t_R FILLER_76_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_757 ();
 FILLER_ASAP7_75t_R FILLER_76_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_773 ();
 DECAPx2_ASAP7_75t_R FILLER_76_781 ();
 FILLER_ASAP7_75t_R FILLER_76_797 ();
 DECAPx2_ASAP7_75t_R FILLER_76_807 ();
 FILLER_ASAP7_75t_R FILLER_76_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_815 ();
 FILLER_ASAP7_75t_R FILLER_76_864 ();
 FILLER_ASAP7_75t_R FILLER_76_894 ();
 FILLER_ASAP7_75t_R FILLER_76_910 ();
 DECAPx2_ASAP7_75t_R FILLER_76_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_924 ();
 DECAPx2_ASAP7_75t_R FILLER_76_932 ();
 DECAPx6_ASAP7_75t_R FILLER_76_945 ();
 FILLER_ASAP7_75t_R FILLER_76_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_961 ();
 DECAPx6_ASAP7_75t_R FILLER_76_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_989 ();
 DECAPx2_ASAP7_75t_R FILLER_76_996 ();
 FILLER_ASAP7_75t_R FILLER_76_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1066 ();
 FILLER_ASAP7_75t_R FILLER_76_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1112 ();
 FILLER_ASAP7_75t_R FILLER_76_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1377 ();
 FILLER_ASAP7_75t_R FILLER_76_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1388 ();
 FILLER_ASAP7_75t_R FILLER_76_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_77_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_23 ();
 FILLER_ASAP7_75t_R FILLER_77_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_73 ();
 DECAPx2_ASAP7_75t_R FILLER_77_80 ();
 FILLER_ASAP7_75t_R FILLER_77_92 ();
 DECAPx2_ASAP7_75t_R FILLER_77_97 ();
 DECAPx4_ASAP7_75t_R FILLER_77_106 ();
 FILLER_ASAP7_75t_R FILLER_77_116 ();
 FILLER_ASAP7_75t_R FILLER_77_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_137 ();
 DECAPx1_ASAP7_75t_R FILLER_77_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_200 ();
 DECAPx10_ASAP7_75t_R FILLER_77_207 ();
 DECAPx1_ASAP7_75t_R FILLER_77_229 ();
 FILLER_ASAP7_75t_R FILLER_77_255 ();
 FILLER_ASAP7_75t_R FILLER_77_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_265 ();
 DECAPx4_ASAP7_75t_R FILLER_77_280 ();
 DECAPx1_ASAP7_75t_R FILLER_77_316 ();
 DECAPx4_ASAP7_75t_R FILLER_77_328 ();
 FILLER_ASAP7_75t_R FILLER_77_338 ();
 FILLER_ASAP7_75t_R FILLER_77_348 ();
 DECAPx2_ASAP7_75t_R FILLER_77_356 ();
 DECAPx10_ASAP7_75t_R FILLER_77_376 ();
 DECAPx2_ASAP7_75t_R FILLER_77_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_404 ();
 DECAPx6_ASAP7_75t_R FILLER_77_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_438 ();
 FILLER_ASAP7_75t_R FILLER_77_458 ();
 DECAPx2_ASAP7_75t_R FILLER_77_478 ();
 FILLER_ASAP7_75t_R FILLER_77_484 ();
 DECAPx6_ASAP7_75t_R FILLER_77_492 ();
 DECAPx2_ASAP7_75t_R FILLER_77_506 ();
 DECAPx2_ASAP7_75t_R FILLER_77_526 ();
 FILLER_ASAP7_75t_R FILLER_77_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_545 ();
 DECAPx10_ASAP7_75t_R FILLER_77_562 ();
 DECAPx1_ASAP7_75t_R FILLER_77_584 ();
 DECAPx1_ASAP7_75t_R FILLER_77_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_625 ();
 FILLER_ASAP7_75t_R FILLER_77_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_631 ();
 DECAPx1_ASAP7_75t_R FILLER_77_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_642 ();
 DECAPx6_ASAP7_75t_R FILLER_77_678 ();
 FILLER_ASAP7_75t_R FILLER_77_692 ();
 DECAPx6_ASAP7_75t_R FILLER_77_706 ();
 DECAPx1_ASAP7_75t_R FILLER_77_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_741 ();
 DECAPx4_ASAP7_75t_R FILLER_77_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_759 ();
 FILLER_ASAP7_75t_R FILLER_77_768 ();
 DECAPx2_ASAP7_75t_R FILLER_77_788 ();
 FILLER_ASAP7_75t_R FILLER_77_794 ();
 DECAPx4_ASAP7_75t_R FILLER_77_816 ();
 FILLER_ASAP7_75t_R FILLER_77_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_828 ();
 DECAPx10_ASAP7_75t_R FILLER_77_839 ();
 DECAPx2_ASAP7_75t_R FILLER_77_867 ();
 FILLER_ASAP7_75t_R FILLER_77_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_875 ();
 DECAPx1_ASAP7_75t_R FILLER_77_882 ();
 DECAPx4_ASAP7_75t_R FILLER_77_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_910 ();
 DECAPx1_ASAP7_75t_R FILLER_77_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_923 ();
 DECAPx6_ASAP7_75t_R FILLER_77_934 ();
 FILLER_ASAP7_75t_R FILLER_77_948 ();
 DECAPx6_ASAP7_75t_R FILLER_77_970 ();
 DECAPx1_ASAP7_75t_R FILLER_77_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_988 ();
 FILLER_ASAP7_75t_R FILLER_77_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1040 ();
 FILLER_ASAP7_75t_R FILLER_77_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1348 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1370 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1392 ();
 FILLER_ASAP7_75t_R FILLER_77_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_78_2 ();
 DECAPx10_ASAP7_75t_R FILLER_78_24 ();
 DECAPx2_ASAP7_75t_R FILLER_78_55 ();
 FILLER_ASAP7_75t_R FILLER_78_61 ();
 DECAPx2_ASAP7_75t_R FILLER_78_89 ();
 DECAPx1_ASAP7_75t_R FILLER_78_101 ();
 FILLER_ASAP7_75t_R FILLER_78_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_137 ();
 DECAPx2_ASAP7_75t_R FILLER_78_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_147 ();
 FILLER_ASAP7_75t_R FILLER_78_155 ();
 DECAPx6_ASAP7_75t_R FILLER_78_160 ();
 DECAPx1_ASAP7_75t_R FILLER_78_174 ();
 DECAPx4_ASAP7_75t_R FILLER_78_181 ();
 FILLER_ASAP7_75t_R FILLER_78_191 ();
 DECAPx6_ASAP7_75t_R FILLER_78_199 ();
 DECAPx1_ASAP7_75t_R FILLER_78_213 ();
 DECAPx1_ASAP7_75t_R FILLER_78_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_271 ();
 FILLER_ASAP7_75t_R FILLER_78_280 ();
 DECAPx6_ASAP7_75t_R FILLER_78_288 ();
 FILLER_ASAP7_75t_R FILLER_78_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_304 ();
 DECAPx1_ASAP7_75t_R FILLER_78_308 ();
 DECAPx6_ASAP7_75t_R FILLER_78_318 ();
 DECAPx2_ASAP7_75t_R FILLER_78_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_338 ();
 DECAPx10_ASAP7_75t_R FILLER_78_345 ();
 FILLER_ASAP7_75t_R FILLER_78_367 ();
 DECAPx4_ASAP7_75t_R FILLER_78_375 ();
 FILLER_ASAP7_75t_R FILLER_78_399 ();
 DECAPx4_ASAP7_75t_R FILLER_78_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_442 ();
 DECAPx2_ASAP7_75t_R FILLER_78_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_461 ();
 DECAPx1_ASAP7_75t_R FILLER_78_464 ();
 FILLER_ASAP7_75t_R FILLER_78_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_478 ();
 DECAPx2_ASAP7_75t_R FILLER_78_496 ();
 DECAPx10_ASAP7_75t_R FILLER_78_508 ();
 DECAPx4_ASAP7_75t_R FILLER_78_530 ();
 FILLER_ASAP7_75t_R FILLER_78_540 ();
 DECAPx2_ASAP7_75t_R FILLER_78_554 ();
 FILLER_ASAP7_75t_R FILLER_78_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_562 ();
 FILLER_ASAP7_75t_R FILLER_78_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_584 ();
 DECAPx1_ASAP7_75t_R FILLER_78_588 ();
 DECAPx2_ASAP7_75t_R FILLER_78_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_604 ();
 DECAPx2_ASAP7_75t_R FILLER_78_637 ();
 FILLER_ASAP7_75t_R FILLER_78_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_645 ();
 FILLER_ASAP7_75t_R FILLER_78_653 ();
 DECAPx2_ASAP7_75t_R FILLER_78_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_667 ();
 DECAPx1_ASAP7_75t_R FILLER_78_684 ();
 FILLER_ASAP7_75t_R FILLER_78_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_710 ();
 DECAPx4_ASAP7_75t_R FILLER_78_725 ();
 FILLER_ASAP7_75t_R FILLER_78_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_744 ();
 DECAPx4_ASAP7_75t_R FILLER_78_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_768 ();
 DECAPx4_ASAP7_75t_R FILLER_78_781 ();
 FILLER_ASAP7_75t_R FILLER_78_791 ();
 DECAPx2_ASAP7_75t_R FILLER_78_799 ();
 FILLER_ASAP7_75t_R FILLER_78_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_807 ();
 FILLER_ASAP7_75t_R FILLER_78_813 ();
 DECAPx10_ASAP7_75t_R FILLER_78_838 ();
 DECAPx1_ASAP7_75t_R FILLER_78_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_864 ();
 DECAPx10_ASAP7_75t_R FILLER_78_879 ();
 DECAPx2_ASAP7_75t_R FILLER_78_901 ();
 FILLER_ASAP7_75t_R FILLER_78_907 ();
 DECAPx2_ASAP7_75t_R FILLER_78_913 ();
 FILLER_ASAP7_75t_R FILLER_78_919 ();
 FILLER_ASAP7_75t_R FILLER_78_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_956 ();
 FILLER_ASAP7_75t_R FILLER_78_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_963 ();
 FILLER_ASAP7_75t_R FILLER_78_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_972 ();
 DECAPx6_ASAP7_75t_R FILLER_78_987 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1011 ();
 FILLER_ASAP7_75t_R FILLER_78_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1025 ();
 FILLER_ASAP7_75t_R FILLER_78_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1039 ();
 FILLER_ASAP7_75t_R FILLER_78_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1069 ();
 FILLER_ASAP7_75t_R FILLER_78_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1083 ();
 FILLER_ASAP7_75t_R FILLER_78_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1128 ();
 FILLER_ASAP7_75t_R FILLER_78_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1160 ();
 FILLER_ASAP7_75t_R FILLER_78_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1188 ();
 FILLER_ASAP7_75t_R FILLER_78_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_78_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1388 ();
 FILLER_ASAP7_75t_R FILLER_78_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_79_2 ();
 FILLER_ASAP7_75t_R FILLER_79_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_18 ();
 FILLER_ASAP7_75t_R FILLER_79_33 ();
 DECAPx4_ASAP7_75t_R FILLER_79_64 ();
 FILLER_ASAP7_75t_R FILLER_79_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_76 ();
 FILLER_ASAP7_75t_R FILLER_79_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_116 ();
 DECAPx2_ASAP7_75t_R FILLER_79_123 ();
 FILLER_ASAP7_75t_R FILLER_79_129 ();
 DECAPx4_ASAP7_75t_R FILLER_79_176 ();
 FILLER_ASAP7_75t_R FILLER_79_186 ();
 FILLER_ASAP7_75t_R FILLER_79_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_204 ();
 DECAPx2_ASAP7_75t_R FILLER_79_212 ();
 DECAPx1_ASAP7_75t_R FILLER_79_232 ();
 DECAPx4_ASAP7_75t_R FILLER_79_242 ();
 DECAPx4_ASAP7_75t_R FILLER_79_258 ();
 DECAPx2_ASAP7_75t_R FILLER_79_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_280 ();
 DECAPx10_ASAP7_75t_R FILLER_79_287 ();
 DECAPx2_ASAP7_75t_R FILLER_79_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_315 ();
 DECAPx10_ASAP7_75t_R FILLER_79_330 ();
 DECAPx10_ASAP7_75t_R FILLER_79_352 ();
 DECAPx10_ASAP7_75t_R FILLER_79_374 ();
 DECAPx10_ASAP7_75t_R FILLER_79_396 ();
 DECAPx10_ASAP7_75t_R FILLER_79_418 ();
 DECAPx1_ASAP7_75t_R FILLER_79_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_444 ();
 DECAPx10_ASAP7_75t_R FILLER_79_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_473 ();
 DECAPx10_ASAP7_75t_R FILLER_79_482 ();
 DECAPx10_ASAP7_75t_R FILLER_79_504 ();
 FILLER_ASAP7_75t_R FILLER_79_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_528 ();
 FILLER_ASAP7_75t_R FILLER_79_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_562 ();
 DECAPx2_ASAP7_75t_R FILLER_79_606 ();
 DECAPx10_ASAP7_75t_R FILLER_79_618 ();
 DECAPx4_ASAP7_75t_R FILLER_79_640 ();
 FILLER_ASAP7_75t_R FILLER_79_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_652 ();
 FILLER_ASAP7_75t_R FILLER_79_656 ();
 FILLER_ASAP7_75t_R FILLER_79_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_663 ();
 DECAPx6_ASAP7_75t_R FILLER_79_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_688 ();
 DECAPx1_ASAP7_75t_R FILLER_79_709 ();
 DECAPx6_ASAP7_75t_R FILLER_79_725 ();
 FILLER_ASAP7_75t_R FILLER_79_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_749 ();
 DECAPx6_ASAP7_75t_R FILLER_79_770 ();
 DECAPx1_ASAP7_75t_R FILLER_79_797 ();
 FILLER_ASAP7_75t_R FILLER_79_809 ();
 DECAPx6_ASAP7_75t_R FILLER_79_814 ();
 DECAPx1_ASAP7_75t_R FILLER_79_828 ();
 DECAPx2_ASAP7_75t_R FILLER_79_837 ();
 DECAPx6_ASAP7_75t_R FILLER_79_846 ();
 FILLER_ASAP7_75t_R FILLER_79_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_862 ();
 DECAPx10_ASAP7_75t_R FILLER_79_869 ();
 DECAPx10_ASAP7_75t_R FILLER_79_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_913 ();
 FILLER_ASAP7_75t_R FILLER_79_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_968 ();
 DECAPx6_ASAP7_75t_R FILLER_79_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_991 ();
 DECAPx10_ASAP7_75t_R FILLER_79_998 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1020 ();
 FILLER_ASAP7_75t_R FILLER_79_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1045 ();
 FILLER_ASAP7_75t_R FILLER_79_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1165 ();
 FILLER_ASAP7_75t_R FILLER_79_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1192 ();
 FILLER_ASAP7_75t_R FILLER_79_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1358 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1380 ();
 FILLER_ASAP7_75t_R FILLER_79_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_80_2 ();
 FILLER_ASAP7_75t_R FILLER_80_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_10 ();
 DECAPx4_ASAP7_75t_R FILLER_80_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_43 ();
 DECAPx2_ASAP7_75t_R FILLER_80_53 ();
 FILLER_ASAP7_75t_R FILLER_80_88 ();
 DECAPx4_ASAP7_75t_R FILLER_80_96 ();
 FILLER_ASAP7_75t_R FILLER_80_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_108 ();
 DECAPx2_ASAP7_75t_R FILLER_80_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_121 ();
 FILLER_ASAP7_75t_R FILLER_80_131 ();
 DECAPx1_ASAP7_75t_R FILLER_80_211 ();
 DECAPx2_ASAP7_75t_R FILLER_80_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_243 ();
 DECAPx10_ASAP7_75t_R FILLER_80_250 ();
 DECAPx2_ASAP7_75t_R FILLER_80_272 ();
 DECAPx10_ASAP7_75t_R FILLER_80_292 ();
 FILLER_ASAP7_75t_R FILLER_80_314 ();
 DECAPx10_ASAP7_75t_R FILLER_80_348 ();
 DECAPx6_ASAP7_75t_R FILLER_80_370 ();
 DECAPx1_ASAP7_75t_R FILLER_80_384 ();
 DECAPx6_ASAP7_75t_R FILLER_80_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_408 ();
 DECAPx10_ASAP7_75t_R FILLER_80_415 ();
 DECAPx2_ASAP7_75t_R FILLER_80_437 ();
 FILLER_ASAP7_75t_R FILLER_80_443 ();
 DECAPx1_ASAP7_75t_R FILLER_80_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_461 ();
 DECAPx6_ASAP7_75t_R FILLER_80_464 ();
 DECAPx4_ASAP7_75t_R FILLER_80_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_497 ();
 DECAPx2_ASAP7_75t_R FILLER_80_506 ();
 DECAPx4_ASAP7_75t_R FILLER_80_529 ();
 FILLER_ASAP7_75t_R FILLER_80_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_541 ();
 DECAPx2_ASAP7_75t_R FILLER_80_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_558 ();
 DECAPx1_ASAP7_75t_R FILLER_80_568 ();
 DECAPx2_ASAP7_75t_R FILLER_80_598 ();
 FILLER_ASAP7_75t_R FILLER_80_604 ();
 DECAPx6_ASAP7_75t_R FILLER_80_670 ();
 DECAPx2_ASAP7_75t_R FILLER_80_684 ();
 FILLER_ASAP7_75t_R FILLER_80_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_733 ();
 DECAPx2_ASAP7_75t_R FILLER_80_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_746 ();
 DECAPx6_ASAP7_75t_R FILLER_80_753 ();
 FILLER_ASAP7_75t_R FILLER_80_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_769 ();
 DECAPx2_ASAP7_75t_R FILLER_80_787 ();
 FILLER_ASAP7_75t_R FILLER_80_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_795 ();
 DECAPx2_ASAP7_75t_R FILLER_80_822 ();
 FILLER_ASAP7_75t_R FILLER_80_880 ();
 DECAPx4_ASAP7_75t_R FILLER_80_912 ();
 DECAPx1_ASAP7_75t_R FILLER_80_933 ();
 DECAPx10_ASAP7_75t_R FILLER_80_940 ();
 DECAPx4_ASAP7_75t_R FILLER_80_962 ();
 FILLER_ASAP7_75t_R FILLER_80_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_982 ();
 FILLER_ASAP7_75t_R FILLER_80_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_991 ();
 FILLER_ASAP7_75t_R FILLER_80_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1023 ();
 FILLER_ASAP7_75t_R FILLER_80_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1077 ();
 FILLER_ASAP7_75t_R FILLER_80_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1154 ();
 FILLER_ASAP7_75t_R FILLER_80_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1388 ();
 FILLER_ASAP7_75t_R FILLER_80_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_81_2 ();
 FILLER_ASAP7_75t_R FILLER_81_8 ();
 FILLER_ASAP7_75t_R FILLER_81_45 ();
 FILLER_ASAP7_75t_R FILLER_81_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_55 ();
 DECAPx1_ASAP7_75t_R FILLER_81_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_63 ();
 FILLER_ASAP7_75t_R FILLER_81_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_78 ();
 DECAPx1_ASAP7_75t_R FILLER_81_105 ();
 DECAPx6_ASAP7_75t_R FILLER_81_115 ();
 DECAPx1_ASAP7_75t_R FILLER_81_129 ();
 FILLER_ASAP7_75t_R FILLER_81_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_149 ();
 DECAPx6_ASAP7_75t_R FILLER_81_156 ();
 DECAPx1_ASAP7_75t_R FILLER_81_170 ();
 DECAPx4_ASAP7_75t_R FILLER_81_177 ();
 DECAPx1_ASAP7_75t_R FILLER_81_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_231 ();
 DECAPx10_ASAP7_75t_R FILLER_81_254 ();
 DECAPx10_ASAP7_75t_R FILLER_81_276 ();
 DECAPx2_ASAP7_75t_R FILLER_81_298 ();
 DECAPx4_ASAP7_75t_R FILLER_81_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_320 ();
 FILLER_ASAP7_75t_R FILLER_81_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_361 ();
 FILLER_ASAP7_75t_R FILLER_81_368 ();
 DECAPx2_ASAP7_75t_R FILLER_81_376 ();
 DECAPx6_ASAP7_75t_R FILLER_81_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_434 ();
 FILLER_ASAP7_75t_R FILLER_81_460 ();
 DECAPx10_ASAP7_75t_R FILLER_81_468 ();
 FILLER_ASAP7_75t_R FILLER_81_496 ();
 FILLER_ASAP7_75t_R FILLER_81_504 ();
 DECAPx6_ASAP7_75t_R FILLER_81_513 ();
 FILLER_ASAP7_75t_R FILLER_81_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_529 ();
 DECAPx10_ASAP7_75t_R FILLER_81_537 ();
 DECAPx10_ASAP7_75t_R FILLER_81_559 ();
 DECAPx2_ASAP7_75t_R FILLER_81_581 ();
 DECAPx6_ASAP7_75t_R FILLER_81_590 ();
 DECAPx1_ASAP7_75t_R FILLER_81_604 ();
 DECAPx6_ASAP7_75t_R FILLER_81_658 ();
 DECAPx1_ASAP7_75t_R FILLER_81_672 ();
 FILLER_ASAP7_75t_R FILLER_81_682 ();
 DECAPx4_ASAP7_75t_R FILLER_81_705 ();
 FILLER_ASAP7_75t_R FILLER_81_715 ();
 DECAPx1_ASAP7_75t_R FILLER_81_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_734 ();
 DECAPx6_ASAP7_75t_R FILLER_81_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_765 ();
 DECAPx4_ASAP7_75t_R FILLER_81_785 ();
 FILLER_ASAP7_75t_R FILLER_81_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_797 ();
 DECAPx2_ASAP7_75t_R FILLER_81_812 ();
 FILLER_ASAP7_75t_R FILLER_81_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_820 ();
 DECAPx6_ASAP7_75t_R FILLER_81_829 ();
 FILLER_ASAP7_75t_R FILLER_81_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_901 ();
 DECAPx4_ASAP7_75t_R FILLER_81_914 ();
 DECAPx4_ASAP7_75t_R FILLER_81_926 ();
 FILLER_ASAP7_75t_R FILLER_81_936 ();
 DECAPx4_ASAP7_75t_R FILLER_81_941 ();
 FILLER_ASAP7_75t_R FILLER_81_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_953 ();
 DECAPx2_ASAP7_75t_R FILLER_81_962 ();
 FILLER_ASAP7_75t_R FILLER_81_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1060 ();
 FILLER_ASAP7_75t_R FILLER_81_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1088 ();
 FILLER_ASAP7_75t_R FILLER_81_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1113 ();
 FILLER_ASAP7_75t_R FILLER_81_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1145 ();
 FILLER_ASAP7_75t_R FILLER_81_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1163 ();
 FILLER_ASAP7_75t_R FILLER_81_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_82_2 ();
 DECAPx1_ASAP7_75t_R FILLER_82_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_31 ();
 FILLER_ASAP7_75t_R FILLER_82_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_40 ();
 DECAPx2_ASAP7_75t_R FILLER_82_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_73 ();
 DECAPx6_ASAP7_75t_R FILLER_82_77 ();
 FILLER_ASAP7_75t_R FILLER_82_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_93 ();
 DECAPx1_ASAP7_75t_R FILLER_82_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_101 ();
 DECAPx2_ASAP7_75t_R FILLER_82_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_134 ();
 DECAPx6_ASAP7_75t_R FILLER_82_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_175 ();
 DECAPx10_ASAP7_75t_R FILLER_82_183 ();
 DECAPx10_ASAP7_75t_R FILLER_82_205 ();
 DECAPx2_ASAP7_75t_R FILLER_82_255 ();
 FILLER_ASAP7_75t_R FILLER_82_261 ();
 DECAPx1_ASAP7_75t_R FILLER_82_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_281 ();
 DECAPx4_ASAP7_75t_R FILLER_82_290 ();
 FILLER_ASAP7_75t_R FILLER_82_300 ();
 DECAPx10_ASAP7_75t_R FILLER_82_316 ();
 DECAPx10_ASAP7_75t_R FILLER_82_338 ();
 DECAPx10_ASAP7_75t_R FILLER_82_374 ();
 DECAPx10_ASAP7_75t_R FILLER_82_396 ();
 FILLER_ASAP7_75t_R FILLER_82_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_441 ();
 DECAPx1_ASAP7_75t_R FILLER_82_458 ();
 FILLER_ASAP7_75t_R FILLER_82_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_466 ();
 DECAPx4_ASAP7_75t_R FILLER_82_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_492 ();
 DECAPx1_ASAP7_75t_R FILLER_82_501 ();
 DECAPx2_ASAP7_75t_R FILLER_82_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_563 ();
 DECAPx10_ASAP7_75t_R FILLER_82_590 ();
 DECAPx6_ASAP7_75t_R FILLER_82_612 ();
 DECAPx1_ASAP7_75t_R FILLER_82_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_633 ();
 DECAPx2_ASAP7_75t_R FILLER_82_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_694 ();
 DECAPx10_ASAP7_75t_R FILLER_82_702 ();
 FILLER_ASAP7_75t_R FILLER_82_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_726 ();
 DECAPx4_ASAP7_75t_R FILLER_82_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_762 ();
 DECAPx10_ASAP7_75t_R FILLER_82_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_791 ();
 FILLER_ASAP7_75t_R FILLER_82_795 ();
 DECAPx6_ASAP7_75t_R FILLER_82_803 ();
 DECAPx1_ASAP7_75t_R FILLER_82_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_821 ();
 FILLER_ASAP7_75t_R FILLER_82_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_840 ();
 FILLER_ASAP7_75t_R FILLER_82_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_911 ();
 FILLER_ASAP7_75t_R FILLER_82_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_940 ();
 DECAPx1_ASAP7_75t_R FILLER_82_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_955 ();
 DECAPx6_ASAP7_75t_R FILLER_82_966 ();
 DECAPx2_ASAP7_75t_R FILLER_82_980 ();
 DECAPx6_ASAP7_75t_R FILLER_82_992 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1006 ();
 FILLER_ASAP7_75t_R FILLER_82_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_82_1041 ();
 FILLER_ASAP7_75t_R FILLER_82_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1164 ();
 FILLER_ASAP7_75t_R FILLER_82_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1179 ();
 FILLER_ASAP7_75t_R FILLER_82_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1388 ();
 FILLER_ASAP7_75t_R FILLER_82_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1404 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_28 ();
 DECAPx4_ASAP7_75t_R FILLER_83_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_42 ();
 DECAPx6_ASAP7_75t_R FILLER_83_49 ();
 DECAPx2_ASAP7_75t_R FILLER_83_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_69 ();
 DECAPx10_ASAP7_75t_R FILLER_83_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_104 ();
 DECAPx1_ASAP7_75t_R FILLER_83_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_121 ();
 DECAPx4_ASAP7_75t_R FILLER_83_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_138 ();
 DECAPx4_ASAP7_75t_R FILLER_83_152 ();
 FILLER_ASAP7_75t_R FILLER_83_162 ();
 DECAPx6_ASAP7_75t_R FILLER_83_190 ();
 DECAPx1_ASAP7_75t_R FILLER_83_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_208 ();
 DECAPx6_ASAP7_75t_R FILLER_83_215 ();
 DECAPx2_ASAP7_75t_R FILLER_83_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_235 ();
 FILLER_ASAP7_75t_R FILLER_83_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_244 ();
 DECAPx10_ASAP7_75t_R FILLER_83_251 ();
 DECAPx2_ASAP7_75t_R FILLER_83_273 ();
 FILLER_ASAP7_75t_R FILLER_83_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_281 ();
 DECAPx10_ASAP7_75t_R FILLER_83_288 ();
 DECAPx6_ASAP7_75t_R FILLER_83_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_324 ();
 DECAPx10_ASAP7_75t_R FILLER_83_333 ();
 DECAPx10_ASAP7_75t_R FILLER_83_355 ();
 DECAPx1_ASAP7_75t_R FILLER_83_377 ();
 DECAPx6_ASAP7_75t_R FILLER_83_387 ();
 FILLER_ASAP7_75t_R FILLER_83_401 ();
 DECAPx2_ASAP7_75t_R FILLER_83_412 ();
 FILLER_ASAP7_75t_R FILLER_83_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_443 ();
 DECAPx1_ASAP7_75t_R FILLER_83_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_454 ();
 DECAPx4_ASAP7_75t_R FILLER_83_461 ();
 FILLER_ASAP7_75t_R FILLER_83_483 ();
 DECAPx6_ASAP7_75t_R FILLER_83_491 ();
 FILLER_ASAP7_75t_R FILLER_83_505 ();
 DECAPx4_ASAP7_75t_R FILLER_83_513 ();
 FILLER_ASAP7_75t_R FILLER_83_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_528 ();
 DECAPx4_ASAP7_75t_R FILLER_83_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_545 ();
 DECAPx2_ASAP7_75t_R FILLER_83_555 ();
 FILLER_ASAP7_75t_R FILLER_83_561 ();
 FILLER_ASAP7_75t_R FILLER_83_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_598 ();
 DECAPx4_ASAP7_75t_R FILLER_83_625 ();
 FILLER_ASAP7_75t_R FILLER_83_635 ();
 FILLER_ASAP7_75t_R FILLER_83_670 ();
 DECAPx1_ASAP7_75t_R FILLER_83_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_688 ();
 DECAPx1_ASAP7_75t_R FILLER_83_705 ();
 DECAPx2_ASAP7_75t_R FILLER_83_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_727 ();
 DECAPx1_ASAP7_75t_R FILLER_83_759 ();
 DECAPx2_ASAP7_75t_R FILLER_83_769 ();
 FILLER_ASAP7_75t_R FILLER_83_775 ();
 DECAPx10_ASAP7_75t_R FILLER_83_843 ();
 DECAPx1_ASAP7_75t_R FILLER_83_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_869 ();
 DECAPx1_ASAP7_75t_R FILLER_83_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_880 ();
 FILLER_ASAP7_75t_R FILLER_83_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_909 ();
 FILLER_ASAP7_75t_R FILLER_83_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_955 ();
 DECAPx1_ASAP7_75t_R FILLER_83_966 ();
 DECAPx2_ASAP7_75t_R FILLER_83_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_982 ();
 DECAPx1_ASAP7_75t_R FILLER_83_995 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1030 ();
 FILLER_ASAP7_75t_R FILLER_83_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1097 ();
 FILLER_ASAP7_75t_R FILLER_83_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1197 ();
 FILLER_ASAP7_75t_R FILLER_83_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1363 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1399 ();
 DECAPx2_ASAP7_75t_R FILLER_84_2 ();
 FILLER_ASAP7_75t_R FILLER_84_8 ();
 FILLER_ASAP7_75t_R FILLER_84_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_53 ();
 DECAPx2_ASAP7_75t_R FILLER_84_60 ();
 FILLER_ASAP7_75t_R FILLER_84_66 ();
 DECAPx4_ASAP7_75t_R FILLER_84_94 ();
 FILLER_ASAP7_75t_R FILLER_84_104 ();
 DECAPx6_ASAP7_75t_R FILLER_84_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_182 ();
 DECAPx2_ASAP7_75t_R FILLER_84_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_209 ();
 DECAPx10_ASAP7_75t_R FILLER_84_230 ();
 DECAPx10_ASAP7_75t_R FILLER_84_252 ();
 DECAPx4_ASAP7_75t_R FILLER_84_274 ();
 DECAPx2_ASAP7_75t_R FILLER_84_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_298 ();
 DECAPx6_ASAP7_75t_R FILLER_84_319 ();
 FILLER_ASAP7_75t_R FILLER_84_333 ();
 DECAPx10_ASAP7_75t_R FILLER_84_341 ();
 DECAPx6_ASAP7_75t_R FILLER_84_363 ();
 DECAPx1_ASAP7_75t_R FILLER_84_377 ();
 DECAPx4_ASAP7_75t_R FILLER_84_389 ();
 FILLER_ASAP7_75t_R FILLER_84_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_409 ();
 DECAPx6_ASAP7_75t_R FILLER_84_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_437 ();
 DECAPx6_ASAP7_75t_R FILLER_84_444 ();
 DECAPx1_ASAP7_75t_R FILLER_84_458 ();
 DECAPx1_ASAP7_75t_R FILLER_84_464 ();
 DECAPx10_ASAP7_75t_R FILLER_84_488 ();
 DECAPx10_ASAP7_75t_R FILLER_84_510 ();
 DECAPx4_ASAP7_75t_R FILLER_84_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_542 ();
 DECAPx1_ASAP7_75t_R FILLER_84_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_570 ();
 FILLER_ASAP7_75t_R FILLER_84_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_592 ();
 DECAPx2_ASAP7_75t_R FILLER_84_606 ();
 FILLER_ASAP7_75t_R FILLER_84_612 ();
 DECAPx10_ASAP7_75t_R FILLER_84_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_639 ();
 FILLER_ASAP7_75t_R FILLER_84_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_664 ();
 DECAPx2_ASAP7_75t_R FILLER_84_682 ();
 FILLER_ASAP7_75t_R FILLER_84_688 ();
 DECAPx2_ASAP7_75t_R FILLER_84_696 ();
 FILLER_ASAP7_75t_R FILLER_84_702 ();
 DECAPx4_ASAP7_75t_R FILLER_84_730 ();
 FILLER_ASAP7_75t_R FILLER_84_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_742 ();
 DECAPx4_ASAP7_75t_R FILLER_84_749 ();
 FILLER_ASAP7_75t_R FILLER_84_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_761 ();
 DECAPx4_ASAP7_75t_R FILLER_84_774 ();
 FILLER_ASAP7_75t_R FILLER_84_784 ();
 DECAPx1_ASAP7_75t_R FILLER_84_789 ();
 FILLER_ASAP7_75t_R FILLER_84_801 ();
 DECAPx1_ASAP7_75t_R FILLER_84_839 ();
 DECAPx4_ASAP7_75t_R FILLER_84_881 ();
 DECAPx1_ASAP7_75t_R FILLER_84_921 ();
 DECAPx1_ASAP7_75t_R FILLER_84_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_947 ();
 DECAPx1_ASAP7_75t_R FILLER_84_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_956 ();
 DECAPx6_ASAP7_75t_R FILLER_84_961 ();
 DECAPx1_ASAP7_75t_R FILLER_84_975 ();
 FILLER_ASAP7_75t_R FILLER_84_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_989 ();
 DECAPx1_ASAP7_75t_R FILLER_84_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1016 ();
 FILLER_ASAP7_75t_R FILLER_84_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1040 ();
 FILLER_ASAP7_75t_R FILLER_84_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1060 ();
 FILLER_ASAP7_75t_R FILLER_84_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1117 ();
 FILLER_ASAP7_75t_R FILLER_84_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1125 ();
 FILLER_ASAP7_75t_R FILLER_84_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1168 ();
 FILLER_ASAP7_75t_R FILLER_84_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1388 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1394 ();
 FILLER_ASAP7_75t_R FILLER_85_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_39 ();
 DECAPx4_ASAP7_75t_R FILLER_85_69 ();
 FILLER_ASAP7_75t_R FILLER_85_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_81 ();
 FILLER_ASAP7_75t_R FILLER_85_85 ();
 DECAPx10_ASAP7_75t_R FILLER_85_119 ();
 DECAPx6_ASAP7_75t_R FILLER_85_141 ();
 FILLER_ASAP7_75t_R FILLER_85_155 ();
 DECAPx6_ASAP7_75t_R FILLER_85_177 ();
 DECAPx1_ASAP7_75t_R FILLER_85_199 ();
 FILLER_ASAP7_75t_R FILLER_85_211 ();
 FILLER_ASAP7_75t_R FILLER_85_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_247 ();
 FILLER_ASAP7_75t_R FILLER_85_260 ();
 DECAPx4_ASAP7_75t_R FILLER_85_276 ();
 DECAPx10_ASAP7_75t_R FILLER_85_292 ();
 DECAPx4_ASAP7_75t_R FILLER_85_314 ();
 FILLER_ASAP7_75t_R FILLER_85_324 ();
 FILLER_ASAP7_75t_R FILLER_85_357 ();
 FILLER_ASAP7_75t_R FILLER_85_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_369 ();
 DECAPx6_ASAP7_75t_R FILLER_85_392 ();
 DECAPx10_ASAP7_75t_R FILLER_85_432 ();
 DECAPx2_ASAP7_75t_R FILLER_85_462 ();
 FILLER_ASAP7_75t_R FILLER_85_468 ();
 DECAPx4_ASAP7_75t_R FILLER_85_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_497 ();
 FILLER_ASAP7_75t_R FILLER_85_508 ();
 DECAPx2_ASAP7_75t_R FILLER_85_526 ();
 DECAPx1_ASAP7_75t_R FILLER_85_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_548 ();
 DECAPx10_ASAP7_75t_R FILLER_85_555 ();
 DECAPx10_ASAP7_75t_R FILLER_85_577 ();
 DECAPx4_ASAP7_75t_R FILLER_85_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_609 ();
 DECAPx6_ASAP7_75t_R FILLER_85_662 ();
 FILLER_ASAP7_75t_R FILLER_85_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_678 ();
 DECAPx4_ASAP7_75t_R FILLER_85_686 ();
 FILLER_ASAP7_75t_R FILLER_85_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_705 ();
 FILLER_ASAP7_75t_R FILLER_85_742 ();
 DECAPx4_ASAP7_75t_R FILLER_85_751 ();
 FILLER_ASAP7_75t_R FILLER_85_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_763 ();
 FILLER_ASAP7_75t_R FILLER_85_770 ();
 DECAPx1_ASAP7_75t_R FILLER_85_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_836 ();
 FILLER_ASAP7_75t_R FILLER_85_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_864 ();
 DECAPx6_ASAP7_75t_R FILLER_85_871 ();
 DECAPx2_ASAP7_75t_R FILLER_85_885 ();
 FILLER_ASAP7_75t_R FILLER_85_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_923 ();
 DECAPx6_ASAP7_75t_R FILLER_85_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_948 ();
 DECAPx2_ASAP7_75t_R FILLER_85_959 ();
 FILLER_ASAP7_75t_R FILLER_85_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_967 ();
 DECAPx6_ASAP7_75t_R FILLER_85_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_992 ();
 DECAPx2_ASAP7_75t_R FILLER_85_996 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1062 ();
 FILLER_ASAP7_75t_R FILLER_85_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1360 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1396 ();
 DECAPx6_ASAP7_75t_R FILLER_86_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_16 ();
 DECAPx1_ASAP7_75t_R FILLER_86_35 ();
 DECAPx2_ASAP7_75t_R FILLER_86_42 ();
 DECAPx1_ASAP7_75t_R FILLER_86_54 ();
 DECAPx4_ASAP7_75t_R FILLER_86_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_81 ();
 DECAPx2_ASAP7_75t_R FILLER_86_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_91 ();
 DECAPx2_ASAP7_75t_R FILLER_86_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_113 ();
 DECAPx1_ASAP7_75t_R FILLER_86_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_144 ();
 DECAPx1_ASAP7_75t_R FILLER_86_161 ();
 DECAPx2_ASAP7_75t_R FILLER_86_181 ();
 FILLER_ASAP7_75t_R FILLER_86_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_189 ();
 DECAPx1_ASAP7_75t_R FILLER_86_202 ();
 DECAPx1_ASAP7_75t_R FILLER_86_213 ();
 DECAPx10_ASAP7_75t_R FILLER_86_223 ();
 DECAPx6_ASAP7_75t_R FILLER_86_245 ();
 DECAPx1_ASAP7_75t_R FILLER_86_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_263 ();
 DECAPx10_ASAP7_75t_R FILLER_86_272 ();
 DECAPx6_ASAP7_75t_R FILLER_86_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_308 ();
 DECAPx10_ASAP7_75t_R FILLER_86_321 ();
 DECAPx10_ASAP7_75t_R FILLER_86_343 ();
 DECAPx6_ASAP7_75t_R FILLER_86_365 ();
 FILLER_ASAP7_75t_R FILLER_86_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_381 ();
 DECAPx4_ASAP7_75t_R FILLER_86_408 ();
 FILLER_ASAP7_75t_R FILLER_86_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_429 ();
 DECAPx2_ASAP7_75t_R FILLER_86_438 ();
 FILLER_ASAP7_75t_R FILLER_86_444 ();
 FILLER_ASAP7_75t_R FILLER_86_460 ();
 DECAPx6_ASAP7_75t_R FILLER_86_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_478 ();
 DECAPx4_ASAP7_75t_R FILLER_86_485 ();
 FILLER_ASAP7_75t_R FILLER_86_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_497 ();
 FILLER_ASAP7_75t_R FILLER_86_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_516 ();
 DECAPx2_ASAP7_75t_R FILLER_86_542 ();
 FILLER_ASAP7_75t_R FILLER_86_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_550 ();
 DECAPx4_ASAP7_75t_R FILLER_86_557 ();
 DECAPx2_ASAP7_75t_R FILLER_86_574 ();
 FILLER_ASAP7_75t_R FILLER_86_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_582 ();
 DECAPx1_ASAP7_75t_R FILLER_86_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_590 ();
 DECAPx1_ASAP7_75t_R FILLER_86_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_611 ();
 DECAPx4_ASAP7_75t_R FILLER_86_665 ();
 FILLER_ASAP7_75t_R FILLER_86_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_677 ();
 DECAPx1_ASAP7_75t_R FILLER_86_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_689 ();
 DECAPx10_ASAP7_75t_R FILLER_86_702 ();
 DECAPx1_ASAP7_75t_R FILLER_86_724 ();
 DECAPx2_ASAP7_75t_R FILLER_86_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_740 ();
 DECAPx1_ASAP7_75t_R FILLER_86_759 ();
 FILLER_ASAP7_75t_R FILLER_86_788 ();
 DECAPx4_ASAP7_75t_R FILLER_86_796 ();
 DECAPx4_ASAP7_75t_R FILLER_86_830 ();
 FILLER_ASAP7_75t_R FILLER_86_843 ();
 DECAPx4_ASAP7_75t_R FILLER_86_851 ();
 FILLER_ASAP7_75t_R FILLER_86_861 ();
 DECAPx6_ASAP7_75t_R FILLER_86_869 ();
 DECAPx1_ASAP7_75t_R FILLER_86_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_887 ();
 FILLER_ASAP7_75t_R FILLER_86_899 ();
 DECAPx2_ASAP7_75t_R FILLER_86_907 ();
 DECAPx1_ASAP7_75t_R FILLER_86_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_951 ();
 FILLER_ASAP7_75t_R FILLER_86_965 ();
 FILLER_ASAP7_75t_R FILLER_86_977 ();
 FILLER_ASAP7_75t_R FILLER_86_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_988 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1021 ();
 FILLER_ASAP7_75t_R FILLER_86_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1101 ();
 FILLER_ASAP7_75t_R FILLER_86_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1124 ();
 FILLER_ASAP7_75t_R FILLER_86_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1198 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1362 ();
 FILLER_ASAP7_75t_R FILLER_86_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1388 ();
 FILLER_ASAP7_75t_R FILLER_86_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_87_2 ();
 DECAPx1_ASAP7_75t_R FILLER_87_16 ();
 DECAPx10_ASAP7_75t_R FILLER_87_26 ();
 FILLER_ASAP7_75t_R FILLER_87_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_50 ();
 DECAPx2_ASAP7_75t_R FILLER_87_60 ();
 FILLER_ASAP7_75t_R FILLER_87_66 ();
 DECAPx4_ASAP7_75t_R FILLER_87_103 ();
 FILLER_ASAP7_75t_R FILLER_87_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_159 ();
 DECAPx1_ASAP7_75t_R FILLER_87_172 ();
 DECAPx2_ASAP7_75t_R FILLER_87_182 ();
 DECAPx1_ASAP7_75t_R FILLER_87_196 ();
 FILLER_ASAP7_75t_R FILLER_87_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_208 ();
 DECAPx1_ASAP7_75t_R FILLER_87_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_240 ();
 DECAPx10_ASAP7_75t_R FILLER_87_249 ();
 DECAPx4_ASAP7_75t_R FILLER_87_271 ();
 DECAPx10_ASAP7_75t_R FILLER_87_309 ();
 DECAPx2_ASAP7_75t_R FILLER_87_331 ();
 FILLER_ASAP7_75t_R FILLER_87_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_339 ();
 DECAPx4_ASAP7_75t_R FILLER_87_346 ();
 DECAPx10_ASAP7_75t_R FILLER_87_362 ();
 DECAPx10_ASAP7_75t_R FILLER_87_384 ();
 DECAPx6_ASAP7_75t_R FILLER_87_406 ();
 DECAPx1_ASAP7_75t_R FILLER_87_420 ();
 DECAPx10_ASAP7_75t_R FILLER_87_438 ();
 DECAPx2_ASAP7_75t_R FILLER_87_460 ();
 FILLER_ASAP7_75t_R FILLER_87_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_468 ();
 FILLER_ASAP7_75t_R FILLER_87_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_477 ();
 DECAPx2_ASAP7_75t_R FILLER_87_495 ();
 DECAPx2_ASAP7_75t_R FILLER_87_519 ();
 FILLER_ASAP7_75t_R FILLER_87_525 ();
 DECAPx6_ASAP7_75t_R FILLER_87_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_561 ();
 DECAPx2_ASAP7_75t_R FILLER_87_594 ();
 FILLER_ASAP7_75t_R FILLER_87_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_602 ();
 DECAPx1_ASAP7_75t_R FILLER_87_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_636 ();
 DECAPx1_ASAP7_75t_R FILLER_87_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_659 ();
 DECAPx4_ASAP7_75t_R FILLER_87_664 ();
 FILLER_ASAP7_75t_R FILLER_87_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_692 ();
 DECAPx10_ASAP7_75t_R FILLER_87_713 ();
 DECAPx1_ASAP7_75t_R FILLER_87_741 ();
 DECAPx4_ASAP7_75t_R FILLER_87_752 ();
 DECAPx6_ASAP7_75t_R FILLER_87_776 ();
 FILLER_ASAP7_75t_R FILLER_87_790 ();
 DECAPx2_ASAP7_75t_R FILLER_87_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_812 ();
 DECAPx2_ASAP7_75t_R FILLER_87_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_825 ();
 FILLER_ASAP7_75t_R FILLER_87_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_870 ();
 DECAPx2_ASAP7_75t_R FILLER_87_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_889 ();
 DECAPx6_ASAP7_75t_R FILLER_87_908 ();
 FILLER_ASAP7_75t_R FILLER_87_922 ();
 FILLER_ASAP7_75t_R FILLER_87_926 ();
 DECAPx4_ASAP7_75t_R FILLER_87_931 ();
 DECAPx2_ASAP7_75t_R FILLER_87_955 ();
 FILLER_ASAP7_75t_R FILLER_87_961 ();
 DECAPx6_ASAP7_75t_R FILLER_87_999 ();
 FILLER_ASAP7_75t_R FILLER_87_1013 ();
 FILLER_ASAP7_75t_R FILLER_87_1034 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1062 ();
 FILLER_ASAP7_75t_R FILLER_87_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1122 ();
 FILLER_ASAP7_75t_R FILLER_87_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1190 ();
 FILLER_ASAP7_75t_R FILLER_87_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1348 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1370 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1392 ();
 FILLER_ASAP7_75t_R FILLER_87_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_88_37 ();
 DECAPx4_ASAP7_75t_R FILLER_88_69 ();
 FILLER_ASAP7_75t_R FILLER_88_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_81 ();
 DECAPx6_ASAP7_75t_R FILLER_88_88 ();
 DECAPx1_ASAP7_75t_R FILLER_88_102 ();
 DECAPx6_ASAP7_75t_R FILLER_88_112 ();
 FILLER_ASAP7_75t_R FILLER_88_126 ();
 DECAPx6_ASAP7_75t_R FILLER_88_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_153 ();
 DECAPx2_ASAP7_75t_R FILLER_88_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_166 ();
 DECAPx4_ASAP7_75t_R FILLER_88_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_221 ();
 DECAPx2_ASAP7_75t_R FILLER_88_230 ();
 FILLER_ASAP7_75t_R FILLER_88_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_238 ();
 DECAPx2_ASAP7_75t_R FILLER_88_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_253 ();
 DECAPx1_ASAP7_75t_R FILLER_88_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_264 ();
 DECAPx1_ASAP7_75t_R FILLER_88_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_272 ();
 DECAPx4_ASAP7_75t_R FILLER_88_327 ();
 FILLER_ASAP7_75t_R FILLER_88_337 ();
 DECAPx2_ASAP7_75t_R FILLER_88_347 ();
 FILLER_ASAP7_75t_R FILLER_88_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_355 ();
 DECAPx2_ASAP7_75t_R FILLER_88_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_370 ();
 DECAPx10_ASAP7_75t_R FILLER_88_377 ();
 DECAPx6_ASAP7_75t_R FILLER_88_399 ();
 FILLER_ASAP7_75t_R FILLER_88_413 ();
 DECAPx10_ASAP7_75t_R FILLER_88_421 ();
 FILLER_ASAP7_75t_R FILLER_88_443 ();
 DECAPx4_ASAP7_75t_R FILLER_88_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_461 ();
 DECAPx1_ASAP7_75t_R FILLER_88_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_468 ();
 DECAPx4_ASAP7_75t_R FILLER_88_483 ();
 FILLER_ASAP7_75t_R FILLER_88_493 ();
 DECAPx10_ASAP7_75t_R FILLER_88_503 ();
 DECAPx2_ASAP7_75t_R FILLER_88_525 ();
 FILLER_ASAP7_75t_R FILLER_88_531 ();
 DECAPx4_ASAP7_75t_R FILLER_88_539 ();
 FILLER_ASAP7_75t_R FILLER_88_549 ();
 DECAPx4_ASAP7_75t_R FILLER_88_570 ();
 FILLER_ASAP7_75t_R FILLER_88_580 ();
 DECAPx4_ASAP7_75t_R FILLER_88_585 ();
 FILLER_ASAP7_75t_R FILLER_88_595 ();
 FILLER_ASAP7_75t_R FILLER_88_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_602 ();
 DECAPx2_ASAP7_75t_R FILLER_88_609 ();
 FILLER_ASAP7_75t_R FILLER_88_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_617 ();
 DECAPx10_ASAP7_75t_R FILLER_88_621 ();
 DECAPx6_ASAP7_75t_R FILLER_88_643 ();
 DECAPx1_ASAP7_75t_R FILLER_88_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_661 ();
 FILLER_ASAP7_75t_R FILLER_88_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_680 ();
 DECAPx1_ASAP7_75t_R FILLER_88_697 ();
 DECAPx1_ASAP7_75t_R FILLER_88_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_715 ();
 DECAPx4_ASAP7_75t_R FILLER_88_752 ();
 FILLER_ASAP7_75t_R FILLER_88_762 ();
 FILLER_ASAP7_75t_R FILLER_88_777 ();
 DECAPx4_ASAP7_75t_R FILLER_88_817 ();
 DECAPx6_ASAP7_75t_R FILLER_88_836 ();
 DECAPx6_ASAP7_75t_R FILLER_88_853 ();
 DECAPx4_ASAP7_75t_R FILLER_88_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_895 ();
 DECAPx6_ASAP7_75t_R FILLER_88_902 ();
 FILLER_ASAP7_75t_R FILLER_88_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_924 ();
 DECAPx4_ASAP7_75t_R FILLER_88_937 ();
 FILLER_ASAP7_75t_R FILLER_88_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_949 ();
 DECAPx1_ASAP7_75t_R FILLER_88_964 ();
 DECAPx4_ASAP7_75t_R FILLER_88_972 ();
 FILLER_ASAP7_75t_R FILLER_88_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1145 ();
 FILLER_ASAP7_75t_R FILLER_88_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1162 ();
 FILLER_ASAP7_75t_R FILLER_88_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1388 ();
 FILLER_ASAP7_75t_R FILLER_88_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1404 ();
 FILLER_ASAP7_75t_R FILLER_89_34 ();
 FILLER_ASAP7_75t_R FILLER_89_45 ();
 DECAPx1_ASAP7_75t_R FILLER_89_62 ();
 DECAPx1_ASAP7_75t_R FILLER_89_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_125 ();
 DECAPx2_ASAP7_75t_R FILLER_89_132 ();
 DECAPx4_ASAP7_75t_R FILLER_89_164 ();
 FILLER_ASAP7_75t_R FILLER_89_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_240 ();
 DECAPx4_ASAP7_75t_R FILLER_89_247 ();
 FILLER_ASAP7_75t_R FILLER_89_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_259 ();
 DECAPx2_ASAP7_75t_R FILLER_89_274 ();
 FILLER_ASAP7_75t_R FILLER_89_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_282 ();
 DECAPx6_ASAP7_75t_R FILLER_89_293 ();
 FILLER_ASAP7_75t_R FILLER_89_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_309 ();
 DECAPx10_ASAP7_75t_R FILLER_89_318 ();
 DECAPx10_ASAP7_75t_R FILLER_89_340 ();
 DECAPx2_ASAP7_75t_R FILLER_89_362 ();
 DECAPx1_ASAP7_75t_R FILLER_89_375 ();
 DECAPx1_ASAP7_75t_R FILLER_89_393 ();
 FILLER_ASAP7_75t_R FILLER_89_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_420 ();
 DECAPx4_ASAP7_75t_R FILLER_89_433 ();
 FILLER_ASAP7_75t_R FILLER_89_457 ();
 DECAPx2_ASAP7_75t_R FILLER_89_473 ();
 DECAPx2_ASAP7_75t_R FILLER_89_501 ();
 FILLER_ASAP7_75t_R FILLER_89_507 ();
 DECAPx2_ASAP7_75t_R FILLER_89_535 ();
 FILLER_ASAP7_75t_R FILLER_89_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_553 ();
 DECAPx2_ASAP7_75t_R FILLER_89_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_600 ();
 DECAPx2_ASAP7_75t_R FILLER_89_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_613 ();
 DECAPx6_ASAP7_75t_R FILLER_89_617 ();
 FILLER_ASAP7_75t_R FILLER_89_631 ();
 DECAPx6_ASAP7_75t_R FILLER_89_665 ();
 DECAPx1_ASAP7_75t_R FILLER_89_679 ();
 DECAPx6_ASAP7_75t_R FILLER_89_689 ();
 FILLER_ASAP7_75t_R FILLER_89_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_705 ();
 DECAPx6_ASAP7_75t_R FILLER_89_730 ();
 DECAPx2_ASAP7_75t_R FILLER_89_744 ();
 FILLER_ASAP7_75t_R FILLER_89_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_762 ();
 DECAPx1_ASAP7_75t_R FILLER_89_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_804 ();
 FILLER_ASAP7_75t_R FILLER_89_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_810 ();
 FILLER_ASAP7_75t_R FILLER_89_817 ();
 DECAPx6_ASAP7_75t_R FILLER_89_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_867 ();
 DECAPx1_ASAP7_75t_R FILLER_89_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_917 ();
 DECAPx2_ASAP7_75t_R FILLER_89_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_932 ();
 DECAPx6_ASAP7_75t_R FILLER_89_945 ();
 DECAPx2_ASAP7_75t_R FILLER_89_959 ();
 DECAPx10_ASAP7_75t_R FILLER_89_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_999 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1017 ();
 FILLER_ASAP7_75t_R FILLER_89_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1040 ();
 FILLER_ASAP7_75t_R FILLER_89_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1055 ();
 FILLER_ASAP7_75t_R FILLER_89_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1136 ();
 FILLER_ASAP7_75t_R FILLER_89_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1195 ();
 FILLER_ASAP7_75t_R FILLER_89_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1218 ();
 FILLER_ASAP7_75t_R FILLER_89_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1361 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1383 ();
 DECAPx4_ASAP7_75t_R FILLER_90_2 ();
 FILLER_ASAP7_75t_R FILLER_90_18 ();
 DECAPx2_ASAP7_75t_R FILLER_90_81 ();
 FILLER_ASAP7_75t_R FILLER_90_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_89 ();
 DECAPx1_ASAP7_75t_R FILLER_90_99 ();
 DECAPx6_ASAP7_75t_R FILLER_90_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_152 ();
 DECAPx2_ASAP7_75t_R FILLER_90_156 ();
 FILLER_ASAP7_75t_R FILLER_90_162 ();
 DECAPx6_ASAP7_75t_R FILLER_90_171 ();
 FILLER_ASAP7_75t_R FILLER_90_185 ();
 DECAPx1_ASAP7_75t_R FILLER_90_194 ();
 DECAPx6_ASAP7_75t_R FILLER_90_204 ();
 FILLER_ASAP7_75t_R FILLER_90_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_220 ();
 DECAPx4_ASAP7_75t_R FILLER_90_227 ();
 DECAPx6_ASAP7_75t_R FILLER_90_245 ();
 DECAPx2_ASAP7_75t_R FILLER_90_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_283 ();
 DECAPx2_ASAP7_75t_R FILLER_90_308 ();
 DECAPx1_ASAP7_75t_R FILLER_90_330 ();
 DECAPx10_ASAP7_75t_R FILLER_90_352 ();
 DECAPx2_ASAP7_75t_R FILLER_90_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_380 ();
 DECAPx10_ASAP7_75t_R FILLER_90_387 ();
 FILLER_ASAP7_75t_R FILLER_90_427 ();
 DECAPx1_ASAP7_75t_R FILLER_90_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_439 ();
 DECAPx6_ASAP7_75t_R FILLER_90_448 ();
 DECAPx4_ASAP7_75t_R FILLER_90_464 ();
 FILLER_ASAP7_75t_R FILLER_90_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_476 ();
 DECAPx2_ASAP7_75t_R FILLER_90_483 ();
 FILLER_ASAP7_75t_R FILLER_90_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_491 ();
 FILLER_ASAP7_75t_R FILLER_90_498 ();
 DECAPx4_ASAP7_75t_R FILLER_90_506 ();
 FILLER_ASAP7_75t_R FILLER_90_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_518 ();
 DECAPx4_ASAP7_75t_R FILLER_90_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_564 ();
 DECAPx10_ASAP7_75t_R FILLER_90_572 ();
 DECAPx2_ASAP7_75t_R FILLER_90_594 ();
 FILLER_ASAP7_75t_R FILLER_90_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_676 ();
 DECAPx1_ASAP7_75t_R FILLER_90_690 ();
 DECAPx2_ASAP7_75t_R FILLER_90_702 ();
 FILLER_ASAP7_75t_R FILLER_90_708 ();
 DECAPx2_ASAP7_75t_R FILLER_90_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_734 ();
 FILLER_ASAP7_75t_R FILLER_90_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_743 ();
 DECAPx4_ASAP7_75t_R FILLER_90_751 ();
 FILLER_ASAP7_75t_R FILLER_90_761 ();
 DECAPx2_ASAP7_75t_R FILLER_90_771 ();
 DECAPx10_ASAP7_75t_R FILLER_90_780 ();
 DECAPx4_ASAP7_75t_R FILLER_90_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_812 ();
 DECAPx1_ASAP7_75t_R FILLER_90_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_823 ();
 FILLER_ASAP7_75t_R FILLER_90_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_840 ();
 DECAPx10_ASAP7_75t_R FILLER_90_844 ();
 DECAPx10_ASAP7_75t_R FILLER_90_866 ();
 DECAPx10_ASAP7_75t_R FILLER_90_888 ();
 FILLER_ASAP7_75t_R FILLER_90_910 ();
 FILLER_ASAP7_75t_R FILLER_90_918 ();
 DECAPx6_ASAP7_75t_R FILLER_90_926 ();
 FILLER_ASAP7_75t_R FILLER_90_940 ();
 DECAPx4_ASAP7_75t_R FILLER_90_948 ();
 FILLER_ASAP7_75t_R FILLER_90_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_967 ();
 DECAPx6_ASAP7_75t_R FILLER_90_976 ();
 DECAPx4_ASAP7_75t_R FILLER_90_996 ();
 FILLER_ASAP7_75t_R FILLER_90_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1008 ();
 FILLER_ASAP7_75t_R FILLER_90_1023 ();
 FILLER_ASAP7_75t_R FILLER_90_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1058 ();
 FILLER_ASAP7_75t_R FILLER_90_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1089 ();
 FILLER_ASAP7_75t_R FILLER_90_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1164 ();
 FILLER_ASAP7_75t_R FILLER_90_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1186 ();
 FILLER_ASAP7_75t_R FILLER_90_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1348 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1370 ();
 FILLER_ASAP7_75t_R FILLER_90_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1388 ();
 FILLER_ASAP7_75t_R FILLER_90_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_91_2 ();
 DECAPx2_ASAP7_75t_R FILLER_91_24 ();
 FILLER_ASAP7_75t_R FILLER_91_30 ();
 DECAPx10_ASAP7_75t_R FILLER_91_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_67 ();
 DECAPx10_ASAP7_75t_R FILLER_91_94 ();
 FILLER_ASAP7_75t_R FILLER_91_116 ();
 FILLER_ASAP7_75t_R FILLER_91_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_126 ();
 DECAPx4_ASAP7_75t_R FILLER_91_130 ();
 DECAPx2_ASAP7_75t_R FILLER_91_156 ();
 DECAPx2_ASAP7_75t_R FILLER_91_188 ();
 FILLER_ASAP7_75t_R FILLER_91_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_196 ();
 DECAPx4_ASAP7_75t_R FILLER_91_209 ();
 FILLER_ASAP7_75t_R FILLER_91_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_236 ();
 FILLER_ASAP7_75t_R FILLER_91_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_247 ();
 FILLER_ASAP7_75t_R FILLER_91_264 ();
 DECAPx2_ASAP7_75t_R FILLER_91_284 ();
 FILLER_ASAP7_75t_R FILLER_91_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_292 ();
 DECAPx2_ASAP7_75t_R FILLER_91_311 ();
 DECAPx2_ASAP7_75t_R FILLER_91_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_333 ();
 DECAPx2_ASAP7_75t_R FILLER_91_350 ();
 FILLER_ASAP7_75t_R FILLER_91_356 ();
 DECAPx2_ASAP7_75t_R FILLER_91_364 ();
 FILLER_ASAP7_75t_R FILLER_91_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_372 ();
 DECAPx2_ASAP7_75t_R FILLER_91_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_405 ();
 DECAPx1_ASAP7_75t_R FILLER_91_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_416 ();
 DECAPx10_ASAP7_75t_R FILLER_91_423 ();
 DECAPx10_ASAP7_75t_R FILLER_91_445 ();
 DECAPx2_ASAP7_75t_R FILLER_91_467 ();
 FILLER_ASAP7_75t_R FILLER_91_473 ();
 FILLER_ASAP7_75t_R FILLER_91_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_513 ();
 DECAPx6_ASAP7_75t_R FILLER_91_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_568 ();
 DECAPx2_ASAP7_75t_R FILLER_91_595 ();
 FILLER_ASAP7_75t_R FILLER_91_607 ();
 FILLER_ASAP7_75t_R FILLER_91_647 ();
 FILLER_ASAP7_75t_R FILLER_91_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_654 ();
 DECAPx10_ASAP7_75t_R FILLER_91_662 ();
 FILLER_ASAP7_75t_R FILLER_91_684 ();
 FILLER_ASAP7_75t_R FILLER_91_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_700 ();
 FILLER_ASAP7_75t_R FILLER_91_709 ();
 DECAPx2_ASAP7_75t_R FILLER_91_725 ();
 FILLER_ASAP7_75t_R FILLER_91_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_733 ();
 DECAPx2_ASAP7_75t_R FILLER_91_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_758 ();
 DECAPx6_ASAP7_75t_R FILLER_91_765 ();
 DECAPx2_ASAP7_75t_R FILLER_91_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_785 ();
 FILLER_ASAP7_75t_R FILLER_91_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_805 ();
 DECAPx4_ASAP7_75t_R FILLER_91_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_819 ();
 FILLER_ASAP7_75t_R FILLER_91_826 ();
 DECAPx2_ASAP7_75t_R FILLER_91_834 ();
 DECAPx4_ASAP7_75t_R FILLER_91_848 ();
 FILLER_ASAP7_75t_R FILLER_91_858 ();
 DECAPx1_ASAP7_75t_R FILLER_91_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_885 ();
 FILLER_ASAP7_75t_R FILLER_91_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_896 ();
 DECAPx10_ASAP7_75t_R FILLER_91_900 ();
 FILLER_ASAP7_75t_R FILLER_91_922 ();
 FILLER_ASAP7_75t_R FILLER_91_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1017 ();
 FILLER_ASAP7_75t_R FILLER_91_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1042 ();
 FILLER_ASAP7_75t_R FILLER_91_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1118 ();
 FILLER_ASAP7_75t_R FILLER_91_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1369 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_92_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_24 ();
 FILLER_ASAP7_75t_R FILLER_92_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_42 ();
 DECAPx6_ASAP7_75t_R FILLER_92_46 ();
 DECAPx2_ASAP7_75t_R FILLER_92_60 ();
 DECAPx1_ASAP7_75t_R FILLER_92_69 ();
 FILLER_ASAP7_75t_R FILLER_92_85 ();
 FILLER_ASAP7_75t_R FILLER_92_113 ();
 FILLER_ASAP7_75t_R FILLER_92_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_126 ();
 DECAPx2_ASAP7_75t_R FILLER_92_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_136 ();
 DECAPx2_ASAP7_75t_R FILLER_92_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_176 ();
 DECAPx4_ASAP7_75t_R FILLER_92_180 ();
 FILLER_ASAP7_75t_R FILLER_92_190 ();
 FILLER_ASAP7_75t_R FILLER_92_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_235 ();
 DECAPx10_ASAP7_75t_R FILLER_92_248 ();
 DECAPx4_ASAP7_75t_R FILLER_92_270 ();
 FILLER_ASAP7_75t_R FILLER_92_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_282 ();
 FILLER_ASAP7_75t_R FILLER_92_301 ();
 DECAPx4_ASAP7_75t_R FILLER_92_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_319 ();
 DECAPx2_ASAP7_75t_R FILLER_92_329 ();
 FILLER_ASAP7_75t_R FILLER_92_335 ();
 DECAPx2_ASAP7_75t_R FILLER_92_349 ();
 DECAPx1_ASAP7_75t_R FILLER_92_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_373 ();
 DECAPx2_ASAP7_75t_R FILLER_92_381 ();
 FILLER_ASAP7_75t_R FILLER_92_390 ();
 FILLER_ASAP7_75t_R FILLER_92_418 ();
 DECAPx4_ASAP7_75t_R FILLER_92_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_461 ();
 DECAPx2_ASAP7_75t_R FILLER_92_464 ();
 DECAPx10_ASAP7_75t_R FILLER_92_484 ();
 DECAPx6_ASAP7_75t_R FILLER_92_506 ();
 DECAPx1_ASAP7_75t_R FILLER_92_520 ();
 DECAPx6_ASAP7_75t_R FILLER_92_533 ();
 DECAPx1_ASAP7_75t_R FILLER_92_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_551 ();
 DECAPx4_ASAP7_75t_R FILLER_92_561 ();
 FILLER_ASAP7_75t_R FILLER_92_577 ();
 DECAPx6_ASAP7_75t_R FILLER_92_598 ();
 DECAPx10_ASAP7_75t_R FILLER_92_627 ();
 FILLER_ASAP7_75t_R FILLER_92_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_651 ();
 DECAPx2_ASAP7_75t_R FILLER_92_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_664 ();
 DECAPx4_ASAP7_75t_R FILLER_92_668 ();
 FILLER_ASAP7_75t_R FILLER_92_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_680 ();
 DECAPx6_ASAP7_75t_R FILLER_92_691 ();
 DECAPx1_ASAP7_75t_R FILLER_92_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_709 ();
 DECAPx4_ASAP7_75t_R FILLER_92_724 ();
 FILLER_ASAP7_75t_R FILLER_92_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_736 ();
 FILLER_ASAP7_75t_R FILLER_92_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_748 ();
 FILLER_ASAP7_75t_R FILLER_92_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_757 ();
 DECAPx1_ASAP7_75t_R FILLER_92_771 ();
 FILLER_ASAP7_75t_R FILLER_92_817 ();
 FILLER_ASAP7_75t_R FILLER_92_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_922 ();
 DECAPx10_ASAP7_75t_R FILLER_92_937 ();
 DECAPx4_ASAP7_75t_R FILLER_92_959 ();
 FILLER_ASAP7_75t_R FILLER_92_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_971 ();
 DECAPx4_ASAP7_75t_R FILLER_92_980 ();
 FILLER_ASAP7_75t_R FILLER_92_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_992 ();
 DECAPx10_ASAP7_75t_R FILLER_92_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1021 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1056 ();
 FILLER_ASAP7_75t_R FILLER_92_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1090 ();
 FILLER_ASAP7_75t_R FILLER_92_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1126 ();
 FILLER_ASAP7_75t_R FILLER_92_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1141 ();
 FILLER_ASAP7_75t_R FILLER_92_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1169 ();
 FILLER_ASAP7_75t_R FILLER_92_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1188 ();
 FILLER_ASAP7_75t_R FILLER_92_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1352 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1374 ();
 FILLER_ASAP7_75t_R FILLER_92_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1388 ();
 FILLER_ASAP7_75t_R FILLER_92_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_93_60 ();
 FILLER_ASAP7_75t_R FILLER_93_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_87 ();
 DECAPx6_ASAP7_75t_R FILLER_93_132 ();
 DECAPx2_ASAP7_75t_R FILLER_93_146 ();
 DECAPx2_ASAP7_75t_R FILLER_93_155 ();
 FILLER_ASAP7_75t_R FILLER_93_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_163 ();
 DECAPx6_ASAP7_75t_R FILLER_93_171 ();
 DECAPx2_ASAP7_75t_R FILLER_93_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_191 ();
 FILLER_ASAP7_75t_R FILLER_93_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_202 ();
 DECAPx1_ASAP7_75t_R FILLER_93_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_215 ();
 DECAPx2_ASAP7_75t_R FILLER_93_223 ();
 FILLER_ASAP7_75t_R FILLER_93_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_231 ();
 DECAPx6_ASAP7_75t_R FILLER_93_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_252 ();
 DECAPx1_ASAP7_75t_R FILLER_93_263 ();
 DECAPx10_ASAP7_75t_R FILLER_93_275 ();
 DECAPx4_ASAP7_75t_R FILLER_93_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_307 ();
 DECAPx6_ASAP7_75t_R FILLER_93_318 ();
 FILLER_ASAP7_75t_R FILLER_93_332 ();
 DECAPx1_ASAP7_75t_R FILLER_93_354 ();
 FILLER_ASAP7_75t_R FILLER_93_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_366 ();
 DECAPx6_ASAP7_75t_R FILLER_93_377 ();
 DECAPx1_ASAP7_75t_R FILLER_93_391 ();
 DECAPx1_ASAP7_75t_R FILLER_93_402 ();
 DECAPx4_ASAP7_75t_R FILLER_93_409 ();
 DECAPx10_ASAP7_75t_R FILLER_93_427 ();
 DECAPx10_ASAP7_75t_R FILLER_93_449 ();
 DECAPx10_ASAP7_75t_R FILLER_93_471 ();
 DECAPx10_ASAP7_75t_R FILLER_93_493 ();
 DECAPx4_ASAP7_75t_R FILLER_93_515 ();
 DECAPx2_ASAP7_75t_R FILLER_93_531 ();
 FILLER_ASAP7_75t_R FILLER_93_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_539 ();
 DECAPx1_ASAP7_75t_R FILLER_93_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_547 ();
 FILLER_ASAP7_75t_R FILLER_93_580 ();
 DECAPx6_ASAP7_75t_R FILLER_93_608 ();
 DECAPx2_ASAP7_75t_R FILLER_93_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_628 ();
 DECAPx6_ASAP7_75t_R FILLER_93_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_649 ();
 FILLER_ASAP7_75t_R FILLER_93_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_678 ();
 DECAPx1_ASAP7_75t_R FILLER_93_692 ();
 DECAPx2_ASAP7_75t_R FILLER_93_712 ();
 FILLER_ASAP7_75t_R FILLER_93_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_720 ();
 DECAPx1_ASAP7_75t_R FILLER_93_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_729 ();
 FILLER_ASAP7_75t_R FILLER_93_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_741 ();
 DECAPx6_ASAP7_75t_R FILLER_93_761 ();
 DECAPx1_ASAP7_75t_R FILLER_93_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_779 ();
 FILLER_ASAP7_75t_R FILLER_93_798 ();
 DECAPx6_ASAP7_75t_R FILLER_93_813 ();
 DECAPx1_ASAP7_75t_R FILLER_93_837 ();
 DECAPx6_ASAP7_75t_R FILLER_93_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_861 ();
 DECAPx4_ASAP7_75t_R FILLER_93_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_880 ();
 DECAPx1_ASAP7_75t_R FILLER_93_895 ();
 DECAPx4_ASAP7_75t_R FILLER_93_911 ();
 FILLER_ASAP7_75t_R FILLER_93_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_923 ();
 DECAPx6_ASAP7_75t_R FILLER_93_926 ();
 FILLER_ASAP7_75t_R FILLER_93_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_942 ();
 DECAPx6_ASAP7_75t_R FILLER_93_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_969 ();
 DECAPx10_ASAP7_75t_R FILLER_93_973 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1044 ();
 FILLER_ASAP7_75t_R FILLER_93_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1217 ();
 FILLER_ASAP7_75t_R FILLER_93_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1363 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1399 ();
 DECAPx4_ASAP7_75t_R FILLER_94_2 ();
 FILLER_ASAP7_75t_R FILLER_94_18 ();
 DECAPx1_ASAP7_75t_R FILLER_94_38 ();
 DECAPx1_ASAP7_75t_R FILLER_94_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_75 ();
 DECAPx1_ASAP7_75t_R FILLER_94_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_86 ();
 DECAPx4_ASAP7_75t_R FILLER_94_90 ();
 FILLER_ASAP7_75t_R FILLER_94_100 ();
 DECAPx1_ASAP7_75t_R FILLER_94_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_118 ();
 DECAPx2_ASAP7_75t_R FILLER_94_145 ();
 FILLER_ASAP7_75t_R FILLER_94_151 ();
 FILLER_ASAP7_75t_R FILLER_94_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_161 ();
 FILLER_ASAP7_75t_R FILLER_94_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_190 ();
 DECAPx2_ASAP7_75t_R FILLER_94_199 ();
 DECAPx10_ASAP7_75t_R FILLER_94_211 ();
 FILLER_ASAP7_75t_R FILLER_94_233 ();
 DECAPx6_ASAP7_75t_R FILLER_94_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_255 ();
 DECAPx2_ASAP7_75t_R FILLER_94_266 ();
 DECAPx10_ASAP7_75t_R FILLER_94_280 ();
 DECAPx10_ASAP7_75t_R FILLER_94_308 ();
 DECAPx10_ASAP7_75t_R FILLER_94_330 ();
 DECAPx10_ASAP7_75t_R FILLER_94_352 ();
 DECAPx10_ASAP7_75t_R FILLER_94_374 ();
 DECAPx10_ASAP7_75t_R FILLER_94_396 ();
 DECAPx1_ASAP7_75t_R FILLER_94_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_449 ();
 DECAPx2_ASAP7_75t_R FILLER_94_456 ();
 DECAPx4_ASAP7_75t_R FILLER_94_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_474 ();
 DECAPx4_ASAP7_75t_R FILLER_94_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_491 ();
 DECAPx4_ASAP7_75t_R FILLER_94_506 ();
 FILLER_ASAP7_75t_R FILLER_94_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_518 ();
 FILLER_ASAP7_75t_R FILLER_94_554 ();
 DECAPx2_ASAP7_75t_R FILLER_94_562 ();
 DECAPx4_ASAP7_75t_R FILLER_94_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_595 ();
 DECAPx4_ASAP7_75t_R FILLER_94_599 ();
 FILLER_ASAP7_75t_R FILLER_94_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_611 ();
 DECAPx2_ASAP7_75t_R FILLER_94_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_626 ();
 DECAPx2_ASAP7_75t_R FILLER_94_659 ();
 FILLER_ASAP7_75t_R FILLER_94_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_667 ();
 FILLER_ASAP7_75t_R FILLER_94_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_718 ();
 FILLER_ASAP7_75t_R FILLER_94_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_727 ();
 DECAPx2_ASAP7_75t_R FILLER_94_740 ();
 FILLER_ASAP7_75t_R FILLER_94_746 ();
 DECAPx4_ASAP7_75t_R FILLER_94_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_761 ();
 DECAPx2_ASAP7_75t_R FILLER_94_774 ();
 DECAPx2_ASAP7_75t_R FILLER_94_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_789 ();
 DECAPx10_ASAP7_75t_R FILLER_94_822 ();
 DECAPx10_ASAP7_75t_R FILLER_94_844 ();
 DECAPx6_ASAP7_75t_R FILLER_94_872 ();
 DECAPx2_ASAP7_75t_R FILLER_94_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_892 ();
 DECAPx6_ASAP7_75t_R FILLER_94_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_919 ();
 FILLER_ASAP7_75t_R FILLER_94_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_934 ();
 DECAPx6_ASAP7_75t_R FILLER_94_947 ();
 FILLER_ASAP7_75t_R FILLER_94_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_975 ();
 DECAPx2_ASAP7_75t_R FILLER_94_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_994 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1049 ();
 FILLER_ASAP7_75t_R FILLER_94_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1104 ();
 FILLER_ASAP7_75t_R FILLER_94_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1175 ();
 FILLER_ASAP7_75t_R FILLER_94_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1378 ();
 FILLER_ASAP7_75t_R FILLER_94_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1388 ();
 FILLER_ASAP7_75t_R FILLER_94_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_95_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_40 ();
 DECAPx4_ASAP7_75t_R FILLER_95_53 ();
 DECAPx1_ASAP7_75t_R FILLER_95_69 ();
 DECAPx10_ASAP7_75t_R FILLER_95_99 ();
 DECAPx2_ASAP7_75t_R FILLER_95_121 ();
 FILLER_ASAP7_75t_R FILLER_95_166 ();
 FILLER_ASAP7_75t_R FILLER_95_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_179 ();
 DECAPx1_ASAP7_75t_R FILLER_95_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_243 ();
 DECAPx2_ASAP7_75t_R FILLER_95_258 ();
 FILLER_ASAP7_75t_R FILLER_95_264 ();
 FILLER_ASAP7_75t_R FILLER_95_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_291 ();
 DECAPx6_ASAP7_75t_R FILLER_95_300 ();
 DECAPx2_ASAP7_75t_R FILLER_95_314 ();
 DECAPx10_ASAP7_75t_R FILLER_95_340 ();
 DECAPx10_ASAP7_75t_R FILLER_95_362 ();
 DECAPx2_ASAP7_75t_R FILLER_95_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_390 ();
 DECAPx6_ASAP7_75t_R FILLER_95_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_411 ();
 DECAPx10_ASAP7_75t_R FILLER_95_418 ();
 DECAPx10_ASAP7_75t_R FILLER_95_440 ();
 DECAPx4_ASAP7_75t_R FILLER_95_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_472 ();
 DECAPx1_ASAP7_75t_R FILLER_95_481 ();
 DECAPx6_ASAP7_75t_R FILLER_95_491 ();
 DECAPx6_ASAP7_75t_R FILLER_95_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_525 ();
 DECAPx6_ASAP7_75t_R FILLER_95_532 ();
 DECAPx1_ASAP7_75t_R FILLER_95_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_550 ();
 DECAPx4_ASAP7_75t_R FILLER_95_557 ();
 FILLER_ASAP7_75t_R FILLER_95_567 ();
 DECAPx4_ASAP7_75t_R FILLER_95_572 ();
 FILLER_ASAP7_75t_R FILLER_95_582 ();
 FILLER_ASAP7_75t_R FILLER_95_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_673 ();
 DECAPx6_ASAP7_75t_R FILLER_95_680 ();
 FILLER_ASAP7_75t_R FILLER_95_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_696 ();
 DECAPx4_ASAP7_75t_R FILLER_95_703 ();
 FILLER_ASAP7_75t_R FILLER_95_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_715 ();
 DECAPx4_ASAP7_75t_R FILLER_95_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_746 ();
 DECAPx4_ASAP7_75t_R FILLER_95_753 ();
 FILLER_ASAP7_75t_R FILLER_95_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_765 ();
 FILLER_ASAP7_75t_R FILLER_95_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_774 ();
 DECAPx2_ASAP7_75t_R FILLER_95_789 ();
 DECAPx2_ASAP7_75t_R FILLER_95_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_809 ();
 DECAPx4_ASAP7_75t_R FILLER_95_813 ();
 FILLER_ASAP7_75t_R FILLER_95_823 ();
 DECAPx1_ASAP7_75t_R FILLER_95_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_860 ();
 DECAPx10_ASAP7_75t_R FILLER_95_902 ();
 DECAPx2_ASAP7_75t_R FILLER_95_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_932 ();
 DECAPx1_ASAP7_75t_R FILLER_95_950 ();
 DECAPx6_ASAP7_75t_R FILLER_95_957 ();
 DECAPx1_ASAP7_75t_R FILLER_95_971 ();
 FILLER_ASAP7_75t_R FILLER_95_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1013 ();
 FILLER_ASAP7_75t_R FILLER_95_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1048 ();
 FILLER_ASAP7_75t_R FILLER_95_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1122 ();
 FILLER_ASAP7_75t_R FILLER_95_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1388 ();
 FILLER_ASAP7_75t_R FILLER_95_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_96_2 ();
 FILLER_ASAP7_75t_R FILLER_96_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_14 ();
 DECAPx4_ASAP7_75t_R FILLER_96_18 ();
 DECAPx1_ASAP7_75t_R FILLER_96_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_38 ();
 FILLER_ASAP7_75t_R FILLER_96_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_73 ();
 DECAPx1_ASAP7_75t_R FILLER_96_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_84 ();
 DECAPx2_ASAP7_75t_R FILLER_96_115 ();
 FILLER_ASAP7_75t_R FILLER_96_121 ();
 DECAPx1_ASAP7_75t_R FILLER_96_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_133 ();
 FILLER_ASAP7_75t_R FILLER_96_137 ();
 DECAPx2_ASAP7_75t_R FILLER_96_158 ();
 FILLER_ASAP7_75t_R FILLER_96_164 ();
 DECAPx4_ASAP7_75t_R FILLER_96_169 ();
 FILLER_ASAP7_75t_R FILLER_96_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_181 ();
 DECAPx4_ASAP7_75t_R FILLER_96_210 ();
 FILLER_ASAP7_75t_R FILLER_96_220 ();
 DECAPx4_ASAP7_75t_R FILLER_96_230 ();
 DECAPx10_ASAP7_75t_R FILLER_96_246 ();
 DECAPx2_ASAP7_75t_R FILLER_96_274 ();
 DECAPx2_ASAP7_75t_R FILLER_96_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_298 ();
 FILLER_ASAP7_75t_R FILLER_96_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_315 ();
 DECAPx6_ASAP7_75t_R FILLER_96_350 ();
 DECAPx2_ASAP7_75t_R FILLER_96_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_370 ();
 DECAPx4_ASAP7_75t_R FILLER_96_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_396 ();
 DECAPx1_ASAP7_75t_R FILLER_96_414 ();
 DECAPx10_ASAP7_75t_R FILLER_96_424 ();
 DECAPx2_ASAP7_75t_R FILLER_96_446 ();
 FILLER_ASAP7_75t_R FILLER_96_452 ();
 FILLER_ASAP7_75t_R FILLER_96_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_472 ();
 DECAPx10_ASAP7_75t_R FILLER_96_479 ();
 DECAPx10_ASAP7_75t_R FILLER_96_501 ();
 FILLER_ASAP7_75t_R FILLER_96_523 ();
 DECAPx2_ASAP7_75t_R FILLER_96_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_547 ();
 DECAPx2_ASAP7_75t_R FILLER_96_581 ();
 FILLER_ASAP7_75t_R FILLER_96_587 ();
 DECAPx2_ASAP7_75t_R FILLER_96_595 ();
 FILLER_ASAP7_75t_R FILLER_96_601 ();
 DECAPx1_ASAP7_75t_R FILLER_96_606 ();
 FILLER_ASAP7_75t_R FILLER_96_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_628 ();
 DECAPx4_ASAP7_75t_R FILLER_96_635 ();
 DECAPx2_ASAP7_75t_R FILLER_96_654 ();
 FILLER_ASAP7_75t_R FILLER_96_660 ();
 DECAPx10_ASAP7_75t_R FILLER_96_665 ();
 FILLER_ASAP7_75t_R FILLER_96_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_689 ();
 DECAPx1_ASAP7_75t_R FILLER_96_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_713 ();
 DECAPx2_ASAP7_75t_R FILLER_96_718 ();
 FILLER_ASAP7_75t_R FILLER_96_730 ();
 FILLER_ASAP7_75t_R FILLER_96_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_766 ();
 DECAPx1_ASAP7_75t_R FILLER_96_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_779 ();
 DECAPx6_ASAP7_75t_R FILLER_96_788 ();
 DECAPx1_ASAP7_75t_R FILLER_96_802 ();
 FILLER_ASAP7_75t_R FILLER_96_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_818 ();
 FILLER_ASAP7_75t_R FILLER_96_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_938 ();
 DECAPx10_ASAP7_75t_R FILLER_96_969 ();
 DECAPx2_ASAP7_75t_R FILLER_96_991 ();
 FILLER_ASAP7_75t_R FILLER_96_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_999 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1162 ();
 FILLER_ASAP7_75t_R FILLER_96_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1361 ();
 FILLER_ASAP7_75t_R FILLER_96_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1388 ();
 FILLER_ASAP7_75t_R FILLER_96_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1404 ();
 FILLER_ASAP7_75t_R FILLER_97_42 ();
 FILLER_ASAP7_75t_R FILLER_97_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_52 ();
 FILLER_ASAP7_75t_R FILLER_97_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_58 ();
 FILLER_ASAP7_75t_R FILLER_97_88 ();
 FILLER_ASAP7_75t_R FILLER_97_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_151 ();
 DECAPx4_ASAP7_75t_R FILLER_97_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_188 ();
 DECAPx10_ASAP7_75t_R FILLER_97_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_227 ();
 FILLER_ASAP7_75t_R FILLER_97_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_258 ();
 DECAPx2_ASAP7_75t_R FILLER_97_271 ();
 FILLER_ASAP7_75t_R FILLER_97_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_279 ();
 DECAPx1_ASAP7_75t_R FILLER_97_294 ();
 DECAPx6_ASAP7_75t_R FILLER_97_312 ();
 DECAPx4_ASAP7_75t_R FILLER_97_356 ();
 FILLER_ASAP7_75t_R FILLER_97_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_368 ();
 DECAPx10_ASAP7_75t_R FILLER_97_375 ();
 DECAPx6_ASAP7_75t_R FILLER_97_397 ();
 FILLER_ASAP7_75t_R FILLER_97_411 ();
 DECAPx10_ASAP7_75t_R FILLER_97_419 ();
 DECAPx10_ASAP7_75t_R FILLER_97_459 ();
 DECAPx10_ASAP7_75t_R FILLER_97_481 ();
 DECAPx6_ASAP7_75t_R FILLER_97_503 ();
 DECAPx1_ASAP7_75t_R FILLER_97_517 ();
 DECAPx10_ASAP7_75t_R FILLER_97_537 ();
 DECAPx10_ASAP7_75t_R FILLER_97_559 ();
 DECAPx10_ASAP7_75t_R FILLER_97_581 ();
 DECAPx4_ASAP7_75t_R FILLER_97_603 ();
 DECAPx4_ASAP7_75t_R FILLER_97_619 ();
 FILLER_ASAP7_75t_R FILLER_97_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_631 ();
 DECAPx6_ASAP7_75t_R FILLER_97_635 ();
 DECAPx1_ASAP7_75t_R FILLER_97_649 ();
 DECAPx2_ASAP7_75t_R FILLER_97_659 ();
 FILLER_ASAP7_75t_R FILLER_97_665 ();
 DECAPx2_ASAP7_75t_R FILLER_97_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_676 ();
 DECAPx1_ASAP7_75t_R FILLER_97_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_708 ();
 FILLER_ASAP7_75t_R FILLER_97_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_730 ();
 FILLER_ASAP7_75t_R FILLER_97_746 ();
 FILLER_ASAP7_75t_R FILLER_97_754 ();
 DECAPx4_ASAP7_75t_R FILLER_97_795 ();
 FILLER_ASAP7_75t_R FILLER_97_823 ();
 DECAPx1_ASAP7_75t_R FILLER_97_843 ();
 DECAPx6_ASAP7_75t_R FILLER_97_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_864 ();
 DECAPx2_ASAP7_75t_R FILLER_97_868 ();
 DECAPx4_ASAP7_75t_R FILLER_97_880 ();
 DECAPx2_ASAP7_75t_R FILLER_97_899 ();
 FILLER_ASAP7_75t_R FILLER_97_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_926 ();
 DECAPx6_ASAP7_75t_R FILLER_97_934 ();
 DECAPx1_ASAP7_75t_R FILLER_97_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_961 ();
 DECAPx2_ASAP7_75t_R FILLER_97_974 ();
 DECAPx1_ASAP7_75t_R FILLER_97_986 ();
 FILLER_ASAP7_75t_R FILLER_97_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1015 ();
 FILLER_ASAP7_75t_R FILLER_97_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1081 ();
 FILLER_ASAP7_75t_R FILLER_97_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1114 ();
 FILLER_ASAP7_75t_R FILLER_97_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1404 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_32 ();
 FILLER_ASAP7_75t_R FILLER_98_47 ();
 DECAPx4_ASAP7_75t_R FILLER_98_55 ();
 DECAPx2_ASAP7_75t_R FILLER_98_71 ();
 DECAPx6_ASAP7_75t_R FILLER_98_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_100 ();
 FILLER_ASAP7_75t_R FILLER_98_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_115 ();
 DECAPx1_ASAP7_75t_R FILLER_98_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_129 ();
 FILLER_ASAP7_75t_R FILLER_98_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_135 ();
 DECAPx6_ASAP7_75t_R FILLER_98_143 ();
 DECAPx1_ASAP7_75t_R FILLER_98_157 ();
 DECAPx6_ASAP7_75t_R FILLER_98_174 ();
 DECAPx1_ASAP7_75t_R FILLER_98_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_192 ();
 DECAPx4_ASAP7_75t_R FILLER_98_203 ();
 FILLER_ASAP7_75t_R FILLER_98_213 ();
 DECAPx2_ASAP7_75t_R FILLER_98_225 ();
 FILLER_ASAP7_75t_R FILLER_98_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_233 ();
 DECAPx1_ASAP7_75t_R FILLER_98_262 ();
 DECAPx10_ASAP7_75t_R FILLER_98_272 ();
 DECAPx6_ASAP7_75t_R FILLER_98_294 ();
 DECAPx10_ASAP7_75t_R FILLER_98_317 ();
 FILLER_ASAP7_75t_R FILLER_98_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_341 ();
 DECAPx2_ASAP7_75t_R FILLER_98_350 ();
 DECAPx6_ASAP7_75t_R FILLER_98_369 ();
 DECAPx1_ASAP7_75t_R FILLER_98_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_387 ();
 DECAPx10_ASAP7_75t_R FILLER_98_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_416 ();
 DECAPx1_ASAP7_75t_R FILLER_98_431 ();
 FILLER_ASAP7_75t_R FILLER_98_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_461 ();
 DECAPx2_ASAP7_75t_R FILLER_98_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_485 ();
 DECAPx4_ASAP7_75t_R FILLER_98_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_504 ();
 DECAPx4_ASAP7_75t_R FILLER_98_513 ();
 FILLER_ASAP7_75t_R FILLER_98_529 ();
 DECAPx10_ASAP7_75t_R FILLER_98_553 ();
 DECAPx1_ASAP7_75t_R FILLER_98_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_579 ();
 DECAPx2_ASAP7_75t_R FILLER_98_644 ();
 FILLER_ASAP7_75t_R FILLER_98_650 ();
 DECAPx2_ASAP7_75t_R FILLER_98_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_684 ();
 FILLER_ASAP7_75t_R FILLER_98_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_706 ();
 DECAPx6_ASAP7_75t_R FILLER_98_719 ();
 FILLER_ASAP7_75t_R FILLER_98_733 ();
 DECAPx6_ASAP7_75t_R FILLER_98_748 ();
 DECAPx2_ASAP7_75t_R FILLER_98_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_768 ();
 DECAPx2_ASAP7_75t_R FILLER_98_775 ();
 DECAPx10_ASAP7_75t_R FILLER_98_784 ();
 DECAPx4_ASAP7_75t_R FILLER_98_806 ();
 FILLER_ASAP7_75t_R FILLER_98_816 ();
 DECAPx1_ASAP7_75t_R FILLER_98_821 ();
 DECAPx1_ASAP7_75t_R FILLER_98_837 ();
 DECAPx4_ASAP7_75t_R FILLER_98_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_859 ();
 DECAPx4_ASAP7_75t_R FILLER_98_880 ();
 FILLER_ASAP7_75t_R FILLER_98_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_892 ();
 DECAPx2_ASAP7_75t_R FILLER_98_901 ();
 DECAPx2_ASAP7_75t_R FILLER_98_913 ();
 FILLER_ASAP7_75t_R FILLER_98_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_927 ();
 DECAPx6_ASAP7_75t_R FILLER_98_937 ();
 DECAPx1_ASAP7_75t_R FILLER_98_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_955 ();
 DECAPx4_ASAP7_75t_R FILLER_98_962 ();
 FILLER_ASAP7_75t_R FILLER_98_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_980 ();
 DECAPx4_ASAP7_75t_R FILLER_98_993 ();
 FILLER_ASAP7_75t_R FILLER_98_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1012 ();
 FILLER_ASAP7_75t_R FILLER_98_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1090 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1130 ();
 FILLER_ASAP7_75t_R FILLER_98_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1382 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1388 ();
 FILLER_ASAP7_75t_R FILLER_98_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_99_2 ();
 DECAPx2_ASAP7_75t_R FILLER_99_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_83 ();
 DECAPx2_ASAP7_75t_R FILLER_99_90 ();
 FILLER_ASAP7_75t_R FILLER_99_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_98 ();
 FILLER_ASAP7_75t_R FILLER_99_128 ();
 DECAPx1_ASAP7_75t_R FILLER_99_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_186 ();
 DECAPx1_ASAP7_75t_R FILLER_99_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_215 ();
 DECAPx2_ASAP7_75t_R FILLER_99_226 ();
 FILLER_ASAP7_75t_R FILLER_99_232 ();
 DECAPx2_ASAP7_75t_R FILLER_99_240 ();
 FILLER_ASAP7_75t_R FILLER_99_246 ();
 FILLER_ASAP7_75t_R FILLER_99_254 ();
 DECAPx2_ASAP7_75t_R FILLER_99_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_284 ();
 DECAPx10_ASAP7_75t_R FILLER_99_303 ();
 DECAPx10_ASAP7_75t_R FILLER_99_325 ();
 DECAPx1_ASAP7_75t_R FILLER_99_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_351 ();
 DECAPx4_ASAP7_75t_R FILLER_99_378 ();
 DECAPx10_ASAP7_75t_R FILLER_99_395 ();
 DECAPx6_ASAP7_75t_R FILLER_99_417 ();
 DECAPx1_ASAP7_75t_R FILLER_99_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_435 ();
 DECAPx10_ASAP7_75t_R FILLER_99_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_466 ();
 FILLER_ASAP7_75t_R FILLER_99_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_475 ();
 DECAPx2_ASAP7_75t_R FILLER_99_490 ();
 FILLER_ASAP7_75t_R FILLER_99_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_498 ();
 DECAPx10_ASAP7_75t_R FILLER_99_505 ();
 DECAPx1_ASAP7_75t_R FILLER_99_527 ();
 DECAPx1_ASAP7_75t_R FILLER_99_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_557 ();
 DECAPx2_ASAP7_75t_R FILLER_99_565 ();
 FILLER_ASAP7_75t_R FILLER_99_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_573 ();
 FILLER_ASAP7_75t_R FILLER_99_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_611 ();
 DECAPx2_ASAP7_75t_R FILLER_99_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_624 ();
 DECAPx1_ASAP7_75t_R FILLER_99_654 ();
 FILLER_ASAP7_75t_R FILLER_99_670 ();
 DECAPx10_ASAP7_75t_R FILLER_99_675 ();
 DECAPx4_ASAP7_75t_R FILLER_99_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_707 ();
 DECAPx6_ASAP7_75t_R FILLER_99_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_741 ();
 DECAPx10_ASAP7_75t_R FILLER_99_749 ();
 DECAPx2_ASAP7_75t_R FILLER_99_771 ();
 FILLER_ASAP7_75t_R FILLER_99_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_779 ();
 DECAPx2_ASAP7_75t_R FILLER_99_808 ();
 DECAPx6_ASAP7_75t_R FILLER_99_828 ();
 DECAPx1_ASAP7_75t_R FILLER_99_842 ();
 DECAPx10_ASAP7_75t_R FILLER_99_855 ();
 DECAPx6_ASAP7_75t_R FILLER_99_877 ();
 FILLER_ASAP7_75t_R FILLER_99_891 ();
 DECAPx6_ASAP7_75t_R FILLER_99_899 ();
 FILLER_ASAP7_75t_R FILLER_99_913 ();
 FILLER_ASAP7_75t_R FILLER_99_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_923 ();
 DECAPx2_ASAP7_75t_R FILLER_99_926 ();
 DECAPx2_ASAP7_75t_R FILLER_99_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_950 ();
 DECAPx2_ASAP7_75t_R FILLER_99_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_963 ();
 DECAPx6_ASAP7_75t_R FILLER_99_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_981 ();
 DECAPx4_ASAP7_75t_R FILLER_99_988 ();
 FILLER_ASAP7_75t_R FILLER_99_998 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1150 ();
 FILLER_ASAP7_75t_R FILLER_99_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_100_2 ();
 FILLER_ASAP7_75t_R FILLER_100_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_14 ();
 FILLER_ASAP7_75t_R FILLER_100_18 ();
 FILLER_ASAP7_75t_R FILLER_100_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_45 ();
 DECAPx2_ASAP7_75t_R FILLER_100_52 ();
 DECAPx2_ASAP7_75t_R FILLER_100_61 ();
 FILLER_ASAP7_75t_R FILLER_100_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_69 ();
 FILLER_ASAP7_75t_R FILLER_100_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_104 ();
 DECAPx10_ASAP7_75t_R FILLER_100_111 ();
 DECAPx4_ASAP7_75t_R FILLER_100_133 ();
 DECAPx6_ASAP7_75t_R FILLER_100_152 ();
 DECAPx1_ASAP7_75t_R FILLER_100_166 ();
 DECAPx6_ASAP7_75t_R FILLER_100_173 ();
 FILLER_ASAP7_75t_R FILLER_100_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_189 ();
 DECAPx4_ASAP7_75t_R FILLER_100_200 ();
 FILLER_ASAP7_75t_R FILLER_100_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_212 ();
 DECAPx10_ASAP7_75t_R FILLER_100_231 ();
 DECAPx6_ASAP7_75t_R FILLER_100_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_279 ();
 DECAPx10_ASAP7_75t_R FILLER_100_286 ();
 DECAPx6_ASAP7_75t_R FILLER_100_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_327 ();
 DECAPx10_ASAP7_75t_R FILLER_100_338 ();
 DECAPx2_ASAP7_75t_R FILLER_100_360 ();
 DECAPx6_ASAP7_75t_R FILLER_100_369 ();
 FILLER_ASAP7_75t_R FILLER_100_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_385 ();
 DECAPx1_ASAP7_75t_R FILLER_100_412 ();
 DECAPx10_ASAP7_75t_R FILLER_100_424 ();
 DECAPx6_ASAP7_75t_R FILLER_100_446 ();
 FILLER_ASAP7_75t_R FILLER_100_460 ();
 DECAPx10_ASAP7_75t_R FILLER_100_472 ();
 DECAPx10_ASAP7_75t_R FILLER_100_494 ();
 DECAPx10_ASAP7_75t_R FILLER_100_516 ();
 DECAPx6_ASAP7_75t_R FILLER_100_538 ();
 DECAPx2_ASAP7_75t_R FILLER_100_552 ();
 FILLER_ASAP7_75t_R FILLER_100_584 ();
 FILLER_ASAP7_75t_R FILLER_100_601 ();
 DECAPx4_ASAP7_75t_R FILLER_100_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_619 ();
 DECAPx2_ASAP7_75t_R FILLER_100_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_629 ();
 DECAPx2_ASAP7_75t_R FILLER_100_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_642 ();
 DECAPx4_ASAP7_75t_R FILLER_100_646 ();
 DECAPx1_ASAP7_75t_R FILLER_100_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_716 ();
 DECAPx1_ASAP7_75t_R FILLER_100_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_751 ();
 DECAPx1_ASAP7_75t_R FILLER_100_758 ();
 DECAPx1_ASAP7_75t_R FILLER_100_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_777 ();
 FILLER_ASAP7_75t_R FILLER_100_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_821 ();
 DECAPx4_ASAP7_75t_R FILLER_100_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_838 ();
 DECAPx2_ASAP7_75t_R FILLER_100_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_863 ();
 DECAPx1_ASAP7_75t_R FILLER_100_875 ();
 FILLER_ASAP7_75t_R FILLER_100_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_949 ();
 DECAPx2_ASAP7_75t_R FILLER_100_986 ();
 FILLER_ASAP7_75t_R FILLER_100_992 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1026 ();
 FILLER_ASAP7_75t_R FILLER_100_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1081 ();
 FILLER_ASAP7_75t_R FILLER_100_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1105 ();
 FILLER_ASAP7_75t_R FILLER_100_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1186 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1388 ();
 FILLER_ASAP7_75t_R FILLER_100_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_101_2 ();
 DECAPx1_ASAP7_75t_R FILLER_101_16 ();
 DECAPx2_ASAP7_75t_R FILLER_101_26 ();
 FILLER_ASAP7_75t_R FILLER_101_32 ();
 DECAPx6_ASAP7_75t_R FILLER_101_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_88 ();
 DECAPx2_ASAP7_75t_R FILLER_101_92 ();
 DECAPx1_ASAP7_75t_R FILLER_101_104 ();
 DECAPx6_ASAP7_75t_R FILLER_101_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_130 ();
 DECAPx1_ASAP7_75t_R FILLER_101_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_142 ();
 DECAPx2_ASAP7_75t_R FILLER_101_146 ();
 FILLER_ASAP7_75t_R FILLER_101_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_154 ();
 DECAPx6_ASAP7_75t_R FILLER_101_171 ();
 DECAPx1_ASAP7_75t_R FILLER_101_185 ();
 FILLER_ASAP7_75t_R FILLER_101_199 ();
 DECAPx1_ASAP7_75t_R FILLER_101_221 ();
 DECAPx1_ASAP7_75t_R FILLER_101_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_249 ();
 DECAPx6_ASAP7_75t_R FILLER_101_256 ();
 DECAPx1_ASAP7_75t_R FILLER_101_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_274 ();
 DECAPx2_ASAP7_75t_R FILLER_101_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_307 ();
 DECAPx2_ASAP7_75t_R FILLER_101_313 ();
 FILLER_ASAP7_75t_R FILLER_101_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_321 ();
 DECAPx2_ASAP7_75t_R FILLER_101_336 ();
 FILLER_ASAP7_75t_R FILLER_101_342 ();
 DECAPx10_ASAP7_75t_R FILLER_101_356 ();
 DECAPx6_ASAP7_75t_R FILLER_101_378 ();
 FILLER_ASAP7_75t_R FILLER_101_392 ();
 DECAPx2_ASAP7_75t_R FILLER_101_403 ();
 FILLER_ASAP7_75t_R FILLER_101_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_411 ();
 DECAPx6_ASAP7_75t_R FILLER_101_418 ();
 DECAPx1_ASAP7_75t_R FILLER_101_432 ();
 DECAPx6_ASAP7_75t_R FILLER_101_442 ();
 DECAPx10_ASAP7_75t_R FILLER_101_463 ();
 DECAPx10_ASAP7_75t_R FILLER_101_485 ();
 DECAPx2_ASAP7_75t_R FILLER_101_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_513 ();
 FILLER_ASAP7_75t_R FILLER_101_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_525 ();
 DECAPx10_ASAP7_75t_R FILLER_101_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_560 ();
 DECAPx1_ASAP7_75t_R FILLER_101_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_571 ();
 DECAPx10_ASAP7_75t_R FILLER_101_575 ();
 FILLER_ASAP7_75t_R FILLER_101_627 ();
 DECAPx6_ASAP7_75t_R FILLER_101_635 ();
 FILLER_ASAP7_75t_R FILLER_101_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_657 ();
 DECAPx4_ASAP7_75t_R FILLER_101_664 ();
 FILLER_ASAP7_75t_R FILLER_101_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_676 ();
 DECAPx2_ASAP7_75t_R FILLER_101_685 ();
 FILLER_ASAP7_75t_R FILLER_101_691 ();
 DECAPx6_ASAP7_75t_R FILLER_101_696 ();
 FILLER_ASAP7_75t_R FILLER_101_710 ();
 FILLER_ASAP7_75t_R FILLER_101_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_780 ();
 FILLER_ASAP7_75t_R FILLER_101_789 ();
 FILLER_ASAP7_75t_R FILLER_101_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_799 ();
 DECAPx6_ASAP7_75t_R FILLER_101_841 ();
 FILLER_ASAP7_75t_R FILLER_101_855 ();
 DECAPx2_ASAP7_75t_R FILLER_101_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_873 ();
 DECAPx2_ASAP7_75t_R FILLER_101_882 ();
 FILLER_ASAP7_75t_R FILLER_101_888 ();
 DECAPx1_ASAP7_75t_R FILLER_101_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_923 ();
 DECAPx2_ASAP7_75t_R FILLER_101_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_932 ();
 DECAPx6_ASAP7_75t_R FILLER_101_939 ();
 DECAPx4_ASAP7_75t_R FILLER_101_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_969 ();
 DECAPx2_ASAP7_75t_R FILLER_101_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_994 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1053 ();
 FILLER_ASAP7_75t_R FILLER_101_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1068 ();
 FILLER_ASAP7_75t_R FILLER_101_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1080 ();
 FILLER_ASAP7_75t_R FILLER_101_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1127 ();
 FILLER_ASAP7_75t_R FILLER_101_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1397 ();
 FILLER_ASAP7_75t_R FILLER_101_1403 ();
 DECAPx4_ASAP7_75t_R FILLER_102_2 ();
 FILLER_ASAP7_75t_R FILLER_102_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_36 ();
 DECAPx2_ASAP7_75t_R FILLER_102_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_49 ();
 FILLER_ASAP7_75t_R FILLER_102_59 ();
 DECAPx4_ASAP7_75t_R FILLER_102_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_100 ();
 DECAPx6_ASAP7_75t_R FILLER_102_179 ();
 FILLER_ASAP7_75t_R FILLER_102_193 ();
 FILLER_ASAP7_75t_R FILLER_102_215 ();
 DECAPx2_ASAP7_75t_R FILLER_102_225 ();
 DECAPx1_ASAP7_75t_R FILLER_102_237 ();
 DECAPx6_ASAP7_75t_R FILLER_102_263 ();
 FILLER_ASAP7_75t_R FILLER_102_277 ();
 DECAPx1_ASAP7_75t_R FILLER_102_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_289 ();
 DECAPx4_ASAP7_75t_R FILLER_102_293 ();
 FILLER_ASAP7_75t_R FILLER_102_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_305 ();
 DECAPx10_ASAP7_75t_R FILLER_102_314 ();
 DECAPx6_ASAP7_75t_R FILLER_102_336 ();
 FILLER_ASAP7_75t_R FILLER_102_350 ();
 DECAPx2_ASAP7_75t_R FILLER_102_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_370 ();
 DECAPx6_ASAP7_75t_R FILLER_102_384 ();
 DECAPx1_ASAP7_75t_R FILLER_102_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_402 ();
 FILLER_ASAP7_75t_R FILLER_102_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_421 ();
 DECAPx6_ASAP7_75t_R FILLER_102_436 ();
 DECAPx2_ASAP7_75t_R FILLER_102_456 ();
 DECAPx2_ASAP7_75t_R FILLER_102_498 ();
 DECAPx6_ASAP7_75t_R FILLER_102_512 ();
 DECAPx4_ASAP7_75t_R FILLER_102_536 ();
 FILLER_ASAP7_75t_R FILLER_102_546 ();
 DECAPx10_ASAP7_75t_R FILLER_102_558 ();
 FILLER_ASAP7_75t_R FILLER_102_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_599 ();
 FILLER_ASAP7_75t_R FILLER_102_632 ();
 FILLER_ASAP7_75t_R FILLER_102_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_642 ();
 DECAPx2_ASAP7_75t_R FILLER_102_675 ();
 FILLER_ASAP7_75t_R FILLER_102_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_683 ();
 DECAPx1_ASAP7_75t_R FILLER_102_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_710 ();
 DECAPx10_ASAP7_75t_R FILLER_102_717 ();
 DECAPx6_ASAP7_75t_R FILLER_102_739 ();
 DECAPx1_ASAP7_75t_R FILLER_102_753 ();
 FILLER_ASAP7_75t_R FILLER_102_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_765 ();
 DECAPx1_ASAP7_75t_R FILLER_102_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_776 ();
 DECAPx10_ASAP7_75t_R FILLER_102_780 ();
 DECAPx1_ASAP7_75t_R FILLER_102_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_806 ();
 DECAPx1_ASAP7_75t_R FILLER_102_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_814 ();
 DECAPx10_ASAP7_75t_R FILLER_102_818 ();
 DECAPx10_ASAP7_75t_R FILLER_102_840 ();
 DECAPx10_ASAP7_75t_R FILLER_102_862 ();
 DECAPx10_ASAP7_75t_R FILLER_102_884 ();
 DECAPx10_ASAP7_75t_R FILLER_102_906 ();
 DECAPx6_ASAP7_75t_R FILLER_102_928 ();
 DECAPx2_ASAP7_75t_R FILLER_102_942 ();
 DECAPx1_ASAP7_75t_R FILLER_102_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_958 ();
 DECAPx2_ASAP7_75t_R FILLER_102_962 ();
 FILLER_ASAP7_75t_R FILLER_102_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_970 ();
 DECAPx10_ASAP7_75t_R FILLER_102_983 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1005 ();
 FILLER_ASAP7_75t_R FILLER_102_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1029 ();
 FILLER_ASAP7_75t_R FILLER_102_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1101 ();
 FILLER_ASAP7_75t_R FILLER_102_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1165 ();
 FILLER_ASAP7_75t_R FILLER_102_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1361 ();
 FILLER_ASAP7_75t_R FILLER_102_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1388 ();
 FILLER_ASAP7_75t_R FILLER_102_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_103_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_46 ();
 FILLER_ASAP7_75t_R FILLER_103_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_75 ();
 DECAPx10_ASAP7_75t_R FILLER_103_82 ();
 DECAPx6_ASAP7_75t_R FILLER_103_120 ();
 FILLER_ASAP7_75t_R FILLER_103_134 ();
 DECAPx6_ASAP7_75t_R FILLER_103_142 ();
 DECAPx2_ASAP7_75t_R FILLER_103_156 ();
 FILLER_ASAP7_75t_R FILLER_103_176 ();
 DECAPx4_ASAP7_75t_R FILLER_103_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_208 ();
 DECAPx6_ASAP7_75t_R FILLER_103_229 ();
 DECAPx1_ASAP7_75t_R FILLER_103_243 ();
 DECAPx4_ASAP7_75t_R FILLER_103_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_263 ();
 DECAPx10_ASAP7_75t_R FILLER_103_270 ();
 DECAPx4_ASAP7_75t_R FILLER_103_292 ();
 FILLER_ASAP7_75t_R FILLER_103_302 ();
 DECAPx10_ASAP7_75t_R FILLER_103_310 ();
 DECAPx10_ASAP7_75t_R FILLER_103_332 ();
 DECAPx10_ASAP7_75t_R FILLER_103_354 ();
 DECAPx10_ASAP7_75t_R FILLER_103_376 ();
 DECAPx10_ASAP7_75t_R FILLER_103_398 ();
 DECAPx6_ASAP7_75t_R FILLER_103_420 ();
 DECAPx2_ASAP7_75t_R FILLER_103_434 ();
 DECAPx6_ASAP7_75t_R FILLER_103_462 ();
 DECAPx1_ASAP7_75t_R FILLER_103_476 ();
 DECAPx6_ASAP7_75t_R FILLER_103_486 ();
 FILLER_ASAP7_75t_R FILLER_103_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_502 ();
 DECAPx2_ASAP7_75t_R FILLER_103_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_535 ();
 DECAPx1_ASAP7_75t_R FILLER_103_564 ();
 FILLER_ASAP7_75t_R FILLER_103_575 ();
 DECAPx2_ASAP7_75t_R FILLER_103_655 ();
 FILLER_ASAP7_75t_R FILLER_103_661 ();
 DECAPx10_ASAP7_75t_R FILLER_103_666 ();
 DECAPx1_ASAP7_75t_R FILLER_103_688 ();
 FILLER_ASAP7_75t_R FILLER_103_730 ();
 DECAPx10_ASAP7_75t_R FILLER_103_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_764 ();
 DECAPx6_ASAP7_75t_R FILLER_103_771 ();
 FILLER_ASAP7_75t_R FILLER_103_797 ();
 DECAPx2_ASAP7_75t_R FILLER_103_802 ();
 FILLER_ASAP7_75t_R FILLER_103_808 ();
 DECAPx2_ASAP7_75t_R FILLER_103_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_822 ();
 DECAPx4_ASAP7_75t_R FILLER_103_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_845 ();
 DECAPx4_ASAP7_75t_R FILLER_103_858 ();
 DECAPx2_ASAP7_75t_R FILLER_103_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_884 ();
 DECAPx6_ASAP7_75t_R FILLER_103_891 ();
 FILLER_ASAP7_75t_R FILLER_103_905 ();
 DECAPx1_ASAP7_75t_R FILLER_103_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_923 ();
 DECAPx1_ASAP7_75t_R FILLER_103_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_930 ();
 DECAPx2_ASAP7_75t_R FILLER_103_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_944 ();
 DECAPx6_ASAP7_75t_R FILLER_103_951 ();
 DECAPx1_ASAP7_75t_R FILLER_103_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_981 ();
 DECAPx2_ASAP7_75t_R FILLER_103_989 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1054 ();
 FILLER_ASAP7_75t_R FILLER_103_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1134 ();
 FILLER_ASAP7_75t_R FILLER_103_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1154 ();
 FILLER_ASAP7_75t_R FILLER_103_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1386 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_104_2 ();
 FILLER_ASAP7_75t_R FILLER_104_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_14 ();
 DECAPx10_ASAP7_75t_R FILLER_104_18 ();
 FILLER_ASAP7_75t_R FILLER_104_40 ();
 FILLER_ASAP7_75t_R FILLER_104_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_50 ();
 FILLER_ASAP7_75t_R FILLER_104_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_91 ();
 DECAPx2_ASAP7_75t_R FILLER_104_95 ();
 DECAPx2_ASAP7_75t_R FILLER_104_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_111 ();
 FILLER_ASAP7_75t_R FILLER_104_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_120 ();
 DECAPx2_ASAP7_75t_R FILLER_104_124 ();
 DECAPx6_ASAP7_75t_R FILLER_104_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_151 ();
 FILLER_ASAP7_75t_R FILLER_104_162 ();
 DECAPx10_ASAP7_75t_R FILLER_104_192 ();
 DECAPx2_ASAP7_75t_R FILLER_104_214 ();
 DECAPx1_ASAP7_75t_R FILLER_104_226 ();
 DECAPx6_ASAP7_75t_R FILLER_104_244 ();
 FILLER_ASAP7_75t_R FILLER_104_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_260 ();
 DECAPx2_ASAP7_75t_R FILLER_104_267 ();
 FILLER_ASAP7_75t_R FILLER_104_273 ();
 DECAPx4_ASAP7_75t_R FILLER_104_295 ();
 DECAPx2_ASAP7_75t_R FILLER_104_313 ();
 FILLER_ASAP7_75t_R FILLER_104_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_321 ();
 DECAPx2_ASAP7_75t_R FILLER_104_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_342 ();
 DECAPx6_ASAP7_75t_R FILLER_104_357 ();
 DECAPx4_ASAP7_75t_R FILLER_104_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_388 ();
 DECAPx10_ASAP7_75t_R FILLER_104_414 ();
 DECAPx4_ASAP7_75t_R FILLER_104_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_446 ();
 DECAPx2_ASAP7_75t_R FILLER_104_456 ();
 DECAPx10_ASAP7_75t_R FILLER_104_464 ();
 DECAPx6_ASAP7_75t_R FILLER_104_486 ();
 FILLER_ASAP7_75t_R FILLER_104_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_502 ();
 FILLER_ASAP7_75t_R FILLER_104_516 ();
 DECAPx10_ASAP7_75t_R FILLER_104_521 ();
 DECAPx1_ASAP7_75t_R FILLER_104_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_547 ();
 DECAPx2_ASAP7_75t_R FILLER_104_554 ();
 FILLER_ASAP7_75t_R FILLER_104_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_562 ();
 DECAPx4_ASAP7_75t_R FILLER_104_595 ();
 FILLER_ASAP7_75t_R FILLER_104_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_619 ();
 DECAPx2_ASAP7_75t_R FILLER_104_623 ();
 FILLER_ASAP7_75t_R FILLER_104_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_643 ();
 DECAPx4_ASAP7_75t_R FILLER_104_647 ();
 FILLER_ASAP7_75t_R FILLER_104_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_697 ();
 DECAPx2_ASAP7_75t_R FILLER_104_704 ();
 FILLER_ASAP7_75t_R FILLER_104_710 ();
 DECAPx2_ASAP7_75t_R FILLER_104_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_749 ();
 FILLER_ASAP7_75t_R FILLER_104_768 ();
 FILLER_ASAP7_75t_R FILLER_104_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_778 ();
 FILLER_ASAP7_75t_R FILLER_104_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_784 ();
 FILLER_ASAP7_75t_R FILLER_104_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_868 ();
 DECAPx2_ASAP7_75t_R FILLER_104_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_913 ();
 DECAPx6_ASAP7_75t_R FILLER_104_928 ();
 DECAPx2_ASAP7_75t_R FILLER_104_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_948 ();
 DECAPx10_ASAP7_75t_R FILLER_104_980 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1078 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1116 ();
 FILLER_ASAP7_75t_R FILLER_104_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1388 ();
 FILLER_ASAP7_75t_R FILLER_104_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_105_2 ();
 FILLER_ASAP7_75t_R FILLER_105_8 ();
 DECAPx2_ASAP7_75t_R FILLER_105_16 ();
 FILLER_ASAP7_75t_R FILLER_105_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_57 ();
 DECAPx1_ASAP7_75t_R FILLER_105_73 ();
 DECAPx10_ASAP7_75t_R FILLER_105_155 ();
 FILLER_ASAP7_75t_R FILLER_105_177 ();
 DECAPx6_ASAP7_75t_R FILLER_105_201 ();
 DECAPx2_ASAP7_75t_R FILLER_105_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_221 ();
 DECAPx1_ASAP7_75t_R FILLER_105_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_242 ();
 FILLER_ASAP7_75t_R FILLER_105_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_251 ();
 DECAPx4_ASAP7_75t_R FILLER_105_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_290 ();
 DECAPx4_ASAP7_75t_R FILLER_105_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_321 ();
 DECAPx2_ASAP7_75t_R FILLER_105_334 ();
 DECAPx4_ASAP7_75t_R FILLER_105_346 ();
 FILLER_ASAP7_75t_R FILLER_105_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_358 ();
 DECAPx6_ASAP7_75t_R FILLER_105_373 ();
 DECAPx10_ASAP7_75t_R FILLER_105_393 ();
 DECAPx1_ASAP7_75t_R FILLER_105_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_419 ();
 DECAPx6_ASAP7_75t_R FILLER_105_432 ();
 DECAPx1_ASAP7_75t_R FILLER_105_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_456 ();
 FILLER_ASAP7_75t_R FILLER_105_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_465 ();
 DECAPx1_ASAP7_75t_R FILLER_105_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_484 ();
 DECAPx10_ASAP7_75t_R FILLER_105_491 ();
 DECAPx6_ASAP7_75t_R FILLER_105_513 ();
 FILLER_ASAP7_75t_R FILLER_105_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_529 ();
 DECAPx10_ASAP7_75t_R FILLER_105_540 ();
 DECAPx10_ASAP7_75t_R FILLER_105_562 ();
 DECAPx10_ASAP7_75t_R FILLER_105_587 ();
 DECAPx2_ASAP7_75t_R FILLER_105_609 ();
 DECAPx2_ASAP7_75t_R FILLER_105_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_633 ();
 DECAPx6_ASAP7_75t_R FILLER_105_638 ();
 FILLER_ASAP7_75t_R FILLER_105_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_654 ();
 FILLER_ASAP7_75t_R FILLER_105_661 ();
 DECAPx2_ASAP7_75t_R FILLER_105_672 ();
 FILLER_ASAP7_75t_R FILLER_105_678 ();
 FILLER_ASAP7_75t_R FILLER_105_683 ();
 DECAPx10_ASAP7_75t_R FILLER_105_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_711 ();
 DECAPx10_ASAP7_75t_R FILLER_105_715 ();
 DECAPx2_ASAP7_75t_R FILLER_105_737 ();
 FILLER_ASAP7_75t_R FILLER_105_753 ();
 DECAPx6_ASAP7_75t_R FILLER_105_810 ();
 DECAPx2_ASAP7_75t_R FILLER_105_832 ();
 FILLER_ASAP7_75t_R FILLER_105_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_840 ();
 FILLER_ASAP7_75t_R FILLER_105_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_867 ();
 DECAPx4_ASAP7_75t_R FILLER_105_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_884 ();
 DECAPx10_ASAP7_75t_R FILLER_105_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_923 ();
 DECAPx2_ASAP7_75t_R FILLER_105_926 ();
 DECAPx1_ASAP7_75t_R FILLER_105_945 ();
 DECAPx4_ASAP7_75t_R FILLER_105_956 ();
 FILLER_ASAP7_75t_R FILLER_105_966 ();
 DECAPx6_ASAP7_75t_R FILLER_105_974 ();
 FILLER_ASAP7_75t_R FILLER_105_988 ();
 FILLER_ASAP7_75t_R FILLER_105_999 ();
 DECAPx1_ASAP7_75t_R FILLER_105_1037 ();
 FILLER_ASAP7_75t_R FILLER_105_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_105_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1095 ();
 FILLER_ASAP7_75t_R FILLER_105_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1404 ();
 FILLER_ASAP7_75t_R FILLER_106_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_4 ();
 DECAPx1_ASAP7_75t_R FILLER_106_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_44 ();
 DECAPx10_ASAP7_75t_R FILLER_106_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_70 ();
 DECAPx1_ASAP7_75t_R FILLER_106_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_78 ();
 DECAPx2_ASAP7_75t_R FILLER_106_85 ();
 FILLER_ASAP7_75t_R FILLER_106_91 ();
 DECAPx4_ASAP7_75t_R FILLER_106_99 ();
 DECAPx6_ASAP7_75t_R FILLER_106_115 ();
 DECAPx2_ASAP7_75t_R FILLER_106_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_135 ();
 FILLER_ASAP7_75t_R FILLER_106_142 ();
 DECAPx6_ASAP7_75t_R FILLER_106_147 ();
 DECAPx6_ASAP7_75t_R FILLER_106_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_189 ();
 FILLER_ASAP7_75t_R FILLER_106_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_198 ();
 DECAPx6_ASAP7_75t_R FILLER_106_211 ();
 DECAPx2_ASAP7_75t_R FILLER_106_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_231 ();
 DECAPx1_ASAP7_75t_R FILLER_106_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_242 ();
 DECAPx10_ASAP7_75t_R FILLER_106_256 ();
 FILLER_ASAP7_75t_R FILLER_106_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_280 ();
 DECAPx10_ASAP7_75t_R FILLER_106_287 ();
 DECAPx10_ASAP7_75t_R FILLER_106_309 ();
 DECAPx4_ASAP7_75t_R FILLER_106_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_341 ();
 DECAPx10_ASAP7_75t_R FILLER_106_348 ();
 DECAPx10_ASAP7_75t_R FILLER_106_370 ();
 DECAPx10_ASAP7_75t_R FILLER_106_392 ();
 FILLER_ASAP7_75t_R FILLER_106_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_416 ();
 DECAPx2_ASAP7_75t_R FILLER_106_425 ();
 DECAPx4_ASAP7_75t_R FILLER_106_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_449 ();
 DECAPx1_ASAP7_75t_R FILLER_106_458 ();
 DECAPx2_ASAP7_75t_R FILLER_106_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_470 ();
 FILLER_ASAP7_75t_R FILLER_106_491 ();
 DECAPx10_ASAP7_75t_R FILLER_106_499 ();
 DECAPx2_ASAP7_75t_R FILLER_106_521 ();
 FILLER_ASAP7_75t_R FILLER_106_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_529 ();
 FILLER_ASAP7_75t_R FILLER_106_536 ();
 FILLER_ASAP7_75t_R FILLER_106_565 ();
 DECAPx4_ASAP7_75t_R FILLER_106_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_647 ();
 DECAPx6_ASAP7_75t_R FILLER_106_680 ();
 FILLER_ASAP7_75t_R FILLER_106_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_714 ();
 DECAPx6_ASAP7_75t_R FILLER_106_741 ();
 FILLER_ASAP7_75t_R FILLER_106_755 ();
 DECAPx2_ASAP7_75t_R FILLER_106_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_769 ();
 DECAPx6_ASAP7_75t_R FILLER_106_773 ();
 FILLER_ASAP7_75t_R FILLER_106_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_789 ();
 DECAPx4_ASAP7_75t_R FILLER_106_799 ();
 FILLER_ASAP7_75t_R FILLER_106_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_811 ();
 DECAPx2_ASAP7_75t_R FILLER_106_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_828 ();
 DECAPx10_ASAP7_75t_R FILLER_106_843 ();
 DECAPx2_ASAP7_75t_R FILLER_106_865 ();
 FILLER_ASAP7_75t_R FILLER_106_871 ();
 FILLER_ASAP7_75t_R FILLER_106_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_885 ();
 FILLER_ASAP7_75t_R FILLER_106_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_902 ();
 FILLER_ASAP7_75t_R FILLER_106_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_917 ();
 DECAPx2_ASAP7_75t_R FILLER_106_939 ();
 DECAPx6_ASAP7_75t_R FILLER_106_951 ();
 FILLER_ASAP7_75t_R FILLER_106_981 ();
 DECAPx6_ASAP7_75t_R FILLER_106_998 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1097 ();
 FILLER_ASAP7_75t_R FILLER_106_1104 ();
 FILLER_ASAP7_75t_R FILLER_106_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1114 ();
 FILLER_ASAP7_75t_R FILLER_106_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1388 ();
 FILLER_ASAP7_75t_R FILLER_106_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1404 ();
 FILLER_ASAP7_75t_R FILLER_107_28 ();
 DECAPx10_ASAP7_75t_R FILLER_107_34 ();
 DECAPx4_ASAP7_75t_R FILLER_107_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_72 ();
 FILLER_ASAP7_75t_R FILLER_107_79 ();
 DECAPx6_ASAP7_75t_R FILLER_107_113 ();
 DECAPx2_ASAP7_75t_R FILLER_107_127 ();
 DECAPx2_ASAP7_75t_R FILLER_107_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_146 ();
 DECAPx2_ASAP7_75t_R FILLER_107_150 ();
 FILLER_ASAP7_75t_R FILLER_107_156 ();
 DECAPx2_ASAP7_75t_R FILLER_107_186 ();
 FILLER_ASAP7_75t_R FILLER_107_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_194 ();
 DECAPx10_ASAP7_75t_R FILLER_107_223 ();
 DECAPx1_ASAP7_75t_R FILLER_107_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_249 ();
 DECAPx1_ASAP7_75t_R FILLER_107_264 ();
 DECAPx4_ASAP7_75t_R FILLER_107_282 ();
 DECAPx6_ASAP7_75t_R FILLER_107_305 ();
 DECAPx2_ASAP7_75t_R FILLER_107_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_325 ();
 DECAPx6_ASAP7_75t_R FILLER_107_334 ();
 DECAPx2_ASAP7_75t_R FILLER_107_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_354 ();
 DECAPx6_ASAP7_75t_R FILLER_107_363 ();
 FILLER_ASAP7_75t_R FILLER_107_377 ();
 DECAPx1_ASAP7_75t_R FILLER_107_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_399 ();
 DECAPx1_ASAP7_75t_R FILLER_107_412 ();
 DECAPx10_ASAP7_75t_R FILLER_107_422 ();
 DECAPx10_ASAP7_75t_R FILLER_107_444 ();
 DECAPx4_ASAP7_75t_R FILLER_107_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_476 ();
 DECAPx1_ASAP7_75t_R FILLER_107_485 ();
 DECAPx2_ASAP7_75t_R FILLER_107_495 ();
 FILLER_ASAP7_75t_R FILLER_107_501 ();
 DECAPx1_ASAP7_75t_R FILLER_107_520 ();
 FILLER_ASAP7_75t_R FILLER_107_546 ();
 DECAPx4_ASAP7_75t_R FILLER_107_554 ();
 FILLER_ASAP7_75t_R FILLER_107_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_566 ();
 FILLER_ASAP7_75t_R FILLER_107_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_628 ();
 DECAPx1_ASAP7_75t_R FILLER_107_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_665 ();
 DECAPx1_ASAP7_75t_R FILLER_107_698 ();
 FILLER_ASAP7_75t_R FILLER_107_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_746 ();
 FILLER_ASAP7_75t_R FILLER_107_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_759 ();
 DECAPx6_ASAP7_75t_R FILLER_107_788 ();
 DECAPx4_ASAP7_75t_R FILLER_107_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_822 ();
 DECAPx6_ASAP7_75t_R FILLER_107_839 ();
 DECAPx1_ASAP7_75t_R FILLER_107_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_857 ();
 DECAPx2_ASAP7_75t_R FILLER_107_874 ();
 DECAPx6_ASAP7_75t_R FILLER_107_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_901 ();
 DECAPx4_ASAP7_75t_R FILLER_107_914 ();
 DECAPx6_ASAP7_75t_R FILLER_107_926 ();
 DECAPx1_ASAP7_75t_R FILLER_107_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_944 ();
 DECAPx6_ASAP7_75t_R FILLER_107_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_966 ();
 DECAPx1_ASAP7_75t_R FILLER_107_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_977 ();
 DECAPx2_ASAP7_75t_R FILLER_107_992 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_107_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1055 ();
 FILLER_ASAP7_75t_R FILLER_107_1061 ();
 FILLER_ASAP7_75t_R FILLER_107_1072 ();
 FILLER_ASAP7_75t_R FILLER_107_1086 ();
 FILLER_ASAP7_75t_R FILLER_107_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1133 ();
 FILLER_ASAP7_75t_R FILLER_107_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1256 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1369 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1391 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_7 ();
 FILLER_ASAP7_75t_R FILLER_108_14 ();
 FILLER_ASAP7_75t_R FILLER_108_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_30 ();
 FILLER_ASAP7_75t_R FILLER_108_37 ();
 DECAPx2_ASAP7_75t_R FILLER_108_42 ();
 FILLER_ASAP7_75t_R FILLER_108_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_59 ();
 DECAPx1_ASAP7_75t_R FILLER_108_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_93 ();
 FILLER_ASAP7_75t_R FILLER_108_129 ();
 DECAPx2_ASAP7_75t_R FILLER_108_183 ();
 FILLER_ASAP7_75t_R FILLER_108_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_191 ();
 DECAPx4_ASAP7_75t_R FILLER_108_200 ();
 DECAPx10_ASAP7_75t_R FILLER_108_236 ();
 DECAPx2_ASAP7_75t_R FILLER_108_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_264 ();
 DECAPx1_ASAP7_75t_R FILLER_108_313 ();
 FILLER_ASAP7_75t_R FILLER_108_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_329 ();
 DECAPx6_ASAP7_75t_R FILLER_108_339 ();
 DECAPx1_ASAP7_75t_R FILLER_108_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_357 ();
 DECAPx1_ASAP7_75t_R FILLER_108_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_370 ();
 DECAPx2_ASAP7_75t_R FILLER_108_384 ();
 DECAPx1_ASAP7_75t_R FILLER_108_416 ();
 DECAPx6_ASAP7_75t_R FILLER_108_432 ();
 FILLER_ASAP7_75t_R FILLER_108_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_448 ();
 DECAPx2_ASAP7_75t_R FILLER_108_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_461 ();
 DECAPx10_ASAP7_75t_R FILLER_108_464 ();
 DECAPx4_ASAP7_75t_R FILLER_108_486 ();
 FILLER_ASAP7_75t_R FILLER_108_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_498 ();
 DECAPx10_ASAP7_75t_R FILLER_108_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_529 ();
 DECAPx4_ASAP7_75t_R FILLER_108_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_546 ();
 FILLER_ASAP7_75t_R FILLER_108_579 ();
 FILLER_ASAP7_75t_R FILLER_108_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_602 ();
 FILLER_ASAP7_75t_R FILLER_108_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_615 ();
 DECAPx4_ASAP7_75t_R FILLER_108_619 ();
 FILLER_ASAP7_75t_R FILLER_108_632 ();
 DECAPx4_ASAP7_75t_R FILLER_108_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_650 ();
 DECAPx2_ASAP7_75t_R FILLER_108_657 ();
 DECAPx1_ASAP7_75t_R FILLER_108_669 ();
 DECAPx2_ASAP7_75t_R FILLER_108_679 ();
 FILLER_ASAP7_75t_R FILLER_108_685 ();
 FILLER_ASAP7_75t_R FILLER_108_690 ();
 DECAPx1_ASAP7_75t_R FILLER_108_724 ();
 DECAPx10_ASAP7_75t_R FILLER_108_734 ();
 DECAPx10_ASAP7_75t_R FILLER_108_756 ();
 FILLER_ASAP7_75t_R FILLER_108_778 ();
 FILLER_ASAP7_75t_R FILLER_108_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_789 ();
 DECAPx1_ASAP7_75t_R FILLER_108_808 ();
 DECAPx2_ASAP7_75t_R FILLER_108_836 ();
 FILLER_ASAP7_75t_R FILLER_108_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_960 ();
 DECAPx6_ASAP7_75t_R FILLER_108_977 ();
 DECAPx1_ASAP7_75t_R FILLER_108_991 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1090 ();
 FILLER_ASAP7_75t_R FILLER_108_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1102 ();
 FILLER_ASAP7_75t_R FILLER_108_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1130 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1202 ();
 FILLER_ASAP7_75t_R FILLER_108_1208 ();
 FILLER_ASAP7_75t_R FILLER_108_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1294 ();
 FILLER_ASAP7_75t_R FILLER_108_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1377 ();
 FILLER_ASAP7_75t_R FILLER_108_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1388 ();
 FILLER_ASAP7_75t_R FILLER_108_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_109_2 ();
 FILLER_ASAP7_75t_R FILLER_109_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_18 ();
 DECAPx2_ASAP7_75t_R FILLER_109_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_77 ();
 DECAPx6_ASAP7_75t_R FILLER_109_81 ();
 DECAPx2_ASAP7_75t_R FILLER_109_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_101 ();
 FILLER_ASAP7_75t_R FILLER_109_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_113 ();
 DECAPx6_ASAP7_75t_R FILLER_109_117 ();
 DECAPx6_ASAP7_75t_R FILLER_109_144 ();
 DECAPx2_ASAP7_75t_R FILLER_109_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_170 ();
 DECAPx2_ASAP7_75t_R FILLER_109_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_201 ();
 DECAPx1_ASAP7_75t_R FILLER_109_214 ();
 DECAPx10_ASAP7_75t_R FILLER_109_241 ();
 DECAPx2_ASAP7_75t_R FILLER_109_263 ();
 FILLER_ASAP7_75t_R FILLER_109_269 ();
 DECAPx1_ASAP7_75t_R FILLER_109_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_283 ();
 DECAPx2_ASAP7_75t_R FILLER_109_294 ();
 FILLER_ASAP7_75t_R FILLER_109_300 ();
 DECAPx2_ASAP7_75t_R FILLER_109_305 ();
 DECAPx2_ASAP7_75t_R FILLER_109_329 ();
 FILLER_ASAP7_75t_R FILLER_109_335 ();
 FILLER_ASAP7_75t_R FILLER_109_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_351 ();
 DECAPx10_ASAP7_75t_R FILLER_109_366 ();
 DECAPx4_ASAP7_75t_R FILLER_109_388 ();
 FILLER_ASAP7_75t_R FILLER_109_398 ();
 DECAPx2_ASAP7_75t_R FILLER_109_409 ();
 FILLER_ASAP7_75t_R FILLER_109_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_417 ();
 DECAPx2_ASAP7_75t_R FILLER_109_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_462 ();
 FILLER_ASAP7_75t_R FILLER_109_471 ();
 DECAPx10_ASAP7_75t_R FILLER_109_479 ();
 DECAPx10_ASAP7_75t_R FILLER_109_501 ();
 DECAPx10_ASAP7_75t_R FILLER_109_523 ();
 FILLER_ASAP7_75t_R FILLER_109_545 ();
 DECAPx2_ASAP7_75t_R FILLER_109_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_560 ();
 DECAPx10_ASAP7_75t_R FILLER_109_564 ();
 DECAPx10_ASAP7_75t_R FILLER_109_586 ();
 DECAPx10_ASAP7_75t_R FILLER_109_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_630 ();
 DECAPx4_ASAP7_75t_R FILLER_109_673 ();
 FILLER_ASAP7_75t_R FILLER_109_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_688 ();
 DECAPx10_ASAP7_75t_R FILLER_109_693 ();
 DECAPx10_ASAP7_75t_R FILLER_109_715 ();
 DECAPx2_ASAP7_75t_R FILLER_109_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_743 ();
 DECAPx4_ASAP7_75t_R FILLER_109_753 ();
 FILLER_ASAP7_75t_R FILLER_109_782 ();
 FILLER_ASAP7_75t_R FILLER_109_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_819 ();
 DECAPx1_ASAP7_75t_R FILLER_109_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_867 ();
 DECAPx2_ASAP7_75t_R FILLER_109_876 ();
 DECAPx4_ASAP7_75t_R FILLER_109_894 ();
 FILLER_ASAP7_75t_R FILLER_109_904 ();
 DECAPx2_ASAP7_75t_R FILLER_109_918 ();
 DECAPx4_ASAP7_75t_R FILLER_109_926 ();
 FILLER_ASAP7_75t_R FILLER_109_936 ();
 DECAPx6_ASAP7_75t_R FILLER_109_962 ();
 DECAPx1_ASAP7_75t_R FILLER_109_986 ();
 DECAPx4_ASAP7_75t_R FILLER_109_998 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1020 ();
 FILLER_ASAP7_75t_R FILLER_109_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1061 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1235 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1361 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_7 ();
 DECAPx1_ASAP7_75t_R FILLER_110_23 ();
 DECAPx6_ASAP7_75t_R FILLER_110_33 ();
 FILLER_ASAP7_75t_R FILLER_110_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_49 ();
 DECAPx2_ASAP7_75t_R FILLER_110_56 ();
 FILLER_ASAP7_75t_R FILLER_110_62 ();
 DECAPx4_ASAP7_75t_R FILLER_110_67 ();
 FILLER_ASAP7_75t_R FILLER_110_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_79 ();
 DECAPx1_ASAP7_75t_R FILLER_110_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_90 ();
 DECAPx1_ASAP7_75t_R FILLER_110_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_101 ();
 DECAPx10_ASAP7_75t_R FILLER_110_105 ();
 FILLER_ASAP7_75t_R FILLER_110_127 ();
 DECAPx10_ASAP7_75t_R FILLER_110_162 ();
 FILLER_ASAP7_75t_R FILLER_110_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_186 ();
 DECAPx2_ASAP7_75t_R FILLER_110_201 ();
 FILLER_ASAP7_75t_R FILLER_110_226 ();
 FILLER_ASAP7_75t_R FILLER_110_234 ();
 DECAPx4_ASAP7_75t_R FILLER_110_258 ();
 FILLER_ASAP7_75t_R FILLER_110_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_270 ();
 DECAPx4_ASAP7_75t_R FILLER_110_281 ();
 DECAPx10_ASAP7_75t_R FILLER_110_301 ();
 DECAPx10_ASAP7_75t_R FILLER_110_323 ();
 DECAPx10_ASAP7_75t_R FILLER_110_345 ();
 DECAPx1_ASAP7_75t_R FILLER_110_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_371 ();
 DECAPx10_ASAP7_75t_R FILLER_110_384 ();
 DECAPx10_ASAP7_75t_R FILLER_110_406 ();
 DECAPx2_ASAP7_75t_R FILLER_110_438 ();
 FILLER_ASAP7_75t_R FILLER_110_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_446 ();
 DECAPx2_ASAP7_75t_R FILLER_110_453 ();
 FILLER_ASAP7_75t_R FILLER_110_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_478 ();
 FILLER_ASAP7_75t_R FILLER_110_485 ();
 DECAPx1_ASAP7_75t_R FILLER_110_493 ();
 DECAPx10_ASAP7_75t_R FILLER_110_503 ();
 DECAPx6_ASAP7_75t_R FILLER_110_525 ();
 DECAPx2_ASAP7_75t_R FILLER_110_539 ();
 DECAPx10_ASAP7_75t_R FILLER_110_553 ();
 DECAPx2_ASAP7_75t_R FILLER_110_575 ();
 FILLER_ASAP7_75t_R FILLER_110_581 ();
 DECAPx4_ASAP7_75t_R FILLER_110_589 ();
 DECAPx1_ASAP7_75t_R FILLER_110_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_613 ();
 FILLER_ASAP7_75t_R FILLER_110_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_631 ();
 DECAPx10_ASAP7_75t_R FILLER_110_635 ();
 DECAPx4_ASAP7_75t_R FILLER_110_657 ();
 FILLER_ASAP7_75t_R FILLER_110_667 ();
 FILLER_ASAP7_75t_R FILLER_110_705 ();
 DECAPx10_ASAP7_75t_R FILLER_110_733 ();
 DECAPx1_ASAP7_75t_R FILLER_110_755 ();
 DECAPx1_ASAP7_75t_R FILLER_110_765 ();
 FILLER_ASAP7_75t_R FILLER_110_781 ();
 DECAPx6_ASAP7_75t_R FILLER_110_790 ();
 FILLER_ASAP7_75t_R FILLER_110_804 ();
 DECAPx2_ASAP7_75t_R FILLER_110_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_819 ();
 DECAPx6_ASAP7_75t_R FILLER_110_826 ();
 FILLER_ASAP7_75t_R FILLER_110_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_842 ();
 DECAPx6_ASAP7_75t_R FILLER_110_851 ();
 DECAPx1_ASAP7_75t_R FILLER_110_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_869 ();
 DECAPx2_ASAP7_75t_R FILLER_110_886 ();
 FILLER_ASAP7_75t_R FILLER_110_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_894 ();
 DECAPx10_ASAP7_75t_R FILLER_110_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_936 ();
 DECAPx10_ASAP7_75t_R FILLER_110_951 ();
 FILLER_ASAP7_75t_R FILLER_110_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_975 ();
 FILLER_ASAP7_75t_R FILLER_110_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1004 ();
 FILLER_ASAP7_75t_R FILLER_110_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1042 ();
 FILLER_ASAP7_75t_R FILLER_110_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1216 ();
 FILLER_ASAP7_75t_R FILLER_110_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1243 ();
 FILLER_ASAP7_75t_R FILLER_110_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1249 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1253 ();
 FILLER_ASAP7_75t_R FILLER_110_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1269 ();
 FILLER_ASAP7_75t_R FILLER_110_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1277 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1352 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1374 ();
 FILLER_ASAP7_75t_R FILLER_110_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1388 ();
 FILLER_ASAP7_75t_R FILLER_110_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1404 ();
 DECAPx1_ASAP7_75t_R FILLER_111_28 ();
 DECAPx1_ASAP7_75t_R FILLER_111_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_39 ();
 DECAPx1_ASAP7_75t_R FILLER_111_46 ();
 DECAPx1_ASAP7_75t_R FILLER_111_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_70 ();
 FILLER_ASAP7_75t_R FILLER_111_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_141 ();
 FILLER_ASAP7_75t_R FILLER_111_151 ();
 DECAPx2_ASAP7_75t_R FILLER_111_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_185 ();
 FILLER_ASAP7_75t_R FILLER_111_200 ();
 DECAPx2_ASAP7_75t_R FILLER_111_218 ();
 FILLER_ASAP7_75t_R FILLER_111_224 ();
 DECAPx1_ASAP7_75t_R FILLER_111_234 ();
 FILLER_ASAP7_75t_R FILLER_111_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_254 ();
 DECAPx6_ASAP7_75t_R FILLER_111_275 ();
 DECAPx2_ASAP7_75t_R FILLER_111_289 ();
 DECAPx10_ASAP7_75t_R FILLER_111_313 ();
 DECAPx10_ASAP7_75t_R FILLER_111_335 ();
 DECAPx6_ASAP7_75t_R FILLER_111_357 ();
 FILLER_ASAP7_75t_R FILLER_111_371 ();
 DECAPx4_ASAP7_75t_R FILLER_111_395 ();
 DECAPx4_ASAP7_75t_R FILLER_111_413 ();
 DECAPx2_ASAP7_75t_R FILLER_111_431 ();
 FILLER_ASAP7_75t_R FILLER_111_437 ();
 DECAPx10_ASAP7_75t_R FILLER_111_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_469 ();
 FILLER_ASAP7_75t_R FILLER_111_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_495 ();
 FILLER_ASAP7_75t_R FILLER_111_526 ();
 DECAPx2_ASAP7_75t_R FILLER_111_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_540 ();
 DECAPx1_ASAP7_75t_R FILLER_111_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_563 ();
 DECAPx1_ASAP7_75t_R FILLER_111_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_575 ();
 DECAPx4_ASAP7_75t_R FILLER_111_646 ();
 DECAPx1_ASAP7_75t_R FILLER_111_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_666 ();
 DECAPx1_ASAP7_75t_R FILLER_111_679 ();
 DECAPx1_ASAP7_75t_R FILLER_111_686 ();
 DECAPx10_ASAP7_75t_R FILLER_111_738 ();
 DECAPx2_ASAP7_75t_R FILLER_111_760 ();
 FILLER_ASAP7_75t_R FILLER_111_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_768 ();
 FILLER_ASAP7_75t_R FILLER_111_775 ();
 DECAPx6_ASAP7_75t_R FILLER_111_783 ();
 FILLER_ASAP7_75t_R FILLER_111_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_799 ();
 DECAPx10_ASAP7_75t_R FILLER_111_816 ();
 DECAPx10_ASAP7_75t_R FILLER_111_838 ();
 FILLER_ASAP7_75t_R FILLER_111_860 ();
 DECAPx6_ASAP7_75t_R FILLER_111_870 ();
 DECAPx1_ASAP7_75t_R FILLER_111_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_926 ();
 FILLER_ASAP7_75t_R FILLER_111_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_941 ();
 DECAPx6_ASAP7_75t_R FILLER_111_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_975 ();
 DECAPx10_ASAP7_75t_R FILLER_111_983 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1061 ();
 FILLER_ASAP7_75t_R FILLER_111_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1088 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1171 ();
 FILLER_ASAP7_75t_R FILLER_111_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1179 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1250 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1260 ();
 FILLER_ASAP7_75t_R FILLER_111_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1295 ();
 FILLER_ASAP7_75t_R FILLER_111_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1351 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1373 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1395 ();
 DECAPx1_ASAP7_75t_R FILLER_112_2 ();
 FILLER_ASAP7_75t_R FILLER_112_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_89 ();
 FILLER_ASAP7_75t_R FILLER_112_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_95 ();
 FILLER_ASAP7_75t_R FILLER_112_128 ();
 DECAPx1_ASAP7_75t_R FILLER_112_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_176 ();
 DECAPx1_ASAP7_75t_R FILLER_112_184 ();
 FILLER_ASAP7_75t_R FILLER_112_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_196 ();
 DECAPx4_ASAP7_75t_R FILLER_112_203 ();
 FILLER_ASAP7_75t_R FILLER_112_213 ();
 DECAPx6_ASAP7_75t_R FILLER_112_221 ();
 FILLER_ASAP7_75t_R FILLER_112_235 ();
 FILLER_ASAP7_75t_R FILLER_112_243 ();
 DECAPx10_ASAP7_75t_R FILLER_112_263 ();
 DECAPx4_ASAP7_75t_R FILLER_112_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_295 ();
 DECAPx2_ASAP7_75t_R FILLER_112_306 ();
 FILLER_ASAP7_75t_R FILLER_112_312 ();
 DECAPx4_ASAP7_75t_R FILLER_112_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_332 ();
 DECAPx6_ASAP7_75t_R FILLER_112_339 ();
 DECAPx2_ASAP7_75t_R FILLER_112_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_359 ();
 DECAPx2_ASAP7_75t_R FILLER_112_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_372 ();
 DECAPx1_ASAP7_75t_R FILLER_112_417 ();
 DECAPx1_ASAP7_75t_R FILLER_112_441 ();
 FILLER_ASAP7_75t_R FILLER_112_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_461 ();
 DECAPx6_ASAP7_75t_R FILLER_112_464 ();
 DECAPx2_ASAP7_75t_R FILLER_112_478 ();
 FILLER_ASAP7_75t_R FILLER_112_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_492 ();
 DECAPx4_ASAP7_75t_R FILLER_112_499 ();
 FILLER_ASAP7_75t_R FILLER_112_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_511 ();
 FILLER_ASAP7_75t_R FILLER_112_518 ();
 FILLER_ASAP7_75t_R FILLER_112_532 ();
 DECAPx10_ASAP7_75t_R FILLER_112_540 ();
 FILLER_ASAP7_75t_R FILLER_112_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_564 ();
 DECAPx2_ASAP7_75t_R FILLER_112_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_600 ();
 FILLER_ASAP7_75t_R FILLER_112_604 ();
 FILLER_ASAP7_75t_R FILLER_112_638 ();
 DECAPx2_ASAP7_75t_R FILLER_112_695 ();
 FILLER_ASAP7_75t_R FILLER_112_701 ();
 DECAPx2_ASAP7_75t_R FILLER_112_715 ();
 FILLER_ASAP7_75t_R FILLER_112_721 ();
 DECAPx2_ASAP7_75t_R FILLER_112_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_735 ();
 DECAPx6_ASAP7_75t_R FILLER_112_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_759 ();
 DECAPx1_ASAP7_75t_R FILLER_112_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_783 ();
 DECAPx1_ASAP7_75t_R FILLER_112_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_795 ();
 DECAPx10_ASAP7_75t_R FILLER_112_804 ();
 DECAPx1_ASAP7_75t_R FILLER_112_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_850 ();
 DECAPx4_ASAP7_75t_R FILLER_112_859 ();
 DECAPx6_ASAP7_75t_R FILLER_112_881 ();
 FILLER_ASAP7_75t_R FILLER_112_895 ();
 DECAPx6_ASAP7_75t_R FILLER_112_929 ();
 DECAPx2_ASAP7_75t_R FILLER_112_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_949 ();
 DECAPx1_ASAP7_75t_R FILLER_112_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_974 ();
 DECAPx1_ASAP7_75t_R FILLER_112_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_986 ();
 DECAPx2_ASAP7_75t_R FILLER_112_996 ();
 FILLER_ASAP7_75t_R FILLER_112_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_112_1021 ();
 FILLER_ASAP7_75t_R FILLER_112_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1042 ();
 FILLER_ASAP7_75t_R FILLER_112_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1161 ();
 FILLER_ASAP7_75t_R FILLER_112_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1388 ();
 FILLER_ASAP7_75t_R FILLER_112_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1404 ();
 DECAPx1_ASAP7_75t_R FILLER_113_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_11 ();
 DECAPx1_ASAP7_75t_R FILLER_113_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_25 ();
 FILLER_ASAP7_75t_R FILLER_113_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_41 ();
 DECAPx4_ASAP7_75t_R FILLER_113_48 ();
 FILLER_ASAP7_75t_R FILLER_113_58 ();
 DECAPx2_ASAP7_75t_R FILLER_113_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_72 ();
 DECAPx6_ASAP7_75t_R FILLER_113_76 ();
 FILLER_ASAP7_75t_R FILLER_113_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_115 ();
 FILLER_ASAP7_75t_R FILLER_113_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_121 ();
 DECAPx4_ASAP7_75t_R FILLER_113_125 ();
 FILLER_ASAP7_75t_R FILLER_113_135 ();
 DECAPx6_ASAP7_75t_R FILLER_113_147 ();
 DECAPx1_ASAP7_75t_R FILLER_113_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_165 ();
 DECAPx6_ASAP7_75t_R FILLER_113_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_208 ();
 DECAPx6_ASAP7_75t_R FILLER_113_225 ();
 DECAPx10_ASAP7_75t_R FILLER_113_247 ();
 DECAPx4_ASAP7_75t_R FILLER_113_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_279 ();
 DECAPx6_ASAP7_75t_R FILLER_113_292 ();
 DECAPx2_ASAP7_75t_R FILLER_113_306 ();
 DECAPx1_ASAP7_75t_R FILLER_113_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_322 ();
 DECAPx2_ASAP7_75t_R FILLER_113_337 ();
 FILLER_ASAP7_75t_R FILLER_113_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_345 ();
 DECAPx2_ASAP7_75t_R FILLER_113_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_374 ();
 DECAPx10_ASAP7_75t_R FILLER_113_396 ();
 DECAPx2_ASAP7_75t_R FILLER_113_418 ();
 DECAPx10_ASAP7_75t_R FILLER_113_432 ();
 DECAPx10_ASAP7_75t_R FILLER_113_454 ();
 DECAPx10_ASAP7_75t_R FILLER_113_476 ();
 DECAPx10_ASAP7_75t_R FILLER_113_498 ();
 DECAPx4_ASAP7_75t_R FILLER_113_520 ();
 DECAPx4_ASAP7_75t_R FILLER_113_552 ();
 FILLER_ASAP7_75t_R FILLER_113_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_564 ();
 DECAPx2_ASAP7_75t_R FILLER_113_571 ();
 FILLER_ASAP7_75t_R FILLER_113_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_579 ();
 DECAPx10_ASAP7_75t_R FILLER_113_583 ();
 DECAPx6_ASAP7_75t_R FILLER_113_605 ();
 DECAPx2_ASAP7_75t_R FILLER_113_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_625 ();
 DECAPx4_ASAP7_75t_R FILLER_113_629 ();
 FILLER_ASAP7_75t_R FILLER_113_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_641 ();
 DECAPx6_ASAP7_75t_R FILLER_113_680 ();
 DECAPx2_ASAP7_75t_R FILLER_113_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_700 ();
 DECAPx10_ASAP7_75t_R FILLER_113_727 ();
 DECAPx6_ASAP7_75t_R FILLER_113_749 ();
 DECAPx2_ASAP7_75t_R FILLER_113_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_775 ();
 DECAPx1_ASAP7_75t_R FILLER_113_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_832 ();
 FILLER_ASAP7_75t_R FILLER_113_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_867 ();
 DECAPx2_ASAP7_75t_R FILLER_113_900 ();
 DECAPx2_ASAP7_75t_R FILLER_113_918 ();
 DECAPx4_ASAP7_75t_R FILLER_113_926 ();
 FILLER_ASAP7_75t_R FILLER_113_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_938 ();
 DECAPx2_ASAP7_75t_R FILLER_113_969 ();
 FILLER_ASAP7_75t_R FILLER_113_975 ();
 DECAPx6_ASAP7_75t_R FILLER_113_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_998 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1057 ();
 FILLER_ASAP7_75t_R FILLER_113_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1109 ();
 FILLER_ASAP7_75t_R FILLER_113_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1202 ();
 FILLER_ASAP7_75t_R FILLER_113_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1214 ();
 FILLER_ASAP7_75t_R FILLER_113_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1272 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1291 ();
 FILLER_ASAP7_75t_R FILLER_113_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1316 ();
 FILLER_ASAP7_75t_R FILLER_113_1322 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1327 ();
 FILLER_ASAP7_75t_R FILLER_113_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1365 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1387 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1401 ();
 DECAPx10_ASAP7_75t_R FILLER_114_7 ();
 FILLER_ASAP7_75t_R FILLER_114_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_31 ();
 DECAPx6_ASAP7_75t_R FILLER_114_58 ();
 DECAPx1_ASAP7_75t_R FILLER_114_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_76 ();
 FILLER_ASAP7_75t_R FILLER_114_83 ();
 DECAPx10_ASAP7_75t_R FILLER_114_88 ();
 DECAPx10_ASAP7_75t_R FILLER_114_110 ();
 DECAPx10_ASAP7_75t_R FILLER_114_132 ();
 DECAPx10_ASAP7_75t_R FILLER_114_154 ();
 DECAPx1_ASAP7_75t_R FILLER_114_176 ();
 FILLER_ASAP7_75t_R FILLER_114_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_189 ();
 DECAPx2_ASAP7_75t_R FILLER_114_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_202 ();
 DECAPx2_ASAP7_75t_R FILLER_114_209 ();
 FILLER_ASAP7_75t_R FILLER_114_215 ();
 DECAPx6_ASAP7_75t_R FILLER_114_231 ();
 DECAPx1_ASAP7_75t_R FILLER_114_245 ();
 FILLER_ASAP7_75t_R FILLER_114_255 ();
 DECAPx2_ASAP7_75t_R FILLER_114_263 ();
 DECAPx6_ASAP7_75t_R FILLER_114_277 ();
 FILLER_ASAP7_75t_R FILLER_114_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_293 ();
 DECAPx10_ASAP7_75t_R FILLER_114_304 ();
 DECAPx6_ASAP7_75t_R FILLER_114_326 ();
 DECAPx2_ASAP7_75t_R FILLER_114_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_346 ();
 DECAPx10_ASAP7_75t_R FILLER_114_353 ();
 DECAPx2_ASAP7_75t_R FILLER_114_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_381 ();
 DECAPx2_ASAP7_75t_R FILLER_114_394 ();
 DECAPx6_ASAP7_75t_R FILLER_114_414 ();
 DECAPx1_ASAP7_75t_R FILLER_114_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_432 ();
 DECAPx2_ASAP7_75t_R FILLER_114_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_448 ();
 DECAPx2_ASAP7_75t_R FILLER_114_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_461 ();
 FILLER_ASAP7_75t_R FILLER_114_464 ();
 DECAPx10_ASAP7_75t_R FILLER_114_472 ();
 DECAPx6_ASAP7_75t_R FILLER_114_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_508 ();
 DECAPx6_ASAP7_75t_R FILLER_114_517 ();
 DECAPx2_ASAP7_75t_R FILLER_114_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_537 ();
 FILLER_ASAP7_75t_R FILLER_114_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_558 ();
 DECAPx10_ASAP7_75t_R FILLER_114_566 ();
 DECAPx2_ASAP7_75t_R FILLER_114_588 ();
 FILLER_ASAP7_75t_R FILLER_114_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_596 ();
 DECAPx2_ASAP7_75t_R FILLER_114_609 ();
 FILLER_ASAP7_75t_R FILLER_114_615 ();
 DECAPx10_ASAP7_75t_R FILLER_114_627 ();
 DECAPx1_ASAP7_75t_R FILLER_114_649 ();
 DECAPx2_ASAP7_75t_R FILLER_114_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_668 ();
 DECAPx10_ASAP7_75t_R FILLER_114_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_694 ();
 DECAPx10_ASAP7_75t_R FILLER_114_735 ();
 DECAPx2_ASAP7_75t_R FILLER_114_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_763 ();
 DECAPx6_ASAP7_75t_R FILLER_114_780 ();
 DECAPx1_ASAP7_75t_R FILLER_114_794 ();
 DECAPx1_ASAP7_75t_R FILLER_114_818 ();
 DECAPx2_ASAP7_75t_R FILLER_114_838 ();
 FILLER_ASAP7_75t_R FILLER_114_860 ();
 DECAPx10_ASAP7_75t_R FILLER_114_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_900 ();
 DECAPx6_ASAP7_75t_R FILLER_114_908 ();
 DECAPx2_ASAP7_75t_R FILLER_114_930 ();
 FILLER_ASAP7_75t_R FILLER_114_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_974 ();
 DECAPx1_ASAP7_75t_R FILLER_114_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_986 ();
 DECAPx1_ASAP7_75t_R FILLER_114_996 ();
 FILLER_ASAP7_75t_R FILLER_114_1029 ();
 FILLER_ASAP7_75t_R FILLER_114_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1153 ();
 FILLER_ASAP7_75t_R FILLER_114_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1182 ();
 FILLER_ASAP7_75t_R FILLER_114_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1251 ();
 FILLER_ASAP7_75t_R FILLER_114_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1280 ();
 FILLER_ASAP7_75t_R FILLER_114_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1301 ();
 FILLER_ASAP7_75t_R FILLER_114_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1351 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1373 ();
 FILLER_ASAP7_75t_R FILLER_114_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1388 ();
 FILLER_ASAP7_75t_R FILLER_114_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_115_37 ();
 DECAPx2_ASAP7_75t_R FILLER_115_50 ();
 FILLER_ASAP7_75t_R FILLER_115_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_64 ();
 FILLER_ASAP7_75t_R FILLER_115_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_105 ();
 DECAPx1_ASAP7_75t_R FILLER_115_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_113 ();
 DECAPx1_ASAP7_75t_R FILLER_115_123 ();
 DECAPx4_ASAP7_75t_R FILLER_115_134 ();
 FILLER_ASAP7_75t_R FILLER_115_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_146 ();
 DECAPx2_ASAP7_75t_R FILLER_115_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_166 ();
 DECAPx1_ASAP7_75t_R FILLER_115_183 ();
 DECAPx4_ASAP7_75t_R FILLER_115_201 ();
 FILLER_ASAP7_75t_R FILLER_115_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_213 ();
 DECAPx4_ASAP7_75t_R FILLER_115_228 ();
 FILLER_ASAP7_75t_R FILLER_115_238 ();
 DECAPx10_ASAP7_75t_R FILLER_115_268 ();
 FILLER_ASAP7_75t_R FILLER_115_290 ();
 DECAPx10_ASAP7_75t_R FILLER_115_312 ();
 DECAPx10_ASAP7_75t_R FILLER_115_334 ();
 DECAPx6_ASAP7_75t_R FILLER_115_356 ();
 DECAPx1_ASAP7_75t_R FILLER_115_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_374 ();
 DECAPx4_ASAP7_75t_R FILLER_115_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_422 ();
 DECAPx10_ASAP7_75t_R FILLER_115_431 ();
 DECAPx10_ASAP7_75t_R FILLER_115_453 ();
 DECAPx2_ASAP7_75t_R FILLER_115_475 ();
 FILLER_ASAP7_75t_R FILLER_115_481 ();
 DECAPx4_ASAP7_75t_R FILLER_115_497 ();
 FILLER_ASAP7_75t_R FILLER_115_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_515 ();
 DECAPx10_ASAP7_75t_R FILLER_115_522 ();
 DECAPx1_ASAP7_75t_R FILLER_115_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_548 ();
 DECAPx2_ASAP7_75t_R FILLER_115_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_591 ();
 DECAPx1_ASAP7_75t_R FILLER_115_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_648 ();
 DECAPx6_ASAP7_75t_R FILLER_115_653 ();
 DECAPx1_ASAP7_75t_R FILLER_115_667 ();
 FILLER_ASAP7_75t_R FILLER_115_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_738 ();
 DECAPx10_ASAP7_75t_R FILLER_115_755 ();
 DECAPx4_ASAP7_75t_R FILLER_115_777 ();
 FILLER_ASAP7_75t_R FILLER_115_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_789 ();
 DECAPx6_ASAP7_75t_R FILLER_115_818 ();
 DECAPx2_ASAP7_75t_R FILLER_115_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_838 ();
 DECAPx10_ASAP7_75t_R FILLER_115_847 ();
 DECAPx10_ASAP7_75t_R FILLER_115_869 ();
 DECAPx2_ASAP7_75t_R FILLER_115_891 ();
 FILLER_ASAP7_75t_R FILLER_115_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_899 ();
 FILLER_ASAP7_75t_R FILLER_115_922 ();
 DECAPx1_ASAP7_75t_R FILLER_115_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_942 ();
 DECAPx6_ASAP7_75t_R FILLER_115_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_986 ();
 DECAPx6_ASAP7_75t_R FILLER_115_996 ();
 FILLER_ASAP7_75t_R FILLER_115_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1040 ();
 FILLER_ASAP7_75t_R FILLER_115_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1065 ();
 FILLER_ASAP7_75t_R FILLER_115_1075 ();
 FILLER_ASAP7_75t_R FILLER_115_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1112 ();
 FILLER_ASAP7_75t_R FILLER_115_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1145 ();
 FILLER_ASAP7_75t_R FILLER_115_1151 ();
 FILLER_ASAP7_75t_R FILLER_115_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1185 ();
 FILLER_ASAP7_75t_R FILLER_115_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1205 ();
 FILLER_ASAP7_75t_R FILLER_115_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1284 ();
 FILLER_ASAP7_75t_R FILLER_115_1290 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1315 ();
 FILLER_ASAP7_75t_R FILLER_115_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1404 ();
 FILLER_ASAP7_75t_R FILLER_116_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_4 ();
 DECAPx1_ASAP7_75t_R FILLER_116_37 ();
 FILLER_ASAP7_75t_R FILLER_116_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_49 ();
 DECAPx2_ASAP7_75t_R FILLER_116_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_117 ();
 DECAPx1_ASAP7_75t_R FILLER_116_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_174 ();
 DECAPx6_ASAP7_75t_R FILLER_116_195 ();
 DECAPx1_ASAP7_75t_R FILLER_116_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_213 ();
 DECAPx2_ASAP7_75t_R FILLER_116_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_232 ();
 FILLER_ASAP7_75t_R FILLER_116_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_257 ();
 FILLER_ASAP7_75t_R FILLER_116_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_266 ();
 DECAPx10_ASAP7_75t_R FILLER_116_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_295 ();
 DECAPx1_ASAP7_75t_R FILLER_116_306 ();
 DECAPx2_ASAP7_75t_R FILLER_116_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_322 ();
 DECAPx10_ASAP7_75t_R FILLER_116_329 ();
 DECAPx1_ASAP7_75t_R FILLER_116_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_355 ();
 DECAPx10_ASAP7_75t_R FILLER_116_362 ();
 DECAPx6_ASAP7_75t_R FILLER_116_384 ();
 DECAPx1_ASAP7_75t_R FILLER_116_398 ();
 FILLER_ASAP7_75t_R FILLER_116_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_410 ();
 DECAPx2_ASAP7_75t_R FILLER_116_417 ();
 FILLER_ASAP7_75t_R FILLER_116_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_425 ();
 DECAPx4_ASAP7_75t_R FILLER_116_450 ();
 FILLER_ASAP7_75t_R FILLER_116_460 ();
 DECAPx6_ASAP7_75t_R FILLER_116_464 ();
 FILLER_ASAP7_75t_R FILLER_116_478 ();
 DECAPx1_ASAP7_75t_R FILLER_116_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_498 ();
 DECAPx1_ASAP7_75t_R FILLER_116_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_520 ();
 DECAPx10_ASAP7_75t_R FILLER_116_535 ();
 FILLER_ASAP7_75t_R FILLER_116_557 ();
 FILLER_ASAP7_75t_R FILLER_116_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_567 ();
 FILLER_ASAP7_75t_R FILLER_116_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_609 ();
 DECAPx1_ASAP7_75t_R FILLER_116_613 ();
 FILLER_ASAP7_75t_R FILLER_116_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_695 ();
 DECAPx1_ASAP7_75t_R FILLER_116_740 ();
 DECAPx6_ASAP7_75t_R FILLER_116_760 ();
 DECAPx1_ASAP7_75t_R FILLER_116_774 ();
 DECAPx1_ASAP7_75t_R FILLER_116_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_805 ();
 DECAPx2_ASAP7_75t_R FILLER_116_821 ();
 FILLER_ASAP7_75t_R FILLER_116_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_829 ();
 DECAPx2_ASAP7_75t_R FILLER_116_842 ();
 FILLER_ASAP7_75t_R FILLER_116_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_850 ();
 DECAPx10_ASAP7_75t_R FILLER_116_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_882 ();
 DECAPx2_ASAP7_75t_R FILLER_116_903 ();
 FILLER_ASAP7_75t_R FILLER_116_909 ();
 DECAPx2_ASAP7_75t_R FILLER_116_926 ();
 FILLER_ASAP7_75t_R FILLER_116_932 ();
 DECAPx4_ASAP7_75t_R FILLER_116_946 ();
 DECAPx10_ASAP7_75t_R FILLER_116_975 ();
 DECAPx1_ASAP7_75t_R FILLER_116_997 ();
 FILLER_ASAP7_75t_R FILLER_116_1018 ();
 FILLER_ASAP7_75t_R FILLER_116_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1061 ();
 FILLER_ASAP7_75t_R FILLER_116_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1083 ();
 FILLER_ASAP7_75t_R FILLER_116_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1187 ();
 FILLER_ASAP7_75t_R FILLER_116_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1236 ();
 FILLER_ASAP7_75t_R FILLER_116_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1303 ();
 FILLER_ASAP7_75t_R FILLER_116_1309 ();
 FILLER_ASAP7_75t_R FILLER_116_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1353 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1388 ();
 FILLER_ASAP7_75t_R FILLER_116_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1404 ();
 FILLER_ASAP7_75t_R FILLER_117_2 ();
 DECAPx4_ASAP7_75t_R FILLER_117_25 ();
 FILLER_ASAP7_75t_R FILLER_117_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_72 ();
 DECAPx6_ASAP7_75t_R FILLER_117_77 ();
 DECAPx1_ASAP7_75t_R FILLER_117_91 ();
 DECAPx4_ASAP7_75t_R FILLER_117_121 ();
 FILLER_ASAP7_75t_R FILLER_117_131 ();
 DECAPx6_ASAP7_75t_R FILLER_117_142 ();
 FILLER_ASAP7_75t_R FILLER_117_156 ();
 DECAPx2_ASAP7_75t_R FILLER_117_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_174 ();
 DECAPx6_ASAP7_75t_R FILLER_117_181 ();
 DECAPx2_ASAP7_75t_R FILLER_117_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_201 ();
 DECAPx1_ASAP7_75t_R FILLER_117_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_212 ();
 DECAPx10_ASAP7_75t_R FILLER_117_225 ();
 DECAPx10_ASAP7_75t_R FILLER_117_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_269 ();
 DECAPx6_ASAP7_75t_R FILLER_117_278 ();
 FILLER_ASAP7_75t_R FILLER_117_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_294 ();
 DECAPx2_ASAP7_75t_R FILLER_117_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_311 ();
 DECAPx2_ASAP7_75t_R FILLER_117_320 ();
 DECAPx2_ASAP7_75t_R FILLER_117_340 ();
 FILLER_ASAP7_75t_R FILLER_117_368 ();
 FILLER_ASAP7_75t_R FILLER_117_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_379 ();
 DECAPx1_ASAP7_75t_R FILLER_117_386 ();
 DECAPx4_ASAP7_75t_R FILLER_117_424 ();
 FILLER_ASAP7_75t_R FILLER_117_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_436 ();
 FILLER_ASAP7_75t_R FILLER_117_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_448 ();
 DECAPx2_ASAP7_75t_R FILLER_117_455 ();
 FILLER_ASAP7_75t_R FILLER_117_461 ();
 DECAPx10_ASAP7_75t_R FILLER_117_471 ();
 DECAPx6_ASAP7_75t_R FILLER_117_493 ();
 DECAPx2_ASAP7_75t_R FILLER_117_507 ();
 DECAPx6_ASAP7_75t_R FILLER_117_519 ();
 FILLER_ASAP7_75t_R FILLER_117_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_535 ();
 DECAPx4_ASAP7_75t_R FILLER_117_546 ();
 FILLER_ASAP7_75t_R FILLER_117_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_558 ();
 DECAPx2_ASAP7_75t_R FILLER_117_569 ();
 FILLER_ASAP7_75t_R FILLER_117_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_577 ();
 DECAPx2_ASAP7_75t_R FILLER_117_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_590 ();
 DECAPx10_ASAP7_75t_R FILLER_117_594 ();
 DECAPx4_ASAP7_75t_R FILLER_117_616 ();
 FILLER_ASAP7_75t_R FILLER_117_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_628 ();
 DECAPx2_ASAP7_75t_R FILLER_117_638 ();
 DECAPx2_ASAP7_75t_R FILLER_117_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_653 ();
 DECAPx2_ASAP7_75t_R FILLER_117_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_666 ();
 DECAPx1_ASAP7_75t_R FILLER_117_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_683 ();
 DECAPx2_ASAP7_75t_R FILLER_117_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_699 ();
 FILLER_ASAP7_75t_R FILLER_117_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_708 ();
 DECAPx2_ASAP7_75t_R FILLER_117_715 ();
 DECAPx1_ASAP7_75t_R FILLER_117_724 ();
 DECAPx6_ASAP7_75t_R FILLER_117_732 ();
 FILLER_ASAP7_75t_R FILLER_117_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_770 ();
 DECAPx1_ASAP7_75t_R FILLER_117_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_785 ();
 DECAPx2_ASAP7_75t_R FILLER_117_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_804 ();
 DECAPx1_ASAP7_75t_R FILLER_117_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_826 ();
 FILLER_ASAP7_75t_R FILLER_117_864 ();
 DECAPx2_ASAP7_75t_R FILLER_117_890 ();
 FILLER_ASAP7_75t_R FILLER_117_896 ();
 DECAPx1_ASAP7_75t_R FILLER_117_907 ();
 DECAPx1_ASAP7_75t_R FILLER_117_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_920 ();
 DECAPx4_ASAP7_75t_R FILLER_117_926 ();
 FILLER_ASAP7_75t_R FILLER_117_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_947 ();
 DECAPx4_ASAP7_75t_R FILLER_117_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_978 ();
 FILLER_ASAP7_75t_R FILLER_117_996 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1006 ();
 FILLER_ASAP7_75t_R FILLER_117_1028 ();
 FILLER_ASAP7_75t_R FILLER_117_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1071 ();
 FILLER_ASAP7_75t_R FILLER_117_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1079 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1122 ();
 FILLER_ASAP7_75t_R FILLER_117_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1221 ();
 FILLER_ASAP7_75t_R FILLER_117_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1242 ();
 FILLER_ASAP7_75t_R FILLER_117_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1354 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1398 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_118_7 ();
 DECAPx2_ASAP7_75t_R FILLER_118_29 ();
 FILLER_ASAP7_75t_R FILLER_118_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_37 ();
 DECAPx2_ASAP7_75t_R FILLER_118_44 ();
 DECAPx4_ASAP7_75t_R FILLER_118_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_70 ();
 DECAPx6_ASAP7_75t_R FILLER_118_77 ();
 DECAPx1_ASAP7_75t_R FILLER_118_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_95 ();
 FILLER_ASAP7_75t_R FILLER_118_108 ();
 DECAPx10_ASAP7_75t_R FILLER_118_113 ();
 DECAPx10_ASAP7_75t_R FILLER_118_135 ();
 DECAPx4_ASAP7_75t_R FILLER_118_157 ();
 FILLER_ASAP7_75t_R FILLER_118_179 ();
 DECAPx6_ASAP7_75t_R FILLER_118_187 ();
 DECAPx4_ASAP7_75t_R FILLER_118_223 ();
 DECAPx10_ASAP7_75t_R FILLER_118_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_269 ();
 DECAPx6_ASAP7_75t_R FILLER_118_276 ();
 FILLER_ASAP7_75t_R FILLER_118_290 ();
 DECAPx10_ASAP7_75t_R FILLER_118_302 ();
 DECAPx2_ASAP7_75t_R FILLER_118_324 ();
 FILLER_ASAP7_75t_R FILLER_118_330 ();
 DECAPx4_ASAP7_75t_R FILLER_118_341 ();
 DECAPx4_ASAP7_75t_R FILLER_118_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_393 ();
 FILLER_ASAP7_75t_R FILLER_118_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_403 ();
 DECAPx10_ASAP7_75t_R FILLER_118_407 ();
 DECAPx4_ASAP7_75t_R FILLER_118_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_439 ();
 DECAPx6_ASAP7_75t_R FILLER_118_446 ();
 FILLER_ASAP7_75t_R FILLER_118_460 ();
 DECAPx1_ASAP7_75t_R FILLER_118_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_482 ();
 DECAPx4_ASAP7_75t_R FILLER_118_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_499 ();
 DECAPx10_ASAP7_75t_R FILLER_118_508 ();
 DECAPx2_ASAP7_75t_R FILLER_118_530 ();
 DECAPx10_ASAP7_75t_R FILLER_118_548 ();
 FILLER_ASAP7_75t_R FILLER_118_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_572 ();
 DECAPx10_ASAP7_75t_R FILLER_118_579 ();
 FILLER_ASAP7_75t_R FILLER_118_601 ();
 FILLER_ASAP7_75t_R FILLER_118_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_617 ();
 DECAPx1_ASAP7_75t_R FILLER_118_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_628 ();
 FILLER_ASAP7_75t_R FILLER_118_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_643 ();
 DECAPx10_ASAP7_75t_R FILLER_118_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_704 ();
 DECAPx10_ASAP7_75t_R FILLER_118_711 ();
 DECAPx4_ASAP7_75t_R FILLER_118_733 ();
 FILLER_ASAP7_75t_R FILLER_118_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_769 ();
 FILLER_ASAP7_75t_R FILLER_118_828 ();
 FILLER_ASAP7_75t_R FILLER_118_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_852 ();
 DECAPx1_ASAP7_75t_R FILLER_118_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_873 ();
 DECAPx2_ASAP7_75t_R FILLER_118_890 ();
 FILLER_ASAP7_75t_R FILLER_118_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_898 ();
 FILLER_ASAP7_75t_R FILLER_118_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_932 ();
 DECAPx4_ASAP7_75t_R FILLER_118_957 ();
 FILLER_ASAP7_75t_R FILLER_118_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_969 ();
 DECAPx2_ASAP7_75t_R FILLER_118_976 ();
 FILLER_ASAP7_75t_R FILLER_118_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1063 ();
 FILLER_ASAP7_75t_R FILLER_118_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1087 ();
 FILLER_ASAP7_75t_R FILLER_118_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1150 ();
 FILLER_ASAP7_75t_R FILLER_118_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1217 ();
 FILLER_ASAP7_75t_R FILLER_118_1223 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1259 ();
 FILLER_ASAP7_75t_R FILLER_118_1269 ();
 FILLER_ASAP7_75t_R FILLER_118_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1290 ();
 FILLER_ASAP7_75t_R FILLER_118_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1312 ();
 FILLER_ASAP7_75t_R FILLER_118_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1388 ();
 FILLER_ASAP7_75t_R FILLER_118_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_119_2 ();
 FILLER_ASAP7_75t_R FILLER_119_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_10 ();
 FILLER_ASAP7_75t_R FILLER_119_17 ();
 DECAPx2_ASAP7_75t_R FILLER_119_33 ();
 FILLER_ASAP7_75t_R FILLER_119_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_50 ();
 DECAPx1_ASAP7_75t_R FILLER_119_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_90 ();
 DECAPx4_ASAP7_75t_R FILLER_119_103 ();
 FILLER_ASAP7_75t_R FILLER_119_113 ();
 DECAPx2_ASAP7_75t_R FILLER_119_118 ();
 FILLER_ASAP7_75t_R FILLER_119_124 ();
 DECAPx2_ASAP7_75t_R FILLER_119_161 ();
 DECAPx1_ASAP7_75t_R FILLER_119_175 ();
 DECAPx2_ASAP7_75t_R FILLER_119_195 ();
 FILLER_ASAP7_75t_R FILLER_119_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_203 ();
 DECAPx2_ASAP7_75t_R FILLER_119_226 ();
 FILLER_ASAP7_75t_R FILLER_119_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_240 ();
 DECAPx1_ASAP7_75t_R FILLER_119_249 ();
 DECAPx10_ASAP7_75t_R FILLER_119_265 ();
 DECAPx2_ASAP7_75t_R FILLER_119_287 ();
 DECAPx10_ASAP7_75t_R FILLER_119_303 ();
 FILLER_ASAP7_75t_R FILLER_119_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_327 ();
 DECAPx2_ASAP7_75t_R FILLER_119_336 ();
 FILLER_ASAP7_75t_R FILLER_119_342 ();
 DECAPx10_ASAP7_75t_R FILLER_119_350 ();
 DECAPx2_ASAP7_75t_R FILLER_119_372 ();
 FILLER_ASAP7_75t_R FILLER_119_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_380 ();
 DECAPx2_ASAP7_75t_R FILLER_119_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_390 ();
 DECAPx6_ASAP7_75t_R FILLER_119_398 ();
 DECAPx2_ASAP7_75t_R FILLER_119_412 ();
 DECAPx6_ASAP7_75t_R FILLER_119_424 ();
 DECAPx2_ASAP7_75t_R FILLER_119_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_444 ();
 DECAPx6_ASAP7_75t_R FILLER_119_451 ();
 DECAPx4_ASAP7_75t_R FILLER_119_471 ();
 DECAPx6_ASAP7_75t_R FILLER_119_509 ();
 DECAPx2_ASAP7_75t_R FILLER_119_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_529 ();
 DECAPx2_ASAP7_75t_R FILLER_119_552 ();
 FILLER_ASAP7_75t_R FILLER_119_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_570 ();
 FILLER_ASAP7_75t_R FILLER_119_597 ();
 DECAPx1_ASAP7_75t_R FILLER_119_625 ();
 DECAPx1_ASAP7_75t_R FILLER_119_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_663 ();
 DECAPx2_ASAP7_75t_R FILLER_119_673 ();
 FILLER_ASAP7_75t_R FILLER_119_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_681 ();
 FILLER_ASAP7_75t_R FILLER_119_685 ();
 FILLER_ASAP7_75t_R FILLER_119_725 ();
 DECAPx2_ASAP7_75t_R FILLER_119_731 ();
 FILLER_ASAP7_75t_R FILLER_119_737 ();
 DECAPx6_ASAP7_75t_R FILLER_119_748 ();
 DECAPx1_ASAP7_75t_R FILLER_119_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_766 ();
 DECAPx4_ASAP7_75t_R FILLER_119_773 ();
 FILLER_ASAP7_75t_R FILLER_119_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_785 ();
 DECAPx6_ASAP7_75t_R FILLER_119_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_842 ();
 DECAPx4_ASAP7_75t_R FILLER_119_852 ();
 FILLER_ASAP7_75t_R FILLER_119_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_864 ();
 DECAPx2_ASAP7_75t_R FILLER_119_871 ();
 FILLER_ASAP7_75t_R FILLER_119_877 ();
 DECAPx1_ASAP7_75t_R FILLER_119_885 ();
 DECAPx4_ASAP7_75t_R FILLER_119_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_923 ();
 DECAPx6_ASAP7_75t_R FILLER_119_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_940 ();
 DECAPx4_ASAP7_75t_R FILLER_119_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_961 ();
 DECAPx2_ASAP7_75t_R FILLER_119_974 ();
 FILLER_ASAP7_75t_R FILLER_119_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_982 ();
 DECAPx4_ASAP7_75t_R FILLER_119_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1042 ();
 FILLER_ASAP7_75t_R FILLER_119_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1067 ();
 FILLER_ASAP7_75t_R FILLER_119_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1121 ();
 FILLER_ASAP7_75t_R FILLER_119_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1148 ();
 FILLER_ASAP7_75t_R FILLER_119_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1181 ();
 FILLER_ASAP7_75t_R FILLER_119_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1227 ();
 FILLER_ASAP7_75t_R FILLER_119_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1297 ();
 FILLER_ASAP7_75t_R FILLER_119_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1319 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1339 ();
 FILLER_ASAP7_75t_R FILLER_119_1369 ();
 FILLER_ASAP7_75t_R FILLER_119_1374 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1399 ();
 FILLER_ASAP7_75t_R FILLER_120_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_4 ();
 FILLER_ASAP7_75t_R FILLER_120_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_143 ();
 DECAPx2_ASAP7_75t_R FILLER_120_170 ();
 FILLER_ASAP7_75t_R FILLER_120_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_187 ();
 DECAPx6_ASAP7_75t_R FILLER_120_194 ();
 FILLER_ASAP7_75t_R FILLER_120_208 ();
 DECAPx2_ASAP7_75t_R FILLER_120_216 ();
 FILLER_ASAP7_75t_R FILLER_120_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_224 ();
 DECAPx2_ASAP7_75t_R FILLER_120_259 ();
 DECAPx2_ASAP7_75t_R FILLER_120_279 ();
 DECAPx6_ASAP7_75t_R FILLER_120_291 ();
 DECAPx1_ASAP7_75t_R FILLER_120_305 ();
 DECAPx2_ASAP7_75t_R FILLER_120_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_321 ();
 DECAPx2_ASAP7_75t_R FILLER_120_330 ();
 FILLER_ASAP7_75t_R FILLER_120_336 ();
 DECAPx6_ASAP7_75t_R FILLER_120_354 ();
 FILLER_ASAP7_75t_R FILLER_120_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_370 ();
 DECAPx4_ASAP7_75t_R FILLER_120_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_387 ();
 FILLER_ASAP7_75t_R FILLER_120_414 ();
 DECAPx1_ASAP7_75t_R FILLER_120_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_426 ();
 DECAPx2_ASAP7_75t_R FILLER_120_435 ();
 FILLER_ASAP7_75t_R FILLER_120_441 ();
 DECAPx4_ASAP7_75t_R FILLER_120_449 ();
 FILLER_ASAP7_75t_R FILLER_120_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_461 ();
 DECAPx6_ASAP7_75t_R FILLER_120_464 ();
 FILLER_ASAP7_75t_R FILLER_120_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_480 ();
 FILLER_ASAP7_75t_R FILLER_120_495 ();
 DECAPx4_ASAP7_75t_R FILLER_120_503 ();
 DECAPx10_ASAP7_75t_R FILLER_120_523 ();
 DECAPx1_ASAP7_75t_R FILLER_120_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_613 ();
 DECAPx2_ASAP7_75t_R FILLER_120_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_626 ();
 FILLER_ASAP7_75t_R FILLER_120_704 ();
 DECAPx10_ASAP7_75t_R FILLER_120_732 ();
 DECAPx6_ASAP7_75t_R FILLER_120_754 ();
 DECAPx1_ASAP7_75t_R FILLER_120_768 ();
 FILLER_ASAP7_75t_R FILLER_120_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_784 ();
 FILLER_ASAP7_75t_R FILLER_120_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_808 ();
 DECAPx1_ASAP7_75t_R FILLER_120_817 ();
 FILLER_ASAP7_75t_R FILLER_120_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_833 ();
 DECAPx10_ASAP7_75t_R FILLER_120_856 ();
 FILLER_ASAP7_75t_R FILLER_120_878 ();
 DECAPx4_ASAP7_75t_R FILLER_120_888 ();
 DECAPx10_ASAP7_75t_R FILLER_120_931 ();
 DECAPx2_ASAP7_75t_R FILLER_120_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_959 ();
 DECAPx4_ASAP7_75t_R FILLER_120_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_973 ();
 DECAPx4_ASAP7_75t_R FILLER_120_997 ();
 FILLER_ASAP7_75t_R FILLER_120_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1079 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1120 ();
 FILLER_ASAP7_75t_R FILLER_120_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1165 ();
 FILLER_ASAP7_75t_R FILLER_120_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1188 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1273 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1286 ();
 FILLER_ASAP7_75t_R FILLER_120_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1302 ();
 FILLER_ASAP7_75t_R FILLER_120_1314 ();
 FILLER_ASAP7_75t_R FILLER_120_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1330 ();
 FILLER_ASAP7_75t_R FILLER_120_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1388 ();
 FILLER_ASAP7_75t_R FILLER_120_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_121_2 ();
 DECAPx2_ASAP7_75t_R FILLER_121_14 ();
 DECAPx1_ASAP7_75t_R FILLER_121_23 ();
 FILLER_ASAP7_75t_R FILLER_121_65 ();
 FILLER_ASAP7_75t_R FILLER_121_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_82 ();
 DECAPx2_ASAP7_75t_R FILLER_121_86 ();
 FILLER_ASAP7_75t_R FILLER_121_92 ();
 DECAPx1_ASAP7_75t_R FILLER_121_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_104 ();
 DECAPx1_ASAP7_75t_R FILLER_121_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_112 ();
 DECAPx2_ASAP7_75t_R FILLER_121_139 ();
 FILLER_ASAP7_75t_R FILLER_121_145 ();
 DECAPx10_ASAP7_75t_R FILLER_121_154 ();
 FILLER_ASAP7_75t_R FILLER_121_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_178 ();
 DECAPx6_ASAP7_75t_R FILLER_121_185 ();
 DECAPx1_ASAP7_75t_R FILLER_121_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_203 ();
 DECAPx1_ASAP7_75t_R FILLER_121_222 ();
 DECAPx1_ASAP7_75t_R FILLER_121_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_236 ();
 DECAPx4_ASAP7_75t_R FILLER_121_255 ();
 FILLER_ASAP7_75t_R FILLER_121_265 ();
 DECAPx1_ASAP7_75t_R FILLER_121_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_277 ();
 DECAPx6_ASAP7_75t_R FILLER_121_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_328 ();
 FILLER_ASAP7_75t_R FILLER_121_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_341 ();
 DECAPx6_ASAP7_75t_R FILLER_121_348 ();
 DECAPx2_ASAP7_75t_R FILLER_121_362 ();
 DECAPx6_ASAP7_75t_R FILLER_121_380 ();
 FILLER_ASAP7_75t_R FILLER_121_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_396 ();
 DECAPx2_ASAP7_75t_R FILLER_121_406 ();
 FILLER_ASAP7_75t_R FILLER_121_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_444 ();
 DECAPx4_ASAP7_75t_R FILLER_121_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_463 ();
 DECAPx10_ASAP7_75t_R FILLER_121_473 ();
 DECAPx4_ASAP7_75t_R FILLER_121_495 ();
 FILLER_ASAP7_75t_R FILLER_121_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_507 ();
 DECAPx4_ASAP7_75t_R FILLER_121_540 ();
 FILLER_ASAP7_75t_R FILLER_121_550 ();
 DECAPx2_ASAP7_75t_R FILLER_121_558 ();
 DECAPx1_ASAP7_75t_R FILLER_121_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_583 ();
 DECAPx1_ASAP7_75t_R FILLER_121_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_597 ();
 DECAPx2_ASAP7_75t_R FILLER_121_601 ();
 FILLER_ASAP7_75t_R FILLER_121_607 ();
 DECAPx2_ASAP7_75t_R FILLER_121_615 ();
 FILLER_ASAP7_75t_R FILLER_121_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_626 ();
 FILLER_ASAP7_75t_R FILLER_121_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_635 ();
 FILLER_ASAP7_75t_R FILLER_121_654 ();
 DECAPx6_ASAP7_75t_R FILLER_121_660 ();
 DECAPx2_ASAP7_75t_R FILLER_121_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_680 ();
 DECAPx10_ASAP7_75t_R FILLER_121_685 ();
 DECAPx2_ASAP7_75t_R FILLER_121_707 ();
 DECAPx1_ASAP7_75t_R FILLER_121_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_720 ();
 DECAPx4_ASAP7_75t_R FILLER_121_724 ();
 FILLER_ASAP7_75t_R FILLER_121_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_755 ();
 FILLER_ASAP7_75t_R FILLER_121_788 ();
 DECAPx2_ASAP7_75t_R FILLER_121_793 ();
 FILLER_ASAP7_75t_R FILLER_121_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_801 ();
 FILLER_ASAP7_75t_R FILLER_121_808 ();
 DECAPx10_ASAP7_75t_R FILLER_121_817 ();
 DECAPx2_ASAP7_75t_R FILLER_121_839 ();
 DECAPx1_ASAP7_75t_R FILLER_121_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_864 ();
 DECAPx2_ASAP7_75t_R FILLER_121_874 ();
 FILLER_ASAP7_75t_R FILLER_121_880 ();
 DECAPx10_ASAP7_75t_R FILLER_121_888 ();
 DECAPx6_ASAP7_75t_R FILLER_121_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_953 ();
 DECAPx2_ASAP7_75t_R FILLER_121_978 ();
 DECAPx1_ASAP7_75t_R FILLER_121_993 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_121_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1067 ();
 FILLER_ASAP7_75t_R FILLER_121_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1075 ();
 FILLER_ASAP7_75t_R FILLER_121_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1086 ();
 FILLER_ASAP7_75t_R FILLER_121_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_121_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1265 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1318 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1404 ();
 FILLER_ASAP7_75t_R FILLER_122_28 ();
 FILLER_ASAP7_75t_R FILLER_122_63 ();
 DECAPx4_ASAP7_75t_R FILLER_122_71 ();
 DECAPx1_ASAP7_75t_R FILLER_122_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_91 ();
 DECAPx6_ASAP7_75t_R FILLER_122_98 ();
 FILLER_ASAP7_75t_R FILLER_122_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_114 ();
 DECAPx6_ASAP7_75t_R FILLER_122_131 ();
 DECAPx1_ASAP7_75t_R FILLER_122_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_149 ();
 DECAPx10_ASAP7_75t_R FILLER_122_160 ();
 DECAPx10_ASAP7_75t_R FILLER_122_182 ();
 FILLER_ASAP7_75t_R FILLER_122_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_206 ();
 DECAPx1_ASAP7_75t_R FILLER_122_221 ();
 DECAPx4_ASAP7_75t_R FILLER_122_260 ();
 DECAPx6_ASAP7_75t_R FILLER_122_276 ();
 DECAPx10_ASAP7_75t_R FILLER_122_296 ();
 DECAPx10_ASAP7_75t_R FILLER_122_318 ();
 DECAPx6_ASAP7_75t_R FILLER_122_340 ();
 FILLER_ASAP7_75t_R FILLER_122_368 ();
 DECAPx10_ASAP7_75t_R FILLER_122_384 ();
 DECAPx10_ASAP7_75t_R FILLER_122_406 ();
 DECAPx6_ASAP7_75t_R FILLER_122_428 ();
 FILLER_ASAP7_75t_R FILLER_122_442 ();
 DECAPx1_ASAP7_75t_R FILLER_122_458 ();
 DECAPx2_ASAP7_75t_R FILLER_122_464 ();
 FILLER_ASAP7_75t_R FILLER_122_470 ();
 DECAPx2_ASAP7_75t_R FILLER_122_478 ();
 DECAPx6_ASAP7_75t_R FILLER_122_491 ();
 FILLER_ASAP7_75t_R FILLER_122_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_507 ();
 DECAPx2_ASAP7_75t_R FILLER_122_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_521 ();
 DECAPx2_ASAP7_75t_R FILLER_122_525 ();
 FILLER_ASAP7_75t_R FILLER_122_531 ();
 DECAPx10_ASAP7_75t_R FILLER_122_541 ();
 DECAPx2_ASAP7_75t_R FILLER_122_563 ();
 FILLER_ASAP7_75t_R FILLER_122_569 ();
 DECAPx10_ASAP7_75t_R FILLER_122_577 ();
 FILLER_ASAP7_75t_R FILLER_122_634 ();
 DECAPx2_ASAP7_75t_R FILLER_122_662 ();
 DECAPx4_ASAP7_75t_R FILLER_122_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_684 ();
 DECAPx10_ASAP7_75t_R FILLER_122_688 ();
 DECAPx4_ASAP7_75t_R FILLER_122_710 ();
 FILLER_ASAP7_75t_R FILLER_122_720 ();
 DECAPx10_ASAP7_75t_R FILLER_122_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_749 ();
 DECAPx6_ASAP7_75t_R FILLER_122_760 ();
 DECAPx1_ASAP7_75t_R FILLER_122_774 ();
 FILLER_ASAP7_75t_R FILLER_122_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_805 ();
 DECAPx2_ASAP7_75t_R FILLER_122_833 ();
 FILLER_ASAP7_75t_R FILLER_122_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_841 ();
 DECAPx4_ASAP7_75t_R FILLER_122_848 ();
 DECAPx2_ASAP7_75t_R FILLER_122_913 ();
 FILLER_ASAP7_75t_R FILLER_122_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_932 ();
 DECAPx1_ASAP7_75t_R FILLER_122_955 ();
 DECAPx2_ASAP7_75t_R FILLER_122_975 ();
 FILLER_ASAP7_75t_R FILLER_122_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1018 ();
 FILLER_ASAP7_75t_R FILLER_122_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1063 ();
 FILLER_ASAP7_75t_R FILLER_122_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1103 ();
 FILLER_ASAP7_75t_R FILLER_122_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_122_1199 ();
 FILLER_ASAP7_75t_R FILLER_122_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1226 ();
 FILLER_ASAP7_75t_R FILLER_122_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_122_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1347 ();
 FILLER_ASAP7_75t_R FILLER_122_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1355 ();
 FILLER_ASAP7_75t_R FILLER_122_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1391 ();
 DECAPx2_ASAP7_75t_R FILLER_123_2 ();
 FILLER_ASAP7_75t_R FILLER_123_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_32 ();
 DECAPx1_ASAP7_75t_R FILLER_123_49 ();
 DECAPx6_ASAP7_75t_R FILLER_123_56 ();
 DECAPx2_ASAP7_75t_R FILLER_123_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_76 ();
 DECAPx10_ASAP7_75t_R FILLER_123_106 ();
 DECAPx10_ASAP7_75t_R FILLER_123_128 ();
 FILLER_ASAP7_75t_R FILLER_123_150 ();
 DECAPx4_ASAP7_75t_R FILLER_123_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_216 ();
 DECAPx1_ASAP7_75t_R FILLER_123_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_229 ();
 DECAPx2_ASAP7_75t_R FILLER_123_274 ();
 FILLER_ASAP7_75t_R FILLER_123_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_282 ();
 DECAPx10_ASAP7_75t_R FILLER_123_291 ();
 DECAPx4_ASAP7_75t_R FILLER_123_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_323 ();
 DECAPx1_ASAP7_75t_R FILLER_123_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_360 ();
 DECAPx4_ASAP7_75t_R FILLER_123_367 ();
 FILLER_ASAP7_75t_R FILLER_123_377 ();
 DECAPx2_ASAP7_75t_R FILLER_123_385 ();
 FILLER_ASAP7_75t_R FILLER_123_391 ();
 FILLER_ASAP7_75t_R FILLER_123_399 ();
 DECAPx2_ASAP7_75t_R FILLER_123_409 ();
 DECAPx4_ASAP7_75t_R FILLER_123_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_433 ();
 DECAPx1_ASAP7_75t_R FILLER_123_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_462 ();
 DECAPx6_ASAP7_75t_R FILLER_123_511 ();
 FILLER_ASAP7_75t_R FILLER_123_525 ();
 DECAPx1_ASAP7_75t_R FILLER_123_537 ();
 DECAPx4_ASAP7_75t_R FILLER_123_560 ();
 FILLER_ASAP7_75t_R FILLER_123_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_598 ();
 DECAPx1_ASAP7_75t_R FILLER_123_602 ();
 DECAPx4_ASAP7_75t_R FILLER_123_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_648 ();
 DECAPx2_ASAP7_75t_R FILLER_123_655 ();
 FILLER_ASAP7_75t_R FILLER_123_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_663 ();
 DECAPx2_ASAP7_75t_R FILLER_123_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_712 ();
 DECAPx4_ASAP7_75t_R FILLER_123_716 ();
 FILLER_ASAP7_75t_R FILLER_123_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_728 ();
 DECAPx2_ASAP7_75t_R FILLER_123_732 ();
 DECAPx2_ASAP7_75t_R FILLER_123_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_753 ();
 DECAPx10_ASAP7_75t_R FILLER_123_770 ();
 DECAPx1_ASAP7_75t_R FILLER_123_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_801 ();
 DECAPx2_ASAP7_75t_R FILLER_123_821 ();
 FILLER_ASAP7_75t_R FILLER_123_827 ();
 DECAPx10_ASAP7_75t_R FILLER_123_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_863 ();
 DECAPx1_ASAP7_75t_R FILLER_123_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_884 ();
 FILLER_ASAP7_75t_R FILLER_123_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_897 ();
 DECAPx2_ASAP7_75t_R FILLER_123_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_926 ();
 FILLER_ASAP7_75t_R FILLER_123_939 ();
 DECAPx2_ASAP7_75t_R FILLER_123_956 ();
 DECAPx10_ASAP7_75t_R FILLER_123_968 ();
 DECAPx1_ASAP7_75t_R FILLER_123_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_994 ();
 FILLER_ASAP7_75t_R FILLER_123_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1085 ();
 FILLER_ASAP7_75t_R FILLER_123_1095 ();
 FILLER_ASAP7_75t_R FILLER_123_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1138 ();
 FILLER_ASAP7_75t_R FILLER_123_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1224 ();
 FILLER_ASAP7_75t_R FILLER_123_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1294 ();
 FILLER_ASAP7_75t_R FILLER_123_1300 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1319 ();
 FILLER_ASAP7_75t_R FILLER_123_1334 ();
 FILLER_ASAP7_75t_R FILLER_123_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1341 ();
 FILLER_ASAP7_75t_R FILLER_123_1376 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_124_2 ();
 FILLER_ASAP7_75t_R FILLER_124_58 ();
 DECAPx1_ASAP7_75t_R FILLER_124_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_74 ();
 DECAPx4_ASAP7_75t_R FILLER_124_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_88 ();
 DECAPx2_ASAP7_75t_R FILLER_124_95 ();
 DECAPx4_ASAP7_75t_R FILLER_124_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_131 ();
 DECAPx10_ASAP7_75t_R FILLER_124_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_166 ();
 DECAPx6_ASAP7_75t_R FILLER_124_170 ();
 DECAPx1_ASAP7_75t_R FILLER_124_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_220 ();
 DECAPx1_ASAP7_75t_R FILLER_124_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_233 ();
 DECAPx4_ASAP7_75t_R FILLER_124_298 ();
 FILLER_ASAP7_75t_R FILLER_124_374 ();
 DECAPx6_ASAP7_75t_R FILLER_124_428 ();
 DECAPx1_ASAP7_75t_R FILLER_124_458 ();
 DECAPx6_ASAP7_75t_R FILLER_124_464 ();
 DECAPx2_ASAP7_75t_R FILLER_124_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_484 ();
 DECAPx1_ASAP7_75t_R FILLER_124_491 ();
 DECAPx6_ASAP7_75t_R FILLER_124_534 ();
 FILLER_ASAP7_75t_R FILLER_124_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_577 ();
 DECAPx4_ASAP7_75t_R FILLER_124_616 ();
 DECAPx6_ASAP7_75t_R FILLER_124_629 ();
 DECAPx1_ASAP7_75t_R FILLER_124_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_647 ();
 DECAPx2_ASAP7_75t_R FILLER_124_682 ();
 DECAPx10_ASAP7_75t_R FILLER_124_756 ();
 DECAPx10_ASAP7_75t_R FILLER_124_778 ();
 DECAPx4_ASAP7_75t_R FILLER_124_800 ();
 DECAPx6_ASAP7_75t_R FILLER_124_817 ();
 DECAPx2_ASAP7_75t_R FILLER_124_831 ();
 FILLER_ASAP7_75t_R FILLER_124_845 ();
 DECAPx10_ASAP7_75t_R FILLER_124_857 ();
 DECAPx2_ASAP7_75t_R FILLER_124_879 ();
 DECAPx1_ASAP7_75t_R FILLER_124_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_905 ();
 DECAPx10_ASAP7_75t_R FILLER_124_921 ();
 DECAPx6_ASAP7_75t_R FILLER_124_943 ();
 FILLER_ASAP7_75t_R FILLER_124_957 ();
 DECAPx6_ASAP7_75t_R FILLER_124_994 ();
 FILLER_ASAP7_75t_R FILLER_124_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1025 ();
 FILLER_ASAP7_75t_R FILLER_124_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1058 ();
 FILLER_ASAP7_75t_R FILLER_124_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1078 ();
 FILLER_ASAP7_75t_R FILLER_124_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1086 ();
 FILLER_ASAP7_75t_R FILLER_124_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1150 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1170 ();
 FILLER_ASAP7_75t_R FILLER_124_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1236 ();
 FILLER_ASAP7_75t_R FILLER_124_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1300 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1322 ();
 FILLER_ASAP7_75t_R FILLER_124_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1388 ();
 FILLER_ASAP7_75t_R FILLER_124_1403 ();
 DECAPx6_ASAP7_75t_R FILLER_125_2 ();
 DECAPx1_ASAP7_75t_R FILLER_125_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_20 ();
 DECAPx2_ASAP7_75t_R FILLER_125_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_34 ();
 DECAPx2_ASAP7_75t_R FILLER_125_51 ();
 FILLER_ASAP7_75t_R FILLER_125_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_59 ();
 DECAPx2_ASAP7_75t_R FILLER_125_86 ();
 FILLER_ASAP7_75t_R FILLER_125_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_94 ();
 DECAPx10_ASAP7_75t_R FILLER_125_166 ();
 DECAPx1_ASAP7_75t_R FILLER_125_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_192 ();
 DECAPx2_ASAP7_75t_R FILLER_125_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_202 ();
 DECAPx1_ASAP7_75t_R FILLER_125_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_219 ();
 DECAPx4_ASAP7_75t_R FILLER_125_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_236 ();
 DECAPx10_ASAP7_75t_R FILLER_125_243 ();
 DECAPx6_ASAP7_75t_R FILLER_125_265 ();
 FILLER_ASAP7_75t_R FILLER_125_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_281 ();
 DECAPx4_ASAP7_75t_R FILLER_125_288 ();
 FILLER_ASAP7_75t_R FILLER_125_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_314 ();
 DECAPx2_ASAP7_75t_R FILLER_125_330 ();
 FILLER_ASAP7_75t_R FILLER_125_336 ();
 FILLER_ASAP7_75t_R FILLER_125_341 ();
 DECAPx2_ASAP7_75t_R FILLER_125_349 ();
 FILLER_ASAP7_75t_R FILLER_125_355 ();
 DECAPx4_ASAP7_75t_R FILLER_125_366 ();
 FILLER_ASAP7_75t_R FILLER_125_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_378 ();
 FILLER_ASAP7_75t_R FILLER_125_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_387 ();
 DECAPx1_ASAP7_75t_R FILLER_125_394 ();
 DECAPx10_ASAP7_75t_R FILLER_125_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_426 ();
 DECAPx6_ASAP7_75t_R FILLER_125_433 ();
 DECAPx10_ASAP7_75t_R FILLER_125_453 ();
 DECAPx10_ASAP7_75t_R FILLER_125_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_508 ();
 DECAPx2_ASAP7_75t_R FILLER_125_527 ();
 FILLER_ASAP7_75t_R FILLER_125_533 ();
 DECAPx1_ASAP7_75t_R FILLER_125_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_553 ();
 DECAPx1_ASAP7_75t_R FILLER_125_582 ();
 DECAPx2_ASAP7_75t_R FILLER_125_595 ();
 FILLER_ASAP7_75t_R FILLER_125_601 ();
 DECAPx10_ASAP7_75t_R FILLER_125_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_631 ();
 FILLER_ASAP7_75t_R FILLER_125_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_648 ();
 DECAPx2_ASAP7_75t_R FILLER_125_655 ();
 FILLER_ASAP7_75t_R FILLER_125_661 ();
 DECAPx1_ASAP7_75t_R FILLER_125_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_670 ();
 DECAPx6_ASAP7_75t_R FILLER_125_706 ();
 FILLER_ASAP7_75t_R FILLER_125_720 ();
 FILLER_ASAP7_75t_R FILLER_125_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_786 ();
 DECAPx4_ASAP7_75t_R FILLER_125_790 ();
 FILLER_ASAP7_75t_R FILLER_125_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_802 ();
 DECAPx6_ASAP7_75t_R FILLER_125_809 ();
 FILLER_ASAP7_75t_R FILLER_125_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_835 ();
 DECAPx2_ASAP7_75t_R FILLER_125_845 ();
 FILLER_ASAP7_75t_R FILLER_125_851 ();
 DECAPx6_ASAP7_75t_R FILLER_125_867 ();
 DECAPx2_ASAP7_75t_R FILLER_125_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_887 ();
 DECAPx4_ASAP7_75t_R FILLER_125_891 ();
 FILLER_ASAP7_75t_R FILLER_125_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_903 ();
 DECAPx6_ASAP7_75t_R FILLER_125_907 ();
 DECAPx1_ASAP7_75t_R FILLER_125_935 ();
 DECAPx4_ASAP7_75t_R FILLER_125_953 ();
 DECAPx2_ASAP7_75t_R FILLER_125_979 ();
 FILLER_ASAP7_75t_R FILLER_125_985 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1021 ();
 FILLER_ASAP7_75t_R FILLER_125_1027 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1050 ();
 FILLER_ASAP7_75t_R FILLER_125_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1147 ();
 FILLER_ASAP7_75t_R FILLER_125_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1179 ();
 FILLER_ASAP7_75t_R FILLER_125_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1208 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1356 ();
 FILLER_ASAP7_75t_R FILLER_125_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1368 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_126_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_6 ();
 DECAPx10_ASAP7_75t_R FILLER_126_29 ();
 DECAPx6_ASAP7_75t_R FILLER_126_51 ();
 FILLER_ASAP7_75t_R FILLER_126_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_73 ();
 DECAPx6_ASAP7_75t_R FILLER_126_84 ();
 FILLER_ASAP7_75t_R FILLER_126_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_100 ();
 DECAPx2_ASAP7_75t_R FILLER_126_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_110 ();
 DECAPx2_ASAP7_75t_R FILLER_126_114 ();
 FILLER_ASAP7_75t_R FILLER_126_120 ();
 DECAPx1_ASAP7_75t_R FILLER_126_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_178 ();
 DECAPx4_ASAP7_75t_R FILLER_126_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_204 ();
 DECAPx10_ASAP7_75t_R FILLER_126_217 ();
 DECAPx6_ASAP7_75t_R FILLER_126_239 ();
 DECAPx1_ASAP7_75t_R FILLER_126_253 ();
 FILLER_ASAP7_75t_R FILLER_126_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_266 ();
 DECAPx6_ASAP7_75t_R FILLER_126_273 ();
 DECAPx1_ASAP7_75t_R FILLER_126_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_305 ();
 DECAPx10_ASAP7_75t_R FILLER_126_312 ();
 DECAPx2_ASAP7_75t_R FILLER_126_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_340 ();
 DECAPx10_ASAP7_75t_R FILLER_126_347 ();
 DECAPx10_ASAP7_75t_R FILLER_126_377 ();
 DECAPx6_ASAP7_75t_R FILLER_126_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_413 ();
 DECAPx1_ASAP7_75t_R FILLER_126_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_424 ();
 DECAPx4_ASAP7_75t_R FILLER_126_443 ();
 FILLER_ASAP7_75t_R FILLER_126_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_455 ();
 DECAPx6_ASAP7_75t_R FILLER_126_470 ();
 FILLER_ASAP7_75t_R FILLER_126_484 ();
 DECAPx10_ASAP7_75t_R FILLER_126_498 ();
 DECAPx10_ASAP7_75t_R FILLER_126_520 ();
 DECAPx10_ASAP7_75t_R FILLER_126_542 ();
 DECAPx2_ASAP7_75t_R FILLER_126_564 ();
 FILLER_ASAP7_75t_R FILLER_126_570 ();
 DECAPx4_ASAP7_75t_R FILLER_126_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_588 ();
 DECAPx1_ASAP7_75t_R FILLER_126_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_603 ();
 FILLER_ASAP7_75t_R FILLER_126_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_632 ();
 DECAPx2_ASAP7_75t_R FILLER_126_668 ();
 FILLER_ASAP7_75t_R FILLER_126_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_676 ();
 DECAPx2_ASAP7_75t_R FILLER_126_683 ();
 FILLER_ASAP7_75t_R FILLER_126_689 ();
 DECAPx2_ASAP7_75t_R FILLER_126_694 ();
 FILLER_ASAP7_75t_R FILLER_126_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_702 ();
 DECAPx6_ASAP7_75t_R FILLER_126_715 ();
 FILLER_ASAP7_75t_R FILLER_126_729 ();
 DECAPx6_ASAP7_75t_R FILLER_126_747 ();
 DECAPx2_ASAP7_75t_R FILLER_126_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_798 ();
 DECAPx2_ASAP7_75t_R FILLER_126_814 ();
 DECAPx2_ASAP7_75t_R FILLER_126_861 ();
 FILLER_ASAP7_75t_R FILLER_126_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_869 ();
 FILLER_ASAP7_75t_R FILLER_126_902 ();
 DECAPx10_ASAP7_75t_R FILLER_126_939 ();
 FILLER_ASAP7_75t_R FILLER_126_961 ();
 DECAPx10_ASAP7_75t_R FILLER_126_969 ();
 DECAPx1_ASAP7_75t_R FILLER_126_991 ();
 FILLER_ASAP7_75t_R FILLER_126_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1094 ();
 FILLER_ASAP7_75t_R FILLER_126_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1103 ();
 FILLER_ASAP7_75t_R FILLER_126_1110 ();
 FILLER_ASAP7_75t_R FILLER_126_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1183 ();
 FILLER_ASAP7_75t_R FILLER_126_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1195 ();
 FILLER_ASAP7_75t_R FILLER_126_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1217 ();
 FILLER_ASAP7_75t_R FILLER_126_1233 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1253 ();
 FILLER_ASAP7_75t_R FILLER_126_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1276 ();
 FILLER_ASAP7_75t_R FILLER_126_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1320 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1382 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_127_2 ();
 FILLER_ASAP7_75t_R FILLER_127_16 ();
 DECAPx1_ASAP7_75t_R FILLER_127_28 ();
 DECAPx1_ASAP7_75t_R FILLER_127_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_58 ();
 DECAPx2_ASAP7_75t_R FILLER_127_62 ();
 DECAPx2_ASAP7_75t_R FILLER_127_120 ();
 FILLER_ASAP7_75t_R FILLER_127_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_200 ();
 FILLER_ASAP7_75t_R FILLER_127_215 ();
 DECAPx4_ASAP7_75t_R FILLER_127_231 ();
 DECAPx1_ASAP7_75t_R FILLER_127_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_251 ();
 DECAPx4_ASAP7_75t_R FILLER_127_278 ();
 FILLER_ASAP7_75t_R FILLER_127_288 ();
 DECAPx10_ASAP7_75t_R FILLER_127_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_318 ();
 DECAPx4_ASAP7_75t_R FILLER_127_325 ();
 DECAPx2_ASAP7_75t_R FILLER_127_347 ();
 DECAPx6_ASAP7_75t_R FILLER_127_359 ();
 DECAPx6_ASAP7_75t_R FILLER_127_385 ();
 DECAPx1_ASAP7_75t_R FILLER_127_399 ();
 DECAPx4_ASAP7_75t_R FILLER_127_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_433 ();
 DECAPx1_ASAP7_75t_R FILLER_127_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_452 ();
 DECAPx10_ASAP7_75t_R FILLER_127_495 ();
 DECAPx4_ASAP7_75t_R FILLER_127_517 ();
 DECAPx4_ASAP7_75t_R FILLER_127_545 ();
 DECAPx2_ASAP7_75t_R FILLER_127_561 ();
 FILLER_ASAP7_75t_R FILLER_127_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_569 ();
 DECAPx6_ASAP7_75t_R FILLER_127_580 ();
 FILLER_ASAP7_75t_R FILLER_127_594 ();
 DECAPx2_ASAP7_75t_R FILLER_127_644 ();
 FILLER_ASAP7_75t_R FILLER_127_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_652 ();
 DECAPx4_ASAP7_75t_R FILLER_127_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_731 ();
 DECAPx10_ASAP7_75t_R FILLER_127_738 ();
 DECAPx6_ASAP7_75t_R FILLER_127_760 ();
 DECAPx2_ASAP7_75t_R FILLER_127_786 ();
 FILLER_ASAP7_75t_R FILLER_127_792 ();
 DECAPx4_ASAP7_75t_R FILLER_127_817 ();
 FILLER_ASAP7_75t_R FILLER_127_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_832 ();
 FILLER_ASAP7_75t_R FILLER_127_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_841 ();
 FILLER_ASAP7_75t_R FILLER_127_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_884 ();
 DECAPx1_ASAP7_75t_R FILLER_127_899 ();
 FILLER_ASAP7_75t_R FILLER_127_922 ();
 DECAPx6_ASAP7_75t_R FILLER_127_932 ();
 DECAPx2_ASAP7_75t_R FILLER_127_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_961 ();
 DECAPx10_ASAP7_75t_R FILLER_127_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1051 ();
 FILLER_ASAP7_75t_R FILLER_127_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1074 ();
 FILLER_ASAP7_75t_R FILLER_127_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1148 ();
 FILLER_ASAP7_75t_R FILLER_127_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1169 ();
 FILLER_ASAP7_75t_R FILLER_127_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1225 ();
 FILLER_ASAP7_75t_R FILLER_127_1232 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1237 ();
 FILLER_ASAP7_75t_R FILLER_127_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1278 ();
 FILLER_ASAP7_75t_R FILLER_127_1293 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1321 ();
 FILLER_ASAP7_75t_R FILLER_127_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1370 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1390 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1399 ();
 DECAPx2_ASAP7_75t_R FILLER_128_2 ();
 DECAPx1_ASAP7_75t_R FILLER_128_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_78 ();
 FILLER_ASAP7_75t_R FILLER_128_85 ();
 DECAPx1_ASAP7_75t_R FILLER_128_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_94 ();
 FILLER_ASAP7_75t_R FILLER_128_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_156 ();
 FILLER_ASAP7_75t_R FILLER_128_170 ();
 DECAPx1_ASAP7_75t_R FILLER_128_179 ();
 DECAPx1_ASAP7_75t_R FILLER_128_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_190 ();
 DECAPx1_ASAP7_75t_R FILLER_128_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_221 ();
 FILLER_ASAP7_75t_R FILLER_128_241 ();
 DECAPx6_ASAP7_75t_R FILLER_128_251 ();
 FILLER_ASAP7_75t_R FILLER_128_265 ();
 DECAPx1_ASAP7_75t_R FILLER_128_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_274 ();
 DECAPx1_ASAP7_75t_R FILLER_128_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_305 ();
 FILLER_ASAP7_75t_R FILLER_128_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_336 ();
 FILLER_ASAP7_75t_R FILLER_128_349 ();
 DECAPx1_ASAP7_75t_R FILLER_128_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_371 ();
 DECAPx10_ASAP7_75t_R FILLER_128_380 ();
 DECAPx2_ASAP7_75t_R FILLER_128_410 ();
 FILLER_ASAP7_75t_R FILLER_128_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_418 ();
 FILLER_ASAP7_75t_R FILLER_128_433 ();
 DECAPx2_ASAP7_75t_R FILLER_128_447 ();
 FILLER_ASAP7_75t_R FILLER_128_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_461 ();
 DECAPx2_ASAP7_75t_R FILLER_128_470 ();
 FILLER_ASAP7_75t_R FILLER_128_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_478 ();
 DECAPx4_ASAP7_75t_R FILLER_128_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_549 ();
 DECAPx2_ASAP7_75t_R FILLER_128_592 ();
 FILLER_ASAP7_75t_R FILLER_128_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_603 ();
 DECAPx2_ASAP7_75t_R FILLER_128_610 ();
 FILLER_ASAP7_75t_R FILLER_128_616 ();
 FILLER_ASAP7_75t_R FILLER_128_621 ();
 DECAPx2_ASAP7_75t_R FILLER_128_626 ();
 FILLER_ASAP7_75t_R FILLER_128_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_704 ();
 DECAPx1_ASAP7_75t_R FILLER_128_711 ();
 DECAPx4_ASAP7_75t_R FILLER_128_718 ();
 FILLER_ASAP7_75t_R FILLER_128_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_730 ();
 DECAPx2_ASAP7_75t_R FILLER_128_746 ();
 FILLER_ASAP7_75t_R FILLER_128_752 ();
 DECAPx6_ASAP7_75t_R FILLER_128_778 ();
 DECAPx1_ASAP7_75t_R FILLER_128_792 ();
 DECAPx10_ASAP7_75t_R FILLER_128_807 ();
 DECAPx6_ASAP7_75t_R FILLER_128_829 ();
 DECAPx2_ASAP7_75t_R FILLER_128_843 ();
 DECAPx4_ASAP7_75t_R FILLER_128_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_865 ();
 DECAPx2_ASAP7_75t_R FILLER_128_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_881 ();
 DECAPx10_ASAP7_75t_R FILLER_128_888 ();
 DECAPx10_ASAP7_75t_R FILLER_128_910 ();
 DECAPx4_ASAP7_75t_R FILLER_128_932 ();
 FILLER_ASAP7_75t_R FILLER_128_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_944 ();
 DECAPx2_ASAP7_75t_R FILLER_128_957 ();
 FILLER_ASAP7_75t_R FILLER_128_963 ();
 DECAPx10_ASAP7_75t_R FILLER_128_988 ();
 FILLER_ASAP7_75t_R FILLER_128_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1020 ();
 FILLER_ASAP7_75t_R FILLER_128_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1053 ();
 FILLER_ASAP7_75t_R FILLER_128_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1070 ();
 FILLER_ASAP7_75t_R FILLER_128_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1234 ();
 FILLER_ASAP7_75t_R FILLER_128_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1281 ();
 FILLER_ASAP7_75t_R FILLER_128_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1313 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1369 ();
 FILLER_ASAP7_75t_R FILLER_128_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1388 ();
 FILLER_ASAP7_75t_R FILLER_128_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_129_2 ();
 DECAPx2_ASAP7_75t_R FILLER_129_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_22 ();
 DECAPx4_ASAP7_75t_R FILLER_129_26 ();
 DECAPx1_ASAP7_75t_R FILLER_129_72 ();
 FILLER_ASAP7_75t_R FILLER_129_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_90 ();
 DECAPx6_ASAP7_75t_R FILLER_129_103 ();
 DECAPx6_ASAP7_75t_R FILLER_129_182 ();
 DECAPx1_ASAP7_75t_R FILLER_129_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_200 ();
 FILLER_ASAP7_75t_R FILLER_129_209 ();
 DECAPx1_ASAP7_75t_R FILLER_129_239 ();
 DECAPx10_ASAP7_75t_R FILLER_129_251 ();
 DECAPx1_ASAP7_75t_R FILLER_129_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_284 ();
 DECAPx1_ASAP7_75t_R FILLER_129_301 ();
 DECAPx1_ASAP7_75t_R FILLER_129_333 ();
 FILLER_ASAP7_75t_R FILLER_129_351 ();
 DECAPx6_ASAP7_75t_R FILLER_129_359 ();
 FILLER_ASAP7_75t_R FILLER_129_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_375 ();
 DECAPx1_ASAP7_75t_R FILLER_129_394 ();
 DECAPx1_ASAP7_75t_R FILLER_129_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_408 ();
 DECAPx1_ASAP7_75t_R FILLER_129_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_419 ();
 DECAPx6_ASAP7_75t_R FILLER_129_429 ();
 DECAPx2_ASAP7_75t_R FILLER_129_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_472 ();
 DECAPx1_ASAP7_75t_R FILLER_129_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_494 ();
 FILLER_ASAP7_75t_R FILLER_129_502 ();
 FILLER_ASAP7_75t_R FILLER_129_559 ();
 FILLER_ASAP7_75t_R FILLER_129_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_576 ();
 DECAPx10_ASAP7_75t_R FILLER_129_609 ();
 DECAPx10_ASAP7_75t_R FILLER_129_631 ();
 DECAPx1_ASAP7_75t_R FILLER_129_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_657 ();
 DECAPx2_ASAP7_75t_R FILLER_129_664 ();
 FILLER_ASAP7_75t_R FILLER_129_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_672 ();
 DECAPx1_ASAP7_75t_R FILLER_129_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_692 ();
 FILLER_ASAP7_75t_R FILLER_129_696 ();
 DECAPx10_ASAP7_75t_R FILLER_129_702 ();
 DECAPx2_ASAP7_75t_R FILLER_129_724 ();
 FILLER_ASAP7_75t_R FILLER_129_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_732 ();
 DECAPx6_ASAP7_75t_R FILLER_129_745 ();
 DECAPx1_ASAP7_75t_R FILLER_129_759 ();
 DECAPx10_ASAP7_75t_R FILLER_129_779 ();
 DECAPx2_ASAP7_75t_R FILLER_129_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_807 ();
 DECAPx6_ASAP7_75t_R FILLER_129_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_830 ();
 DECAPx10_ASAP7_75t_R FILLER_129_847 ();
 DECAPx4_ASAP7_75t_R FILLER_129_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_879 ();
 DECAPx4_ASAP7_75t_R FILLER_129_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_897 ();
 DECAPx2_ASAP7_75t_R FILLER_129_907 ();
 DECAPx1_ASAP7_75t_R FILLER_129_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_923 ();
 DECAPx1_ASAP7_75t_R FILLER_129_926 ();
 DECAPx2_ASAP7_75t_R FILLER_129_967 ();
 FILLER_ASAP7_75t_R FILLER_129_973 ();
 DECAPx1_ASAP7_75t_R FILLER_129_984 ();
 FILLER_ASAP7_75t_R FILLER_129_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_129_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1113 ();
 FILLER_ASAP7_75t_R FILLER_129_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1190 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1211 ();
 FILLER_ASAP7_75t_R FILLER_129_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1250 ();
 FILLER_ASAP7_75t_R FILLER_129_1264 ();
 FILLER_ASAP7_75t_R FILLER_129_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1293 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_129_1333 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1355 ();
 FILLER_ASAP7_75t_R FILLER_129_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1367 ();
 DECAPx2_ASAP7_75t_R FILLER_130_2 ();
 DECAPx6_ASAP7_75t_R FILLER_130_20 ();
 DECAPx2_ASAP7_75t_R FILLER_130_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_40 ();
 DECAPx1_ASAP7_75t_R FILLER_130_57 ();
 DECAPx6_ASAP7_75t_R FILLER_130_113 ();
 FILLER_ASAP7_75t_R FILLER_130_127 ();
 DECAPx1_ASAP7_75t_R FILLER_130_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_136 ();
 DECAPx6_ASAP7_75t_R FILLER_130_153 ();
 DECAPx1_ASAP7_75t_R FILLER_130_167 ();
 DECAPx6_ASAP7_75t_R FILLER_130_174 ();
 DECAPx6_ASAP7_75t_R FILLER_130_202 ();
 DECAPx2_ASAP7_75t_R FILLER_130_216 ();
 DECAPx4_ASAP7_75t_R FILLER_130_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_240 ();
 DECAPx2_ASAP7_75t_R FILLER_130_247 ();
 FILLER_ASAP7_75t_R FILLER_130_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_255 ();
 DECAPx2_ASAP7_75t_R FILLER_130_259 ();
 DECAPx4_ASAP7_75t_R FILLER_130_271 ();
 FILLER_ASAP7_75t_R FILLER_130_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_283 ();
 DECAPx2_ASAP7_75t_R FILLER_130_310 ();
 FILLER_ASAP7_75t_R FILLER_130_316 ();
 DECAPx10_ASAP7_75t_R FILLER_130_324 ();
 DECAPx2_ASAP7_75t_R FILLER_130_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_352 ();
 FILLER_ASAP7_75t_R FILLER_130_360 ();
 DECAPx1_ASAP7_75t_R FILLER_130_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_381 ();
 DECAPx6_ASAP7_75t_R FILLER_130_396 ();
 DECAPx2_ASAP7_75t_R FILLER_130_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_443 ();
 DECAPx1_ASAP7_75t_R FILLER_130_458 ();
 DECAPx4_ASAP7_75t_R FILLER_130_470 ();
 FILLER_ASAP7_75t_R FILLER_130_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_482 ();
 DECAPx4_ASAP7_75t_R FILLER_130_512 ();
 FILLER_ASAP7_75t_R FILLER_130_522 ();
 DECAPx10_ASAP7_75t_R FILLER_130_536 ();
 DECAPx10_ASAP7_75t_R FILLER_130_558 ();
 DECAPx2_ASAP7_75t_R FILLER_130_580 ();
 DECAPx2_ASAP7_75t_R FILLER_130_592 ();
 FILLER_ASAP7_75t_R FILLER_130_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_600 ();
 FILLER_ASAP7_75t_R FILLER_130_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_609 ();
 DECAPx2_ASAP7_75t_R FILLER_130_616 ();
 DECAPx1_ASAP7_75t_R FILLER_130_628 ();
 FILLER_ASAP7_75t_R FILLER_130_650 ();
 DECAPx4_ASAP7_75t_R FILLER_130_687 ();
 FILLER_ASAP7_75t_R FILLER_130_697 ();
 DECAPx2_ASAP7_75t_R FILLER_130_705 ();
 FILLER_ASAP7_75t_R FILLER_130_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_713 ();
 DECAPx6_ASAP7_75t_R FILLER_130_718 ();
 DECAPx1_ASAP7_75t_R FILLER_130_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_736 ();
 DECAPx1_ASAP7_75t_R FILLER_130_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_748 ();
 DECAPx2_ASAP7_75t_R FILLER_130_759 ();
 FILLER_ASAP7_75t_R FILLER_130_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_767 ();
 FILLER_ASAP7_75t_R FILLER_130_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_776 ();
 DECAPx2_ASAP7_75t_R FILLER_130_787 ();
 FILLER_ASAP7_75t_R FILLER_130_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_795 ();
 FILLER_ASAP7_75t_R FILLER_130_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_806 ();
 DECAPx1_ASAP7_75t_R FILLER_130_835 ();
 DECAPx2_ASAP7_75t_R FILLER_130_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_857 ();
 DECAPx1_ASAP7_75t_R FILLER_130_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_884 ();
 DECAPx1_ASAP7_75t_R FILLER_130_895 ();
 FILLER_ASAP7_75t_R FILLER_130_915 ();
 FILLER_ASAP7_75t_R FILLER_130_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_929 ();
 DECAPx10_ASAP7_75t_R FILLER_130_940 ();
 DECAPx10_ASAP7_75t_R FILLER_130_962 ();
 DECAPx2_ASAP7_75t_R FILLER_130_984 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1021 ();
 FILLER_ASAP7_75t_R FILLER_130_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1138 ();
 FILLER_ASAP7_75t_R FILLER_130_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1171 ();
 FILLER_ASAP7_75t_R FILLER_130_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1245 ();
 FILLER_ASAP7_75t_R FILLER_130_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1303 ();
 FILLER_ASAP7_75t_R FILLER_130_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1385 ();
 FILLER_ASAP7_75t_R FILLER_130_1394 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1399 ();
 FILLER_ASAP7_75t_R FILLER_131_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_4 ();
 FILLER_ASAP7_75t_R FILLER_131_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_33 ();
 DECAPx10_ASAP7_75t_R FILLER_131_37 ();
 FILLER_ASAP7_75t_R FILLER_131_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_75 ();
 DECAPx4_ASAP7_75t_R FILLER_131_106 ();
 DECAPx10_ASAP7_75t_R FILLER_131_122 ();
 DECAPx6_ASAP7_75t_R FILLER_131_144 ();
 FILLER_ASAP7_75t_R FILLER_131_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_160 ();
 DECAPx1_ASAP7_75t_R FILLER_131_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_174 ();
 DECAPx6_ASAP7_75t_R FILLER_131_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_218 ();
 DECAPx10_ASAP7_75t_R FILLER_131_225 ();
 DECAPx6_ASAP7_75t_R FILLER_131_279 ();
 DECAPx2_ASAP7_75t_R FILLER_131_293 ();
 DECAPx2_ASAP7_75t_R FILLER_131_302 ();
 DECAPx2_ASAP7_75t_R FILLER_131_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_317 ();
 DECAPx2_ASAP7_75t_R FILLER_131_321 ();
 FILLER_ASAP7_75t_R FILLER_131_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_329 ();
 DECAPx1_ASAP7_75t_R FILLER_131_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_376 ();
 DECAPx6_ASAP7_75t_R FILLER_131_380 ();
 DECAPx2_ASAP7_75t_R FILLER_131_394 ();
 DECAPx2_ASAP7_75t_R FILLER_131_409 ();
 FILLER_ASAP7_75t_R FILLER_131_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_417 ();
 DECAPx6_ASAP7_75t_R FILLER_131_434 ();
 FILLER_ASAP7_75t_R FILLER_131_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_450 ();
 DECAPx6_ASAP7_75t_R FILLER_131_465 ();
 DECAPx1_ASAP7_75t_R FILLER_131_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_483 ();
 DECAPx10_ASAP7_75t_R FILLER_131_500 ();
 DECAPx6_ASAP7_75t_R FILLER_131_522 ();
 DECAPx1_ASAP7_75t_R FILLER_131_536 ();
 DECAPx6_ASAP7_75t_R FILLER_131_550 ();
 FILLER_ASAP7_75t_R FILLER_131_564 ();
 DECAPx2_ASAP7_75t_R FILLER_131_572 ();
 DECAPx1_ASAP7_75t_R FILLER_131_636 ();
 FILLER_ASAP7_75t_R FILLER_131_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_724 ();
 DECAPx2_ASAP7_75t_R FILLER_131_764 ();
 DECAPx2_ASAP7_75t_R FILLER_131_806 ();
 DECAPx4_ASAP7_75t_R FILLER_131_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_825 ();
 DECAPx1_ASAP7_75t_R FILLER_131_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_857 ();
 FILLER_ASAP7_75t_R FILLER_131_880 ();
 DECAPx1_ASAP7_75t_R FILLER_131_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_905 ();
 DECAPx2_ASAP7_75t_R FILLER_131_915 ();
 FILLER_ASAP7_75t_R FILLER_131_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_923 ();
 DECAPx10_ASAP7_75t_R FILLER_131_932 ();
 DECAPx4_ASAP7_75t_R FILLER_131_954 ();
 FILLER_ASAP7_75t_R FILLER_131_964 ();
 DECAPx10_ASAP7_75t_R FILLER_131_982 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1061 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1077 ();
 FILLER_ASAP7_75t_R FILLER_131_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1172 ();
 FILLER_ASAP7_75t_R FILLER_131_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1212 ();
 FILLER_ASAP7_75t_R FILLER_131_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1270 ();
 FILLER_ASAP7_75t_R FILLER_131_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1296 ();
 FILLER_ASAP7_75t_R FILLER_131_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1314 ();
 FILLER_ASAP7_75t_R FILLER_131_1320 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1348 ();
 FILLER_ASAP7_75t_R FILLER_131_1358 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1360 ();
 FILLER_ASAP7_75t_R FILLER_131_1376 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_132_2 ();
 FILLER_ASAP7_75t_R FILLER_132_8 ();
 FILLER_ASAP7_75t_R FILLER_132_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_87 ();
 FILLER_ASAP7_75t_R FILLER_132_123 ();
 DECAPx1_ASAP7_75t_R FILLER_132_132 ();
 DECAPx6_ASAP7_75t_R FILLER_132_139 ();
 DECAPx1_ASAP7_75t_R FILLER_132_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_183 ();
 DECAPx6_ASAP7_75t_R FILLER_132_212 ();
 FILLER_ASAP7_75t_R FILLER_132_226 ();
 FILLER_ASAP7_75t_R FILLER_132_234 ();
 DECAPx6_ASAP7_75t_R FILLER_132_242 ();
 DECAPx2_ASAP7_75t_R FILLER_132_256 ();
 DECAPx6_ASAP7_75t_R FILLER_132_265 ();
 DECAPx1_ASAP7_75t_R FILLER_132_279 ();
 DECAPx2_ASAP7_75t_R FILLER_132_290 ();
 DECAPx2_ASAP7_75t_R FILLER_132_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_305 ();
 DECAPx2_ASAP7_75t_R FILLER_132_319 ();
 DECAPx4_ASAP7_75t_R FILLER_132_355 ();
 DECAPx10_ASAP7_75t_R FILLER_132_368 ();
 DECAPx2_ASAP7_75t_R FILLER_132_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_405 ();
 FILLER_ASAP7_75t_R FILLER_132_414 ();
 DECAPx2_ASAP7_75t_R FILLER_132_448 ();
 DECAPx1_ASAP7_75t_R FILLER_132_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_461 ();
 DECAPx6_ASAP7_75t_R FILLER_132_464 ();
 DECAPx2_ASAP7_75t_R FILLER_132_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_494 ();
 DECAPx6_ASAP7_75t_R FILLER_132_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_589 ();
 DECAPx2_ASAP7_75t_R FILLER_132_602 ();
 FILLER_ASAP7_75t_R FILLER_132_608 ();
 FILLER_ASAP7_75t_R FILLER_132_616 ();
 DECAPx1_ASAP7_75t_R FILLER_132_683 ();
 DECAPx2_ASAP7_75t_R FILLER_132_704 ();
 DECAPx4_ASAP7_75t_R FILLER_132_713 ();
 FILLER_ASAP7_75t_R FILLER_132_723 ();
 DECAPx4_ASAP7_75t_R FILLER_132_751 ();
 DECAPx2_ASAP7_75t_R FILLER_132_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_780 ();
 DECAPx10_ASAP7_75t_R FILLER_132_787 ();
 FILLER_ASAP7_75t_R FILLER_132_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_811 ();
 DECAPx4_ASAP7_75t_R FILLER_132_815 ();
 DECAPx4_ASAP7_75t_R FILLER_132_834 ();
 FILLER_ASAP7_75t_R FILLER_132_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_846 ();
 DECAPx6_ASAP7_75t_R FILLER_132_856 ();
 FILLER_ASAP7_75t_R FILLER_132_870 ();
 DECAPx4_ASAP7_75t_R FILLER_132_878 ();
 FILLER_ASAP7_75t_R FILLER_132_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_890 ();
 DECAPx2_ASAP7_75t_R FILLER_132_897 ();
 FILLER_ASAP7_75t_R FILLER_132_903 ();
 DECAPx10_ASAP7_75t_R FILLER_132_914 ();
 DECAPx6_ASAP7_75t_R FILLER_132_936 ();
 DECAPx1_ASAP7_75t_R FILLER_132_950 ();
 FILLER_ASAP7_75t_R FILLER_132_963 ();
 DECAPx2_ASAP7_75t_R FILLER_132_974 ();
 FILLER_ASAP7_75t_R FILLER_132_980 ();
 DECAPx4_ASAP7_75t_R FILLER_132_991 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1038 ();
 FILLER_ASAP7_75t_R FILLER_132_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1133 ();
 FILLER_ASAP7_75t_R FILLER_132_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1288 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1307 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1318 ();
 FILLER_ASAP7_75t_R FILLER_132_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1326 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1361 ();
 FILLER_ASAP7_75t_R FILLER_132_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1401 ();
 DECAPx4_ASAP7_75t_R FILLER_133_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_19 ();
 FILLER_ASAP7_75t_R FILLER_133_23 ();
 DECAPx2_ASAP7_75t_R FILLER_133_28 ();
 FILLER_ASAP7_75t_R FILLER_133_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_36 ();
 DECAPx4_ASAP7_75t_R FILLER_133_63 ();
 FILLER_ASAP7_75t_R FILLER_133_73 ();
 FILLER_ASAP7_75t_R FILLER_133_78 ();
 DECAPx2_ASAP7_75t_R FILLER_133_83 ();
 FILLER_ASAP7_75t_R FILLER_133_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_91 ();
 FILLER_ASAP7_75t_R FILLER_133_98 ();
 DECAPx4_ASAP7_75t_R FILLER_133_112 ();
 DECAPx10_ASAP7_75t_R FILLER_133_171 ();
 FILLER_ASAP7_75t_R FILLER_133_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_195 ();
 FILLER_ASAP7_75t_R FILLER_133_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_204 ();
 DECAPx6_ASAP7_75t_R FILLER_133_212 ();
 FILLER_ASAP7_75t_R FILLER_133_248 ();
 FILLER_ASAP7_75t_R FILLER_133_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_266 ();
 DECAPx2_ASAP7_75t_R FILLER_133_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_276 ();
 DECAPx4_ASAP7_75t_R FILLER_133_329 ();
 DECAPx2_ASAP7_75t_R FILLER_133_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_354 ();
 DECAPx2_ASAP7_75t_R FILLER_133_361 ();
 FILLER_ASAP7_75t_R FILLER_133_375 ();
 DECAPx10_ASAP7_75t_R FILLER_133_383 ();
 DECAPx1_ASAP7_75t_R FILLER_133_405 ();
 DECAPx1_ASAP7_75t_R FILLER_133_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_429 ();
 FILLER_ASAP7_75t_R FILLER_133_459 ();
 FILLER_ASAP7_75t_R FILLER_133_474 ();
 DECAPx1_ASAP7_75t_R FILLER_133_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_493 ();
 DECAPx4_ASAP7_75t_R FILLER_133_533 ();
 FILLER_ASAP7_75t_R FILLER_133_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_576 ();
 DECAPx4_ASAP7_75t_R FILLER_133_580 ();
 DECAPx2_ASAP7_75t_R FILLER_133_616 ();
 FILLER_ASAP7_75t_R FILLER_133_622 ();
 DECAPx4_ASAP7_75t_R FILLER_133_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_637 ();
 DECAPx6_ASAP7_75t_R FILLER_133_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_655 ();
 DECAPx4_ASAP7_75t_R FILLER_133_662 ();
 DECAPx10_ASAP7_75t_R FILLER_133_698 ();
 DECAPx2_ASAP7_75t_R FILLER_133_720 ();
 FILLER_ASAP7_75t_R FILLER_133_726 ();
 DECAPx4_ASAP7_75t_R FILLER_133_737 ();
 FILLER_ASAP7_75t_R FILLER_133_747 ();
 DECAPx6_ASAP7_75t_R FILLER_133_778 ();
 DECAPx1_ASAP7_75t_R FILLER_133_792 ();
 DECAPx6_ASAP7_75t_R FILLER_133_805 ();
 DECAPx1_ASAP7_75t_R FILLER_133_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_823 ();
 FILLER_ASAP7_75t_R FILLER_133_827 ();
 DECAPx2_ASAP7_75t_R FILLER_133_838 ();
 FILLER_ASAP7_75t_R FILLER_133_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_846 ();
 DECAPx10_ASAP7_75t_R FILLER_133_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_882 ();
 DECAPx6_ASAP7_75t_R FILLER_133_889 ();
 FILLER_ASAP7_75t_R FILLER_133_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_905 ();
 DECAPx2_ASAP7_75t_R FILLER_133_916 ();
 FILLER_ASAP7_75t_R FILLER_133_922 ();
 DECAPx2_ASAP7_75t_R FILLER_133_926 ();
 FILLER_ASAP7_75t_R FILLER_133_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_934 ();
 DECAPx2_ASAP7_75t_R FILLER_133_941 ();
 DECAPx4_ASAP7_75t_R FILLER_133_966 ();
 FILLER_ASAP7_75t_R FILLER_133_999 ();
 FILLER_ASAP7_75t_R FILLER_133_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1021 ();
 FILLER_ASAP7_75t_R FILLER_133_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1068 ();
 FILLER_ASAP7_75t_R FILLER_133_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1086 ();
 FILLER_ASAP7_75t_R FILLER_133_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1131 ();
 FILLER_ASAP7_75t_R FILLER_133_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1143 ();
 FILLER_ASAP7_75t_R FILLER_133_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1199 ();
 FILLER_ASAP7_75t_R FILLER_133_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1227 ();
 FILLER_ASAP7_75t_R FILLER_133_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1251 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1280 ();
 FILLER_ASAP7_75t_R FILLER_133_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1304 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1326 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1342 ();
 FILLER_ASAP7_75t_R FILLER_133_1368 ();
 FILLER_ASAP7_75t_R FILLER_133_1377 ();
 DECAPx4_ASAP7_75t_R FILLER_134_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_12 ();
 DECAPx2_ASAP7_75t_R FILLER_134_19 ();
 DECAPx2_ASAP7_75t_R FILLER_134_31 ();
 FILLER_ASAP7_75t_R FILLER_134_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_39 ();
 DECAPx2_ASAP7_75t_R FILLER_134_46 ();
 FILLER_ASAP7_75t_R FILLER_134_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_57 ();
 DECAPx10_ASAP7_75t_R FILLER_134_84 ();
 DECAPx4_ASAP7_75t_R FILLER_134_106 ();
 DECAPx1_ASAP7_75t_R FILLER_134_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_128 ();
 DECAPx1_ASAP7_75t_R FILLER_134_135 ();
 DECAPx6_ASAP7_75t_R FILLER_134_165 ();
 FILLER_ASAP7_75t_R FILLER_134_179 ();
 DECAPx6_ASAP7_75t_R FILLER_134_203 ();
 DECAPx1_ASAP7_75t_R FILLER_134_217 ();
 DECAPx1_ASAP7_75t_R FILLER_134_243 ();
 FILLER_ASAP7_75t_R FILLER_134_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_304 ();
 DECAPx2_ASAP7_75t_R FILLER_134_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_317 ();
 DECAPx10_ASAP7_75t_R FILLER_134_321 ();
 DECAPx1_ASAP7_75t_R FILLER_134_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_392 ();
 DECAPx10_ASAP7_75t_R FILLER_134_410 ();
 FILLER_ASAP7_75t_R FILLER_134_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_434 ();
 DECAPx1_ASAP7_75t_R FILLER_134_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_446 ();
 DECAPx4_ASAP7_75t_R FILLER_134_450 ();
 FILLER_ASAP7_75t_R FILLER_134_460 ();
 DECAPx1_ASAP7_75t_R FILLER_134_490 ();
 DECAPx2_ASAP7_75t_R FILLER_134_501 ();
 FILLER_ASAP7_75t_R FILLER_134_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_509 ();
 FILLER_ASAP7_75t_R FILLER_134_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_515 ();
 DECAPx2_ASAP7_75t_R FILLER_134_525 ();
 FILLER_ASAP7_75t_R FILLER_134_531 ();
 DECAPx10_ASAP7_75t_R FILLER_134_539 ();
 DECAPx4_ASAP7_75t_R FILLER_134_561 ();
 DECAPx6_ASAP7_75t_R FILLER_134_584 ();
 DECAPx2_ASAP7_75t_R FILLER_134_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_604 ();
 DECAPx4_ASAP7_75t_R FILLER_134_608 ();
 FILLER_ASAP7_75t_R FILLER_134_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_620 ();
 DECAPx6_ASAP7_75t_R FILLER_134_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_648 ();
 DECAPx4_ASAP7_75t_R FILLER_134_681 ();
 FILLER_ASAP7_75t_R FILLER_134_691 ();
 DECAPx2_ASAP7_75t_R FILLER_134_699 ();
 FILLER_ASAP7_75t_R FILLER_134_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_710 ();
 DECAPx10_ASAP7_75t_R FILLER_134_715 ();
 DECAPx10_ASAP7_75t_R FILLER_134_737 ();
 DECAPx2_ASAP7_75t_R FILLER_134_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_797 ();
 DECAPx2_ASAP7_75t_R FILLER_134_811 ();
 DECAPx4_ASAP7_75t_R FILLER_134_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_849 ();
 DECAPx4_ASAP7_75t_R FILLER_134_859 ();
 FILLER_ASAP7_75t_R FILLER_134_869 ();
 DECAPx2_ASAP7_75t_R FILLER_134_889 ();
 FILLER_ASAP7_75t_R FILLER_134_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_897 ();
 FILLER_ASAP7_75t_R FILLER_134_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_909 ();
 DECAPx2_ASAP7_75t_R FILLER_134_928 ();
 DECAPx2_ASAP7_75t_R FILLER_134_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_946 ();
 FILLER_ASAP7_75t_R FILLER_134_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_955 ();
 DECAPx1_ASAP7_75t_R FILLER_134_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_969 ();
 DECAPx10_ASAP7_75t_R FILLER_134_985 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1038 ();
 FILLER_ASAP7_75t_R FILLER_134_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1095 ();
 FILLER_ASAP7_75t_R FILLER_134_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1117 ();
 FILLER_ASAP7_75t_R FILLER_134_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1125 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1237 ();
 FILLER_ASAP7_75t_R FILLER_134_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1319 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1329 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1333 ();
 FILLER_ASAP7_75t_R FILLER_134_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1382 ();
 FILLER_ASAP7_75t_R FILLER_134_1394 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1399 ();
 DECAPx2_ASAP7_75t_R FILLER_135_2 ();
 FILLER_ASAP7_75t_R FILLER_135_8 ();
 FILLER_ASAP7_75t_R FILLER_135_39 ();
 DECAPx6_ASAP7_75t_R FILLER_135_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_104 ();
 DECAPx2_ASAP7_75t_R FILLER_135_118 ();
 DECAPx4_ASAP7_75t_R FILLER_135_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_153 ();
 DECAPx6_ASAP7_75t_R FILLER_135_157 ();
 DECAPx2_ASAP7_75t_R FILLER_135_171 ();
 DECAPx1_ASAP7_75t_R FILLER_135_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_193 ();
 DECAPx2_ASAP7_75t_R FILLER_135_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_212 ();
 DECAPx4_ASAP7_75t_R FILLER_135_244 ();
 DECAPx6_ASAP7_75t_R FILLER_135_270 ();
 FILLER_ASAP7_75t_R FILLER_135_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_286 ();
 FILLER_ASAP7_75t_R FILLER_135_290 ();
 DECAPx10_ASAP7_75t_R FILLER_135_298 ();
 DECAPx2_ASAP7_75t_R FILLER_135_320 ();
 DECAPx2_ASAP7_75t_R FILLER_135_329 ();
 DECAPx2_ASAP7_75t_R FILLER_135_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_350 ();
 FILLER_ASAP7_75t_R FILLER_135_357 ();
 DECAPx4_ASAP7_75t_R FILLER_135_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_417 ();
 DECAPx6_ASAP7_75t_R FILLER_135_431 ();
 FILLER_ASAP7_75t_R FILLER_135_445 ();
 DECAPx10_ASAP7_75t_R FILLER_135_473 ();
 DECAPx10_ASAP7_75t_R FILLER_135_495 ();
 DECAPx4_ASAP7_75t_R FILLER_135_517 ();
 FILLER_ASAP7_75t_R FILLER_135_527 ();
 DECAPx2_ASAP7_75t_R FILLER_135_545 ();
 FILLER_ASAP7_75t_R FILLER_135_551 ();
 DECAPx1_ASAP7_75t_R FILLER_135_575 ();
 DECAPx1_ASAP7_75t_R FILLER_135_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_620 ();
 DECAPx1_ASAP7_75t_R FILLER_135_666 ();
 DECAPx2_ASAP7_75t_R FILLER_135_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_691 ();
 DECAPx1_ASAP7_75t_R FILLER_135_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_722 ();
 DECAPx2_ASAP7_75t_R FILLER_135_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_744 ();
 FILLER_ASAP7_75t_R FILLER_135_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_754 ();
 DECAPx4_ASAP7_75t_R FILLER_135_762 ();
 FILLER_ASAP7_75t_R FILLER_135_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_829 ();
 DECAPx4_ASAP7_75t_R FILLER_135_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_849 ();
 DECAPx10_ASAP7_75t_R FILLER_135_859 ();
 DECAPx2_ASAP7_75t_R FILLER_135_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_887 ();
 DECAPx2_ASAP7_75t_R FILLER_135_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_900 ();
 DECAPx6_ASAP7_75t_R FILLER_135_907 ();
 FILLER_ASAP7_75t_R FILLER_135_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_923 ();
 DECAPx1_ASAP7_75t_R FILLER_135_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_936 ();
 DECAPx10_ASAP7_75t_R FILLER_135_945 ();
 DECAPx6_ASAP7_75t_R FILLER_135_967 ();
 DECAPx6_ASAP7_75t_R FILLER_135_984 ();
 DECAPx1_ASAP7_75t_R FILLER_135_998 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1078 ();
 FILLER_ASAP7_75t_R FILLER_135_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1164 ();
 FILLER_ASAP7_75t_R FILLER_135_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1220 ();
 FILLER_ASAP7_75t_R FILLER_135_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1274 ();
 FILLER_ASAP7_75t_R FILLER_135_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1289 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1367 ();
 FILLER_ASAP7_75t_R FILLER_135_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1388 ();
 FILLER_ASAP7_75t_R FILLER_135_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1404 ();
 DECAPx4_ASAP7_75t_R FILLER_136_2 ();
 FILLER_ASAP7_75t_R FILLER_136_12 ();
 DECAPx1_ASAP7_75t_R FILLER_136_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_24 ();
 DECAPx4_ASAP7_75t_R FILLER_136_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_70 ();
 FILLER_ASAP7_75t_R FILLER_136_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_82 ();
 FILLER_ASAP7_75t_R FILLER_136_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_101 ();
 DECAPx2_ASAP7_75t_R FILLER_136_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_162 ();
 DECAPx2_ASAP7_75t_R FILLER_136_175 ();
 FILLER_ASAP7_75t_R FILLER_136_181 ();
 DECAPx4_ASAP7_75t_R FILLER_136_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_221 ();
 DECAPx10_ASAP7_75t_R FILLER_136_236 ();
 DECAPx4_ASAP7_75t_R FILLER_136_258 ();
 FILLER_ASAP7_75t_R FILLER_136_268 ();
 DECAPx2_ASAP7_75t_R FILLER_136_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_292 ();
 DECAPx4_ASAP7_75t_R FILLER_136_296 ();
 FILLER_ASAP7_75t_R FILLER_136_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_308 ();
 DECAPx1_ASAP7_75t_R FILLER_136_316 ();
 FILLER_ASAP7_75t_R FILLER_136_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_357 ();
 DECAPx1_ASAP7_75t_R FILLER_136_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_390 ();
 DECAPx6_ASAP7_75t_R FILLER_136_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_414 ();
 DECAPx2_ASAP7_75t_R FILLER_136_441 ();
 FILLER_ASAP7_75t_R FILLER_136_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_461 ();
 DECAPx2_ASAP7_75t_R FILLER_136_470 ();
 FILLER_ASAP7_75t_R FILLER_136_476 ();
 DECAPx4_ASAP7_75t_R FILLER_136_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_503 ();
 DECAPx2_ASAP7_75t_R FILLER_136_510 ();
 FILLER_ASAP7_75t_R FILLER_136_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_518 ();
 FILLER_ASAP7_75t_R FILLER_136_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_530 ();
 DECAPx6_ASAP7_75t_R FILLER_136_543 ();
 DECAPx1_ASAP7_75t_R FILLER_136_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_561 ();
 DECAPx4_ASAP7_75t_R FILLER_136_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_608 ();
 DECAPx4_ASAP7_75t_R FILLER_136_629 ();
 DECAPx10_ASAP7_75t_R FILLER_136_642 ();
 DECAPx6_ASAP7_75t_R FILLER_136_664 ();
 DECAPx2_ASAP7_75t_R FILLER_136_678 ();
 FILLER_ASAP7_75t_R FILLER_136_690 ();
 DECAPx10_ASAP7_75t_R FILLER_136_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_757 ();
 DECAPx1_ASAP7_75t_R FILLER_136_764 ();
 DECAPx6_ASAP7_75t_R FILLER_136_775 ();
 FILLER_ASAP7_75t_R FILLER_136_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_791 ();
 DECAPx1_ASAP7_75t_R FILLER_136_802 ();
 DECAPx10_ASAP7_75t_R FILLER_136_809 ();
 FILLER_ASAP7_75t_R FILLER_136_831 ();
 DECAPx4_ASAP7_75t_R FILLER_136_853 ();
 FILLER_ASAP7_75t_R FILLER_136_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_865 ();
 DECAPx4_ASAP7_75t_R FILLER_136_878 ();
 DECAPx10_ASAP7_75t_R FILLER_136_902 ();
 DECAPx4_ASAP7_75t_R FILLER_136_932 ();
 DECAPx10_ASAP7_75t_R FILLER_136_948 ();
 DECAPx2_ASAP7_75t_R FILLER_136_970 ();
 DECAPx10_ASAP7_75t_R FILLER_136_996 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1018 ();
 FILLER_ASAP7_75t_R FILLER_136_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1045 ();
 FILLER_ASAP7_75t_R FILLER_136_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1069 ();
 FILLER_ASAP7_75t_R FILLER_136_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1080 ();
 FILLER_ASAP7_75t_R FILLER_136_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1186 ();
 FILLER_ASAP7_75t_R FILLER_136_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1222 ();
 FILLER_ASAP7_75t_R FILLER_136_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1257 ();
 FILLER_ASAP7_75t_R FILLER_136_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1281 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1297 ();
 FILLER_ASAP7_75t_R FILLER_136_1303 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1317 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1342 ();
 FILLER_ASAP7_75t_R FILLER_136_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1365 ();
 FILLER_ASAP7_75t_R FILLER_136_1375 ();
 FILLER_ASAP7_75t_R FILLER_136_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1396 ();
 FILLER_ASAP7_75t_R FILLER_136_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1404 ();
 DECAPx2_ASAP7_75t_R FILLER_137_2 ();
 FILLER_ASAP7_75t_R FILLER_137_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_10 ();
 DECAPx2_ASAP7_75t_R FILLER_137_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_52 ();
 DECAPx2_ASAP7_75t_R FILLER_137_56 ();
 DECAPx6_ASAP7_75t_R FILLER_137_65 ();
 FILLER_ASAP7_75t_R FILLER_137_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_108 ();
 DECAPx1_ASAP7_75t_R FILLER_137_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_119 ();
 DECAPx1_ASAP7_75t_R FILLER_137_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_159 ();
 DECAPx1_ASAP7_75t_R FILLER_137_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_190 ();
 DECAPx10_ASAP7_75t_R FILLER_137_211 ();
 DECAPx2_ASAP7_75t_R FILLER_137_233 ();
 FILLER_ASAP7_75t_R FILLER_137_239 ();
 DECAPx1_ASAP7_75t_R FILLER_137_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_267 ();
 DECAPx2_ASAP7_75t_R FILLER_137_294 ();
 FILLER_ASAP7_75t_R FILLER_137_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_302 ();
 DECAPx1_ASAP7_75t_R FILLER_137_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_355 ();
 DECAPx2_ASAP7_75t_R FILLER_137_394 ();
 FILLER_ASAP7_75t_R FILLER_137_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_402 ();
 DECAPx4_ASAP7_75t_R FILLER_137_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_423 ();
 DECAPx2_ASAP7_75t_R FILLER_137_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_441 ();
 DECAPx10_ASAP7_75t_R FILLER_137_449 ();
 DECAPx1_ASAP7_75t_R FILLER_137_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_475 ();
 DECAPx6_ASAP7_75t_R FILLER_137_550 ();
 FILLER_ASAP7_75t_R FILLER_137_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_566 ();
 DECAPx4_ASAP7_75t_R FILLER_137_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_583 ();
 DECAPx10_ASAP7_75t_R FILLER_137_587 ();
 DECAPx6_ASAP7_75t_R FILLER_137_609 ();
 DECAPx1_ASAP7_75t_R FILLER_137_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_627 ();
 DECAPx6_ASAP7_75t_R FILLER_137_638 ();
 DECAPx1_ASAP7_75t_R FILLER_137_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_656 ();
 DECAPx6_ASAP7_75t_R FILLER_137_709 ();
 FILLER_ASAP7_75t_R FILLER_137_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_725 ();
 DECAPx4_ASAP7_75t_R FILLER_137_736 ();
 DECAPx4_ASAP7_75t_R FILLER_137_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_759 ();
 DECAPx6_ASAP7_75t_R FILLER_137_792 ();
 FILLER_ASAP7_75t_R FILLER_137_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_808 ();
 DECAPx6_ASAP7_75t_R FILLER_137_828 ();
 FILLER_ASAP7_75t_R FILLER_137_842 ();
 FILLER_ASAP7_75t_R FILLER_137_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_852 ();
 DECAPx10_ASAP7_75t_R FILLER_137_863 ();
 FILLER_ASAP7_75t_R FILLER_137_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_887 ();
 DECAPx1_ASAP7_75t_R FILLER_137_896 ();
 DECAPx1_ASAP7_75t_R FILLER_137_910 ();
 DECAPx10_ASAP7_75t_R FILLER_137_926 ();
 FILLER_ASAP7_75t_R FILLER_137_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_956 ();
 DECAPx4_ASAP7_75t_R FILLER_137_970 ();
 FILLER_ASAP7_75t_R FILLER_137_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_982 ();
 DECAPx2_ASAP7_75t_R FILLER_137_989 ();
 FILLER_ASAP7_75t_R FILLER_137_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_997 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1020 ();
 FILLER_ASAP7_75t_R FILLER_137_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1044 ();
 FILLER_ASAP7_75t_R FILLER_137_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1100 ();
 FILLER_ASAP7_75t_R FILLER_137_1110 ();
 FILLER_ASAP7_75t_R FILLER_137_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1152 ();
 FILLER_ASAP7_75t_R FILLER_137_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1186 ();
 FILLER_ASAP7_75t_R FILLER_137_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1238 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1312 ();
 FILLER_ASAP7_75t_R FILLER_137_1318 ();
 FILLER_ASAP7_75t_R FILLER_137_1326 ();
 FILLER_ASAP7_75t_R FILLER_137_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1358 ();
 FILLER_ASAP7_75t_R FILLER_137_1368 ();
 DECAPx10_ASAP7_75t_R FILLER_138_2 ();
 FILLER_ASAP7_75t_R FILLER_138_24 ();
 DECAPx4_ASAP7_75t_R FILLER_138_29 ();
 FILLER_ASAP7_75t_R FILLER_138_39 ();
 DECAPx1_ASAP7_75t_R FILLER_138_48 ();
 DECAPx2_ASAP7_75t_R FILLER_138_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_64 ();
 DECAPx6_ASAP7_75t_R FILLER_138_68 ();
 DECAPx1_ASAP7_75t_R FILLER_138_82 ();
 DECAPx1_ASAP7_75t_R FILLER_138_92 ();
 DECAPx10_ASAP7_75t_R FILLER_138_99 ();
 DECAPx1_ASAP7_75t_R FILLER_138_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_125 ();
 DECAPx6_ASAP7_75t_R FILLER_138_133 ();
 FILLER_ASAP7_75t_R FILLER_138_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_156 ();
 DECAPx4_ASAP7_75t_R FILLER_138_164 ();
 DECAPx1_ASAP7_75t_R FILLER_138_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_181 ();
 FILLER_ASAP7_75t_R FILLER_138_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_187 ();
 DECAPx6_ASAP7_75t_R FILLER_138_196 ();
 FILLER_ASAP7_75t_R FILLER_138_210 ();
 DECAPx2_ASAP7_75t_R FILLER_138_230 ();
 DECAPx1_ASAP7_75t_R FILLER_138_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_319 ();
 DECAPx6_ASAP7_75t_R FILLER_138_323 ();
 FILLER_ASAP7_75t_R FILLER_138_337 ();
 DECAPx1_ASAP7_75t_R FILLER_138_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_369 ();
 DECAPx2_ASAP7_75t_R FILLER_138_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_382 ();
 DECAPx1_ASAP7_75t_R FILLER_138_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_423 ();
 FILLER_ASAP7_75t_R FILLER_138_434 ();
 DECAPx4_ASAP7_75t_R FILLER_138_468 ();
 FILLER_ASAP7_75t_R FILLER_138_478 ();
 DECAPx10_ASAP7_75t_R FILLER_138_486 ();
 DECAPx6_ASAP7_75t_R FILLER_138_508 ();
 DECAPx6_ASAP7_75t_R FILLER_138_526 ();
 DECAPx10_ASAP7_75t_R FILLER_138_558 ();
 FILLER_ASAP7_75t_R FILLER_138_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_582 ();
 DECAPx4_ASAP7_75t_R FILLER_138_593 ();
 DECAPx2_ASAP7_75t_R FILLER_138_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_619 ();
 DECAPx6_ASAP7_75t_R FILLER_138_626 ();
 DECAPx2_ASAP7_75t_R FILLER_138_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_646 ();
 DECAPx10_ASAP7_75t_R FILLER_138_661 ();
 DECAPx2_ASAP7_75t_R FILLER_138_689 ();
 FILLER_ASAP7_75t_R FILLER_138_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_697 ();
 DECAPx10_ASAP7_75t_R FILLER_138_701 ();
 DECAPx10_ASAP7_75t_R FILLER_138_723 ();
 DECAPx10_ASAP7_75t_R FILLER_138_745 ();
 DECAPx1_ASAP7_75t_R FILLER_138_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_771 ();
 FILLER_ASAP7_75t_R FILLER_138_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_784 ();
 FILLER_ASAP7_75t_R FILLER_138_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_817 ();
 FILLER_ASAP7_75t_R FILLER_138_824 ();
 DECAPx6_ASAP7_75t_R FILLER_138_834 ();
 DECAPx2_ASAP7_75t_R FILLER_138_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_854 ();
 DECAPx10_ASAP7_75t_R FILLER_138_868 ();
 DECAPx4_ASAP7_75t_R FILLER_138_890 ();
 DECAPx4_ASAP7_75t_R FILLER_138_906 ();
 FILLER_ASAP7_75t_R FILLER_138_916 ();
 DECAPx10_ASAP7_75t_R FILLER_138_924 ();
 DECAPx2_ASAP7_75t_R FILLER_138_946 ();
 FILLER_ASAP7_75t_R FILLER_138_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_954 ();
 DECAPx1_ASAP7_75t_R FILLER_138_962 ();
 DECAPx10_ASAP7_75t_R FILLER_138_973 ();
 DECAPx6_ASAP7_75t_R FILLER_138_995 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1013 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1184 ();
 FILLER_ASAP7_75t_R FILLER_138_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1199 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1221 ();
 FILLER_ASAP7_75t_R FILLER_138_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1252 ();
 FILLER_ASAP7_75t_R FILLER_138_1263 ();
 FILLER_ASAP7_75t_R FILLER_138_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1308 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1336 ();
 FILLER_ASAP7_75t_R FILLER_138_1366 ();
 FILLER_ASAP7_75t_R FILLER_138_1384 ();
 FILLER_ASAP7_75t_R FILLER_138_1394 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_139_2 ();
 DECAPx6_ASAP7_75t_R FILLER_139_24 ();
 DECAPx4_ASAP7_75t_R FILLER_139_64 ();
 DECAPx1_ASAP7_75t_R FILLER_139_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_84 ();
 DECAPx2_ASAP7_75t_R FILLER_139_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_122 ();
 DECAPx2_ASAP7_75t_R FILLER_139_149 ();
 DECAPx6_ASAP7_75t_R FILLER_139_181 ();
 FILLER_ASAP7_75t_R FILLER_139_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_197 ();
 DECAPx6_ASAP7_75t_R FILLER_139_204 ();
 FILLER_ASAP7_75t_R FILLER_139_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_220 ();
 FILLER_ASAP7_75t_R FILLER_139_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_247 ();
 DECAPx4_ASAP7_75t_R FILLER_139_261 ();
 FILLER_ASAP7_75t_R FILLER_139_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_287 ();
 DECAPx4_ASAP7_75t_R FILLER_139_291 ();
 FILLER_ASAP7_75t_R FILLER_139_301 ();
 DECAPx10_ASAP7_75t_R FILLER_139_329 ();
 FILLER_ASAP7_75t_R FILLER_139_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_353 ();
 DECAPx2_ASAP7_75t_R FILLER_139_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_363 ();
 FILLER_ASAP7_75t_R FILLER_139_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_372 ();
 DECAPx10_ASAP7_75t_R FILLER_139_413 ();
 DECAPx2_ASAP7_75t_R FILLER_139_435 ();
 FILLER_ASAP7_75t_R FILLER_139_441 ();
 DECAPx2_ASAP7_75t_R FILLER_139_449 ();
 FILLER_ASAP7_75t_R FILLER_139_458 ();
 DECAPx1_ASAP7_75t_R FILLER_139_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_496 ();
 DECAPx10_ASAP7_75t_R FILLER_139_529 ();
 FILLER_ASAP7_75t_R FILLER_139_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_553 ();
 DECAPx4_ASAP7_75t_R FILLER_139_582 ();
 DECAPx1_ASAP7_75t_R FILLER_139_598 ();
 DECAPx6_ASAP7_75t_R FILLER_139_605 ();
 DECAPx1_ASAP7_75t_R FILLER_139_645 ();
 DECAPx10_ASAP7_75t_R FILLER_139_689 ();
 DECAPx6_ASAP7_75t_R FILLER_139_711 ();
 DECAPx1_ASAP7_75t_R FILLER_139_725 ();
 DECAPx2_ASAP7_75t_R FILLER_139_736 ();
 FILLER_ASAP7_75t_R FILLER_139_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_744 ();
 FILLER_ASAP7_75t_R FILLER_139_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_757 ();
 DECAPx10_ASAP7_75t_R FILLER_139_761 ();
 DECAPx10_ASAP7_75t_R FILLER_139_783 ();
 DECAPx2_ASAP7_75t_R FILLER_139_805 ();
 FILLER_ASAP7_75t_R FILLER_139_811 ();
 FILLER_ASAP7_75t_R FILLER_139_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_845 ();
 DECAPx2_ASAP7_75t_R FILLER_139_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_857 ();
 DECAPx2_ASAP7_75t_R FILLER_139_866 ();
 DECAPx2_ASAP7_75t_R FILLER_139_885 ();
 DECAPx10_ASAP7_75t_R FILLER_139_897 ();
 DECAPx1_ASAP7_75t_R FILLER_139_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_923 ();
 DECAPx2_ASAP7_75t_R FILLER_139_926 ();
 FILLER_ASAP7_75t_R FILLER_139_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_934 ();
 DECAPx10_ASAP7_75t_R FILLER_139_949 ();
 DECAPx4_ASAP7_75t_R FILLER_139_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_981 ();
 DECAPx1_ASAP7_75t_R FILLER_139_999 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1040 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1239 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1293 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_140_2 ();
 DECAPx1_ASAP7_75t_R FILLER_140_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_20 ();
 DECAPx1_ASAP7_75t_R FILLER_140_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_51 ();
 DECAPx2_ASAP7_75t_R FILLER_140_55 ();
 FILLER_ASAP7_75t_R FILLER_140_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_137 ();
 FILLER_ASAP7_75t_R FILLER_140_141 ();
 DECAPx2_ASAP7_75t_R FILLER_140_150 ();
 FILLER_ASAP7_75t_R FILLER_140_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_158 ();
 DECAPx1_ASAP7_75t_R FILLER_140_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_169 ();
 FILLER_ASAP7_75t_R FILLER_140_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_182 ();
 DECAPx2_ASAP7_75t_R FILLER_140_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_203 ();
 FILLER_ASAP7_75t_R FILLER_140_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_212 ();
 DECAPx1_ASAP7_75t_R FILLER_140_227 ();
 DECAPx6_ASAP7_75t_R FILLER_140_245 ();
 FILLER_ASAP7_75t_R FILLER_140_259 ();
 DECAPx4_ASAP7_75t_R FILLER_140_279 ();
 FILLER_ASAP7_75t_R FILLER_140_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_291 ();
 FILLER_ASAP7_75t_R FILLER_140_302 ();
 DECAPx2_ASAP7_75t_R FILLER_140_311 ();
 FILLER_ASAP7_75t_R FILLER_140_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_322 ();
 DECAPx2_ASAP7_75t_R FILLER_140_329 ();
 FILLER_ASAP7_75t_R FILLER_140_335 ();
 DECAPx2_ASAP7_75t_R FILLER_140_343 ();
 FILLER_ASAP7_75t_R FILLER_140_349 ();
 DECAPx2_ASAP7_75t_R FILLER_140_363 ();
 FILLER_ASAP7_75t_R FILLER_140_369 ();
 FILLER_ASAP7_75t_R FILLER_140_379 ();
 DECAPx4_ASAP7_75t_R FILLER_140_409 ();
 FILLER_ASAP7_75t_R FILLER_140_419 ();
 FILLER_ASAP7_75t_R FILLER_140_456 ();
 DECAPx4_ASAP7_75t_R FILLER_140_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_474 ();
 DECAPx6_ASAP7_75t_R FILLER_140_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_492 ();
 DECAPx4_ASAP7_75t_R FILLER_140_509 ();
 FILLER_ASAP7_75t_R FILLER_140_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_521 ();
 DECAPx6_ASAP7_75t_R FILLER_140_548 ();
 DECAPx2_ASAP7_75t_R FILLER_140_562 ();
 DECAPx1_ASAP7_75t_R FILLER_140_578 ();
 DECAPx2_ASAP7_75t_R FILLER_140_614 ();
 FILLER_ASAP7_75t_R FILLER_140_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_622 ();
 DECAPx1_ASAP7_75t_R FILLER_140_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_633 ();
 DECAPx6_ASAP7_75t_R FILLER_140_637 ();
 DECAPx4_ASAP7_75t_R FILLER_140_667 ();
 FILLER_ASAP7_75t_R FILLER_140_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_679 ();
 DECAPx6_ASAP7_75t_R FILLER_140_712 ();
 DECAPx4_ASAP7_75t_R FILLER_140_734 ();
 DECAPx10_ASAP7_75t_R FILLER_140_752 ();
 DECAPx6_ASAP7_75t_R FILLER_140_774 ();
 DECAPx1_ASAP7_75t_R FILLER_140_788 ();
 DECAPx6_ASAP7_75t_R FILLER_140_802 ();
 FILLER_ASAP7_75t_R FILLER_140_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_836 ();
 DECAPx6_ASAP7_75t_R FILLER_140_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_869 ();
 DECAPx6_ASAP7_75t_R FILLER_140_886 ();
 DECAPx2_ASAP7_75t_R FILLER_140_908 ();
 FILLER_ASAP7_75t_R FILLER_140_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_916 ();
 DECAPx2_ASAP7_75t_R FILLER_140_927 ();
 DECAPx6_ASAP7_75t_R FILLER_140_951 ();
 FILLER_ASAP7_75t_R FILLER_140_965 ();
 DECAPx10_ASAP7_75t_R FILLER_140_973 ();
 DECAPx10_ASAP7_75t_R FILLER_140_995 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1049 ();
 FILLER_ASAP7_75t_R FILLER_140_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1153 ();
 FILLER_ASAP7_75t_R FILLER_140_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1198 ();
 FILLER_ASAP7_75t_R FILLER_140_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1251 ();
 FILLER_ASAP7_75t_R FILLER_140_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1269 ();
 FILLER_ASAP7_75t_R FILLER_140_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1345 ();
 FILLER_ASAP7_75t_R FILLER_140_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1396 ();
 FILLER_ASAP7_75t_R FILLER_140_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_141_2 ();
 DECAPx1_ASAP7_75t_R FILLER_141_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_20 ();
 FILLER_ASAP7_75t_R FILLER_141_39 ();
 DECAPx1_ASAP7_75t_R FILLER_141_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_97 ();
 DECAPx10_ASAP7_75t_R FILLER_141_101 ();
 DECAPx6_ASAP7_75t_R FILLER_141_123 ();
 DECAPx1_ASAP7_75t_R FILLER_141_137 ();
 DECAPx2_ASAP7_75t_R FILLER_141_167 ();
 FILLER_ASAP7_75t_R FILLER_141_173 ();
 FILLER_ASAP7_75t_R FILLER_141_181 ();
 DECAPx2_ASAP7_75t_R FILLER_141_207 ();
 DECAPx1_ASAP7_75t_R FILLER_141_227 ();
 DECAPx10_ASAP7_75t_R FILLER_141_241 ();
 DECAPx2_ASAP7_75t_R FILLER_141_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_269 ();
 DECAPx2_ASAP7_75t_R FILLER_141_286 ();
 FILLER_ASAP7_75t_R FILLER_141_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_294 ();
 DECAPx2_ASAP7_75t_R FILLER_141_308 ();
 FILLER_ASAP7_75t_R FILLER_141_342 ();
 FILLER_ASAP7_75t_R FILLER_141_373 ();
 DECAPx1_ASAP7_75t_R FILLER_141_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_419 ();
 FILLER_ASAP7_75t_R FILLER_141_464 ();
 DECAPx1_ASAP7_75t_R FILLER_141_476 ();
 DECAPx2_ASAP7_75t_R FILLER_141_498 ();
 FILLER_ASAP7_75t_R FILLER_141_504 ();
 FILLER_ASAP7_75t_R FILLER_141_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_530 ();
 DECAPx4_ASAP7_75t_R FILLER_141_563 ();
 FILLER_ASAP7_75t_R FILLER_141_573 ();
 FILLER_ASAP7_75t_R FILLER_141_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_612 ();
 DECAPx4_ASAP7_75t_R FILLER_141_651 ();
 DECAPx10_ASAP7_75t_R FILLER_141_687 ();
 DECAPx10_ASAP7_75t_R FILLER_141_709 ();
 DECAPx10_ASAP7_75t_R FILLER_141_731 ();
 DECAPx6_ASAP7_75t_R FILLER_141_753 ();
 FILLER_ASAP7_75t_R FILLER_141_786 ();
 DECAPx4_ASAP7_75t_R FILLER_141_810 ();
 DECAPx10_ASAP7_75t_R FILLER_141_832 ();
 FILLER_ASAP7_75t_R FILLER_141_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_874 ();
 DECAPx10_ASAP7_75t_R FILLER_141_881 ();
 DECAPx6_ASAP7_75t_R FILLER_141_903 ();
 DECAPx2_ASAP7_75t_R FILLER_141_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_923 ();
 DECAPx4_ASAP7_75t_R FILLER_141_926 ();
 FILLER_ASAP7_75t_R FILLER_141_936 ();
 DECAPx4_ASAP7_75t_R FILLER_141_945 ();
 FILLER_ASAP7_75t_R FILLER_141_955 ();
 DECAPx4_ASAP7_75t_R FILLER_141_963 ();
 FILLER_ASAP7_75t_R FILLER_141_973 ();
 FILLER_ASAP7_75t_R FILLER_141_981 ();
 DECAPx2_ASAP7_75t_R FILLER_141_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1010 ();
 FILLER_ASAP7_75t_R FILLER_141_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1078 ();
 FILLER_ASAP7_75t_R FILLER_141_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1115 ();
 FILLER_ASAP7_75t_R FILLER_141_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1148 ();
 FILLER_ASAP7_75t_R FILLER_141_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1250 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1272 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1288 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1308 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1341 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1351 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1374 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1395 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1399 ();
 DECAPx2_ASAP7_75t_R FILLER_142_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_8 ();
 FILLER_ASAP7_75t_R FILLER_142_47 ();
 DECAPx1_ASAP7_75t_R FILLER_142_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_59 ();
 DECAPx1_ASAP7_75t_R FILLER_142_63 ();
 DECAPx2_ASAP7_75t_R FILLER_142_73 ();
 FILLER_ASAP7_75t_R FILLER_142_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_81 ();
 DECAPx10_ASAP7_75t_R FILLER_142_85 ();
 FILLER_ASAP7_75t_R FILLER_142_120 ();
 DECAPx10_ASAP7_75t_R FILLER_142_125 ();
 FILLER_ASAP7_75t_R FILLER_142_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_155 ();
 DECAPx6_ASAP7_75t_R FILLER_142_159 ();
 FILLER_ASAP7_75t_R FILLER_142_173 ();
 DECAPx2_ASAP7_75t_R FILLER_142_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_187 ();
 DECAPx4_ASAP7_75t_R FILLER_142_200 ();
 FILLER_ASAP7_75t_R FILLER_142_210 ();
 DECAPx2_ASAP7_75t_R FILLER_142_228 ();
 FILLER_ASAP7_75t_R FILLER_142_234 ();
 FILLER_ASAP7_75t_R FILLER_142_246 ();
 FILLER_ASAP7_75t_R FILLER_142_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_341 ();
 DECAPx4_ASAP7_75t_R FILLER_142_348 ();
 FILLER_ASAP7_75t_R FILLER_142_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_363 ();
 DECAPx1_ASAP7_75t_R FILLER_142_378 ();
 FILLER_ASAP7_75t_R FILLER_142_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_390 ();
 DECAPx10_ASAP7_75t_R FILLER_142_424 ();
 DECAPx6_ASAP7_75t_R FILLER_142_446 ();
 FILLER_ASAP7_75t_R FILLER_142_460 ();
 DECAPx6_ASAP7_75t_R FILLER_142_464 ();
 DECAPx6_ASAP7_75t_R FILLER_142_492 ();
 DECAPx2_ASAP7_75t_R FILLER_142_516 ();
 FILLER_ASAP7_75t_R FILLER_142_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_524 ();
 DECAPx2_ASAP7_75t_R FILLER_142_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_549 ();
 DECAPx1_ASAP7_75t_R FILLER_142_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_568 ();
 FILLER_ASAP7_75t_R FILLER_142_581 ();
 DECAPx2_ASAP7_75t_R FILLER_142_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_599 ();
 DECAPx1_ASAP7_75t_R FILLER_142_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_639 ();
 DECAPx6_ASAP7_75t_R FILLER_142_643 ();
 DECAPx1_ASAP7_75t_R FILLER_142_657 ();
 DECAPx2_ASAP7_75t_R FILLER_142_667 ();
 FILLER_ASAP7_75t_R FILLER_142_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_675 ();
 FILLER_ASAP7_75t_R FILLER_142_679 ();
 FILLER_ASAP7_75t_R FILLER_142_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_693 ();
 DECAPx10_ASAP7_75t_R FILLER_142_697 ();
 DECAPx2_ASAP7_75t_R FILLER_142_719 ();
 FILLER_ASAP7_75t_R FILLER_142_725 ();
 DECAPx4_ASAP7_75t_R FILLER_142_741 ();
 FILLER_ASAP7_75t_R FILLER_142_751 ();
 DECAPx6_ASAP7_75t_R FILLER_142_769 ();
 DECAPx1_ASAP7_75t_R FILLER_142_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_787 ();
 DECAPx6_ASAP7_75t_R FILLER_142_815 ();
 FILLER_ASAP7_75t_R FILLER_142_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_853 ();
 DECAPx10_ASAP7_75t_R FILLER_142_866 ();
 DECAPx10_ASAP7_75t_R FILLER_142_888 ();
 FILLER_ASAP7_75t_R FILLER_142_910 ();
 DECAPx4_ASAP7_75t_R FILLER_142_922 ();
 FILLER_ASAP7_75t_R FILLER_142_932 ();
 DECAPx10_ASAP7_75t_R FILLER_142_946 ();
 DECAPx10_ASAP7_75t_R FILLER_142_968 ();
 FILLER_ASAP7_75t_R FILLER_142_990 ();
 DECAPx1_ASAP7_75t_R FILLER_142_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1079 ();
 FILLER_ASAP7_75t_R FILLER_142_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1115 ();
 FILLER_ASAP7_75t_R FILLER_142_1121 ();
 FILLER_ASAP7_75t_R FILLER_142_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1225 ();
 FILLER_ASAP7_75t_R FILLER_142_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1259 ();
 FILLER_ASAP7_75t_R FILLER_142_1280 ();
 FILLER_ASAP7_75t_R FILLER_142_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1305 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1327 ();
 FILLER_ASAP7_75t_R FILLER_142_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1388 ();
 FILLER_ASAP7_75t_R FILLER_142_1394 ();
 FILLER_ASAP7_75t_R FILLER_142_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_143_2 ();
 DECAPx2_ASAP7_75t_R FILLER_143_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_22 ();
 DECAPx6_ASAP7_75t_R FILLER_143_26 ();
 DECAPx6_ASAP7_75t_R FILLER_143_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_91 ();
 DECAPx4_ASAP7_75t_R FILLER_143_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_142 ();
 DECAPx10_ASAP7_75t_R FILLER_143_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_182 ();
 DECAPx10_ASAP7_75t_R FILLER_143_191 ();
 DECAPx10_ASAP7_75t_R FILLER_143_213 ();
 FILLER_ASAP7_75t_R FILLER_143_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_237 ();
 DECAPx2_ASAP7_75t_R FILLER_143_268 ();
 DECAPx1_ASAP7_75t_R FILLER_143_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_285 ();
 DECAPx4_ASAP7_75t_R FILLER_143_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_335 ();
 DECAPx1_ASAP7_75t_R FILLER_143_350 ();
 DECAPx2_ASAP7_75t_R FILLER_143_362 ();
 FILLER_ASAP7_75t_R FILLER_143_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_370 ();
 FILLER_ASAP7_75t_R FILLER_143_392 ();
 DECAPx1_ASAP7_75t_R FILLER_143_400 ();
 DECAPx2_ASAP7_75t_R FILLER_143_418 ();
 FILLER_ASAP7_75t_R FILLER_143_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_426 ();
 DECAPx4_ASAP7_75t_R FILLER_143_437 ();
 DECAPx2_ASAP7_75t_R FILLER_143_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_481 ();
 DECAPx10_ASAP7_75t_R FILLER_143_500 ();
 DECAPx10_ASAP7_75t_R FILLER_143_522 ();
 DECAPx1_ASAP7_75t_R FILLER_143_544 ();
 DECAPx2_ASAP7_75t_R FILLER_143_564 ();
 FILLER_ASAP7_75t_R FILLER_143_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_572 ();
 DECAPx10_ASAP7_75t_R FILLER_143_576 ();
 DECAPx2_ASAP7_75t_R FILLER_143_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_604 ();
 DECAPx4_ASAP7_75t_R FILLER_143_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_621 ();
 DECAPx4_ASAP7_75t_R FILLER_143_631 ();
 FILLER_ASAP7_75t_R FILLER_143_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_643 ();
 DECAPx4_ASAP7_75t_R FILLER_143_670 ();
 DECAPx2_ASAP7_75t_R FILLER_143_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_734 ();
 DECAPx10_ASAP7_75t_R FILLER_143_742 ();
 DECAPx10_ASAP7_75t_R FILLER_143_764 ();
 DECAPx1_ASAP7_75t_R FILLER_143_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_790 ();
 DECAPx10_ASAP7_75t_R FILLER_143_817 ();
 DECAPx6_ASAP7_75t_R FILLER_143_839 ();
 DECAPx1_ASAP7_75t_R FILLER_143_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_857 ();
 DECAPx10_ASAP7_75t_R FILLER_143_865 ();
 DECAPx2_ASAP7_75t_R FILLER_143_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_893 ();
 DECAPx6_ASAP7_75t_R FILLER_143_904 ();
 DECAPx2_ASAP7_75t_R FILLER_143_918 ();
 FILLER_ASAP7_75t_R FILLER_143_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_934 ();
 DECAPx4_ASAP7_75t_R FILLER_143_951 ();
 DECAPx10_ASAP7_75t_R FILLER_143_967 ();
 DECAPx10_ASAP7_75t_R FILLER_143_989 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1101 ();
 FILLER_ASAP7_75t_R FILLER_143_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1305 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1331 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1358 ();
 FILLER_ASAP7_75t_R FILLER_143_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_144_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_30 ();
 DECAPx2_ASAP7_75t_R FILLER_144_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_43 ();
 FILLER_ASAP7_75t_R FILLER_144_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_52 ();
 DECAPx2_ASAP7_75t_R FILLER_144_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_114 ();
 DECAPx4_ASAP7_75t_R FILLER_144_131 ();
 FILLER_ASAP7_75t_R FILLER_144_141 ();
 FILLER_ASAP7_75t_R FILLER_144_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_181 ();
 DECAPx2_ASAP7_75t_R FILLER_144_202 ();
 FILLER_ASAP7_75t_R FILLER_144_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_210 ();
 DECAPx1_ASAP7_75t_R FILLER_144_225 ();
 DECAPx4_ASAP7_75t_R FILLER_144_239 ();
 FILLER_ASAP7_75t_R FILLER_144_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_251 ();
 DECAPx1_ASAP7_75t_R FILLER_144_268 ();
 DECAPx10_ASAP7_75t_R FILLER_144_282 ();
 FILLER_ASAP7_75t_R FILLER_144_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_306 ();
 FILLER_ASAP7_75t_R FILLER_144_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_312 ();
 DECAPx6_ASAP7_75t_R FILLER_144_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_400 ();
 DECAPx1_ASAP7_75t_R FILLER_144_407 ();
 FILLER_ASAP7_75t_R FILLER_144_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_442 ();
 DECAPx1_ASAP7_75t_R FILLER_144_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_461 ();
 DECAPx1_ASAP7_75t_R FILLER_144_464 ();
 DECAPx6_ASAP7_75t_R FILLER_144_478 ();
 DECAPx4_ASAP7_75t_R FILLER_144_514 ();
 FILLER_ASAP7_75t_R FILLER_144_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_526 ();
 FILLER_ASAP7_75t_R FILLER_144_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_545 ();
 DECAPx2_ASAP7_75t_R FILLER_144_556 ();
 FILLER_ASAP7_75t_R FILLER_144_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_564 ();
 DECAPx2_ASAP7_75t_R FILLER_144_568 ();
 FILLER_ASAP7_75t_R FILLER_144_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_576 ();
 DECAPx10_ASAP7_75t_R FILLER_144_592 ();
 DECAPx2_ASAP7_75t_R FILLER_144_614 ();
 FILLER_ASAP7_75t_R FILLER_144_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_622 ();
 DECAPx1_ASAP7_75t_R FILLER_144_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_636 ();
 DECAPx4_ASAP7_75t_R FILLER_144_669 ();
 FILLER_ASAP7_75t_R FILLER_144_679 ();
 DECAPx10_ASAP7_75t_R FILLER_144_687 ();
 DECAPx10_ASAP7_75t_R FILLER_144_709 ();
 DECAPx10_ASAP7_75t_R FILLER_144_731 ();
 DECAPx1_ASAP7_75t_R FILLER_144_753 ();
 DECAPx2_ASAP7_75t_R FILLER_144_765 ();
 FILLER_ASAP7_75t_R FILLER_144_771 ();
 DECAPx2_ASAP7_75t_R FILLER_144_780 ();
 FILLER_ASAP7_75t_R FILLER_144_786 ();
 DECAPx2_ASAP7_75t_R FILLER_144_794 ();
 FILLER_ASAP7_75t_R FILLER_144_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_814 ();
 DECAPx1_ASAP7_75t_R FILLER_144_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_825 ();
 DECAPx1_ASAP7_75t_R FILLER_144_838 ();
 DECAPx4_ASAP7_75t_R FILLER_144_859 ();
 FILLER_ASAP7_75t_R FILLER_144_869 ();
 FILLER_ASAP7_75t_R FILLER_144_891 ();
 DECAPx4_ASAP7_75t_R FILLER_144_925 ();
 FILLER_ASAP7_75t_R FILLER_144_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_937 ();
 DECAPx6_ASAP7_75t_R FILLER_144_944 ();
 DECAPx2_ASAP7_75t_R FILLER_144_973 ();
 DECAPx6_ASAP7_75t_R FILLER_144_993 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1020 ();
 FILLER_ASAP7_75t_R FILLER_144_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_144_1270 ();
 FILLER_ASAP7_75t_R FILLER_144_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1292 ();
 FILLER_ASAP7_75t_R FILLER_144_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1300 ();
 FILLER_ASAP7_75t_R FILLER_144_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1330 ();
 DECAPx4_ASAP7_75t_R FILLER_145_2 ();
 FILLER_ASAP7_75t_R FILLER_145_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_14 ();
 DECAPx2_ASAP7_75t_R FILLER_145_45 ();
 DECAPx4_ASAP7_75t_R FILLER_145_57 ();
 FILLER_ASAP7_75t_R FILLER_145_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_69 ();
 FILLER_ASAP7_75t_R FILLER_145_85 ();
 DECAPx1_ASAP7_75t_R FILLER_145_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_143 ();
 DECAPx10_ASAP7_75t_R FILLER_145_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_173 ();
 DECAPx2_ASAP7_75t_R FILLER_145_197 ();
 FILLER_ASAP7_75t_R FILLER_145_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_205 ();
 DECAPx10_ASAP7_75t_R FILLER_145_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_274 ();
 DECAPx1_ASAP7_75t_R FILLER_145_285 ();
 DECAPx6_ASAP7_75t_R FILLER_145_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_313 ();
 DECAPx1_ASAP7_75t_R FILLER_145_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_348 ();
 DECAPx10_ASAP7_75t_R FILLER_145_359 ();
 FILLER_ASAP7_75t_R FILLER_145_381 ();
 DECAPx6_ASAP7_75t_R FILLER_145_389 ();
 DECAPx2_ASAP7_75t_R FILLER_145_403 ();
 DECAPx10_ASAP7_75t_R FILLER_145_415 ();
 DECAPx2_ASAP7_75t_R FILLER_145_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_443 ();
 DECAPx10_ASAP7_75t_R FILLER_145_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_502 ();
 DECAPx1_ASAP7_75t_R FILLER_145_529 ();
 DECAPx2_ASAP7_75t_R FILLER_145_538 ();
 DECAPx6_ASAP7_75t_R FILLER_145_582 ();
 DECAPx1_ASAP7_75t_R FILLER_145_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_616 ();
 DECAPx1_ASAP7_75t_R FILLER_145_638 ();
 DECAPx4_ASAP7_75t_R FILLER_145_648 ();
 FILLER_ASAP7_75t_R FILLER_145_664 ();
 DECAPx10_ASAP7_75t_R FILLER_145_672 ();
 DECAPx10_ASAP7_75t_R FILLER_145_694 ();
 DECAPx10_ASAP7_75t_R FILLER_145_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_738 ();
 DECAPx1_ASAP7_75t_R FILLER_145_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_749 ();
 FILLER_ASAP7_75t_R FILLER_145_778 ();
 DECAPx1_ASAP7_75t_R FILLER_145_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_809 ();
 DECAPx6_ASAP7_75t_R FILLER_145_822 ();
 DECAPx1_ASAP7_75t_R FILLER_145_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_840 ();
 FILLER_ASAP7_75t_R FILLER_145_852 ();
 FILLER_ASAP7_75t_R FILLER_145_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_866 ();
 DECAPx10_ASAP7_75t_R FILLER_145_874 ();
 DECAPx6_ASAP7_75t_R FILLER_145_896 ();
 DECAPx10_ASAP7_75t_R FILLER_145_926 ();
 DECAPx10_ASAP7_75t_R FILLER_145_948 ();
 DECAPx6_ASAP7_75t_R FILLER_145_970 ();
 FILLER_ASAP7_75t_R FILLER_145_984 ();
 DECAPx1_ASAP7_75t_R FILLER_145_996 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1283 ();
 FILLER_ASAP7_75t_R FILLER_145_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1348 ();
 FILLER_ASAP7_75t_R FILLER_145_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_146_2 ();
 DECAPx2_ASAP7_75t_R FILLER_146_24 ();
 FILLER_ASAP7_75t_R FILLER_146_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_41 ();
 DECAPx10_ASAP7_75t_R FILLER_146_68 ();
 FILLER_ASAP7_75t_R FILLER_146_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_106 ();
 DECAPx6_ASAP7_75t_R FILLER_146_110 ();
 DECAPx1_ASAP7_75t_R FILLER_146_124 ();
 FILLER_ASAP7_75t_R FILLER_146_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_176 ();
 DECAPx10_ASAP7_75t_R FILLER_146_191 ();
 FILLER_ASAP7_75t_R FILLER_146_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_215 ();
 DECAPx6_ASAP7_75t_R FILLER_146_232 ();
 FILLER_ASAP7_75t_R FILLER_146_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_248 ();
 DECAPx1_ASAP7_75t_R FILLER_146_265 ();
 DECAPx1_ASAP7_75t_R FILLER_146_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_287 ();
 DECAPx6_ASAP7_75t_R FILLER_146_339 ();
 DECAPx2_ASAP7_75t_R FILLER_146_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_359 ();
 FILLER_ASAP7_75t_R FILLER_146_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_372 ();
 DECAPx6_ASAP7_75t_R FILLER_146_383 ();
 DECAPx1_ASAP7_75t_R FILLER_146_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_401 ();
 DECAPx10_ASAP7_75t_R FILLER_146_412 ();
 FILLER_ASAP7_75t_R FILLER_146_434 ();
 DECAPx1_ASAP7_75t_R FILLER_146_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_461 ();
 DECAPx6_ASAP7_75t_R FILLER_146_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_478 ();
 DECAPx1_ASAP7_75t_R FILLER_146_485 ();
 DECAPx4_ASAP7_75t_R FILLER_146_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_502 ();
 FILLER_ASAP7_75t_R FILLER_146_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_520 ();
 FILLER_ASAP7_75t_R FILLER_146_535 ();
 DECAPx10_ASAP7_75t_R FILLER_146_550 ();
 FILLER_ASAP7_75t_R FILLER_146_572 ();
 FILLER_ASAP7_75t_R FILLER_146_585 ();
 DECAPx2_ASAP7_75t_R FILLER_146_616 ();
 FILLER_ASAP7_75t_R FILLER_146_628 ();
 FILLER_ASAP7_75t_R FILLER_146_639 ();
 DECAPx2_ASAP7_75t_R FILLER_146_647 ();
 FILLER_ASAP7_75t_R FILLER_146_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_655 ();
 DECAPx2_ASAP7_75t_R FILLER_146_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_665 ();
 DECAPx10_ASAP7_75t_R FILLER_146_698 ();
 DECAPx10_ASAP7_75t_R FILLER_146_720 ();
 DECAPx6_ASAP7_75t_R FILLER_146_742 ();
 DECAPx1_ASAP7_75t_R FILLER_146_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_760 ();
 DECAPx10_ASAP7_75t_R FILLER_146_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_813 ();
 DECAPx2_ASAP7_75t_R FILLER_146_820 ();
 FILLER_ASAP7_75t_R FILLER_146_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_828 ();
 DECAPx10_ASAP7_75t_R FILLER_146_836 ();
 DECAPx10_ASAP7_75t_R FILLER_146_858 ();
 DECAPx6_ASAP7_75t_R FILLER_146_880 ();
 DECAPx2_ASAP7_75t_R FILLER_146_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_900 ();
 DECAPx10_ASAP7_75t_R FILLER_146_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_929 ();
 DECAPx10_ASAP7_75t_R FILLER_146_936 ();
 DECAPx10_ASAP7_75t_R FILLER_146_958 ();
 DECAPx10_ASAP7_75t_R FILLER_146_980 ();
 FILLER_ASAP7_75t_R FILLER_146_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1093 ();
 FILLER_ASAP7_75t_R FILLER_146_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1187 ();
 FILLER_ASAP7_75t_R FILLER_146_1220 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1252 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1281 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1312 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1385 ();
 FILLER_ASAP7_75t_R FILLER_146_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_147_2 ();
 FILLER_ASAP7_75t_R FILLER_147_24 ();
 DECAPx4_ASAP7_75t_R FILLER_147_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_45 ();
 DECAPx1_ASAP7_75t_R FILLER_147_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_56 ();
 DECAPx4_ASAP7_75t_R FILLER_147_60 ();
 DECAPx6_ASAP7_75t_R FILLER_147_79 ();
 FILLER_ASAP7_75t_R FILLER_147_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_95 ();
 DECAPx10_ASAP7_75t_R FILLER_147_99 ();
 DECAPx1_ASAP7_75t_R FILLER_147_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_125 ();
 DECAPx4_ASAP7_75t_R FILLER_147_140 ();
 DECAPx1_ASAP7_75t_R FILLER_147_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_160 ();
 DECAPx6_ASAP7_75t_R FILLER_147_164 ();
 FILLER_ASAP7_75t_R FILLER_147_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_180 ();
 DECAPx1_ASAP7_75t_R FILLER_147_187 ();
 FILLER_ASAP7_75t_R FILLER_147_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_199 ();
 DECAPx2_ASAP7_75t_R FILLER_147_214 ();
 FILLER_ASAP7_75t_R FILLER_147_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_222 ();
 DECAPx4_ASAP7_75t_R FILLER_147_239 ();
 FILLER_ASAP7_75t_R FILLER_147_249 ();
 DECAPx2_ASAP7_75t_R FILLER_147_265 ();
 FILLER_ASAP7_75t_R FILLER_147_271 ();
 DECAPx4_ASAP7_75t_R FILLER_147_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_293 ();
 DECAPx4_ASAP7_75t_R FILLER_147_298 ();
 FILLER_ASAP7_75t_R FILLER_147_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_330 ();
 FILLER_ASAP7_75t_R FILLER_147_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_363 ();
 DECAPx1_ASAP7_75t_R FILLER_147_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_388 ();
 DECAPx1_ASAP7_75t_R FILLER_147_433 ();
 DECAPx2_ASAP7_75t_R FILLER_147_463 ();
 DECAPx6_ASAP7_75t_R FILLER_147_501 ();
 DECAPx2_ASAP7_75t_R FILLER_147_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_521 ();
 DECAPx6_ASAP7_75t_R FILLER_147_528 ();
 DECAPx10_ASAP7_75t_R FILLER_147_548 ();
 DECAPx4_ASAP7_75t_R FILLER_147_570 ();
 FILLER_ASAP7_75t_R FILLER_147_580 ();
 FILLER_ASAP7_75t_R FILLER_147_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_611 ();
 DECAPx6_ASAP7_75t_R FILLER_147_626 ();
 FILLER_ASAP7_75t_R FILLER_147_640 ();
 DECAPx1_ASAP7_75t_R FILLER_147_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_672 ();
 DECAPx2_ASAP7_75t_R FILLER_147_702 ();
 DECAPx10_ASAP7_75t_R FILLER_147_718 ();
 DECAPx1_ASAP7_75t_R FILLER_147_740 ();
 DECAPx10_ASAP7_75t_R FILLER_147_752 ();
 DECAPx2_ASAP7_75t_R FILLER_147_774 ();
 DECAPx1_ASAP7_75t_R FILLER_147_818 ();
 DECAPx4_ASAP7_75t_R FILLER_147_842 ();
 DECAPx6_ASAP7_75t_R FILLER_147_860 ();
 FILLER_ASAP7_75t_R FILLER_147_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_876 ();
 DECAPx10_ASAP7_75t_R FILLER_147_881 ();
 DECAPx6_ASAP7_75t_R FILLER_147_903 ();
 DECAPx2_ASAP7_75t_R FILLER_147_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_923 ();
 DECAPx4_ASAP7_75t_R FILLER_147_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_936 ();
 DECAPx2_ASAP7_75t_R FILLER_147_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_953 ();
 DECAPx1_ASAP7_75t_R FILLER_147_960 ();
 DECAPx10_ASAP7_75t_R FILLER_147_971 ();
 DECAPx10_ASAP7_75t_R FILLER_147_993 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1084 ();
 FILLER_ASAP7_75t_R FILLER_147_1099 ();
 FILLER_ASAP7_75t_R FILLER_147_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1146 ();
 FILLER_ASAP7_75t_R FILLER_147_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1169 ();
 FILLER_ASAP7_75t_R FILLER_147_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1193 ();
 FILLER_ASAP7_75t_R FILLER_147_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1233 ();
 FILLER_ASAP7_75t_R FILLER_147_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1253 ();
 FILLER_ASAP7_75t_R FILLER_147_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_148_2 ();
 DECAPx2_ASAP7_75t_R FILLER_148_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_47 ();
 DECAPx2_ASAP7_75t_R FILLER_148_54 ();
 FILLER_ASAP7_75t_R FILLER_148_60 ();
 DECAPx1_ASAP7_75t_R FILLER_148_91 ();
 DECAPx1_ASAP7_75t_R FILLER_148_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_110 ();
 DECAPx6_ASAP7_75t_R FILLER_148_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_135 ();
 DECAPx6_ASAP7_75t_R FILLER_148_150 ();
 DECAPx2_ASAP7_75t_R FILLER_148_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_170 ();
 DECAPx2_ASAP7_75t_R FILLER_148_193 ();
 DECAPx2_ASAP7_75t_R FILLER_148_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_223 ();
 DECAPx1_ASAP7_75t_R FILLER_148_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_238 ();
 DECAPx1_ASAP7_75t_R FILLER_148_257 ();
 DECAPx2_ASAP7_75t_R FILLER_148_264 ();
 FILLER_ASAP7_75t_R FILLER_148_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_272 ();
 DECAPx10_ASAP7_75t_R FILLER_148_281 ();
 FILLER_ASAP7_75t_R FILLER_148_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_305 ();
 DECAPx2_ASAP7_75t_R FILLER_148_342 ();
 FILLER_ASAP7_75t_R FILLER_148_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_350 ();
 DECAPx6_ASAP7_75t_R FILLER_148_361 ();
 DECAPx2_ASAP7_75t_R FILLER_148_375 ();
 DECAPx1_ASAP7_75t_R FILLER_148_391 ();
 DECAPx2_ASAP7_75t_R FILLER_148_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_411 ();
 DECAPx4_ASAP7_75t_R FILLER_148_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_432 ();
 DECAPx2_ASAP7_75t_R FILLER_148_443 ();
 FILLER_ASAP7_75t_R FILLER_148_449 ();
 DECAPx1_ASAP7_75t_R FILLER_148_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_461 ();
 DECAPx2_ASAP7_75t_R FILLER_148_467 ();
 FILLER_ASAP7_75t_R FILLER_148_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_475 ();
 DECAPx4_ASAP7_75t_R FILLER_148_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_492 ();
 DECAPx1_ASAP7_75t_R FILLER_148_504 ();
 DECAPx6_ASAP7_75t_R FILLER_148_515 ();
 DECAPx1_ASAP7_75t_R FILLER_148_529 ();
 DECAPx1_ASAP7_75t_R FILLER_148_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_547 ();
 DECAPx10_ASAP7_75t_R FILLER_148_569 ();
 DECAPx10_ASAP7_75t_R FILLER_148_591 ();
 DECAPx6_ASAP7_75t_R FILLER_148_613 ();
 FILLER_ASAP7_75t_R FILLER_148_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_629 ();
 DECAPx10_ASAP7_75t_R FILLER_148_638 ();
 DECAPx1_ASAP7_75t_R FILLER_148_660 ();
 DECAPx2_ASAP7_75t_R FILLER_148_682 ();
 DECAPx10_ASAP7_75t_R FILLER_148_694 ();
 FILLER_ASAP7_75t_R FILLER_148_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_757 ();
 FILLER_ASAP7_75t_R FILLER_148_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_797 ();
 DECAPx1_ASAP7_75t_R FILLER_148_806 ();
 DECAPx2_ASAP7_75t_R FILLER_148_816 ();
 FILLER_ASAP7_75t_R FILLER_148_822 ();
 DECAPx4_ASAP7_75t_R FILLER_148_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_846 ();
 DECAPx1_ASAP7_75t_R FILLER_148_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_863 ();
 DECAPx1_ASAP7_75t_R FILLER_148_876 ();
 FILLER_ASAP7_75t_R FILLER_148_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_897 ();
 DECAPx10_ASAP7_75t_R FILLER_148_906 ();
 DECAPx2_ASAP7_75t_R FILLER_148_928 ();
 FILLER_ASAP7_75t_R FILLER_148_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_936 ();
 DECAPx10_ASAP7_75t_R FILLER_148_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_980 ();
 FILLER_ASAP7_75t_R FILLER_148_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1016 ();
 FILLER_ASAP7_75t_R FILLER_148_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1079 ();
 FILLER_ASAP7_75t_R FILLER_148_1098 ();
 FILLER_ASAP7_75t_R FILLER_148_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1271 ();
 FILLER_ASAP7_75t_R FILLER_148_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1319 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1357 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1396 ();
 FILLER_ASAP7_75t_R FILLER_148_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_149_2 ();
 FILLER_ASAP7_75t_R FILLER_149_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_26 ();
 DECAPx2_ASAP7_75t_R FILLER_149_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_99 ();
 DECAPx4_ASAP7_75t_R FILLER_149_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_142 ();
 DECAPx10_ASAP7_75t_R FILLER_149_188 ();
 DECAPx10_ASAP7_75t_R FILLER_149_210 ();
 DECAPx2_ASAP7_75t_R FILLER_149_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_305 ();
 DECAPx2_ASAP7_75t_R FILLER_149_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_322 ();
 FILLER_ASAP7_75t_R FILLER_149_329 ();
 DECAPx6_ASAP7_75t_R FILLER_149_334 ();
 FILLER_ASAP7_75t_R FILLER_149_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_350 ();
 DECAPx6_ASAP7_75t_R FILLER_149_365 ();
 FILLER_ASAP7_75t_R FILLER_149_399 ();
 DECAPx2_ASAP7_75t_R FILLER_149_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_431 ();
 DECAPx2_ASAP7_75t_R FILLER_149_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_448 ();
 DECAPx4_ASAP7_75t_R FILLER_149_475 ();
 FILLER_ASAP7_75t_R FILLER_149_485 ();
 DECAPx6_ASAP7_75t_R FILLER_149_509 ();
 DECAPx1_ASAP7_75t_R FILLER_149_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_527 ();
 DECAPx4_ASAP7_75t_R FILLER_149_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_556 ();
 DECAPx4_ASAP7_75t_R FILLER_149_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_575 ();
 DECAPx4_ASAP7_75t_R FILLER_149_584 ();
 DECAPx1_ASAP7_75t_R FILLER_149_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_648 ();
 DECAPx10_ASAP7_75t_R FILLER_149_669 ();
 DECAPx1_ASAP7_75t_R FILLER_149_701 ();
 DECAPx2_ASAP7_75t_R FILLER_149_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_714 ();
 DECAPx1_ASAP7_75t_R FILLER_149_724 ();
 DECAPx1_ASAP7_75t_R FILLER_149_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_745 ();
 DECAPx2_ASAP7_75t_R FILLER_149_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_761 ();
 DECAPx1_ASAP7_75t_R FILLER_149_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_774 ();
 DECAPx1_ASAP7_75t_R FILLER_149_789 ();
 FILLER_ASAP7_75t_R FILLER_149_807 ();
 DECAPx1_ASAP7_75t_R FILLER_149_822 ();
 DECAPx2_ASAP7_75t_R FILLER_149_834 ();
 FILLER_ASAP7_75t_R FILLER_149_840 ();
 DECAPx4_ASAP7_75t_R FILLER_149_845 ();
 FILLER_ASAP7_75t_R FILLER_149_855 ();
 DECAPx2_ASAP7_75t_R FILLER_149_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_871 ();
 DECAPx6_ASAP7_75t_R FILLER_149_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_897 ();
 DECAPx4_ASAP7_75t_R FILLER_149_904 ();
 DECAPx1_ASAP7_75t_R FILLER_149_920 ();
 DECAPx10_ASAP7_75t_R FILLER_149_926 ();
 DECAPx10_ASAP7_75t_R FILLER_149_948 ();
 DECAPx1_ASAP7_75t_R FILLER_149_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_981 ();
 DECAPx6_ASAP7_75t_R FILLER_149_990 ();
 FILLER_ASAP7_75t_R FILLER_149_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1066 ();
 FILLER_ASAP7_75t_R FILLER_149_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1151 ();
 FILLER_ASAP7_75t_R FILLER_149_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1207 ();
 FILLER_ASAP7_75t_R FILLER_149_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1304 ();
 FILLER_ASAP7_75t_R FILLER_149_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1395 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1399 ();
 DECAPx6_ASAP7_75t_R FILLER_150_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_16 ();
 DECAPx1_ASAP7_75t_R FILLER_150_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_53 ();
 DECAPx6_ASAP7_75t_R FILLER_150_57 ();
 DECAPx2_ASAP7_75t_R FILLER_150_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_84 ();
 FILLER_ASAP7_75t_R FILLER_150_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_93 ();
 DECAPx4_ASAP7_75t_R FILLER_150_102 ();
 FILLER_ASAP7_75t_R FILLER_150_112 ();
 FILLER_ASAP7_75t_R FILLER_150_122 ();
 FILLER_ASAP7_75t_R FILLER_150_134 ();
 FILLER_ASAP7_75t_R FILLER_150_156 ();
 DECAPx4_ASAP7_75t_R FILLER_150_161 ();
 FILLER_ASAP7_75t_R FILLER_150_171 ();
 DECAPx10_ASAP7_75t_R FILLER_150_176 ();
 DECAPx1_ASAP7_75t_R FILLER_150_198 ();
 DECAPx1_ASAP7_75t_R FILLER_150_226 ();
 DECAPx4_ASAP7_75t_R FILLER_150_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_254 ();
 DECAPx6_ASAP7_75t_R FILLER_150_262 ();
 DECAPx1_ASAP7_75t_R FILLER_150_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_280 ();
 FILLER_ASAP7_75t_R FILLER_150_295 ();
 DECAPx10_ASAP7_75t_R FILLER_150_307 ();
 DECAPx4_ASAP7_75t_R FILLER_150_329 ();
 FILLER_ASAP7_75t_R FILLER_150_339 ();
 DECAPx1_ASAP7_75t_R FILLER_150_355 ();
 DECAPx1_ASAP7_75t_R FILLER_150_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_393 ();
 FILLER_ASAP7_75t_R FILLER_150_410 ();
 DECAPx4_ASAP7_75t_R FILLER_150_432 ();
 FILLER_ASAP7_75t_R FILLER_150_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_444 ();
 DECAPx4_ASAP7_75t_R FILLER_150_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_461 ();
 DECAPx2_ASAP7_75t_R FILLER_150_464 ();
 FILLER_ASAP7_75t_R FILLER_150_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_472 ();
 DECAPx6_ASAP7_75t_R FILLER_150_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_490 ();
 DECAPx1_ASAP7_75t_R FILLER_150_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_501 ();
 DECAPx4_ASAP7_75t_R FILLER_150_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_525 ();
 DECAPx1_ASAP7_75t_R FILLER_150_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_538 ();
 DECAPx6_ASAP7_75t_R FILLER_150_547 ();
 DECAPx2_ASAP7_75t_R FILLER_150_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_567 ();
 DECAPx6_ASAP7_75t_R FILLER_150_586 ();
 DECAPx2_ASAP7_75t_R FILLER_150_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_606 ();
 DECAPx1_ASAP7_75t_R FILLER_150_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_619 ();
 DECAPx2_ASAP7_75t_R FILLER_150_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_636 ();
 DECAPx1_ASAP7_75t_R FILLER_150_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_662 ();
 DECAPx1_ASAP7_75t_R FILLER_150_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_721 ();
 FILLER_ASAP7_75t_R FILLER_150_729 ();
 DECAPx10_ASAP7_75t_R FILLER_150_737 ();
 DECAPx2_ASAP7_75t_R FILLER_150_759 ();
 DECAPx10_ASAP7_75t_R FILLER_150_773 ();
 FILLER_ASAP7_75t_R FILLER_150_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_813 ();
 DECAPx10_ASAP7_75t_R FILLER_150_829 ();
 DECAPx10_ASAP7_75t_R FILLER_150_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_873 ();
 DECAPx6_ASAP7_75t_R FILLER_150_882 ();
 FILLER_ASAP7_75t_R FILLER_150_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_898 ();
 DECAPx4_ASAP7_75t_R FILLER_150_907 ();
 FILLER_ASAP7_75t_R FILLER_150_917 ();
 DECAPx10_ASAP7_75t_R FILLER_150_931 ();
 DECAPx1_ASAP7_75t_R FILLER_150_953 ();
 FILLER_ASAP7_75t_R FILLER_150_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_978 ();
 DECAPx10_ASAP7_75t_R FILLER_150_985 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1007 ();
 FILLER_ASAP7_75t_R FILLER_150_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1149 ();
 FILLER_ASAP7_75t_R FILLER_150_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1202 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1270 ();
 FILLER_ASAP7_75t_R FILLER_150_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1288 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1299 ();
 FILLER_ASAP7_75t_R FILLER_150_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1307 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1327 ();
 FILLER_ASAP7_75t_R FILLER_150_1341 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1354 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_151_2 ();
 FILLER_ASAP7_75t_R FILLER_151_30 ();
 DECAPx6_ASAP7_75t_R FILLER_151_35 ();
 DECAPx1_ASAP7_75t_R FILLER_151_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_67 ();
 DECAPx2_ASAP7_75t_R FILLER_151_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_94 ();
 FILLER_ASAP7_75t_R FILLER_151_98 ();
 FILLER_ASAP7_75t_R FILLER_151_115 ();
 DECAPx2_ASAP7_75t_R FILLER_151_120 ();
 DECAPx6_ASAP7_75t_R FILLER_151_148 ();
 DECAPx2_ASAP7_75t_R FILLER_151_162 ();
 DECAPx1_ASAP7_75t_R FILLER_151_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_190 ();
 DECAPx4_ASAP7_75t_R FILLER_151_209 ();
 DECAPx2_ASAP7_75t_R FILLER_151_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_287 ();
 DECAPx2_ASAP7_75t_R FILLER_151_314 ();
 FILLER_ASAP7_75t_R FILLER_151_320 ();
 DECAPx4_ASAP7_75t_R FILLER_151_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_350 ();
 DECAPx10_ASAP7_75t_R FILLER_151_365 ();
 DECAPx6_ASAP7_75t_R FILLER_151_387 ();
 DECAPx1_ASAP7_75t_R FILLER_151_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_405 ();
 DECAPx2_ASAP7_75t_R FILLER_151_414 ();
 FILLER_ASAP7_75t_R FILLER_151_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_429 ();
 DECAPx1_ASAP7_75t_R FILLER_151_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_481 ();
 DECAPx4_ASAP7_75t_R FILLER_151_488 ();
 DECAPx2_ASAP7_75t_R FILLER_151_538 ();
 DECAPx10_ASAP7_75t_R FILLER_151_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_573 ();
 FILLER_ASAP7_75t_R FILLER_151_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_590 ();
 DECAPx6_ASAP7_75t_R FILLER_151_599 ();
 DECAPx2_ASAP7_75t_R FILLER_151_613 ();
 DECAPx10_ASAP7_75t_R FILLER_151_629 ();
 DECAPx10_ASAP7_75t_R FILLER_151_651 ();
 DECAPx6_ASAP7_75t_R FILLER_151_673 ();
 FILLER_ASAP7_75t_R FILLER_151_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_689 ();
 DECAPx6_ASAP7_75t_R FILLER_151_699 ();
 DECAPx1_ASAP7_75t_R FILLER_151_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_717 ();
 DECAPx4_ASAP7_75t_R FILLER_151_727 ();
 FILLER_ASAP7_75t_R FILLER_151_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_739 ();
 DECAPx2_ASAP7_75t_R FILLER_151_760 ();
 FILLER_ASAP7_75t_R FILLER_151_783 ();
 DECAPx2_ASAP7_75t_R FILLER_151_817 ();
 DECAPx1_ASAP7_75t_R FILLER_151_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_840 ();
 DECAPx10_ASAP7_75t_R FILLER_151_849 ();
 DECAPx10_ASAP7_75t_R FILLER_151_871 ();
 DECAPx10_ASAP7_75t_R FILLER_151_893 ();
 DECAPx2_ASAP7_75t_R FILLER_151_915 ();
 FILLER_ASAP7_75t_R FILLER_151_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_923 ();
 DECAPx6_ASAP7_75t_R FILLER_151_926 ();
 DECAPx6_ASAP7_75t_R FILLER_151_966 ();
 DECAPx2_ASAP7_75t_R FILLER_151_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_986 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1013 ();
 FILLER_ASAP7_75t_R FILLER_151_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1042 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1053 ();
 FILLER_ASAP7_75t_R FILLER_151_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1134 ();
 FILLER_ASAP7_75t_R FILLER_151_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1150 ();
 FILLER_ASAP7_75t_R FILLER_151_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1292 ();
 FILLER_ASAP7_75t_R FILLER_151_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1340 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1361 ();
 FILLER_ASAP7_75t_R FILLER_151_1377 ();
 DECAPx10_ASAP7_75t_R FILLER_152_2 ();
 DECAPx4_ASAP7_75t_R FILLER_152_34 ();
 FILLER_ASAP7_75t_R FILLER_152_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_56 ();
 FILLER_ASAP7_75t_R FILLER_152_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_117 ();
 DECAPx6_ASAP7_75t_R FILLER_152_128 ();
 DECAPx2_ASAP7_75t_R FILLER_152_142 ();
 FILLER_ASAP7_75t_R FILLER_152_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_160 ();
 DECAPx2_ASAP7_75t_R FILLER_152_193 ();
 FILLER_ASAP7_75t_R FILLER_152_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_201 ();
 DECAPx2_ASAP7_75t_R FILLER_152_212 ();
 FILLER_ASAP7_75t_R FILLER_152_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_220 ();
 FILLER_ASAP7_75t_R FILLER_152_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_261 ();
 DECAPx10_ASAP7_75t_R FILLER_152_265 ();
 DECAPx4_ASAP7_75t_R FILLER_152_287 ();
 FILLER_ASAP7_75t_R FILLER_152_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_299 ();
 DECAPx2_ASAP7_75t_R FILLER_152_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_324 ();
 DECAPx4_ASAP7_75t_R FILLER_152_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_369 ();
 DECAPx4_ASAP7_75t_R FILLER_152_388 ();
 FILLER_ASAP7_75t_R FILLER_152_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_400 ();
 DECAPx1_ASAP7_75t_R FILLER_152_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_415 ();
 FILLER_ASAP7_75t_R FILLER_152_442 ();
 DECAPx2_ASAP7_75t_R FILLER_152_450 ();
 FILLER_ASAP7_75t_R FILLER_152_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_461 ();
 DECAPx1_ASAP7_75t_R FILLER_152_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_468 ();
 DECAPx2_ASAP7_75t_R FILLER_152_475 ();
 DECAPx2_ASAP7_75t_R FILLER_152_529 ();
 FILLER_ASAP7_75t_R FILLER_152_535 ();
 DECAPx1_ASAP7_75t_R FILLER_152_553 ();
 FILLER_ASAP7_75t_R FILLER_152_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_576 ();
 FILLER_ASAP7_75t_R FILLER_152_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_585 ();
 DECAPx1_ASAP7_75t_R FILLER_152_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_616 ();
 DECAPx2_ASAP7_75t_R FILLER_152_658 ();
 FILLER_ASAP7_75t_R FILLER_152_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_666 ();
 DECAPx4_ASAP7_75t_R FILLER_152_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_686 ();
 DECAPx4_ASAP7_75t_R FILLER_152_716 ();
 FILLER_ASAP7_75t_R FILLER_152_726 ();
 DECAPx6_ASAP7_75t_R FILLER_152_738 ();
 DECAPx1_ASAP7_75t_R FILLER_152_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_756 ();
 FILLER_ASAP7_75t_R FILLER_152_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_765 ();
 DECAPx2_ASAP7_75t_R FILLER_152_772 ();
 DECAPx10_ASAP7_75t_R FILLER_152_784 ();
 DECAPx2_ASAP7_75t_R FILLER_152_809 ();
 FILLER_ASAP7_75t_R FILLER_152_815 ();
 DECAPx10_ASAP7_75t_R FILLER_152_825 ();
 DECAPx6_ASAP7_75t_R FILLER_152_847 ();
 DECAPx4_ASAP7_75t_R FILLER_152_868 ();
 DECAPx2_ASAP7_75t_R FILLER_152_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_897 ();
 DECAPx6_ASAP7_75t_R FILLER_152_904 ();
 DECAPx2_ASAP7_75t_R FILLER_152_918 ();
 DECAPx10_ASAP7_75t_R FILLER_152_930 ();
 DECAPx6_ASAP7_75t_R FILLER_152_952 ();
 FILLER_ASAP7_75t_R FILLER_152_966 ();
 DECAPx2_ASAP7_75t_R FILLER_152_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_990 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1029 ();
 FILLER_ASAP7_75t_R FILLER_152_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1104 ();
 FILLER_ASAP7_75t_R FILLER_152_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1223 ();
 FILLER_ASAP7_75t_R FILLER_152_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1270 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1304 ();
 FILLER_ASAP7_75t_R FILLER_152_1314 ();
 FILLER_ASAP7_75t_R FILLER_152_1328 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1396 ();
 FILLER_ASAP7_75t_R FILLER_152_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_153_2 ();
 FILLER_ASAP7_75t_R FILLER_153_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_40 ();
 DECAPx2_ASAP7_75t_R FILLER_153_67 ();
 FILLER_ASAP7_75t_R FILLER_153_73 ();
 FILLER_ASAP7_75t_R FILLER_153_81 ();
 DECAPx6_ASAP7_75t_R FILLER_153_86 ();
 DECAPx1_ASAP7_75t_R FILLER_153_100 ();
 DECAPx1_ASAP7_75t_R FILLER_153_147 ();
 DECAPx4_ASAP7_75t_R FILLER_153_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_179 ();
 DECAPx2_ASAP7_75t_R FILLER_153_196 ();
 FILLER_ASAP7_75t_R FILLER_153_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_204 ();
 DECAPx10_ASAP7_75t_R FILLER_153_215 ();
 DECAPx2_ASAP7_75t_R FILLER_153_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_243 ();
 DECAPx2_ASAP7_75t_R FILLER_153_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_260 ();
 DECAPx4_ASAP7_75t_R FILLER_153_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_277 ();
 DECAPx10_ASAP7_75t_R FILLER_153_294 ();
 DECAPx2_ASAP7_75t_R FILLER_153_316 ();
 FILLER_ASAP7_75t_R FILLER_153_322 ();
 DECAPx2_ASAP7_75t_R FILLER_153_340 ();
 FILLER_ASAP7_75t_R FILLER_153_346 ();
 DECAPx1_ASAP7_75t_R FILLER_153_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_370 ();
 DECAPx1_ASAP7_75t_R FILLER_153_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_393 ();
 DECAPx6_ASAP7_75t_R FILLER_153_414 ();
 FILLER_ASAP7_75t_R FILLER_153_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_430 ();
 DECAPx4_ASAP7_75t_R FILLER_153_434 ();
 FILLER_ASAP7_75t_R FILLER_153_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_446 ();
 DECAPx4_ASAP7_75t_R FILLER_153_479 ();
 DECAPx6_ASAP7_75t_R FILLER_153_525 ();
 DECAPx1_ASAP7_75t_R FILLER_153_539 ();
 DECAPx6_ASAP7_75t_R FILLER_153_549 ();
 DECAPx2_ASAP7_75t_R FILLER_153_563 ();
 DECAPx1_ASAP7_75t_R FILLER_153_577 ();
 FILLER_ASAP7_75t_R FILLER_153_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_595 ();
 DECAPx6_ASAP7_75t_R FILLER_153_628 ();
 DECAPx2_ASAP7_75t_R FILLER_153_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_686 ();
 DECAPx4_ASAP7_75t_R FILLER_153_705 ();
 FILLER_ASAP7_75t_R FILLER_153_715 ();
 DECAPx4_ASAP7_75t_R FILLER_153_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_737 ();
 DECAPx1_ASAP7_75t_R FILLER_153_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_757 ();
 DECAPx1_ASAP7_75t_R FILLER_153_765 ();
 DECAPx1_ASAP7_75t_R FILLER_153_783 ();
 DECAPx1_ASAP7_75t_R FILLER_153_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_797 ();
 DECAPx10_ASAP7_75t_R FILLER_153_829 ();
 DECAPx2_ASAP7_75t_R FILLER_153_851 ();
 FILLER_ASAP7_75t_R FILLER_153_857 ();
 DECAPx1_ASAP7_75t_R FILLER_153_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_867 ();
 FILLER_ASAP7_75t_R FILLER_153_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_878 ();
 DECAPx4_ASAP7_75t_R FILLER_153_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_911 ();
 DECAPx1_ASAP7_75t_R FILLER_153_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_923 ();
 FILLER_ASAP7_75t_R FILLER_153_932 ();
 DECAPx10_ASAP7_75t_R FILLER_153_948 ();
 DECAPx4_ASAP7_75t_R FILLER_153_970 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1052 ();
 FILLER_ASAP7_75t_R FILLER_153_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1111 ();
 FILLER_ASAP7_75t_R FILLER_153_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1160 ();
 FILLER_ASAP7_75t_R FILLER_153_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1180 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1208 ();
 FILLER_ASAP7_75t_R FILLER_153_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1272 ();
 FILLER_ASAP7_75t_R FILLER_153_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1379 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1392 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_154_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_24 ();
 FILLER_ASAP7_75t_R FILLER_154_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_41 ();
 DECAPx2_ASAP7_75t_R FILLER_154_48 ();
 FILLER_ASAP7_75t_R FILLER_154_54 ();
 DECAPx2_ASAP7_75t_R FILLER_154_59 ();
 FILLER_ASAP7_75t_R FILLER_154_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_67 ();
 DECAPx6_ASAP7_75t_R FILLER_154_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_145 ();
 DECAPx6_ASAP7_75t_R FILLER_154_156 ();
 DECAPx2_ASAP7_75t_R FILLER_154_170 ();
 FILLER_ASAP7_75t_R FILLER_154_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_192 ();
 DECAPx4_ASAP7_75t_R FILLER_154_219 ();
 FILLER_ASAP7_75t_R FILLER_154_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_231 ();
 DECAPx6_ASAP7_75t_R FILLER_154_242 ();
 FILLER_ASAP7_75t_R FILLER_154_256 ();
 DECAPx6_ASAP7_75t_R FILLER_154_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_286 ();
 DECAPx4_ASAP7_75t_R FILLER_154_313 ();
 DECAPx6_ASAP7_75t_R FILLER_154_337 ();
 FILLER_ASAP7_75t_R FILLER_154_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_367 ();
 FILLER_ASAP7_75t_R FILLER_154_396 ();
 DECAPx1_ASAP7_75t_R FILLER_154_408 ();
 DECAPx2_ASAP7_75t_R FILLER_154_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_461 ();
 DECAPx2_ASAP7_75t_R FILLER_154_467 ();
 DECAPx6_ASAP7_75t_R FILLER_154_476 ();
 FILLER_ASAP7_75t_R FILLER_154_490 ();
 FILLER_ASAP7_75t_R FILLER_154_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_516 ();
 DECAPx1_ASAP7_75t_R FILLER_154_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_537 ();
 DECAPx6_ASAP7_75t_R FILLER_154_554 ();
 DECAPx2_ASAP7_75t_R FILLER_154_568 ();
 FILLER_ASAP7_75t_R FILLER_154_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_582 ();
 DECAPx4_ASAP7_75t_R FILLER_154_589 ();
 FILLER_ASAP7_75t_R FILLER_154_599 ();
 FILLER_ASAP7_75t_R FILLER_154_604 ();
 DECAPx4_ASAP7_75t_R FILLER_154_612 ();
 DECAPx6_ASAP7_75t_R FILLER_154_625 ();
 DECAPx2_ASAP7_75t_R FILLER_154_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_645 ();
 FILLER_ASAP7_75t_R FILLER_154_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_684 ();
 DECAPx6_ASAP7_75t_R FILLER_154_693 ();
 DECAPx1_ASAP7_75t_R FILLER_154_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_711 ();
 FILLER_ASAP7_75t_R FILLER_154_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_756 ();
 DECAPx1_ASAP7_75t_R FILLER_154_765 ();
 DECAPx1_ASAP7_75t_R FILLER_154_777 ();
 DECAPx10_ASAP7_75t_R FILLER_154_807 ();
 DECAPx6_ASAP7_75t_R FILLER_154_829 ();
 FILLER_ASAP7_75t_R FILLER_154_843 ();
 DECAPx10_ASAP7_75t_R FILLER_154_853 ();
 DECAPx10_ASAP7_75t_R FILLER_154_875 ();
 DECAPx6_ASAP7_75t_R FILLER_154_897 ();
 FILLER_ASAP7_75t_R FILLER_154_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_920 ();
 FILLER_ASAP7_75t_R FILLER_154_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_963 ();
 DECAPx10_ASAP7_75t_R FILLER_154_972 ();
 DECAPx10_ASAP7_75t_R FILLER_154_994 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1038 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1050 ();
 FILLER_ASAP7_75t_R FILLER_154_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1175 ();
 FILLER_ASAP7_75t_R FILLER_154_1186 ();
 FILLER_ASAP7_75t_R FILLER_154_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1277 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1312 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1351 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1373 ();
 FILLER_ASAP7_75t_R FILLER_154_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1396 ();
 FILLER_ASAP7_75t_R FILLER_154_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_155_2 ();
 DECAPx2_ASAP7_75t_R FILLER_155_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_30 ();
 FILLER_ASAP7_75t_R FILLER_155_57 ();
 DECAPx2_ASAP7_75t_R FILLER_155_62 ();
 DECAPx6_ASAP7_75t_R FILLER_155_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_103 ();
 DECAPx6_ASAP7_75t_R FILLER_155_112 ();
 DECAPx1_ASAP7_75t_R FILLER_155_126 ();
 DECAPx4_ASAP7_75t_R FILLER_155_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_153 ();
 DECAPx1_ASAP7_75t_R FILLER_155_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_165 ();
 DECAPx4_ASAP7_75t_R FILLER_155_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_208 ();
 DECAPx4_ASAP7_75t_R FILLER_155_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_241 ();
 DECAPx1_ASAP7_75t_R FILLER_155_248 ();
 DECAPx10_ASAP7_75t_R FILLER_155_258 ();
 DECAPx2_ASAP7_75t_R FILLER_155_280 ();
 FILLER_ASAP7_75t_R FILLER_155_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_295 ();
 DECAPx1_ASAP7_75t_R FILLER_155_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_310 ();
 DECAPx10_ASAP7_75t_R FILLER_155_314 ();
 DECAPx10_ASAP7_75t_R FILLER_155_336 ();
 DECAPx10_ASAP7_75t_R FILLER_155_358 ();
 DECAPx10_ASAP7_75t_R FILLER_155_380 ();
 FILLER_ASAP7_75t_R FILLER_155_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_404 ();
 DECAPx10_ASAP7_75t_R FILLER_155_415 ();
 DECAPx1_ASAP7_75t_R FILLER_155_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_441 ();
 DECAPx6_ASAP7_75t_R FILLER_155_454 ();
 DECAPx1_ASAP7_75t_R FILLER_155_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_472 ();
 DECAPx10_ASAP7_75t_R FILLER_155_497 ();
 DECAPx6_ASAP7_75t_R FILLER_155_519 ();
 DECAPx1_ASAP7_75t_R FILLER_155_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_561 ();
 DECAPx10_ASAP7_75t_R FILLER_155_576 ();
 DECAPx1_ASAP7_75t_R FILLER_155_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_602 ();
 DECAPx2_ASAP7_75t_R FILLER_155_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_619 ();
 DECAPx4_ASAP7_75t_R FILLER_155_623 ();
 FILLER_ASAP7_75t_R FILLER_155_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_659 ();
 DECAPx4_ASAP7_75t_R FILLER_155_673 ();
 FILLER_ASAP7_75t_R FILLER_155_701 ();
 DECAPx4_ASAP7_75t_R FILLER_155_711 ();
 DECAPx6_ASAP7_75t_R FILLER_155_727 ();
 FILLER_ASAP7_75t_R FILLER_155_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_743 ();
 DECAPx1_ASAP7_75t_R FILLER_155_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_758 ();
 DECAPx1_ASAP7_75t_R FILLER_155_778 ();
 FILLER_ASAP7_75t_R FILLER_155_794 ();
 FILLER_ASAP7_75t_R FILLER_155_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_806 ();
 DECAPx6_ASAP7_75t_R FILLER_155_814 ();
 DECAPx6_ASAP7_75t_R FILLER_155_834 ();
 DECAPx10_ASAP7_75t_R FILLER_155_855 ();
 DECAPx2_ASAP7_75t_R FILLER_155_891 ();
 DECAPx6_ASAP7_75t_R FILLER_155_907 ();
 FILLER_ASAP7_75t_R FILLER_155_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_923 ();
 DECAPx4_ASAP7_75t_R FILLER_155_926 ();
 FILLER_ASAP7_75t_R FILLER_155_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_959 ();
 DECAPx2_ASAP7_75t_R FILLER_155_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_980 ();
 DECAPx4_ASAP7_75t_R FILLER_155_988 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1022 ();
 FILLER_ASAP7_75t_R FILLER_155_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1086 ();
 FILLER_ASAP7_75t_R FILLER_155_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1102 ();
 FILLER_ASAP7_75t_R FILLER_155_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1227 ();
 FILLER_ASAP7_75t_R FILLER_155_1238 ();
 FILLER_ASAP7_75t_R FILLER_155_1281 ();
 FILLER_ASAP7_75t_R FILLER_155_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1338 ();
 FILLER_ASAP7_75t_R FILLER_155_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_156_2 ();
 DECAPx6_ASAP7_75t_R FILLER_156_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_45 ();
 DECAPx6_ASAP7_75t_R FILLER_156_49 ();
 DECAPx2_ASAP7_75t_R FILLER_156_63 ();
 DECAPx4_ASAP7_75t_R FILLER_156_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_113 ();
 FILLER_ASAP7_75t_R FILLER_156_117 ();
 DECAPx10_ASAP7_75t_R FILLER_156_126 ();
 FILLER_ASAP7_75t_R FILLER_156_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_150 ();
 DECAPx4_ASAP7_75t_R FILLER_156_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_187 ();
 FILLER_ASAP7_75t_R FILLER_156_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_206 ();
 DECAPx2_ASAP7_75t_R FILLER_156_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_267 ();
 DECAPx1_ASAP7_75t_R FILLER_156_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_280 ();
 DECAPx4_ASAP7_75t_R FILLER_156_287 ();
 DECAPx10_ASAP7_75t_R FILLER_156_323 ();
 DECAPx6_ASAP7_75t_R FILLER_156_345 ();
 DECAPx1_ASAP7_75t_R FILLER_156_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_363 ();
 DECAPx4_ASAP7_75t_R FILLER_156_376 ();
 DECAPx6_ASAP7_75t_R FILLER_156_392 ();
 DECAPx1_ASAP7_75t_R FILLER_156_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_461 ();
 FILLER_ASAP7_75t_R FILLER_156_498 ();
 DECAPx1_ASAP7_75t_R FILLER_156_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_518 ();
 FILLER_ASAP7_75t_R FILLER_156_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_535 ();
 DECAPx4_ASAP7_75t_R FILLER_156_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_549 ();
 DECAPx6_ASAP7_75t_R FILLER_156_576 ();
 DECAPx2_ASAP7_75t_R FILLER_156_590 ();
 FILLER_ASAP7_75t_R FILLER_156_634 ();
 FILLER_ASAP7_75t_R FILLER_156_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_667 ();
 FILLER_ASAP7_75t_R FILLER_156_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_720 ();
 DECAPx10_ASAP7_75t_R FILLER_156_734 ();
 DECAPx10_ASAP7_75t_R FILLER_156_756 ();
 DECAPx6_ASAP7_75t_R FILLER_156_778 ();
 FILLER_ASAP7_75t_R FILLER_156_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_794 ();
 DECAPx4_ASAP7_75t_R FILLER_156_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_857 ();
 DECAPx2_ASAP7_75t_R FILLER_156_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_874 ();
 DECAPx4_ASAP7_75t_R FILLER_156_881 ();
 FILLER_ASAP7_75t_R FILLER_156_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_893 ();
 DECAPx10_ASAP7_75t_R FILLER_156_906 ();
 DECAPx4_ASAP7_75t_R FILLER_156_928 ();
 FILLER_ASAP7_75t_R FILLER_156_938 ();
 DECAPx6_ASAP7_75t_R FILLER_156_948 ();
 DECAPx2_ASAP7_75t_R FILLER_156_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1025 ();
 FILLER_ASAP7_75t_R FILLER_156_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1127 ();
 FILLER_ASAP7_75t_R FILLER_156_1148 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1199 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1255 ();
 FILLER_ASAP7_75t_R FILLER_156_1261 ();
 FILLER_ASAP7_75t_R FILLER_156_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1286 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1310 ();
 FILLER_ASAP7_75t_R FILLER_156_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1359 ();
 FILLER_ASAP7_75t_R FILLER_156_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1396 ();
 DECAPx6_ASAP7_75t_R FILLER_157_2 ();
 DECAPx2_ASAP7_75t_R FILLER_157_16 ();
 DECAPx2_ASAP7_75t_R FILLER_157_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_36 ();
 DECAPx2_ASAP7_75t_R FILLER_157_48 ();
 FILLER_ASAP7_75t_R FILLER_157_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_60 ();
 DECAPx6_ASAP7_75t_R FILLER_157_71 ();
 FILLER_ASAP7_75t_R FILLER_157_85 ();
 FILLER_ASAP7_75t_R FILLER_157_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_98 ();
 DECAPx1_ASAP7_75t_R FILLER_157_125 ();
 DECAPx6_ASAP7_75t_R FILLER_157_161 ();
 FILLER_ASAP7_75t_R FILLER_157_175 ();
 DECAPx10_ASAP7_75t_R FILLER_157_193 ();
 FILLER_ASAP7_75t_R FILLER_157_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_223 ();
 DECAPx2_ASAP7_75t_R FILLER_157_230 ();
 FILLER_ASAP7_75t_R FILLER_157_236 ();
 DECAPx10_ASAP7_75t_R FILLER_157_248 ();
 DECAPx4_ASAP7_75t_R FILLER_157_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_280 ();
 DECAPx4_ASAP7_75t_R FILLER_157_287 ();
 DECAPx4_ASAP7_75t_R FILLER_157_303 ();
 DECAPx2_ASAP7_75t_R FILLER_157_325 ();
 DECAPx1_ASAP7_75t_R FILLER_157_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_360 ();
 DECAPx2_ASAP7_75t_R FILLER_157_375 ();
 FILLER_ASAP7_75t_R FILLER_157_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_383 ();
 DECAPx10_ASAP7_75t_R FILLER_157_410 ();
 DECAPx2_ASAP7_75t_R FILLER_157_432 ();
 FILLER_ASAP7_75t_R FILLER_157_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_440 ();
 DECAPx6_ASAP7_75t_R FILLER_157_449 ();
 DECAPx2_ASAP7_75t_R FILLER_157_463 ();
 FILLER_ASAP7_75t_R FILLER_157_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_474 ();
 DECAPx2_ASAP7_75t_R FILLER_157_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_523 ();
 DECAPx2_ASAP7_75t_R FILLER_157_539 ();
 DECAPx4_ASAP7_75t_R FILLER_157_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_568 ();
 DECAPx10_ASAP7_75t_R FILLER_157_595 ();
 FILLER_ASAP7_75t_R FILLER_157_617 ();
 DECAPx6_ASAP7_75t_R FILLER_157_645 ();
 FILLER_ASAP7_75t_R FILLER_157_659 ();
 FILLER_ASAP7_75t_R FILLER_157_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_684 ();
 DECAPx2_ASAP7_75t_R FILLER_157_695 ();
 FILLER_ASAP7_75t_R FILLER_157_701 ();
 DECAPx1_ASAP7_75t_R FILLER_157_711 ();
 DECAPx1_ASAP7_75t_R FILLER_157_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_725 ();
 DECAPx6_ASAP7_75t_R FILLER_157_731 ();
 DECAPx1_ASAP7_75t_R FILLER_157_745 ();
 DECAPx2_ASAP7_75t_R FILLER_157_755 ();
 DECAPx10_ASAP7_75t_R FILLER_157_781 ();
 DECAPx2_ASAP7_75t_R FILLER_157_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_809 ();
 DECAPx1_ASAP7_75t_R FILLER_157_816 ();
 DECAPx2_ASAP7_75t_R FILLER_157_823 ();
 DECAPx10_ASAP7_75t_R FILLER_157_832 ();
 FILLER_ASAP7_75t_R FILLER_157_854 ();
 DECAPx1_ASAP7_75t_R FILLER_157_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_874 ();
 DECAPx2_ASAP7_75t_R FILLER_157_893 ();
 DECAPx6_ASAP7_75t_R FILLER_157_907 ();
 FILLER_ASAP7_75t_R FILLER_157_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_923 ();
 DECAPx4_ASAP7_75t_R FILLER_157_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_943 ();
 DECAPx2_ASAP7_75t_R FILLER_157_952 ();
 DECAPx1_ASAP7_75t_R FILLER_157_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_977 ();
 DECAPx2_ASAP7_75t_R FILLER_157_990 ();
 FILLER_ASAP7_75t_R FILLER_157_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1045 ();
 FILLER_ASAP7_75t_R FILLER_157_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1082 ();
 FILLER_ASAP7_75t_R FILLER_157_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1195 ();
 FILLER_ASAP7_75t_R FILLER_157_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1203 ();
 FILLER_ASAP7_75t_R FILLER_157_1220 ();
 FILLER_ASAP7_75t_R FILLER_157_1225 ();
 FILLER_ASAP7_75t_R FILLER_157_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1253 ();
 FILLER_ASAP7_75t_R FILLER_157_1275 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1297 ();
 FILLER_ASAP7_75t_R FILLER_157_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1327 ();
 FILLER_ASAP7_75t_R FILLER_157_1365 ();
 FILLER_ASAP7_75t_R FILLER_157_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1378 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1382 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1395 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1399 ();
 DECAPx6_ASAP7_75t_R FILLER_158_2 ();
 FILLER_ASAP7_75t_R FILLER_158_16 ();
 FILLER_ASAP7_75t_R FILLER_158_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_75 ();
 DECAPx2_ASAP7_75t_R FILLER_158_90 ();
 FILLER_ASAP7_75t_R FILLER_158_96 ();
 FILLER_ASAP7_75t_R FILLER_158_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_135 ();
 DECAPx1_ASAP7_75t_R FILLER_158_143 ();
 DECAPx10_ASAP7_75t_R FILLER_158_173 ();
 FILLER_ASAP7_75t_R FILLER_158_195 ();
 DECAPx10_ASAP7_75t_R FILLER_158_221 ();
 DECAPx10_ASAP7_75t_R FILLER_158_243 ();
 DECAPx2_ASAP7_75t_R FILLER_158_265 ();
 DECAPx10_ASAP7_75t_R FILLER_158_279 ();
 DECAPx10_ASAP7_75t_R FILLER_158_301 ();
 DECAPx2_ASAP7_75t_R FILLER_158_323 ();
 FILLER_ASAP7_75t_R FILLER_158_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_331 ();
 DECAPx2_ASAP7_75t_R FILLER_158_338 ();
 FILLER_ASAP7_75t_R FILLER_158_344 ();
 DECAPx1_ASAP7_75t_R FILLER_158_366 ();
 FILLER_ASAP7_75t_R FILLER_158_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_386 ();
 DECAPx1_ASAP7_75t_R FILLER_158_394 ();
 DECAPx4_ASAP7_75t_R FILLER_158_411 ();
 FILLER_ASAP7_75t_R FILLER_158_421 ();
 DECAPx6_ASAP7_75t_R FILLER_158_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_461 ();
 DECAPx6_ASAP7_75t_R FILLER_158_464 ();
 FILLER_ASAP7_75t_R FILLER_158_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_480 ();
 DECAPx2_ASAP7_75t_R FILLER_158_487 ();
 FILLER_ASAP7_75t_R FILLER_158_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_495 ();
 FILLER_ASAP7_75t_R FILLER_158_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_501 ();
 DECAPx6_ASAP7_75t_R FILLER_158_505 ();
 DECAPx2_ASAP7_75t_R FILLER_158_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_525 ();
 DECAPx2_ASAP7_75t_R FILLER_158_532 ();
 FILLER_ASAP7_75t_R FILLER_158_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_550 ();
 DECAPx4_ASAP7_75t_R FILLER_158_557 ();
 FILLER_ASAP7_75t_R FILLER_158_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_569 ();
 FILLER_ASAP7_75t_R FILLER_158_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_578 ();
 DECAPx2_ASAP7_75t_R FILLER_158_614 ();
 DECAPx2_ASAP7_75t_R FILLER_158_626 ();
 FILLER_ASAP7_75t_R FILLER_158_632 ();
 DECAPx10_ASAP7_75t_R FILLER_158_637 ();
 DECAPx10_ASAP7_75t_R FILLER_158_659 ();
 DECAPx10_ASAP7_75t_R FILLER_158_681 ();
 FILLER_ASAP7_75t_R FILLER_158_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_705 ();
 DECAPx2_ASAP7_75t_R FILLER_158_713 ();
 FILLER_ASAP7_75t_R FILLER_158_719 ();
 DECAPx1_ASAP7_75t_R FILLER_158_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_731 ();
 DECAPx2_ASAP7_75t_R FILLER_158_744 ();
 DECAPx2_ASAP7_75t_R FILLER_158_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_763 ();
 FILLER_ASAP7_75t_R FILLER_158_780 ();
 DECAPx6_ASAP7_75t_R FILLER_158_799 ();
 DECAPx2_ASAP7_75t_R FILLER_158_813 ();
 DECAPx6_ASAP7_75t_R FILLER_158_822 ();
 FILLER_ASAP7_75t_R FILLER_158_836 ();
 DECAPx10_ASAP7_75t_R FILLER_158_852 ();
 DECAPx10_ASAP7_75t_R FILLER_158_874 ();
 DECAPx6_ASAP7_75t_R FILLER_158_896 ();
 DECAPx2_ASAP7_75t_R FILLER_158_910 ();
 DECAPx6_ASAP7_75t_R FILLER_158_923 ();
 FILLER_ASAP7_75t_R FILLER_158_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_967 ();
 DECAPx10_ASAP7_75t_R FILLER_158_975 ();
 DECAPx6_ASAP7_75t_R FILLER_158_997 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1037 ();
 FILLER_ASAP7_75t_R FILLER_158_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1068 ();
 FILLER_ASAP7_75t_R FILLER_158_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1117 ();
 FILLER_ASAP7_75t_R FILLER_158_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1168 ();
 FILLER_ASAP7_75t_R FILLER_158_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1203 ();
 FILLER_ASAP7_75t_R FILLER_158_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1238 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1256 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1267 ();
 FILLER_ASAP7_75t_R FILLER_158_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1288 ();
 FILLER_ASAP7_75t_R FILLER_158_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1296 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1372 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_159_2 ();
 DECAPx6_ASAP7_75t_R FILLER_159_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_38 ();
 DECAPx10_ASAP7_75t_R FILLER_159_46 ();
 DECAPx4_ASAP7_75t_R FILLER_159_68 ();
 DECAPx2_ASAP7_75t_R FILLER_159_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_110 ();
 DECAPx4_ASAP7_75t_R FILLER_159_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_149 ();
 DECAPx10_ASAP7_75t_R FILLER_159_166 ();
 FILLER_ASAP7_75t_R FILLER_159_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_190 ();
 DECAPx4_ASAP7_75t_R FILLER_159_201 ();
 DECAPx2_ASAP7_75t_R FILLER_159_225 ();
 FILLER_ASAP7_75t_R FILLER_159_231 ();
 DECAPx4_ASAP7_75t_R FILLER_159_239 ();
 FILLER_ASAP7_75t_R FILLER_159_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_251 ();
 DECAPx10_ASAP7_75t_R FILLER_159_260 ();
 DECAPx4_ASAP7_75t_R FILLER_159_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_292 ();
 DECAPx10_ASAP7_75t_R FILLER_159_299 ();
 DECAPx2_ASAP7_75t_R FILLER_159_321 ();
 FILLER_ASAP7_75t_R FILLER_159_327 ();
 DECAPx10_ASAP7_75t_R FILLER_159_337 ();
 DECAPx10_ASAP7_75t_R FILLER_159_359 ();
 DECAPx10_ASAP7_75t_R FILLER_159_381 ();
 FILLER_ASAP7_75t_R FILLER_159_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_405 ();
 DECAPx2_ASAP7_75t_R FILLER_159_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_429 ();
 DECAPx2_ASAP7_75t_R FILLER_159_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_457 ();
 DECAPx10_ASAP7_75t_R FILLER_159_476 ();
 DECAPx4_ASAP7_75t_R FILLER_159_498 ();
 FILLER_ASAP7_75t_R FILLER_159_508 ();
 DECAPx2_ASAP7_75t_R FILLER_159_520 ();
 FILLER_ASAP7_75t_R FILLER_159_526 ();
 FILLER_ASAP7_75t_R FILLER_159_548 ();
 DECAPx6_ASAP7_75t_R FILLER_159_576 ();
 DECAPx2_ASAP7_75t_R FILLER_159_596 ();
 DECAPx10_ASAP7_75t_R FILLER_159_605 ();
 DECAPx1_ASAP7_75t_R FILLER_159_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_631 ();
 DECAPx1_ASAP7_75t_R FILLER_159_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_666 ();
 FILLER_ASAP7_75t_R FILLER_159_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_727 ();
 DECAPx4_ASAP7_75t_R FILLER_159_756 ();
 FILLER_ASAP7_75t_R FILLER_159_766 ();
 FILLER_ASAP7_75t_R FILLER_159_785 ();
 FILLER_ASAP7_75t_R FILLER_159_804 ();
 DECAPx1_ASAP7_75t_R FILLER_159_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_838 ();
 FILLER_ASAP7_75t_R FILLER_159_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_852 ();
 DECAPx10_ASAP7_75t_R FILLER_159_859 ();
 DECAPx10_ASAP7_75t_R FILLER_159_881 ();
 DECAPx6_ASAP7_75t_R FILLER_159_903 ();
 DECAPx2_ASAP7_75t_R FILLER_159_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_923 ();
 DECAPx6_ASAP7_75t_R FILLER_159_932 ();
 FILLER_ASAP7_75t_R FILLER_159_946 ();
 DECAPx2_ASAP7_75t_R FILLER_159_954 ();
 DECAPx2_ASAP7_75t_R FILLER_159_967 ();
 DECAPx1_ASAP7_75t_R FILLER_159_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_983 ();
 DECAPx4_ASAP7_75t_R FILLER_159_991 ();
 FILLER_ASAP7_75t_R FILLER_159_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1047 ();
 FILLER_ASAP7_75t_R FILLER_159_1069 ();
 FILLER_ASAP7_75t_R FILLER_159_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1104 ();
 FILLER_ASAP7_75t_R FILLER_159_1116 ();
 FILLER_ASAP7_75t_R FILLER_159_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1214 ();
 FILLER_ASAP7_75t_R FILLER_159_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1271 ();
 FILLER_ASAP7_75t_R FILLER_159_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1358 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_160_2 ();
 DECAPx2_ASAP7_75t_R FILLER_160_50 ();
 FILLER_ASAP7_75t_R FILLER_160_56 ();
 DECAPx2_ASAP7_75t_R FILLER_160_61 ();
 DECAPx6_ASAP7_75t_R FILLER_160_75 ();
 DECAPx10_ASAP7_75t_R FILLER_160_105 ();
 DECAPx10_ASAP7_75t_R FILLER_160_127 ();
 DECAPx10_ASAP7_75t_R FILLER_160_149 ();
 DECAPx2_ASAP7_75t_R FILLER_160_181 ();
 DECAPx1_ASAP7_75t_R FILLER_160_213 ();
 DECAPx1_ASAP7_75t_R FILLER_160_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_229 ();
 DECAPx2_ASAP7_75t_R FILLER_160_244 ();
 FILLER_ASAP7_75t_R FILLER_160_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_252 ();
 DECAPx10_ASAP7_75t_R FILLER_160_265 ();
 FILLER_ASAP7_75t_R FILLER_160_287 ();
 DECAPx6_ASAP7_75t_R FILLER_160_295 ();
 DECAPx4_ASAP7_75t_R FILLER_160_317 ();
 FILLER_ASAP7_75t_R FILLER_160_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_329 ();
 DECAPx2_ASAP7_75t_R FILLER_160_336 ();
 FILLER_ASAP7_75t_R FILLER_160_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_344 ();
 DECAPx10_ASAP7_75t_R FILLER_160_363 ();
 DECAPx1_ASAP7_75t_R FILLER_160_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_389 ();
 DECAPx10_ASAP7_75t_R FILLER_160_396 ();
 DECAPx6_ASAP7_75t_R FILLER_160_418 ();
 DECAPx2_ASAP7_75t_R FILLER_160_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_438 ();
 DECAPx6_ASAP7_75t_R FILLER_160_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_461 ();
 DECAPx2_ASAP7_75t_R FILLER_160_474 ();
 DECAPx10_ASAP7_75t_R FILLER_160_498 ();
 DECAPx6_ASAP7_75t_R FILLER_160_520 ();
 FILLER_ASAP7_75t_R FILLER_160_534 ();
 FILLER_ASAP7_75t_R FILLER_160_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_546 ();
 DECAPx4_ASAP7_75t_R FILLER_160_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_563 ();
 DECAPx4_ASAP7_75t_R FILLER_160_567 ();
 DECAPx10_ASAP7_75t_R FILLER_160_587 ();
 DECAPx2_ASAP7_75t_R FILLER_160_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_650 ();
 FILLER_ASAP7_75t_R FILLER_160_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_671 ();
 DECAPx10_ASAP7_75t_R FILLER_160_698 ();
 DECAPx2_ASAP7_75t_R FILLER_160_735 ();
 FILLER_ASAP7_75t_R FILLER_160_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_743 ();
 DECAPx2_ASAP7_75t_R FILLER_160_759 ();
 FILLER_ASAP7_75t_R FILLER_160_765 ();
 DECAPx4_ASAP7_75t_R FILLER_160_781 ();
 DECAPx2_ASAP7_75t_R FILLER_160_798 ();
 FILLER_ASAP7_75t_R FILLER_160_804 ();
 FILLER_ASAP7_75t_R FILLER_160_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_815 ();
 DECAPx4_ASAP7_75t_R FILLER_160_826 ();
 FILLER_ASAP7_75t_R FILLER_160_836 ();
 DECAPx1_ASAP7_75t_R FILLER_160_848 ();
 DECAPx2_ASAP7_75t_R FILLER_160_868 ();
 FILLER_ASAP7_75t_R FILLER_160_874 ();
 DECAPx1_ASAP7_75t_R FILLER_160_888 ();
 FILLER_ASAP7_75t_R FILLER_160_912 ();
 DECAPx6_ASAP7_75t_R FILLER_160_925 ();
 DECAPx1_ASAP7_75t_R FILLER_160_939 ();
 FILLER_ASAP7_75t_R FILLER_160_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_951 ();
 DECAPx4_ASAP7_75t_R FILLER_160_960 ();
 FILLER_ASAP7_75t_R FILLER_160_970 ();
 DECAPx1_ASAP7_75t_R FILLER_160_995 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1035 ();
 FILLER_ASAP7_75t_R FILLER_160_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1163 ();
 FILLER_ASAP7_75t_R FILLER_160_1174 ();
 FILLER_ASAP7_75t_R FILLER_160_1182 ();
 FILLER_ASAP7_75t_R FILLER_160_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1257 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1283 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1294 ();
 FILLER_ASAP7_75t_R FILLER_160_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1302 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1314 ();
 FILLER_ASAP7_75t_R FILLER_160_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1326 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1354 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1358 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1362 ();
 FILLER_ASAP7_75t_R FILLER_160_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_161_2 ();
 DECAPx1_ASAP7_75t_R FILLER_161_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_28 ();
 FILLER_ASAP7_75t_R FILLER_161_35 ();
 DECAPx2_ASAP7_75t_R FILLER_161_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_75 ();
 FILLER_ASAP7_75t_R FILLER_161_82 ();
 DECAPx4_ASAP7_75t_R FILLER_161_90 ();
 FILLER_ASAP7_75t_R FILLER_161_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_116 ();
 DECAPx2_ASAP7_75t_R FILLER_161_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_133 ();
 DECAPx1_ASAP7_75t_R FILLER_161_169 ();
 DECAPx2_ASAP7_75t_R FILLER_161_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_185 ();
 DECAPx2_ASAP7_75t_R FILLER_161_196 ();
 DECAPx1_ASAP7_75t_R FILLER_161_205 ();
 FILLER_ASAP7_75t_R FILLER_161_228 ();
 DECAPx10_ASAP7_75t_R FILLER_161_236 ();
 DECAPx4_ASAP7_75t_R FILLER_161_258 ();
 FILLER_ASAP7_75t_R FILLER_161_268 ();
 DECAPx10_ASAP7_75t_R FILLER_161_278 ();
 FILLER_ASAP7_75t_R FILLER_161_300 ();
 DECAPx6_ASAP7_75t_R FILLER_161_308 ();
 DECAPx1_ASAP7_75t_R FILLER_161_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_326 ();
 DECAPx6_ASAP7_75t_R FILLER_161_333 ();
 DECAPx1_ASAP7_75t_R FILLER_161_358 ();
 FILLER_ASAP7_75t_R FILLER_161_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_374 ();
 DECAPx1_ASAP7_75t_R FILLER_161_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_385 ();
 DECAPx6_ASAP7_75t_R FILLER_161_402 ();
 DECAPx1_ASAP7_75t_R FILLER_161_416 ();
 FILLER_ASAP7_75t_R FILLER_161_426 ();
 FILLER_ASAP7_75t_R FILLER_161_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_444 ();
 DECAPx6_ASAP7_75t_R FILLER_161_448 ();
 DECAPx1_ASAP7_75t_R FILLER_161_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_485 ();
 FILLER_ASAP7_75t_R FILLER_161_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_509 ();
 DECAPx10_ASAP7_75t_R FILLER_161_526 ();
 DECAPx6_ASAP7_75t_R FILLER_161_548 ();
 DECAPx1_ASAP7_75t_R FILLER_161_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_577 ();
 FILLER_ASAP7_75t_R FILLER_161_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_590 ();
 DECAPx4_ASAP7_75t_R FILLER_161_599 ();
 FILLER_ASAP7_75t_R FILLER_161_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_611 ();
 DECAPx4_ASAP7_75t_R FILLER_161_642 ();
 DECAPx4_ASAP7_75t_R FILLER_161_658 ();
 FILLER_ASAP7_75t_R FILLER_161_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_670 ();
 DECAPx10_ASAP7_75t_R FILLER_161_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_707 ();
 DECAPx10_ASAP7_75t_R FILLER_161_718 ();
 DECAPx1_ASAP7_75t_R FILLER_161_740 ();
 DECAPx1_ASAP7_75t_R FILLER_161_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_763 ();
 DECAPx6_ASAP7_75t_R FILLER_161_782 ();
 DECAPx4_ASAP7_75t_R FILLER_161_816 ();
 FILLER_ASAP7_75t_R FILLER_161_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_828 ();
 DECAPx1_ASAP7_75t_R FILLER_161_842 ();
 DECAPx6_ASAP7_75t_R FILLER_161_856 ();
 DECAPx2_ASAP7_75t_R FILLER_161_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_876 ();
 DECAPx2_ASAP7_75t_R FILLER_161_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_912 ();
 DECAPx1_ASAP7_75t_R FILLER_161_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_923 ();
 DECAPx2_ASAP7_75t_R FILLER_161_926 ();
 FILLER_ASAP7_75t_R FILLER_161_939 ();
 DECAPx2_ASAP7_75t_R FILLER_161_992 ();
 FILLER_ASAP7_75t_R FILLER_161_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1007 ();
 FILLER_ASAP7_75t_R FILLER_161_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1095 ();
 FILLER_ASAP7_75t_R FILLER_161_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_161_1148 ();
 FILLER_ASAP7_75t_R FILLER_161_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1177 ();
 FILLER_ASAP7_75t_R FILLER_161_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_161_1255 ();
 FILLER_ASAP7_75t_R FILLER_161_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1318 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1356 ();
 FILLER_ASAP7_75t_R FILLER_161_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1365 ();
 FILLER_ASAP7_75t_R FILLER_161_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1374 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1399 ();
 FILLER_ASAP7_75t_R FILLER_162_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_40 ();
 DECAPx4_ASAP7_75t_R FILLER_162_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_107 ();
 DECAPx6_ASAP7_75t_R FILLER_162_134 ();
 FILLER_ASAP7_75t_R FILLER_162_148 ();
 FILLER_ASAP7_75t_R FILLER_162_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_188 ();
 DECAPx10_ASAP7_75t_R FILLER_162_195 ();
 DECAPx2_ASAP7_75t_R FILLER_162_217 ();
 FILLER_ASAP7_75t_R FILLER_162_223 ();
 DECAPx10_ASAP7_75t_R FILLER_162_231 ();
 DECAPx10_ASAP7_75t_R FILLER_162_253 ();
 DECAPx10_ASAP7_75t_R FILLER_162_275 ();
 DECAPx2_ASAP7_75t_R FILLER_162_297 ();
 FILLER_ASAP7_75t_R FILLER_162_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_305 ();
 FILLER_ASAP7_75t_R FILLER_162_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_314 ();
 DECAPx4_ASAP7_75t_R FILLER_162_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_333 ();
 FILLER_ASAP7_75t_R FILLER_162_360 ();
 DECAPx6_ASAP7_75t_R FILLER_162_397 ();
 DECAPx2_ASAP7_75t_R FILLER_162_411 ();
 DECAPx4_ASAP7_75t_R FILLER_162_433 ();
 FILLER_ASAP7_75t_R FILLER_162_443 ();
 DECAPx2_ASAP7_75t_R FILLER_162_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_461 ();
 DECAPx6_ASAP7_75t_R FILLER_162_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_478 ();
 FILLER_ASAP7_75t_R FILLER_162_489 ();
 FILLER_ASAP7_75t_R FILLER_162_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_519 ();
 DECAPx2_ASAP7_75t_R FILLER_162_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_542 ();
 FILLER_ASAP7_75t_R FILLER_162_559 ();
 FILLER_ASAP7_75t_R FILLER_162_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_570 ();
 FILLER_ASAP7_75t_R FILLER_162_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_591 ();
 DECAPx2_ASAP7_75t_R FILLER_162_600 ();
 DECAPx2_ASAP7_75t_R FILLER_162_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_680 ();
 DECAPx10_ASAP7_75t_R FILLER_162_709 ();
 DECAPx2_ASAP7_75t_R FILLER_162_731 ();
 DECAPx4_ASAP7_75t_R FILLER_162_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_761 ();
 FILLER_ASAP7_75t_R FILLER_162_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_780 ();
 DECAPx10_ASAP7_75t_R FILLER_162_791 ();
 DECAPx2_ASAP7_75t_R FILLER_162_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_819 ();
 DECAPx2_ASAP7_75t_R FILLER_162_826 ();
 FILLER_ASAP7_75t_R FILLER_162_832 ();
 DECAPx2_ASAP7_75t_R FILLER_162_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_852 ();
 FILLER_ASAP7_75t_R FILLER_162_860 ();
 DECAPx10_ASAP7_75t_R FILLER_162_870 ();
 DECAPx10_ASAP7_75t_R FILLER_162_892 ();
 DECAPx10_ASAP7_75t_R FILLER_162_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_936 ();
 DECAPx10_ASAP7_75t_R FILLER_162_949 ();
 FILLER_ASAP7_75t_R FILLER_162_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_973 ();
 DECAPx10_ASAP7_75t_R FILLER_162_980 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1034 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1050 ();
 FILLER_ASAP7_75t_R FILLER_162_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1185 ();
 FILLER_ASAP7_75t_R FILLER_162_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1248 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1300 ();
 FILLER_ASAP7_75t_R FILLER_162_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1312 ();
 FILLER_ASAP7_75t_R FILLER_162_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1365 ();
 FILLER_ASAP7_75t_R FILLER_162_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1377 ();
 FILLER_ASAP7_75t_R FILLER_162_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1388 ();
 FILLER_ASAP7_75t_R FILLER_162_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_163_2 ();
 DECAPx1_ASAP7_75t_R FILLER_163_16 ();
 FILLER_ASAP7_75t_R FILLER_163_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_38 ();
 DECAPx1_ASAP7_75t_R FILLER_163_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_99 ();
 FILLER_ASAP7_75t_R FILLER_163_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_116 ();
 FILLER_ASAP7_75t_R FILLER_163_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_122 ();
 DECAPx1_ASAP7_75t_R FILLER_163_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_146 ();
 DECAPx6_ASAP7_75t_R FILLER_163_150 ();
 DECAPx1_ASAP7_75t_R FILLER_163_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_168 ();
 DECAPx2_ASAP7_75t_R FILLER_163_179 ();
 FILLER_ASAP7_75t_R FILLER_163_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_187 ();
 FILLER_ASAP7_75t_R FILLER_163_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_198 ();
 FILLER_ASAP7_75t_R FILLER_163_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_220 ();
 FILLER_ASAP7_75t_R FILLER_163_235 ();
 DECAPx10_ASAP7_75t_R FILLER_163_257 ();
 DECAPx10_ASAP7_75t_R FILLER_163_279 ();
 DECAPx10_ASAP7_75t_R FILLER_163_301 ();
 DECAPx6_ASAP7_75t_R FILLER_163_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_337 ();
 DECAPx1_ASAP7_75t_R FILLER_163_345 ();
 DECAPx6_ASAP7_75t_R FILLER_163_352 ();
 FILLER_ASAP7_75t_R FILLER_163_366 ();
 FILLER_ASAP7_75t_R FILLER_163_375 ();
 DECAPx6_ASAP7_75t_R FILLER_163_380 ();
 FILLER_ASAP7_75t_R FILLER_163_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_396 ();
 DECAPx1_ASAP7_75t_R FILLER_163_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_418 ();
 DECAPx4_ASAP7_75t_R FILLER_163_431 ();
 FILLER_ASAP7_75t_R FILLER_163_441 ();
 DECAPx10_ASAP7_75t_R FILLER_163_469 ();
 DECAPx2_ASAP7_75t_R FILLER_163_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_504 ();
 DECAPx2_ASAP7_75t_R FILLER_163_508 ();
 FILLER_ASAP7_75t_R FILLER_163_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_516 ();
 DECAPx2_ASAP7_75t_R FILLER_163_529 ();
 DECAPx2_ASAP7_75t_R FILLER_163_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_583 ();
 DECAPx2_ASAP7_75t_R FILLER_163_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_606 ();
 DECAPx4_ASAP7_75t_R FILLER_163_615 ();
 DECAPx10_ASAP7_75t_R FILLER_163_665 ();
 FILLER_ASAP7_75t_R FILLER_163_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_689 ();
 DECAPx6_ASAP7_75t_R FILLER_163_696 ();
 DECAPx2_ASAP7_75t_R FILLER_163_710 ();
 FILLER_ASAP7_75t_R FILLER_163_735 ();
 DECAPx2_ASAP7_75t_R FILLER_163_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_780 ();
 DECAPx1_ASAP7_75t_R FILLER_163_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_791 ();
 DECAPx2_ASAP7_75t_R FILLER_163_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_804 ();
 DECAPx2_ASAP7_75t_R FILLER_163_811 ();
 FILLER_ASAP7_75t_R FILLER_163_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_835 ();
 DECAPx6_ASAP7_75t_R FILLER_163_842 ();
 FILLER_ASAP7_75t_R FILLER_163_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_858 ();
 FILLER_ASAP7_75t_R FILLER_163_875 ();
 DECAPx10_ASAP7_75t_R FILLER_163_887 ();
 DECAPx2_ASAP7_75t_R FILLER_163_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_923 ();
 DECAPx2_ASAP7_75t_R FILLER_163_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_932 ();
 DECAPx1_ASAP7_75t_R FILLER_163_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_955 ();
 DECAPx4_ASAP7_75t_R FILLER_163_962 ();
 DECAPx2_ASAP7_75t_R FILLER_163_979 ();
 FILLER_ASAP7_75t_R FILLER_163_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_987 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1116 ();
 FILLER_ASAP7_75t_R FILLER_163_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1132 ();
 FILLER_ASAP7_75t_R FILLER_163_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1177 ();
 FILLER_ASAP7_75t_R FILLER_163_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1237 ();
 FILLER_ASAP7_75t_R FILLER_163_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1291 ();
 FILLER_ASAP7_75t_R FILLER_163_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1299 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1339 ();
 FILLER_ASAP7_75t_R FILLER_163_1361 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1366 ();
 FILLER_ASAP7_75t_R FILLER_163_1376 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_164_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_8 ();
 FILLER_ASAP7_75t_R FILLER_164_67 ();
 FILLER_ASAP7_75t_R FILLER_164_75 ();
 DECAPx1_ASAP7_75t_R FILLER_164_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_84 ();
 DECAPx2_ASAP7_75t_R FILLER_164_111 ();
 FILLER_ASAP7_75t_R FILLER_164_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_132 ();
 DECAPx6_ASAP7_75t_R FILLER_164_159 ();
 DECAPx1_ASAP7_75t_R FILLER_164_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_177 ();
 DECAPx4_ASAP7_75t_R FILLER_164_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_217 ();
 DECAPx6_ASAP7_75t_R FILLER_164_234 ();
 DECAPx2_ASAP7_75t_R FILLER_164_248 ();
 DECAPx1_ASAP7_75t_R FILLER_164_261 ();
 DECAPx1_ASAP7_75t_R FILLER_164_271 ();
 DECAPx2_ASAP7_75t_R FILLER_164_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_289 ();
 DECAPx10_ASAP7_75t_R FILLER_164_302 ();
 DECAPx6_ASAP7_75t_R FILLER_164_332 ();
 DECAPx2_ASAP7_75t_R FILLER_164_352 ();
 FILLER_ASAP7_75t_R FILLER_164_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_360 ();
 DECAPx10_ASAP7_75t_R FILLER_164_364 ();
 DECAPx4_ASAP7_75t_R FILLER_164_386 ();
 DECAPx10_ASAP7_75t_R FILLER_164_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_427 ();
 FILLER_ASAP7_75t_R FILLER_164_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_433 ();
 DECAPx2_ASAP7_75t_R FILLER_164_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_447 ();
 DECAPx2_ASAP7_75t_R FILLER_164_454 ();
 FILLER_ASAP7_75t_R FILLER_164_460 ();
 DECAPx1_ASAP7_75t_R FILLER_164_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_468 ();
 FILLER_ASAP7_75t_R FILLER_164_479 ();
 FILLER_ASAP7_75t_R FILLER_164_484 ();
 DECAPx4_ASAP7_75t_R FILLER_164_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_504 ();
 DECAPx2_ASAP7_75t_R FILLER_164_518 ();
 DECAPx10_ASAP7_75t_R FILLER_164_534 ();
 DECAPx1_ASAP7_75t_R FILLER_164_556 ();
 DECAPx10_ASAP7_75t_R FILLER_164_563 ();
 DECAPx2_ASAP7_75t_R FILLER_164_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_591 ();
 DECAPx6_ASAP7_75t_R FILLER_164_600 ();
 FILLER_ASAP7_75t_R FILLER_164_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_616 ();
 DECAPx6_ASAP7_75t_R FILLER_164_627 ();
 DECAPx1_ASAP7_75t_R FILLER_164_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_653 ();
 DECAPx6_ASAP7_75t_R FILLER_164_660 ();
 FILLER_ASAP7_75t_R FILLER_164_674 ();
 DECAPx1_ASAP7_75t_R FILLER_164_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_710 ();
 DECAPx4_ASAP7_75t_R FILLER_164_731 ();
 FILLER_ASAP7_75t_R FILLER_164_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_743 ();
 FILLER_ASAP7_75t_R FILLER_164_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_754 ();
 DECAPx10_ASAP7_75t_R FILLER_164_761 ();
 DECAPx6_ASAP7_75t_R FILLER_164_783 ();
 DECAPx1_ASAP7_75t_R FILLER_164_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_801 ();
 DECAPx6_ASAP7_75t_R FILLER_164_805 ();
 FILLER_ASAP7_75t_R FILLER_164_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_821 ();
 FILLER_ASAP7_75t_R FILLER_164_828 ();
 DECAPx2_ASAP7_75t_R FILLER_164_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_916 ();
 DECAPx1_ASAP7_75t_R FILLER_164_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_937 ();
 DECAPx2_ASAP7_75t_R FILLER_164_953 ();
 FILLER_ASAP7_75t_R FILLER_164_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_979 ();
 FILLER_ASAP7_75t_R FILLER_164_995 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1030 ();
 FILLER_ASAP7_75t_R FILLER_164_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1073 ();
 FILLER_ASAP7_75t_R FILLER_164_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1095 ();
 FILLER_ASAP7_75t_R FILLER_164_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1116 ();
 FILLER_ASAP7_75t_R FILLER_164_1126 ();
 FILLER_ASAP7_75t_R FILLER_164_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1158 ();
 FILLER_ASAP7_75t_R FILLER_164_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1164 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1209 ();
 FILLER_ASAP7_75t_R FILLER_164_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1317 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1339 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1401 ();
 DECAPx10_ASAP7_75t_R FILLER_165_2 ();
 DECAPx1_ASAP7_75t_R FILLER_165_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_37 ();
 DECAPx1_ASAP7_75t_R FILLER_165_41 ();
 DECAPx1_ASAP7_75t_R FILLER_165_51 ();
 DECAPx2_ASAP7_75t_R FILLER_165_58 ();
 DECAPx10_ASAP7_75t_R FILLER_165_67 ();
 DECAPx1_ASAP7_75t_R FILLER_165_89 ();
 DECAPx10_ASAP7_75t_R FILLER_165_147 ();
 DECAPx6_ASAP7_75t_R FILLER_165_169 ();
 FILLER_ASAP7_75t_R FILLER_165_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_206 ();
 DECAPx2_ASAP7_75t_R FILLER_165_213 ();
 FILLER_ASAP7_75t_R FILLER_165_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_221 ();
 DECAPx2_ASAP7_75t_R FILLER_165_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_261 ();
 DECAPx4_ASAP7_75t_R FILLER_165_276 ();
 DECAPx4_ASAP7_75t_R FILLER_165_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_308 ();
 DECAPx2_ASAP7_75t_R FILLER_165_335 ();
 DECAPx4_ASAP7_75t_R FILLER_165_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_383 ();
 DECAPx1_ASAP7_75t_R FILLER_165_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_398 ();
 DECAPx2_ASAP7_75t_R FILLER_165_419 ();
 FILLER_ASAP7_75t_R FILLER_165_425 ();
 DECAPx2_ASAP7_75t_R FILLER_165_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_465 ();
 DECAPx2_ASAP7_75t_R FILLER_165_527 ();
 FILLER_ASAP7_75t_R FILLER_165_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_535 ();
 DECAPx4_ASAP7_75t_R FILLER_165_566 ();
 DECAPx4_ASAP7_75t_R FILLER_165_586 ();
 FILLER_ASAP7_75t_R FILLER_165_596 ();
 FILLER_ASAP7_75t_R FILLER_165_605 ();
 DECAPx1_ASAP7_75t_R FILLER_165_614 ();
 DECAPx10_ASAP7_75t_R FILLER_165_628 ();
 DECAPx1_ASAP7_75t_R FILLER_165_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_670 ();
 DECAPx4_ASAP7_75t_R FILLER_165_697 ();
 FILLER_ASAP7_75t_R FILLER_165_707 ();
 DECAPx10_ASAP7_75t_R FILLER_165_714 ();
 DECAPx10_ASAP7_75t_R FILLER_165_736 ();
 DECAPx2_ASAP7_75t_R FILLER_165_758 ();
 DECAPx4_ASAP7_75t_R FILLER_165_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_781 ();
 DECAPx2_ASAP7_75t_R FILLER_165_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_794 ();
 DECAPx2_ASAP7_75t_R FILLER_165_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_817 ();
 DECAPx1_ASAP7_75t_R FILLER_165_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_832 ();
 DECAPx2_ASAP7_75t_R FILLER_165_855 ();
 DECAPx1_ASAP7_75t_R FILLER_165_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_879 ();
 DECAPx2_ASAP7_75t_R FILLER_165_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_896 ();
 DECAPx1_ASAP7_75t_R FILLER_165_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_923 ();
 FILLER_ASAP7_75t_R FILLER_165_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_942 ();
 DECAPx10_ASAP7_75t_R FILLER_165_989 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1023 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1043 ();
 FILLER_ASAP7_75t_R FILLER_165_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1078 ();
 FILLER_ASAP7_75t_R FILLER_165_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1134 ();
 FILLER_ASAP7_75t_R FILLER_165_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1159 ();
 FILLER_ASAP7_75t_R FILLER_165_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1225 ();
 FILLER_ASAP7_75t_R FILLER_165_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1233 ();
 FILLER_ASAP7_75t_R FILLER_165_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1262 ();
 FILLER_ASAP7_75t_R FILLER_165_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1280 ();
 FILLER_ASAP7_75t_R FILLER_165_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1293 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1361 ();
 FILLER_ASAP7_75t_R FILLER_165_1383 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1391 ();
 DECAPx6_ASAP7_75t_R FILLER_166_2 ();
 DECAPx1_ASAP7_75t_R FILLER_166_16 ();
 DECAPx2_ASAP7_75t_R FILLER_166_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_34 ();
 DECAPx6_ASAP7_75t_R FILLER_166_45 ();
 FILLER_ASAP7_75t_R FILLER_166_59 ();
 FILLER_ASAP7_75t_R FILLER_166_71 ();
 DECAPx1_ASAP7_75t_R FILLER_166_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_89 ();
 DECAPx2_ASAP7_75t_R FILLER_166_93 ();
 DECAPx2_ASAP7_75t_R FILLER_166_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_108 ();
 DECAPx2_ASAP7_75t_R FILLER_166_112 ();
 FILLER_ASAP7_75t_R FILLER_166_118 ();
 DECAPx6_ASAP7_75t_R FILLER_166_123 ();
 FILLER_ASAP7_75t_R FILLER_166_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_152 ();
 FILLER_ASAP7_75t_R FILLER_166_156 ();
 FILLER_ASAP7_75t_R FILLER_166_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_177 ();
 DECAPx2_ASAP7_75t_R FILLER_166_181 ();
 FILLER_ASAP7_75t_R FILLER_166_201 ();
 DECAPx10_ASAP7_75t_R FILLER_166_217 ();
 DECAPx4_ASAP7_75t_R FILLER_166_239 ();
 DECAPx1_ASAP7_75t_R FILLER_166_252 ();
 DECAPx10_ASAP7_75t_R FILLER_166_262 ();
 DECAPx4_ASAP7_75t_R FILLER_166_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_294 ();
 DECAPx1_ASAP7_75t_R FILLER_166_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_305 ();
 DECAPx2_ASAP7_75t_R FILLER_166_316 ();
 FILLER_ASAP7_75t_R FILLER_166_322 ();
 DECAPx2_ASAP7_75t_R FILLER_166_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_339 ();
 DECAPx10_ASAP7_75t_R FILLER_166_346 ();
 DECAPx6_ASAP7_75t_R FILLER_166_374 ();
 DECAPx1_ASAP7_75t_R FILLER_166_388 ();
 DECAPx2_ASAP7_75t_R FILLER_166_400 ();
 FILLER_ASAP7_75t_R FILLER_166_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_408 ();
 DECAPx2_ASAP7_75t_R FILLER_166_417 ();
 FILLER_ASAP7_75t_R FILLER_166_423 ();
 DECAPx2_ASAP7_75t_R FILLER_166_439 ();
 FILLER_ASAP7_75t_R FILLER_166_445 ();
 DECAPx4_ASAP7_75t_R FILLER_166_450 ();
 FILLER_ASAP7_75t_R FILLER_166_460 ();
 DECAPx10_ASAP7_75t_R FILLER_166_480 ();
 DECAPx6_ASAP7_75t_R FILLER_166_502 ();
 DECAPx10_ASAP7_75t_R FILLER_166_519 ();
 DECAPx10_ASAP7_75t_R FILLER_166_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_573 ();
 FILLER_ASAP7_75t_R FILLER_166_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_596 ();
 DECAPx6_ASAP7_75t_R FILLER_166_635 ();
 FILLER_ASAP7_75t_R FILLER_166_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_651 ();
 FILLER_ASAP7_75t_R FILLER_166_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_660 ();
 FILLER_ASAP7_75t_R FILLER_166_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_673 ();
 DECAPx10_ASAP7_75t_R FILLER_166_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_706 ();
 DECAPx10_ASAP7_75t_R FILLER_166_717 ();
 DECAPx10_ASAP7_75t_R FILLER_166_739 ();
 FILLER_ASAP7_75t_R FILLER_166_761 ();
 DECAPx4_ASAP7_75t_R FILLER_166_792 ();
 DECAPx10_ASAP7_75t_R FILLER_166_810 ();
 DECAPx1_ASAP7_75t_R FILLER_166_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_836 ();
 DECAPx6_ASAP7_75t_R FILLER_166_843 ();
 DECAPx1_ASAP7_75t_R FILLER_166_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_861 ();
 DECAPx6_ASAP7_75t_R FILLER_166_868 ();
 DECAPx2_ASAP7_75t_R FILLER_166_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_888 ();
 FILLER_ASAP7_75t_R FILLER_166_901 ();
 DECAPx1_ASAP7_75t_R FILLER_166_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_933 ();
 DECAPx6_ASAP7_75t_R FILLER_166_942 ();
 FILLER_ASAP7_75t_R FILLER_166_956 ();
 DECAPx4_ASAP7_75t_R FILLER_166_964 ();
 FILLER_ASAP7_75t_R FILLER_166_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_976 ();
 DECAPx6_ASAP7_75t_R FILLER_166_987 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1045 ();
 FILLER_ASAP7_75t_R FILLER_166_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1079 ();
 FILLER_ASAP7_75t_R FILLER_166_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1131 ();
 FILLER_ASAP7_75t_R FILLER_166_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1200 ();
 FILLER_ASAP7_75t_R FILLER_166_1206 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1302 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1317 ();
 FILLER_ASAP7_75t_R FILLER_166_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1366 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1385 ();
 FILLER_ASAP7_75t_R FILLER_166_1394 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1399 ();
 DECAPx6_ASAP7_75t_R FILLER_167_2 ();
 FILLER_ASAP7_75t_R FILLER_167_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_18 ();
 FILLER_ASAP7_75t_R FILLER_167_33 ();
 FILLER_ASAP7_75t_R FILLER_167_45 ();
 FILLER_ASAP7_75t_R FILLER_167_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_63 ();
 FILLER_ASAP7_75t_R FILLER_167_90 ();
 DECAPx10_ASAP7_75t_R FILLER_167_102 ();
 DECAPx4_ASAP7_75t_R FILLER_167_124 ();
 FILLER_ASAP7_75t_R FILLER_167_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_136 ();
 DECAPx2_ASAP7_75t_R FILLER_167_199 ();
 FILLER_ASAP7_75t_R FILLER_167_205 ();
 DECAPx2_ASAP7_75t_R FILLER_167_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_223 ();
 DECAPx6_ASAP7_75t_R FILLER_167_244 ();
 DECAPx1_ASAP7_75t_R FILLER_167_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_269 ();
 DECAPx1_ASAP7_75t_R FILLER_167_284 ();
 DECAPx10_ASAP7_75t_R FILLER_167_314 ();
 DECAPx2_ASAP7_75t_R FILLER_167_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_342 ();
 DECAPx6_ASAP7_75t_R FILLER_167_351 ();
 DECAPx1_ASAP7_75t_R FILLER_167_365 ();
 DECAPx10_ASAP7_75t_R FILLER_167_377 ();
 DECAPx10_ASAP7_75t_R FILLER_167_399 ();
 FILLER_ASAP7_75t_R FILLER_167_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_423 ();
 DECAPx10_ASAP7_75t_R FILLER_167_440 ();
 DECAPx10_ASAP7_75t_R FILLER_167_462 ();
 DECAPx10_ASAP7_75t_R FILLER_167_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_514 ();
 DECAPx10_ASAP7_75t_R FILLER_167_525 ();
 DECAPx2_ASAP7_75t_R FILLER_167_557 ();
 FILLER_ASAP7_75t_R FILLER_167_563 ();
 DECAPx4_ASAP7_75t_R FILLER_167_573 ();
 FILLER_ASAP7_75t_R FILLER_167_583 ();
 DECAPx6_ASAP7_75t_R FILLER_167_609 ();
 FILLER_ASAP7_75t_R FILLER_167_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_625 ();
 DECAPx1_ASAP7_75t_R FILLER_167_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_640 ();
 DECAPx10_ASAP7_75t_R FILLER_167_671 ();
 DECAPx4_ASAP7_75t_R FILLER_167_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_703 ();
 DECAPx1_ASAP7_75t_R FILLER_167_719 ();
 DECAPx4_ASAP7_75t_R FILLER_167_731 ();
 FILLER_ASAP7_75t_R FILLER_167_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_743 ();
 DECAPx2_ASAP7_75t_R FILLER_167_752 ();
 FILLER_ASAP7_75t_R FILLER_167_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_760 ();
 FILLER_ASAP7_75t_R FILLER_167_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_778 ();
 FILLER_ASAP7_75t_R FILLER_167_786 ();
 DECAPx10_ASAP7_75t_R FILLER_167_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_824 ();
 DECAPx4_ASAP7_75t_R FILLER_167_845 ();
 FILLER_ASAP7_75t_R FILLER_167_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_866 ();
 DECAPx1_ASAP7_75t_R FILLER_167_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_926 ();
 FILLER_ASAP7_75t_R FILLER_167_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_937 ();
 DECAPx6_ASAP7_75t_R FILLER_167_946 ();
 DECAPx2_ASAP7_75t_R FILLER_167_960 ();
 DECAPx6_ASAP7_75t_R FILLER_167_973 ();
 DECAPx1_ASAP7_75t_R FILLER_167_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_998 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1064 ();
 FILLER_ASAP7_75t_R FILLER_167_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1125 ();
 FILLER_ASAP7_75t_R FILLER_167_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1192 ();
 FILLER_ASAP7_75t_R FILLER_167_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1236 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1259 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1315 ();
 FILLER_ASAP7_75t_R FILLER_167_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1323 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1343 ();
 FILLER_ASAP7_75t_R FILLER_167_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1361 ();
 DECAPx6_ASAP7_75t_R FILLER_168_2 ();
 FILLER_ASAP7_75t_R FILLER_168_16 ();
 DECAPx2_ASAP7_75t_R FILLER_168_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_46 ();
 DECAPx2_ASAP7_75t_R FILLER_168_57 ();
 FILLER_ASAP7_75t_R FILLER_168_63 ();
 FILLER_ASAP7_75t_R FILLER_168_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_77 ();
 DECAPx2_ASAP7_75t_R FILLER_168_81 ();
 FILLER_ASAP7_75t_R FILLER_168_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_128 ();
 DECAPx1_ASAP7_75t_R FILLER_168_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_136 ();
 DECAPx6_ASAP7_75t_R FILLER_168_143 ();
 DECAPx1_ASAP7_75t_R FILLER_168_157 ();
 DECAPx10_ASAP7_75t_R FILLER_168_177 ();
 DECAPx6_ASAP7_75t_R FILLER_168_199 ();
 FILLER_ASAP7_75t_R FILLER_168_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_215 ();
 DECAPx4_ASAP7_75t_R FILLER_168_230 ();
 DECAPx2_ASAP7_75t_R FILLER_168_254 ();
 FILLER_ASAP7_75t_R FILLER_168_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_268 ();
 DECAPx10_ASAP7_75t_R FILLER_168_277 ();
 FILLER_ASAP7_75t_R FILLER_168_299 ();
 FILLER_ASAP7_75t_R FILLER_168_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_312 ();
 DECAPx10_ASAP7_75t_R FILLER_168_316 ();
 DECAPx10_ASAP7_75t_R FILLER_168_338 ();
 DECAPx10_ASAP7_75t_R FILLER_168_360 ();
 DECAPx2_ASAP7_75t_R FILLER_168_382 ();
 FILLER_ASAP7_75t_R FILLER_168_388 ();
 FILLER_ASAP7_75t_R FILLER_168_396 ();
 DECAPx10_ASAP7_75t_R FILLER_168_404 ();
 DECAPx6_ASAP7_75t_R FILLER_168_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_440 ();
 FILLER_ASAP7_75t_R FILLER_168_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_461 ();
 DECAPx4_ASAP7_75t_R FILLER_168_467 ();
 FILLER_ASAP7_75t_R FILLER_168_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_483 ();
 DECAPx1_ASAP7_75t_R FILLER_168_490 ();
 DECAPx2_ASAP7_75t_R FILLER_168_530 ();
 FILLER_ASAP7_75t_R FILLER_168_536 ();
 DECAPx2_ASAP7_75t_R FILLER_168_562 ();
 FILLER_ASAP7_75t_R FILLER_168_592 ();
 DECAPx6_ASAP7_75t_R FILLER_168_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_623 ();
 DECAPx4_ASAP7_75t_R FILLER_168_638 ();
 FILLER_ASAP7_75t_R FILLER_168_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_658 ();
 FILLER_ASAP7_75t_R FILLER_168_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_719 ();
 DECAPx1_ASAP7_75t_R FILLER_168_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_730 ();
 DECAPx4_ASAP7_75t_R FILLER_168_739 ();
 FILLER_ASAP7_75t_R FILLER_168_749 ();
 FILLER_ASAP7_75t_R FILLER_168_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_786 ();
 DECAPx6_ASAP7_75t_R FILLER_168_790 ();
 DECAPx1_ASAP7_75t_R FILLER_168_804 ();
 DECAPx2_ASAP7_75t_R FILLER_168_822 ();
 DECAPx6_ASAP7_75t_R FILLER_168_841 ();
 DECAPx10_ASAP7_75t_R FILLER_168_895 ();
 DECAPx10_ASAP7_75t_R FILLER_168_923 ();
 DECAPx4_ASAP7_75t_R FILLER_168_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_955 ();
 FILLER_ASAP7_75t_R FILLER_168_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_964 ();
 DECAPx2_ASAP7_75t_R FILLER_168_980 ();
 FILLER_ASAP7_75t_R FILLER_168_986 ();
 DECAPx1_ASAP7_75t_R FILLER_168_994 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1022 ();
 FILLER_ASAP7_75t_R FILLER_168_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1075 ();
 FILLER_ASAP7_75t_R FILLER_168_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1160 ();
 FILLER_ASAP7_75t_R FILLER_168_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1209 ();
 FILLER_ASAP7_75t_R FILLER_168_1220 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1277 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1292 ();
 FILLER_ASAP7_75t_R FILLER_168_1302 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1310 ();
 FILLER_ASAP7_75t_R FILLER_168_1320 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1328 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1338 ();
 FILLER_ASAP7_75t_R FILLER_168_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1354 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1368 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1398 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_169_2 ();
 DECAPx10_ASAP7_75t_R FILLER_169_24 ();
 DECAPx2_ASAP7_75t_R FILLER_169_46 ();
 FILLER_ASAP7_75t_R FILLER_169_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_54 ();
 DECAPx10_ASAP7_75t_R FILLER_169_65 ();
 DECAPx10_ASAP7_75t_R FILLER_169_87 ();
 DECAPx2_ASAP7_75t_R FILLER_169_109 ();
 DECAPx4_ASAP7_75t_R FILLER_169_156 ();
 FILLER_ASAP7_75t_R FILLER_169_166 ();
 DECAPx1_ASAP7_75t_R FILLER_169_194 ();
 DECAPx6_ASAP7_75t_R FILLER_169_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_263 ();
 FILLER_ASAP7_75t_R FILLER_169_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_281 ();
 DECAPx10_ASAP7_75t_R FILLER_169_288 ();
 FILLER_ASAP7_75t_R FILLER_169_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_312 ();
 DECAPx2_ASAP7_75t_R FILLER_169_341 ();
 FILLER_ASAP7_75t_R FILLER_169_347 ();
 DECAPx2_ASAP7_75t_R FILLER_169_361 ();
 DECAPx1_ASAP7_75t_R FILLER_169_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_392 ();
 DECAPx2_ASAP7_75t_R FILLER_169_422 ();
 FILLER_ASAP7_75t_R FILLER_169_428 ();
 DECAPx2_ASAP7_75t_R FILLER_169_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_529 ();
 DECAPx1_ASAP7_75t_R FILLER_169_544 ();
 DECAPx2_ASAP7_75t_R FILLER_169_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_563 ();
 DECAPx10_ASAP7_75t_R FILLER_169_572 ();
 DECAPx1_ASAP7_75t_R FILLER_169_594 ();
 DECAPx2_ASAP7_75t_R FILLER_169_604 ();
 FILLER_ASAP7_75t_R FILLER_169_610 ();
 DECAPx1_ASAP7_75t_R FILLER_169_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_632 ();
 DECAPx6_ASAP7_75t_R FILLER_169_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_655 ();
 DECAPx1_ASAP7_75t_R FILLER_169_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_680 ();
 DECAPx2_ASAP7_75t_R FILLER_169_701 ();
 FILLER_ASAP7_75t_R FILLER_169_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_712 ();
 DECAPx4_ASAP7_75t_R FILLER_169_723 ();
 FILLER_ASAP7_75t_R FILLER_169_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_743 ();
 DECAPx10_ASAP7_75t_R FILLER_169_766 ();
 DECAPx1_ASAP7_75t_R FILLER_169_788 ();
 DECAPx6_ASAP7_75t_R FILLER_169_820 ();
 DECAPx2_ASAP7_75t_R FILLER_169_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_840 ();
 DECAPx6_ASAP7_75t_R FILLER_169_861 ();
 FILLER_ASAP7_75t_R FILLER_169_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_877 ();
 DECAPx6_ASAP7_75t_R FILLER_169_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_900 ();
 FILLER_ASAP7_75t_R FILLER_169_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_911 ();
 FILLER_ASAP7_75t_R FILLER_169_926 ();
 FILLER_ASAP7_75t_R FILLER_169_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_947 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1008 ();
 FILLER_ASAP7_75t_R FILLER_169_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1032 ();
 FILLER_ASAP7_75t_R FILLER_169_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1066 ();
 FILLER_ASAP7_75t_R FILLER_169_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1075 ();
 FILLER_ASAP7_75t_R FILLER_169_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1221 ();
 FILLER_ASAP7_75t_R FILLER_169_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1292 ();
 FILLER_ASAP7_75t_R FILLER_169_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1347 ();
 FILLER_ASAP7_75t_R FILLER_169_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1368 ();
 DECAPx4_ASAP7_75t_R FILLER_170_2 ();
 FILLER_ASAP7_75t_R FILLER_170_12 ();
 DECAPx10_ASAP7_75t_R FILLER_170_40 ();
 FILLER_ASAP7_75t_R FILLER_170_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_90 ();
 FILLER_ASAP7_75t_R FILLER_170_101 ();
 DECAPx10_ASAP7_75t_R FILLER_170_109 ();
 DECAPx6_ASAP7_75t_R FILLER_170_131 ();
 DECAPx1_ASAP7_75t_R FILLER_170_171 ();
 DECAPx1_ASAP7_75t_R FILLER_170_219 ();
 DECAPx1_ASAP7_75t_R FILLER_170_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_241 ();
 DECAPx2_ASAP7_75t_R FILLER_170_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_261 ();
 DECAPx2_ASAP7_75t_R FILLER_170_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_274 ();
 DECAPx1_ASAP7_75t_R FILLER_170_283 ();
 DECAPx4_ASAP7_75t_R FILLER_170_299 ();
 FILLER_ASAP7_75t_R FILLER_170_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_311 ();
 DECAPx4_ASAP7_75t_R FILLER_170_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_328 ();
 DECAPx6_ASAP7_75t_R FILLER_170_335 ();
 DECAPx2_ASAP7_75t_R FILLER_170_357 ();
 FILLER_ASAP7_75t_R FILLER_170_363 ();
 FILLER_ASAP7_75t_R FILLER_170_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_381 ();
 DECAPx1_ASAP7_75t_R FILLER_170_396 ();
 DECAPx6_ASAP7_75t_R FILLER_170_406 ();
 DECAPx2_ASAP7_75t_R FILLER_170_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_461 ();
 DECAPx2_ASAP7_75t_R FILLER_170_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_479 ();
 DECAPx6_ASAP7_75t_R FILLER_170_489 ();
 DECAPx2_ASAP7_75t_R FILLER_170_503 ();
 DECAPx2_ASAP7_75t_R FILLER_170_515 ();
 DECAPx4_ASAP7_75t_R FILLER_170_529 ();
 FILLER_ASAP7_75t_R FILLER_170_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_541 ();
 DECAPx2_ASAP7_75t_R FILLER_170_557 ();
 FILLER_ASAP7_75t_R FILLER_170_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_565 ();
 DECAPx4_ASAP7_75t_R FILLER_170_574 ();
 FILLER_ASAP7_75t_R FILLER_170_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_586 ();
 DECAPx1_ASAP7_75t_R FILLER_170_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_605 ();
 DECAPx1_ASAP7_75t_R FILLER_170_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_639 ();
 DECAPx1_ASAP7_75t_R FILLER_170_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_659 ();
 DECAPx10_ASAP7_75t_R FILLER_170_705 ();
 DECAPx2_ASAP7_75t_R FILLER_170_727 ();
 FILLER_ASAP7_75t_R FILLER_170_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_735 ();
 DECAPx10_ASAP7_75t_R FILLER_170_742 ();
 DECAPx6_ASAP7_75t_R FILLER_170_764 ();
 FILLER_ASAP7_75t_R FILLER_170_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_780 ();
 DECAPx4_ASAP7_75t_R FILLER_170_795 ();
 DECAPx2_ASAP7_75t_R FILLER_170_815 ();
 DECAPx6_ASAP7_75t_R FILLER_170_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_850 ();
 FILLER_ASAP7_75t_R FILLER_170_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_859 ();
 DECAPx6_ASAP7_75t_R FILLER_170_870 ();
 FILLER_ASAP7_75t_R FILLER_170_884 ();
 FILLER_ASAP7_75t_R FILLER_170_894 ();
 FILLER_ASAP7_75t_R FILLER_170_906 ();
 FILLER_ASAP7_75t_R FILLER_170_914 ();
 DECAPx1_ASAP7_75t_R FILLER_170_922 ();
 DECAPx2_ASAP7_75t_R FILLER_170_929 ();
 FILLER_ASAP7_75t_R FILLER_170_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_953 ();
 DECAPx2_ASAP7_75t_R FILLER_170_960 ();
 FILLER_ASAP7_75t_R FILLER_170_966 ();
 DECAPx4_ASAP7_75t_R FILLER_170_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_991 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1005 ();
 FILLER_ASAP7_75t_R FILLER_170_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1168 ();
 FILLER_ASAP7_75t_R FILLER_170_1194 ();
 FILLER_ASAP7_75t_R FILLER_170_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1204 ();
 FILLER_ASAP7_75t_R FILLER_170_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1224 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1245 ();
 FILLER_ASAP7_75t_R FILLER_170_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1268 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1290 ();
 FILLER_ASAP7_75t_R FILLER_170_1300 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1332 ();
 FILLER_ASAP7_75t_R FILLER_170_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_171_2 ();
 FILLER_ASAP7_75t_R FILLER_171_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_18 ();
 DECAPx2_ASAP7_75t_R FILLER_171_60 ();
 FILLER_ASAP7_75t_R FILLER_171_81 ();
 DECAPx2_ASAP7_75t_R FILLER_171_109 ();
 FILLER_ASAP7_75t_R FILLER_171_115 ();
 DECAPx1_ASAP7_75t_R FILLER_171_125 ();
 DECAPx10_ASAP7_75t_R FILLER_171_132 ();
 DECAPx1_ASAP7_75t_R FILLER_171_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_158 ();
 FILLER_ASAP7_75t_R FILLER_171_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_164 ();
 DECAPx10_ASAP7_75t_R FILLER_171_201 ();
 DECAPx2_ASAP7_75t_R FILLER_171_223 ();
 FILLER_ASAP7_75t_R FILLER_171_229 ();
 DECAPx2_ASAP7_75t_R FILLER_171_247 ();
 DECAPx10_ASAP7_75t_R FILLER_171_261 ();
 DECAPx2_ASAP7_75t_R FILLER_171_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_289 ();
 FILLER_ASAP7_75t_R FILLER_171_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_324 ();
 DECAPx6_ASAP7_75t_R FILLER_171_333 ();
 FILLER_ASAP7_75t_R FILLER_171_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_349 ();
 DECAPx10_ASAP7_75t_R FILLER_171_356 ();
 DECAPx1_ASAP7_75t_R FILLER_171_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_382 ();
 DECAPx2_ASAP7_75t_R FILLER_171_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_395 ();
 DECAPx6_ASAP7_75t_R FILLER_171_402 ();
 DECAPx1_ASAP7_75t_R FILLER_171_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_446 ();
 DECAPx4_ASAP7_75t_R FILLER_171_479 ();
 FILLER_ASAP7_75t_R FILLER_171_489 ();
 DECAPx1_ASAP7_75t_R FILLER_171_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_505 ();
 DECAPx2_ASAP7_75t_R FILLER_171_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_533 ();
 DECAPx1_ASAP7_75t_R FILLER_171_556 ();
 FILLER_ASAP7_75t_R FILLER_171_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_596 ();
 FILLER_ASAP7_75t_R FILLER_171_631 ();
 FILLER_ASAP7_75t_R FILLER_171_647 ();
 DECAPx4_ASAP7_75t_R FILLER_171_673 ();
 FILLER_ASAP7_75t_R FILLER_171_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_685 ();
 DECAPx6_ASAP7_75t_R FILLER_171_696 ();
 DECAPx1_ASAP7_75t_R FILLER_171_710 ();
 DECAPx2_ASAP7_75t_R FILLER_171_728 ();
 FILLER_ASAP7_75t_R FILLER_171_734 ();
 DECAPx2_ASAP7_75t_R FILLER_171_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_754 ();
 DECAPx1_ASAP7_75t_R FILLER_171_775 ();
 DECAPx10_ASAP7_75t_R FILLER_171_786 ();
 DECAPx10_ASAP7_75t_R FILLER_171_808 ();
 DECAPx10_ASAP7_75t_R FILLER_171_830 ();
 DECAPx1_ASAP7_75t_R FILLER_171_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_856 ();
 FILLER_ASAP7_75t_R FILLER_171_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_887 ();
 FILLER_ASAP7_75t_R FILLER_171_944 ();
 DECAPx4_ASAP7_75t_R FILLER_171_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_968 ();
 DECAPx6_ASAP7_75t_R FILLER_171_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_990 ();
 FILLER_ASAP7_75t_R FILLER_171_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_999 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1079 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1248 ();
 FILLER_ASAP7_75t_R FILLER_171_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1267 ();
 FILLER_ASAP7_75t_R FILLER_171_1277 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1293 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1319 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1325 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1378 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_172_2 ();
 DECAPx1_ASAP7_75t_R FILLER_172_24 ();
 FILLER_ASAP7_75t_R FILLER_172_31 ();
 FILLER_ASAP7_75t_R FILLER_172_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_76 ();
 FILLER_ASAP7_75t_R FILLER_172_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_85 ();
 DECAPx10_ASAP7_75t_R FILLER_172_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_114 ();
 FILLER_ASAP7_75t_R FILLER_172_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_143 ();
 DECAPx4_ASAP7_75t_R FILLER_172_153 ();
 DECAPx1_ASAP7_75t_R FILLER_172_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_210 ();
 DECAPx6_ASAP7_75t_R FILLER_172_217 ();
 FILLER_ASAP7_75t_R FILLER_172_241 ();
 FILLER_ASAP7_75t_R FILLER_172_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_251 ();
 DECAPx4_ASAP7_75t_R FILLER_172_284 ();
 FILLER_ASAP7_75t_R FILLER_172_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_303 ();
 DECAPx4_ASAP7_75t_R FILLER_172_307 ();
 FILLER_ASAP7_75t_R FILLER_172_317 ();
 DECAPx1_ASAP7_75t_R FILLER_172_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_346 ();
 FILLER_ASAP7_75t_R FILLER_172_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_375 ();
 DECAPx10_ASAP7_75t_R FILLER_172_382 ();
 DECAPx4_ASAP7_75t_R FILLER_172_404 ();
 FILLER_ASAP7_75t_R FILLER_172_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_426 ();
 DECAPx1_ASAP7_75t_R FILLER_172_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_461 ();
 FILLER_ASAP7_75t_R FILLER_172_467 ();
 DECAPx1_ASAP7_75t_R FILLER_172_477 ();
 DECAPx1_ASAP7_75t_R FILLER_172_487 ();
 DECAPx4_ASAP7_75t_R FILLER_172_530 ();
 FILLER_ASAP7_75t_R FILLER_172_540 ();
 DECAPx2_ASAP7_75t_R FILLER_172_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_563 ();
 DECAPx1_ASAP7_75t_R FILLER_172_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_582 ();
 DECAPx6_ASAP7_75t_R FILLER_172_604 ();
 DECAPx1_ASAP7_75t_R FILLER_172_618 ();
 DECAPx10_ASAP7_75t_R FILLER_172_632 ();
 DECAPx4_ASAP7_75t_R FILLER_172_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_664 ();
 DECAPx4_ASAP7_75t_R FILLER_172_677 ();
 FILLER_ASAP7_75t_R FILLER_172_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_711 ();
 DECAPx2_ASAP7_75t_R FILLER_172_718 ();
 FILLER_ASAP7_75t_R FILLER_172_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_726 ();
 DECAPx1_ASAP7_75t_R FILLER_172_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_741 ();
 DECAPx1_ASAP7_75t_R FILLER_172_770 ();
 DECAPx1_ASAP7_75t_R FILLER_172_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_784 ();
 DECAPx4_ASAP7_75t_R FILLER_172_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_798 ();
 DECAPx6_ASAP7_75t_R FILLER_172_805 ();
 DECAPx1_ASAP7_75t_R FILLER_172_819 ();
 DECAPx10_ASAP7_75t_R FILLER_172_829 ();
 DECAPx2_ASAP7_75t_R FILLER_172_857 ();
 FILLER_ASAP7_75t_R FILLER_172_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_865 ();
 DECAPx4_ASAP7_75t_R FILLER_172_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_886 ();
 DECAPx10_ASAP7_75t_R FILLER_172_903 ();
 DECAPx2_ASAP7_75t_R FILLER_172_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_931 ();
 DECAPx2_ASAP7_75t_R FILLER_172_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_946 ();
 DECAPx2_ASAP7_75t_R FILLER_172_960 ();
 DECAPx4_ASAP7_75t_R FILLER_172_976 ();
 FILLER_ASAP7_75t_R FILLER_172_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1001 ();
 FILLER_ASAP7_75t_R FILLER_172_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1091 ();
 FILLER_ASAP7_75t_R FILLER_172_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1171 ();
 FILLER_ASAP7_75t_R FILLER_172_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1195 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1208 ();
 FILLER_ASAP7_75t_R FILLER_172_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1224 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1307 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1315 ();
 FILLER_ASAP7_75t_R FILLER_172_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1333 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1368 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1385 ();
 FILLER_ASAP7_75t_R FILLER_172_1398 ();
 DECAPx1_ASAP7_75t_R FILLER_173_2 ();
 FILLER_ASAP7_75t_R FILLER_173_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_40 ();
 FILLER_ASAP7_75t_R FILLER_173_44 ();
 DECAPx2_ASAP7_75t_R FILLER_173_49 ();
 DECAPx2_ASAP7_75t_R FILLER_173_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_102 ();
 DECAPx2_ASAP7_75t_R FILLER_173_106 ();
 DECAPx4_ASAP7_75t_R FILLER_173_128 ();
 FILLER_ASAP7_75t_R FILLER_173_138 ();
 FILLER_ASAP7_75t_R FILLER_173_166 ();
 DECAPx4_ASAP7_75t_R FILLER_173_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_242 ();
 DECAPx6_ASAP7_75t_R FILLER_173_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_265 ();
 FILLER_ASAP7_75t_R FILLER_173_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_271 ();
 DECAPx2_ASAP7_75t_R FILLER_173_282 ();
 FILLER_ASAP7_75t_R FILLER_173_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_290 ();
 DECAPx6_ASAP7_75t_R FILLER_173_305 ();
 DECAPx2_ASAP7_75t_R FILLER_173_319 ();
 DECAPx6_ASAP7_75t_R FILLER_173_331 ();
 DECAPx1_ASAP7_75t_R FILLER_173_345 ();
 DECAPx1_ASAP7_75t_R FILLER_173_362 ();
 DECAPx4_ASAP7_75t_R FILLER_173_392 ();
 FILLER_ASAP7_75t_R FILLER_173_402 ();
 DECAPx1_ASAP7_75t_R FILLER_173_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_442 ();
 DECAPx2_ASAP7_75t_R FILLER_173_461 ();
 DECAPx10_ASAP7_75t_R FILLER_173_503 ();
 DECAPx6_ASAP7_75t_R FILLER_173_525 ();
 FILLER_ASAP7_75t_R FILLER_173_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_541 ();
 DECAPx4_ASAP7_75t_R FILLER_173_552 ();
 DECAPx4_ASAP7_75t_R FILLER_173_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_586 ();
 DECAPx10_ASAP7_75t_R FILLER_173_593 ();
 DECAPx1_ASAP7_75t_R FILLER_173_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_619 ();
 DECAPx1_ASAP7_75t_R FILLER_173_626 ();
 DECAPx6_ASAP7_75t_R FILLER_173_636 ();
 DECAPx1_ASAP7_75t_R FILLER_173_650 ();
 DECAPx1_ASAP7_75t_R FILLER_173_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_680 ();
 DECAPx1_ASAP7_75t_R FILLER_173_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_705 ();
 DECAPx2_ASAP7_75t_R FILLER_173_713 ();
 DECAPx10_ASAP7_75t_R FILLER_173_733 ();
 DECAPx1_ASAP7_75t_R FILLER_173_755 ();
 DECAPx1_ASAP7_75t_R FILLER_173_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_769 ();
 DECAPx2_ASAP7_75t_R FILLER_173_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_784 ();
 FILLER_ASAP7_75t_R FILLER_173_801 ();
 DECAPx6_ASAP7_75t_R FILLER_173_822 ();
 DECAPx2_ASAP7_75t_R FILLER_173_836 ();
 DECAPx4_ASAP7_75t_R FILLER_173_854 ();
 FILLER_ASAP7_75t_R FILLER_173_864 ();
 DECAPx10_ASAP7_75t_R FILLER_173_874 ();
 DECAPx4_ASAP7_75t_R FILLER_173_896 ();
 FILLER_ASAP7_75t_R FILLER_173_906 ();
 DECAPx2_ASAP7_75t_R FILLER_173_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_923 ();
 DECAPx2_ASAP7_75t_R FILLER_173_926 ();
 FILLER_ASAP7_75t_R FILLER_173_932 ();
 DECAPx2_ASAP7_75t_R FILLER_173_942 ();
 DECAPx1_ASAP7_75t_R FILLER_173_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_964 ();
 DECAPx1_ASAP7_75t_R FILLER_173_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_985 ();
 DECAPx1_ASAP7_75t_R FILLER_173_996 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_173_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1031 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1142 ();
 FILLER_ASAP7_75t_R FILLER_173_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1207 ();
 FILLER_ASAP7_75t_R FILLER_173_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1274 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1289 ();
 FILLER_ASAP7_75t_R FILLER_173_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1308 ();
 FILLER_ASAP7_75t_R FILLER_173_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_173_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1354 ();
 FILLER_ASAP7_75t_R FILLER_173_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1362 ();
 DECAPx6_ASAP7_75t_R FILLER_174_2 ();
 DECAPx1_ASAP7_75t_R FILLER_174_16 ();
 FILLER_ASAP7_75t_R FILLER_174_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_25 ();
 DECAPx10_ASAP7_75t_R FILLER_174_32 ();
 DECAPx10_ASAP7_75t_R FILLER_174_60 ();
 FILLER_ASAP7_75t_R FILLER_174_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_88 ();
 DECAPx1_ASAP7_75t_R FILLER_174_123 ();
 DECAPx2_ASAP7_75t_R FILLER_174_133 ();
 FILLER_ASAP7_75t_R FILLER_174_139 ();
 DECAPx2_ASAP7_75t_R FILLER_174_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_153 ();
 DECAPx1_ASAP7_75t_R FILLER_174_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_176 ();
 DECAPx6_ASAP7_75t_R FILLER_174_190 ();
 DECAPx1_ASAP7_75t_R FILLER_174_204 ();
 DECAPx10_ASAP7_75t_R FILLER_174_217 ();
 DECAPx2_ASAP7_75t_R FILLER_174_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_245 ();
 DECAPx10_ASAP7_75t_R FILLER_174_252 ();
 DECAPx4_ASAP7_75t_R FILLER_174_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_309 ();
 DECAPx1_ASAP7_75t_R FILLER_174_313 ();
 DECAPx10_ASAP7_75t_R FILLER_174_323 ();
 DECAPx2_ASAP7_75t_R FILLER_174_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_361 ();
 DECAPx1_ASAP7_75t_R FILLER_174_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_369 ();
 DECAPx1_ASAP7_75t_R FILLER_174_422 ();
 FILLER_ASAP7_75t_R FILLER_174_437 ();
 DECAPx2_ASAP7_75t_R FILLER_174_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_461 ();
 DECAPx2_ASAP7_75t_R FILLER_174_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_470 ();
 DECAPx6_ASAP7_75t_R FILLER_174_477 ();
 DECAPx1_ASAP7_75t_R FILLER_174_491 ();
 DECAPx1_ASAP7_75t_R FILLER_174_521 ();
 DECAPx1_ASAP7_75t_R FILLER_174_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_535 ();
 DECAPx6_ASAP7_75t_R FILLER_174_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_583 ();
 FILLER_ASAP7_75t_R FILLER_174_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_600 ();
 DECAPx2_ASAP7_75t_R FILLER_174_610 ();
 FILLER_ASAP7_75t_R FILLER_174_616 ();
 FILLER_ASAP7_75t_R FILLER_174_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_667 ();
 DECAPx1_ASAP7_75t_R FILLER_174_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_678 ();
 DECAPx1_ASAP7_75t_R FILLER_174_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_703 ();
 DECAPx6_ASAP7_75t_R FILLER_174_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_732 ();
 DECAPx2_ASAP7_75t_R FILLER_174_745 ();
 FILLER_ASAP7_75t_R FILLER_174_751 ();
 DECAPx6_ASAP7_75t_R FILLER_174_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_799 ();
 DECAPx10_ASAP7_75t_R FILLER_174_806 ();
 DECAPx10_ASAP7_75t_R FILLER_174_834 ();
 DECAPx2_ASAP7_75t_R FILLER_174_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_862 ();
 DECAPx4_ASAP7_75t_R FILLER_174_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_881 ();
 DECAPx6_ASAP7_75t_R FILLER_174_890 ();
 DECAPx1_ASAP7_75t_R FILLER_174_904 ();
 DECAPx1_ASAP7_75t_R FILLER_174_927 ();
 DECAPx6_ASAP7_75t_R FILLER_174_939 ();
 DECAPx1_ASAP7_75t_R FILLER_174_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_957 ();
 DECAPx2_ASAP7_75t_R FILLER_174_981 ();
 DECAPx10_ASAP7_75t_R FILLER_174_994 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1096 ();
 FILLER_ASAP7_75t_R FILLER_174_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1136 ();
 FILLER_ASAP7_75t_R FILLER_174_1142 ();
 FILLER_ASAP7_75t_R FILLER_174_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1161 ();
 FILLER_ASAP7_75t_R FILLER_174_1167 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1175 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1185 ();
 FILLER_ASAP7_75t_R FILLER_174_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1256 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1263 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1385 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1395 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_175_2 ();
 DECAPx10_ASAP7_75t_R FILLER_175_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_46 ();
 DECAPx6_ASAP7_75t_R FILLER_175_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_93 ();
 DECAPx6_ASAP7_75t_R FILLER_175_97 ();
 DECAPx1_ASAP7_75t_R FILLER_175_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_115 ();
 DECAPx10_ASAP7_75t_R FILLER_175_148 ();
 DECAPx10_ASAP7_75t_R FILLER_175_170 ();
 DECAPx2_ASAP7_75t_R FILLER_175_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_204 ();
 DECAPx2_ASAP7_75t_R FILLER_175_219 ();
 FILLER_ASAP7_75t_R FILLER_175_241 ();
 DECAPx2_ASAP7_75t_R FILLER_175_249 ();
 FILLER_ASAP7_75t_R FILLER_175_261 ();
 DECAPx1_ASAP7_75t_R FILLER_175_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_312 ();
 DECAPx1_ASAP7_75t_R FILLER_175_321 ();
 DECAPx6_ASAP7_75t_R FILLER_175_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_356 ();
 DECAPx10_ASAP7_75t_R FILLER_175_363 ();
 DECAPx1_ASAP7_75t_R FILLER_175_385 ();
 DECAPx6_ASAP7_75t_R FILLER_175_403 ();
 DECAPx2_ASAP7_75t_R FILLER_175_417 ();
 FILLER_ASAP7_75t_R FILLER_175_446 ();
 DECAPx1_ASAP7_75t_R FILLER_175_466 ();
 DECAPx1_ASAP7_75t_R FILLER_175_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_488 ();
 DECAPx1_ASAP7_75t_R FILLER_175_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_507 ();
 DECAPx1_ASAP7_75t_R FILLER_175_548 ();
 DECAPx6_ASAP7_75t_R FILLER_175_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_572 ();
 DECAPx4_ASAP7_75t_R FILLER_175_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_597 ();
 DECAPx1_ASAP7_75t_R FILLER_175_614 ();
 DECAPx10_ASAP7_75t_R FILLER_175_644 ();
 DECAPx4_ASAP7_75t_R FILLER_175_666 ();
 DECAPx6_ASAP7_75t_R FILLER_175_689 ();
 DECAPx2_ASAP7_75t_R FILLER_175_713 ();
 DECAPx2_ASAP7_75t_R FILLER_175_725 ();
 FILLER_ASAP7_75t_R FILLER_175_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_733 ();
 DECAPx10_ASAP7_75t_R FILLER_175_746 ();
 DECAPx6_ASAP7_75t_R FILLER_175_768 ();
 DECAPx10_ASAP7_75t_R FILLER_175_792 ();
 DECAPx2_ASAP7_75t_R FILLER_175_814 ();
 FILLER_ASAP7_75t_R FILLER_175_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_822 ();
 DECAPx1_ASAP7_75t_R FILLER_175_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_850 ();
 FILLER_ASAP7_75t_R FILLER_175_867 ();
 FILLER_ASAP7_75t_R FILLER_175_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_881 ();
 FILLER_ASAP7_75t_R FILLER_175_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_892 ();
 DECAPx2_ASAP7_75t_R FILLER_175_916 ();
 FILLER_ASAP7_75t_R FILLER_175_922 ();
 DECAPx4_ASAP7_75t_R FILLER_175_942 ();
 DECAPx2_ASAP7_75t_R FILLER_175_962 ();
 DECAPx1_ASAP7_75t_R FILLER_175_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_980 ();
 DECAPx10_ASAP7_75t_R FILLER_175_987 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1020 ();
 FILLER_ASAP7_75t_R FILLER_175_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1044 ();
 FILLER_ASAP7_75t_R FILLER_175_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1128 ();
 FILLER_ASAP7_75t_R FILLER_175_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_175_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1179 ();
 DECAPx4_ASAP7_75t_R FILLER_175_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1211 ();
 FILLER_ASAP7_75t_R FILLER_175_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1248 ();
 FILLER_ASAP7_75t_R FILLER_175_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1291 ();
 FILLER_ASAP7_75t_R FILLER_175_1295 ();
 DECAPx4_ASAP7_75t_R FILLER_175_1313 ();
 FILLER_ASAP7_75t_R FILLER_175_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1325 ();
 FILLER_ASAP7_75t_R FILLER_175_1360 ();
 FILLER_ASAP7_75t_R FILLER_175_1365 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1374 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1378 ();
 DECAPx6_ASAP7_75t_R FILLER_176_2 ();
 DECAPx2_ASAP7_75t_R FILLER_176_16 ();
 FILLER_ASAP7_75t_R FILLER_176_25 ();
 DECAPx1_ASAP7_75t_R FILLER_176_33 ();
 FILLER_ASAP7_75t_R FILLER_176_59 ();
 DECAPx6_ASAP7_75t_R FILLER_176_64 ();
 FILLER_ASAP7_75t_R FILLER_176_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_80 ();
 DECAPx1_ASAP7_75t_R FILLER_176_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_97 ();
 FILLER_ASAP7_75t_R FILLER_176_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_126 ();
 FILLER_ASAP7_75t_R FILLER_176_153 ();
 DECAPx2_ASAP7_75t_R FILLER_176_167 ();
 FILLER_ASAP7_75t_R FILLER_176_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_175 ();
 DECAPx1_ASAP7_75t_R FILLER_176_210 ();
 FILLER_ASAP7_75t_R FILLER_176_221 ();
 DECAPx2_ASAP7_75t_R FILLER_176_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_244 ();
 DECAPx1_ASAP7_75t_R FILLER_176_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_257 ();
 DECAPx10_ASAP7_75t_R FILLER_176_274 ();
 DECAPx1_ASAP7_75t_R FILLER_176_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_300 ();
 DECAPx4_ASAP7_75t_R FILLER_176_304 ();
 FILLER_ASAP7_75t_R FILLER_176_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_316 ();
 DECAPx10_ASAP7_75t_R FILLER_176_323 ();
 DECAPx4_ASAP7_75t_R FILLER_176_345 ();
 FILLER_ASAP7_75t_R FILLER_176_355 ();
 DECAPx10_ASAP7_75t_R FILLER_176_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_405 ();
 DECAPx4_ASAP7_75t_R FILLER_176_412 ();
 FILLER_ASAP7_75t_R FILLER_176_422 ();
 DECAPx10_ASAP7_75t_R FILLER_176_430 ();
 DECAPx1_ASAP7_75t_R FILLER_176_452 ();
 DECAPx1_ASAP7_75t_R FILLER_176_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_468 ();
 DECAPx6_ASAP7_75t_R FILLER_176_483 ();
 FILLER_ASAP7_75t_R FILLER_176_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_499 ();
 FILLER_ASAP7_75t_R FILLER_176_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_508 ();
 DECAPx2_ASAP7_75t_R FILLER_176_512 ();
 FILLER_ASAP7_75t_R FILLER_176_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_528 ();
 DECAPx6_ASAP7_75t_R FILLER_176_532 ();
 FILLER_ASAP7_75t_R FILLER_176_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_568 ();
 DECAPx1_ASAP7_75t_R FILLER_176_578 ();
 FILLER_ASAP7_75t_R FILLER_176_596 ();
 FILLER_ASAP7_75t_R FILLER_176_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_618 ();
 DECAPx2_ASAP7_75t_R FILLER_176_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_631 ();
 DECAPx2_ASAP7_75t_R FILLER_176_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_641 ();
 DECAPx4_ASAP7_75t_R FILLER_176_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_658 ();
 DECAPx1_ASAP7_75t_R FILLER_176_673 ();
 DECAPx2_ASAP7_75t_R FILLER_176_685 ();
 FILLER_ASAP7_75t_R FILLER_176_691 ();
 FILLER_ASAP7_75t_R FILLER_176_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_702 ();
 FILLER_ASAP7_75t_R FILLER_176_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_711 ();
 DECAPx6_ASAP7_75t_R FILLER_176_720 ();
 FILLER_ASAP7_75t_R FILLER_176_774 ();
 DECAPx10_ASAP7_75t_R FILLER_176_792 ();
 DECAPx10_ASAP7_75t_R FILLER_176_814 ();
 DECAPx1_ASAP7_75t_R FILLER_176_836 ();
 DECAPx6_ASAP7_75t_R FILLER_176_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_860 ();
 DECAPx1_ASAP7_75t_R FILLER_176_864 ();
 FILLER_ASAP7_75t_R FILLER_176_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_886 ();
 DECAPx2_ASAP7_75t_R FILLER_176_909 ();
 FILLER_ASAP7_75t_R FILLER_176_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_917 ();
 DECAPx4_ASAP7_75t_R FILLER_176_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_948 ();
 DECAPx10_ASAP7_75t_R FILLER_176_963 ();
 FILLER_ASAP7_75t_R FILLER_176_985 ();
 FILLER_ASAP7_75t_R FILLER_176_997 ();
 FILLER_ASAP7_75t_R FILLER_176_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1086 ();
 FILLER_ASAP7_75t_R FILLER_176_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1109 ();
 FILLER_ASAP7_75t_R FILLER_176_1115 ();
 FILLER_ASAP7_75t_R FILLER_176_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1224 ();
 FILLER_ASAP7_75t_R FILLER_176_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1318 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1327 ();
 FILLER_ASAP7_75t_R FILLER_176_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1357 ();
 FILLER_ASAP7_75t_R FILLER_176_1394 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1399 ();
 DECAPx2_ASAP7_75t_R FILLER_177_2 ();
 DECAPx6_ASAP7_75t_R FILLER_177_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_58 ();
 DECAPx1_ASAP7_75t_R FILLER_177_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_66 ();
 FILLER_ASAP7_75t_R FILLER_177_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_120 ();
 DECAPx4_ASAP7_75t_R FILLER_177_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_140 ();
 DECAPx1_ASAP7_75t_R FILLER_177_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_148 ();
 DECAPx2_ASAP7_75t_R FILLER_177_162 ();
 DECAPx2_ASAP7_75t_R FILLER_177_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_200 ();
 FILLER_ASAP7_75t_R FILLER_177_207 ();
 DECAPx6_ASAP7_75t_R FILLER_177_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_235 ();
 DECAPx2_ASAP7_75t_R FILLER_177_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_268 ();
 DECAPx2_ASAP7_75t_R FILLER_177_283 ();
 FILLER_ASAP7_75t_R FILLER_177_289 ();
 DECAPx10_ASAP7_75t_R FILLER_177_301 ();
 DECAPx2_ASAP7_75t_R FILLER_177_323 ();
 FILLER_ASAP7_75t_R FILLER_177_329 ();
 DECAPx6_ASAP7_75t_R FILLER_177_337 ();
 DECAPx2_ASAP7_75t_R FILLER_177_351 ();
 DECAPx2_ASAP7_75t_R FILLER_177_363 ();
 FILLER_ASAP7_75t_R FILLER_177_369 ();
 FILLER_ASAP7_75t_R FILLER_177_374 ();
 DECAPx1_ASAP7_75t_R FILLER_177_393 ();
 FILLER_ASAP7_75t_R FILLER_177_435 ();
 DECAPx6_ASAP7_75t_R FILLER_177_443 ();
 FILLER_ASAP7_75t_R FILLER_177_457 ();
 DECAPx1_ASAP7_75t_R FILLER_177_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_483 ();
 DECAPx6_ASAP7_75t_R FILLER_177_490 ();
 DECAPx1_ASAP7_75t_R FILLER_177_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_508 ();
 DECAPx4_ASAP7_75t_R FILLER_177_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_527 ();
 DECAPx1_ASAP7_75t_R FILLER_177_534 ();
 FILLER_ASAP7_75t_R FILLER_177_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_546 ();
 DECAPx6_ASAP7_75t_R FILLER_177_554 ();
 FILLER_ASAP7_75t_R FILLER_177_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_570 ();
 FILLER_ASAP7_75t_R FILLER_177_595 ();
 DECAPx6_ASAP7_75t_R FILLER_177_609 ();
 DECAPx2_ASAP7_75t_R FILLER_177_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_637 ();
 DECAPx2_ASAP7_75t_R FILLER_177_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_702 ();
 DECAPx2_ASAP7_75t_R FILLER_177_726 ();
 FILLER_ASAP7_75t_R FILLER_177_732 ();
 DECAPx10_ASAP7_75t_R FILLER_177_751 ();
 DECAPx2_ASAP7_75t_R FILLER_177_773 ();
 FILLER_ASAP7_75t_R FILLER_177_779 ();
 DECAPx4_ASAP7_75t_R FILLER_177_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_797 ();
 DECAPx2_ASAP7_75t_R FILLER_177_819 ();
 FILLER_ASAP7_75t_R FILLER_177_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_827 ();
 FILLER_ASAP7_75t_R FILLER_177_836 ();
 DECAPx10_ASAP7_75t_R FILLER_177_844 ();
 DECAPx10_ASAP7_75t_R FILLER_177_866 ();
 DECAPx2_ASAP7_75t_R FILLER_177_888 ();
 FILLER_ASAP7_75t_R FILLER_177_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_896 ();
 DECAPx6_ASAP7_75t_R FILLER_177_907 ();
 FILLER_ASAP7_75t_R FILLER_177_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_923 ();
 DECAPx1_ASAP7_75t_R FILLER_177_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_930 ();
 DECAPx4_ASAP7_75t_R FILLER_177_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_966 ();
 FILLER_ASAP7_75t_R FILLER_177_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_977 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1027 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1042 ();
 FILLER_ASAP7_75t_R FILLER_177_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1066 ();
 FILLER_ASAP7_75t_R FILLER_177_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1082 ();
 FILLER_ASAP7_75t_R FILLER_177_1089 ();
 FILLER_ASAP7_75t_R FILLER_177_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1155 ();
 FILLER_ASAP7_75t_R FILLER_177_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1198 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1208 ();
 FILLER_ASAP7_75t_R FILLER_177_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1251 ();
 FILLER_ASAP7_75t_R FILLER_177_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1273 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1295 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1309 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1327 ();
 FILLER_ASAP7_75t_R FILLER_177_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1339 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1399 ();
 FILLER_ASAP7_75t_R FILLER_178_2 ();
 DECAPx2_ASAP7_75t_R FILLER_178_36 ();
 FILLER_ASAP7_75t_R FILLER_178_42 ();
 DECAPx2_ASAP7_75t_R FILLER_178_83 ();
 FILLER_ASAP7_75t_R FILLER_178_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_118 ();
 DECAPx1_ASAP7_75t_R FILLER_178_122 ();
 DECAPx1_ASAP7_75t_R FILLER_178_134 ();
 DECAPx1_ASAP7_75t_R FILLER_178_141 ();
 DECAPx4_ASAP7_75t_R FILLER_178_171 ();
 DECAPx1_ASAP7_75t_R FILLER_178_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_221 ();
 DECAPx2_ASAP7_75t_R FILLER_178_236 ();
 FILLER_ASAP7_75t_R FILLER_178_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_244 ();
 DECAPx4_ASAP7_75t_R FILLER_178_267 ();
 FILLER_ASAP7_75t_R FILLER_178_277 ();
 DECAPx4_ASAP7_75t_R FILLER_178_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_299 ();
 DECAPx10_ASAP7_75t_R FILLER_178_317 ();
 DECAPx10_ASAP7_75t_R FILLER_178_339 ();
 DECAPx10_ASAP7_75t_R FILLER_178_361 ();
 FILLER_ASAP7_75t_R FILLER_178_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_385 ();
 FILLER_ASAP7_75t_R FILLER_178_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_422 ();
 DECAPx1_ASAP7_75t_R FILLER_178_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_435 ();
 DECAPx4_ASAP7_75t_R FILLER_178_450 ();
 FILLER_ASAP7_75t_R FILLER_178_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_479 ();
 DECAPx2_ASAP7_75t_R FILLER_178_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_512 ();
 FILLER_ASAP7_75t_R FILLER_178_538 ();
 DECAPx4_ASAP7_75t_R FILLER_178_556 ();
 FILLER_ASAP7_75t_R FILLER_178_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_568 ();
 FILLER_ASAP7_75t_R FILLER_178_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_579 ();
 DECAPx2_ASAP7_75t_R FILLER_178_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_598 ();
 FILLER_ASAP7_75t_R FILLER_178_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_618 ();
 FILLER_ASAP7_75t_R FILLER_178_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_660 ();
 DECAPx1_ASAP7_75t_R FILLER_178_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_690 ();
 DECAPx2_ASAP7_75t_R FILLER_178_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_711 ();
 DECAPx10_ASAP7_75t_R FILLER_178_719 ();
 DECAPx4_ASAP7_75t_R FILLER_178_741 ();
 FILLER_ASAP7_75t_R FILLER_178_761 ();
 DECAPx4_ASAP7_75t_R FILLER_178_771 ();
 DECAPx1_ASAP7_75t_R FILLER_178_794 ();
 FILLER_ASAP7_75t_R FILLER_178_814 ();
 FILLER_ASAP7_75t_R FILLER_178_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_847 ();
 DECAPx2_ASAP7_75t_R FILLER_178_858 ();
 FILLER_ASAP7_75t_R FILLER_178_864 ();
 DECAPx10_ASAP7_75t_R FILLER_178_872 ();
 DECAPx1_ASAP7_75t_R FILLER_178_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_898 ();
 DECAPx4_ASAP7_75t_R FILLER_178_915 ();
 DECAPx4_ASAP7_75t_R FILLER_178_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_954 ();
 FILLER_ASAP7_75t_R FILLER_178_963 ();
 FILLER_ASAP7_75t_R FILLER_178_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1129 ();
 FILLER_ASAP7_75t_R FILLER_178_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1149 ();
 FILLER_ASAP7_75t_R FILLER_178_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1225 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1247 ();
 FILLER_ASAP7_75t_R FILLER_178_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1286 ();
 FILLER_ASAP7_75t_R FILLER_178_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1331 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1364 ();
 FILLER_ASAP7_75t_R FILLER_178_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1372 ();
 FILLER_ASAP7_75t_R FILLER_178_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1388 ();
 FILLER_ASAP7_75t_R FILLER_178_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1396 ();
 DECAPx6_ASAP7_75t_R FILLER_179_2 ();
 FILLER_ASAP7_75t_R FILLER_179_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_22 ();
 FILLER_ASAP7_75t_R FILLER_179_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_31 ();
 DECAPx1_ASAP7_75t_R FILLER_179_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_62 ();
 DECAPx10_ASAP7_75t_R FILLER_179_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_100 ();
 DECAPx1_ASAP7_75t_R FILLER_179_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_149 ();
 DECAPx2_ASAP7_75t_R FILLER_179_153 ();
 DECAPx6_ASAP7_75t_R FILLER_179_162 ();
 FILLER_ASAP7_75t_R FILLER_179_176 ();
 DECAPx10_ASAP7_75t_R FILLER_179_184 ();
 DECAPx6_ASAP7_75t_R FILLER_179_206 ();
 DECAPx1_ASAP7_75t_R FILLER_179_220 ();
 DECAPx2_ASAP7_75t_R FILLER_179_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_255 ();
 FILLER_ASAP7_75t_R FILLER_179_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_273 ();
 DECAPx2_ASAP7_75t_R FILLER_179_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_287 ();
 FILLER_ASAP7_75t_R FILLER_179_294 ();
 DECAPx6_ASAP7_75t_R FILLER_179_299 ();
 DECAPx2_ASAP7_75t_R FILLER_179_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_319 ();
 DECAPx10_ASAP7_75t_R FILLER_179_326 ();
 DECAPx2_ASAP7_75t_R FILLER_179_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_354 ();
 DECAPx6_ASAP7_75t_R FILLER_179_361 ();
 FILLER_ASAP7_75t_R FILLER_179_375 ();
 DECAPx2_ASAP7_75t_R FILLER_179_383 ();
 FILLER_ASAP7_75t_R FILLER_179_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_403 ();
 DECAPx6_ASAP7_75t_R FILLER_179_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_421 ();
 DECAPx10_ASAP7_75t_R FILLER_179_464 ();
 DECAPx4_ASAP7_75t_R FILLER_179_502 ();
 DECAPx10_ASAP7_75t_R FILLER_179_526 ();
 DECAPx1_ASAP7_75t_R FILLER_179_548 ();
 DECAPx1_ASAP7_75t_R FILLER_179_560 ();
 DECAPx2_ASAP7_75t_R FILLER_179_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_596 ();
 DECAPx2_ASAP7_75t_R FILLER_179_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_609 ();
 DECAPx2_ASAP7_75t_R FILLER_179_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_641 ();
 DECAPx2_ASAP7_75t_R FILLER_179_650 ();
 DECAPx10_ASAP7_75t_R FILLER_179_664 ();
 DECAPx2_ASAP7_75t_R FILLER_179_686 ();
 FILLER_ASAP7_75t_R FILLER_179_692 ();
 DECAPx6_ASAP7_75t_R FILLER_179_702 ();
 FILLER_ASAP7_75t_R FILLER_179_716 ();
 DECAPx4_ASAP7_75t_R FILLER_179_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_734 ();
 DECAPx1_ASAP7_75t_R FILLER_179_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_765 ();
 DECAPx6_ASAP7_75t_R FILLER_179_782 ();
 FILLER_ASAP7_75t_R FILLER_179_802 ();
 DECAPx2_ASAP7_75t_R FILLER_179_819 ();
 FILLER_ASAP7_75t_R FILLER_179_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_848 ();
 FILLER_ASAP7_75t_R FILLER_179_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_865 ();
 DECAPx1_ASAP7_75t_R FILLER_179_882 ();
 DECAPx4_ASAP7_75t_R FILLER_179_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_906 ();
 DECAPx1_ASAP7_75t_R FILLER_179_920 ();
 DECAPx2_ASAP7_75t_R FILLER_179_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_932 ();
 DECAPx4_ASAP7_75t_R FILLER_179_954 ();
 FILLER_ASAP7_75t_R FILLER_179_964 ();
 DECAPx10_ASAP7_75t_R FILLER_179_974 ();
 DECAPx1_ASAP7_75t_R FILLER_179_996 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1107 ();
 FILLER_ASAP7_75t_R FILLER_179_1113 ();
 FILLER_ASAP7_75t_R FILLER_179_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1182 ();
 FILLER_ASAP7_75t_R FILLER_179_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1190 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1199 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1209 ();
 FILLER_ASAP7_75t_R FILLER_179_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1259 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_180_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_28 ();
 FILLER_ASAP7_75t_R FILLER_180_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_37 ();
 DECAPx1_ASAP7_75t_R FILLER_180_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_45 ();
 FILLER_ASAP7_75t_R FILLER_180_49 ();
 DECAPx2_ASAP7_75t_R FILLER_180_58 ();
 DECAPx2_ASAP7_75t_R FILLER_180_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_73 ();
 DECAPx10_ASAP7_75t_R FILLER_180_80 ();
 DECAPx10_ASAP7_75t_R FILLER_180_102 ();
 DECAPx2_ASAP7_75t_R FILLER_180_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_130 ();
 DECAPx2_ASAP7_75t_R FILLER_180_137 ();
 FILLER_ASAP7_75t_R FILLER_180_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_145 ();
 DECAPx6_ASAP7_75t_R FILLER_180_190 ();
 DECAPx10_ASAP7_75t_R FILLER_180_218 ();
 DECAPx10_ASAP7_75t_R FILLER_180_240 ();
 DECAPx4_ASAP7_75t_R FILLER_180_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_272 ();
 FILLER_ASAP7_75t_R FILLER_180_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_307 ();
 DECAPx4_ASAP7_75t_R FILLER_180_314 ();
 FILLER_ASAP7_75t_R FILLER_180_324 ();
 DECAPx2_ASAP7_75t_R FILLER_180_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_340 ();
 DECAPx1_ASAP7_75t_R FILLER_180_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_353 ();
 FILLER_ASAP7_75t_R FILLER_180_360 ();
 DECAPx4_ASAP7_75t_R FILLER_180_368 ();
 DECAPx6_ASAP7_75t_R FILLER_180_386 ();
 DECAPx2_ASAP7_75t_R FILLER_180_400 ();
 DECAPx10_ASAP7_75t_R FILLER_180_409 ();
 DECAPx1_ASAP7_75t_R FILLER_180_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_435 ();
 DECAPx6_ASAP7_75t_R FILLER_180_443 ();
 DECAPx1_ASAP7_75t_R FILLER_180_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_461 ();
 DECAPx6_ASAP7_75t_R FILLER_180_472 ();
 DECAPx2_ASAP7_75t_R FILLER_180_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_492 ();
 DECAPx2_ASAP7_75t_R FILLER_180_503 ();
 DECAPx2_ASAP7_75t_R FILLER_180_527 ();
 DECAPx10_ASAP7_75t_R FILLER_180_549 ();
 DECAPx2_ASAP7_75t_R FILLER_180_571 ();
 FILLER_ASAP7_75t_R FILLER_180_577 ();
 DECAPx2_ASAP7_75t_R FILLER_180_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_588 ();
 DECAPx10_ASAP7_75t_R FILLER_180_595 ();
 DECAPx2_ASAP7_75t_R FILLER_180_617 ();
 FILLER_ASAP7_75t_R FILLER_180_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_625 ();
 DECAPx4_ASAP7_75t_R FILLER_180_638 ();
 FILLER_ASAP7_75t_R FILLER_180_648 ();
 DECAPx6_ASAP7_75t_R FILLER_180_656 ();
 DECAPx1_ASAP7_75t_R FILLER_180_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_674 ();
 DECAPx2_ASAP7_75t_R FILLER_180_681 ();
 FILLER_ASAP7_75t_R FILLER_180_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_689 ();
 FILLER_ASAP7_75t_R FILLER_180_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_699 ();
 FILLER_ASAP7_75t_R FILLER_180_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_714 ();
 DECAPx6_ASAP7_75t_R FILLER_180_727 ();
 DECAPx1_ASAP7_75t_R FILLER_180_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_745 ();
 DECAPx2_ASAP7_75t_R FILLER_180_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_760 ();
 DECAPx1_ASAP7_75t_R FILLER_180_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_778 ();
 DECAPx2_ASAP7_75t_R FILLER_180_788 ();
 FILLER_ASAP7_75t_R FILLER_180_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_796 ();
 DECAPx4_ASAP7_75t_R FILLER_180_803 ();
 DECAPx10_ASAP7_75t_R FILLER_180_820 ();
 DECAPx2_ASAP7_75t_R FILLER_180_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_848 ();
 DECAPx4_ASAP7_75t_R FILLER_180_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_890 ();
 FILLER_ASAP7_75t_R FILLER_180_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_903 ();
 DECAPx4_ASAP7_75t_R FILLER_180_914 ();
 FILLER_ASAP7_75t_R FILLER_180_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_940 ();
 DECAPx2_ASAP7_75t_R FILLER_180_956 ();
 FILLER_ASAP7_75t_R FILLER_180_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_964 ();
 DECAPx6_ASAP7_75t_R FILLER_180_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_997 ();
 FILLER_ASAP7_75t_R FILLER_180_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1033 ();
 FILLER_ASAP7_75t_R FILLER_180_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1116 ();
 FILLER_ASAP7_75t_R FILLER_180_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1204 ();
 FILLER_ASAP7_75t_R FILLER_180_1223 ();
 FILLER_ASAP7_75t_R FILLER_180_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1293 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1313 ();
 FILLER_ASAP7_75t_R FILLER_180_1324 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1366 ();
 FILLER_ASAP7_75t_R FILLER_180_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1388 ();
 FILLER_ASAP7_75t_R FILLER_180_1394 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1399 ();
 DECAPx2_ASAP7_75t_R FILLER_181_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_8 ();
 DECAPx2_ASAP7_75t_R FILLER_181_67 ();
 FILLER_ASAP7_75t_R FILLER_181_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_101 ();
 DECAPx2_ASAP7_75t_R FILLER_181_105 ();
 FILLER_ASAP7_75t_R FILLER_181_123 ();
 DECAPx6_ASAP7_75t_R FILLER_181_128 ();
 DECAPx2_ASAP7_75t_R FILLER_181_142 ();
 DECAPx2_ASAP7_75t_R FILLER_181_158 ();
 DECAPx6_ASAP7_75t_R FILLER_181_180 ();
 DECAPx1_ASAP7_75t_R FILLER_181_194 ();
 FILLER_ASAP7_75t_R FILLER_181_206 ();
 FILLER_ASAP7_75t_R FILLER_181_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_216 ();
 DECAPx4_ASAP7_75t_R FILLER_181_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_244 ();
 DECAPx2_ASAP7_75t_R FILLER_181_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_257 ();
 DECAPx1_ASAP7_75t_R FILLER_181_265 ();
 DECAPx2_ASAP7_75t_R FILLER_181_272 ();
 FILLER_ASAP7_75t_R FILLER_181_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_286 ();
 DECAPx10_ASAP7_75t_R FILLER_181_290 ();
 DECAPx6_ASAP7_75t_R FILLER_181_312 ();
 DECAPx2_ASAP7_75t_R FILLER_181_326 ();
 DECAPx2_ASAP7_75t_R FILLER_181_339 ();
 FILLER_ASAP7_75t_R FILLER_181_345 ();
 DECAPx1_ASAP7_75t_R FILLER_181_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_357 ();
 DECAPx2_ASAP7_75t_R FILLER_181_374 ();
 FILLER_ASAP7_75t_R FILLER_181_380 ();
 DECAPx2_ASAP7_75t_R FILLER_181_392 ();
 DECAPx4_ASAP7_75t_R FILLER_181_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_428 ();
 FILLER_ASAP7_75t_R FILLER_181_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_437 ();
 DECAPx4_ASAP7_75t_R FILLER_181_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_454 ();
 DECAPx1_ASAP7_75t_R FILLER_181_493 ();
 DECAPx6_ASAP7_75t_R FILLER_181_507 ();
 FILLER_ASAP7_75t_R FILLER_181_521 ();
 DECAPx1_ASAP7_75t_R FILLER_181_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_549 ();
 DECAPx6_ASAP7_75t_R FILLER_181_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_570 ();
 DECAPx2_ASAP7_75t_R FILLER_181_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_587 ();
 DECAPx1_ASAP7_75t_R FILLER_181_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_618 ();
 DECAPx6_ASAP7_75t_R FILLER_181_627 ();
 FILLER_ASAP7_75t_R FILLER_181_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_643 ();
 FILLER_ASAP7_75t_R FILLER_181_658 ();
 FILLER_ASAP7_75t_R FILLER_181_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_700 ();
 DECAPx4_ASAP7_75t_R FILLER_181_717 ();
 FILLER_ASAP7_75t_R FILLER_181_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_737 ();
 DECAPx10_ASAP7_75t_R FILLER_181_745 ();
 DECAPx2_ASAP7_75t_R FILLER_181_767 ();
 FILLER_ASAP7_75t_R FILLER_181_787 ();
 DECAPx2_ASAP7_75t_R FILLER_181_797 ();
 FILLER_ASAP7_75t_R FILLER_181_803 ();
 DECAPx4_ASAP7_75t_R FILLER_181_823 ();
 FILLER_ASAP7_75t_R FILLER_181_833 ();
 DECAPx2_ASAP7_75t_R FILLER_181_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_856 ();
 DECAPx6_ASAP7_75t_R FILLER_181_867 ();
 FILLER_ASAP7_75t_R FILLER_181_881 ();
 DECAPx10_ASAP7_75t_R FILLER_181_902 ();
 FILLER_ASAP7_75t_R FILLER_181_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_936 ();
 DECAPx1_ASAP7_75t_R FILLER_181_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_960 ();
 FILLER_ASAP7_75t_R FILLER_181_979 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1047 ();
 FILLER_ASAP7_75t_R FILLER_181_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1059 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1116 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1133 ();
 FILLER_ASAP7_75t_R FILLER_181_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1153 ();
 FILLER_ASAP7_75t_R FILLER_181_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1288 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1379 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1393 ();
 FILLER_ASAP7_75t_R FILLER_181_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_182_2 ();
 DECAPx6_ASAP7_75t_R FILLER_182_30 ();
 DECAPx2_ASAP7_75t_R FILLER_182_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_53 ();
 DECAPx6_ASAP7_75t_R FILLER_182_60 ();
 DECAPx2_ASAP7_75t_R FILLER_182_80 ();
 FILLER_ASAP7_75t_R FILLER_182_86 ();
 DECAPx4_ASAP7_75t_R FILLER_182_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_109 ();
 FILLER_ASAP7_75t_R FILLER_182_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_138 ();
 DECAPx2_ASAP7_75t_R FILLER_182_142 ();
 DECAPx1_ASAP7_75t_R FILLER_182_155 ();
 DECAPx4_ASAP7_75t_R FILLER_182_162 ();
 DECAPx2_ASAP7_75t_R FILLER_182_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_187 ();
 FILLER_ASAP7_75t_R FILLER_182_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_240 ();
 DECAPx6_ASAP7_75t_R FILLER_182_281 ();
 FILLER_ASAP7_75t_R FILLER_182_295 ();
 DECAPx10_ASAP7_75t_R FILLER_182_313 ();
 DECAPx10_ASAP7_75t_R FILLER_182_335 ();
 DECAPx10_ASAP7_75t_R FILLER_182_357 ();
 DECAPx4_ASAP7_75t_R FILLER_182_379 ();
 FILLER_ASAP7_75t_R FILLER_182_389 ();
 FILLER_ASAP7_75t_R FILLER_182_417 ();
 DECAPx4_ASAP7_75t_R FILLER_182_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_461 ();
 DECAPx6_ASAP7_75t_R FILLER_182_464 ();
 FILLER_ASAP7_75t_R FILLER_182_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_480 ();
 DECAPx4_ASAP7_75t_R FILLER_182_487 ();
 FILLER_ASAP7_75t_R FILLER_182_497 ();
 DECAPx4_ASAP7_75t_R FILLER_182_506 ();
 FILLER_ASAP7_75t_R FILLER_182_516 ();
 FILLER_ASAP7_75t_R FILLER_182_532 ();
 FILLER_ASAP7_75t_R FILLER_182_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_574 ();
 DECAPx2_ASAP7_75t_R FILLER_182_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_601 ();
 FILLER_ASAP7_75t_R FILLER_182_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_607 ();
 FILLER_ASAP7_75t_R FILLER_182_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_620 ();
 DECAPx1_ASAP7_75t_R FILLER_182_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_661 ();
 DECAPx4_ASAP7_75t_R FILLER_182_670 ();
 FILLER_ASAP7_75t_R FILLER_182_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_682 ();
 DECAPx10_ASAP7_75t_R FILLER_182_693 ();
 DECAPx6_ASAP7_75t_R FILLER_182_715 ();
 DECAPx1_ASAP7_75t_R FILLER_182_729 ();
 DECAPx10_ASAP7_75t_R FILLER_182_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_762 ();
 DECAPx4_ASAP7_75t_R FILLER_182_770 ();
 FILLER_ASAP7_75t_R FILLER_182_786 ();
 DECAPx1_ASAP7_75t_R FILLER_182_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_834 ();
 DECAPx4_ASAP7_75t_R FILLER_182_843 ();
 DECAPx10_ASAP7_75t_R FILLER_182_865 ();
 DECAPx6_ASAP7_75t_R FILLER_182_887 ();
 DECAPx1_ASAP7_75t_R FILLER_182_911 ();
 FILLER_ASAP7_75t_R FILLER_182_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_923 ();
 DECAPx2_ASAP7_75t_R FILLER_182_932 ();
 FILLER_ASAP7_75t_R FILLER_182_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_940 ();
 DECAPx10_ASAP7_75t_R FILLER_182_957 ();
 DECAPx10_ASAP7_75t_R FILLER_182_979 ();
 FILLER_ASAP7_75t_R FILLER_182_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1061 ();
 FILLER_ASAP7_75t_R FILLER_182_1071 ();
 FILLER_ASAP7_75t_R FILLER_182_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1214 ();
 FILLER_ASAP7_75t_R FILLER_182_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1236 ();
 FILLER_ASAP7_75t_R FILLER_182_1242 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1257 ();
 FILLER_ASAP7_75t_R FILLER_182_1298 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1339 ();
 FILLER_ASAP7_75t_R FILLER_182_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1388 ();
 FILLER_ASAP7_75t_R FILLER_182_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1396 ();
 DECAPx10_ASAP7_75t_R FILLER_183_2 ();
 DECAPx1_ASAP7_75t_R FILLER_183_24 ();
 DECAPx4_ASAP7_75t_R FILLER_183_34 ();
 FILLER_ASAP7_75t_R FILLER_183_44 ();
 DECAPx1_ASAP7_75t_R FILLER_183_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_82 ();
 DECAPx4_ASAP7_75t_R FILLER_183_109 ();
 DECAPx1_ASAP7_75t_R FILLER_183_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_130 ();
 DECAPx2_ASAP7_75t_R FILLER_183_190 ();
 FILLER_ASAP7_75t_R FILLER_183_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_214 ();
 DECAPx2_ASAP7_75t_R FILLER_183_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_241 ();
 FILLER_ASAP7_75t_R FILLER_183_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_258 ();
 DECAPx4_ASAP7_75t_R FILLER_183_265 ();
 DECAPx1_ASAP7_75t_R FILLER_183_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_286 ();
 DECAPx1_ASAP7_75t_R FILLER_183_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_294 ();
 DECAPx2_ASAP7_75t_R FILLER_183_321 ();
 FILLER_ASAP7_75t_R FILLER_183_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_329 ();
 DECAPx4_ASAP7_75t_R FILLER_183_338 ();
 FILLER_ASAP7_75t_R FILLER_183_348 ();
 DECAPx10_ASAP7_75t_R FILLER_183_356 ();
 DECAPx2_ASAP7_75t_R FILLER_183_378 ();
 FILLER_ASAP7_75t_R FILLER_183_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_386 ();
 DECAPx2_ASAP7_75t_R FILLER_183_393 ();
 FILLER_ASAP7_75t_R FILLER_183_399 ();
 DECAPx10_ASAP7_75t_R FILLER_183_417 ();
 FILLER_ASAP7_75t_R FILLER_183_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_444 ();
 DECAPx6_ASAP7_75t_R FILLER_183_451 ();
 FILLER_ASAP7_75t_R FILLER_183_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_467 ();
 DECAPx4_ASAP7_75t_R FILLER_183_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_494 ();
 DECAPx4_ASAP7_75t_R FILLER_183_506 ();
 FILLER_ASAP7_75t_R FILLER_183_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_518 ();
 DECAPx6_ASAP7_75t_R FILLER_183_533 ();
 FILLER_ASAP7_75t_R FILLER_183_547 ();
 DECAPx1_ASAP7_75t_R FILLER_183_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_559 ();
 DECAPx2_ASAP7_75t_R FILLER_183_563 ();
 FILLER_ASAP7_75t_R FILLER_183_569 ();
 DECAPx2_ASAP7_75t_R FILLER_183_581 ();
 FILLER_ASAP7_75t_R FILLER_183_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_589 ();
 DECAPx4_ASAP7_75t_R FILLER_183_596 ();
 FILLER_ASAP7_75t_R FILLER_183_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_608 ();
 DECAPx1_ASAP7_75t_R FILLER_183_622 ();
 DECAPx6_ASAP7_75t_R FILLER_183_632 ();
 DECAPx10_ASAP7_75t_R FILLER_183_649 ();
 DECAPx4_ASAP7_75t_R FILLER_183_671 ();
 FILLER_ASAP7_75t_R FILLER_183_681 ();
 DECAPx10_ASAP7_75t_R FILLER_183_690 ();
 DECAPx2_ASAP7_75t_R FILLER_183_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_718 ();
 DECAPx6_ASAP7_75t_R FILLER_183_726 ();
 DECAPx1_ASAP7_75t_R FILLER_183_740 ();
 DECAPx6_ASAP7_75t_R FILLER_183_758 ();
 DECAPx1_ASAP7_75t_R FILLER_183_772 ();
 DECAPx10_ASAP7_75t_R FILLER_183_783 ();
 FILLER_ASAP7_75t_R FILLER_183_805 ();
 DECAPx6_ASAP7_75t_R FILLER_183_813 ();
 FILLER_ASAP7_75t_R FILLER_183_827 ();
 FILLER_ASAP7_75t_R FILLER_183_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_853 ();
 DECAPx2_ASAP7_75t_R FILLER_183_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_892 ();
 DECAPx6_ASAP7_75t_R FILLER_183_906 ();
 DECAPx1_ASAP7_75t_R FILLER_183_920 ();
 DECAPx10_ASAP7_75t_R FILLER_183_926 ();
 DECAPx10_ASAP7_75t_R FILLER_183_948 ();
 DECAPx10_ASAP7_75t_R FILLER_183_970 ();
 DECAPx10_ASAP7_75t_R FILLER_183_992 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1036 ();
 FILLER_ASAP7_75t_R FILLER_183_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1101 ();
 FILLER_ASAP7_75t_R FILLER_183_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1188 ();
 FILLER_ASAP7_75t_R FILLER_183_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1229 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1256 ();
 FILLER_ASAP7_75t_R FILLER_183_1270 ();
 FILLER_ASAP7_75t_R FILLER_183_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1277 ();
 FILLER_ASAP7_75t_R FILLER_183_1326 ();
 FILLER_ASAP7_75t_R FILLER_183_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1378 ();
 DECAPx6_ASAP7_75t_R FILLER_184_2 ();
 DECAPx6_ASAP7_75t_R FILLER_184_42 ();
 DECAPx1_ASAP7_75t_R FILLER_184_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_60 ();
 DECAPx2_ASAP7_75t_R FILLER_184_64 ();
 FILLER_ASAP7_75t_R FILLER_184_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_72 ();
 DECAPx4_ASAP7_75t_R FILLER_184_79 ();
 FILLER_ASAP7_75t_R FILLER_184_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_97 ();
 DECAPx1_ASAP7_75t_R FILLER_184_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_105 ();
 DECAPx2_ASAP7_75t_R FILLER_184_138 ();
 FILLER_ASAP7_75t_R FILLER_184_144 ();
 FILLER_ASAP7_75t_R FILLER_184_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_151 ();
 DECAPx6_ASAP7_75t_R FILLER_184_158 ();
 DECAPx1_ASAP7_75t_R FILLER_184_172 ();
 DECAPx1_ASAP7_75t_R FILLER_184_179 ();
 DECAPx6_ASAP7_75t_R FILLER_184_189 ();
 DECAPx1_ASAP7_75t_R FILLER_184_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_213 ();
 FILLER_ASAP7_75t_R FILLER_184_224 ();
 DECAPx4_ASAP7_75t_R FILLER_184_233 ();
 FILLER_ASAP7_75t_R FILLER_184_243 ();
 DECAPx10_ASAP7_75t_R FILLER_184_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_305 ();
 DECAPx4_ASAP7_75t_R FILLER_184_321 ();
 FILLER_ASAP7_75t_R FILLER_184_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_333 ();
 DECAPx4_ASAP7_75t_R FILLER_184_337 ();
 FILLER_ASAP7_75t_R FILLER_184_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_355 ();
 DECAPx1_ASAP7_75t_R FILLER_184_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_374 ();
 FILLER_ASAP7_75t_R FILLER_184_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_383 ();
 DECAPx10_ASAP7_75t_R FILLER_184_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_414 ();
 DECAPx4_ASAP7_75t_R FILLER_184_429 ();
 FILLER_ASAP7_75t_R FILLER_184_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_441 ();
 DECAPx6_ASAP7_75t_R FILLER_184_448 ();
 DECAPx4_ASAP7_75t_R FILLER_184_464 ();
 FILLER_ASAP7_75t_R FILLER_184_474 ();
 DECAPx10_ASAP7_75t_R FILLER_184_482 ();
 DECAPx6_ASAP7_75t_R FILLER_184_504 ();
 DECAPx1_ASAP7_75t_R FILLER_184_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_537 ();
 DECAPx10_ASAP7_75t_R FILLER_184_548 ();
 FILLER_ASAP7_75t_R FILLER_184_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_572 ();
 FILLER_ASAP7_75t_R FILLER_184_583 ();
 DECAPx1_ASAP7_75t_R FILLER_184_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_642 ();
 DECAPx4_ASAP7_75t_R FILLER_184_646 ();
 DECAPx4_ASAP7_75t_R FILLER_184_664 ();
 FILLER_ASAP7_75t_R FILLER_184_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_686 ();
 FILLER_ASAP7_75t_R FILLER_184_696 ();
 DECAPx2_ASAP7_75t_R FILLER_184_704 ();
 FILLER_ASAP7_75t_R FILLER_184_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_712 ();
 DECAPx1_ASAP7_75t_R FILLER_184_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_739 ();
 DECAPx4_ASAP7_75t_R FILLER_184_752 ();
 FILLER_ASAP7_75t_R FILLER_184_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_764 ();
 DECAPx1_ASAP7_75t_R FILLER_184_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_775 ();
 DECAPx10_ASAP7_75t_R FILLER_184_794 ();
 DECAPx2_ASAP7_75t_R FILLER_184_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_856 ();
 DECAPx1_ASAP7_75t_R FILLER_184_867 ();
 DECAPx2_ASAP7_75t_R FILLER_184_887 ();
 FILLER_ASAP7_75t_R FILLER_184_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_908 ();
 DECAPx2_ASAP7_75t_R FILLER_184_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_957 ();
 FILLER_ASAP7_75t_R FILLER_184_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_966 ();
 DECAPx4_ASAP7_75t_R FILLER_184_973 ();
 FILLER_ASAP7_75t_R FILLER_184_983 ();
 DECAPx4_ASAP7_75t_R FILLER_184_999 ();
 FILLER_ASAP7_75t_R FILLER_184_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1082 ();
 FILLER_ASAP7_75t_R FILLER_184_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1114 ();
 FILLER_ASAP7_75t_R FILLER_184_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_184_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1236 ();
 FILLER_ASAP7_75t_R FILLER_184_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1303 ();
 FILLER_ASAP7_75t_R FILLER_184_1309 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1359 ();
 FILLER_ASAP7_75t_R FILLER_184_1373 ();
 FILLER_ASAP7_75t_R FILLER_184_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1385 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1388 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1404 ();
 DECAPx6_ASAP7_75t_R FILLER_185_2 ();
 DECAPx2_ASAP7_75t_R FILLER_185_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_22 ();
 FILLER_ASAP7_75t_R FILLER_185_29 ();
 FILLER_ASAP7_75t_R FILLER_185_34 ();
 DECAPx4_ASAP7_75t_R FILLER_185_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_62 ();
 DECAPx6_ASAP7_75t_R FILLER_185_95 ();
 FILLER_ASAP7_75t_R FILLER_185_109 ();
 DECAPx1_ASAP7_75t_R FILLER_185_114 ();
 FILLER_ASAP7_75t_R FILLER_185_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_130 ();
 DECAPx6_ASAP7_75t_R FILLER_185_147 ();
 DECAPx1_ASAP7_75t_R FILLER_185_194 ();
 FILLER_ASAP7_75t_R FILLER_185_212 ();
 FILLER_ASAP7_75t_R FILLER_185_236 ();
 DECAPx6_ASAP7_75t_R FILLER_185_244 ();
 FILLER_ASAP7_75t_R FILLER_185_258 ();
 DECAPx1_ASAP7_75t_R FILLER_185_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_276 ();
 DECAPx10_ASAP7_75t_R FILLER_185_283 ();
 DECAPx10_ASAP7_75t_R FILLER_185_305 ();
 DECAPx10_ASAP7_75t_R FILLER_185_327 ();
 DECAPx2_ASAP7_75t_R FILLER_185_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_355 ();
 FILLER_ASAP7_75t_R FILLER_185_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_366 ();
 DECAPx10_ASAP7_75t_R FILLER_185_399 ();
 DECAPx6_ASAP7_75t_R FILLER_185_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_435 ();
 DECAPx4_ASAP7_75t_R FILLER_185_450 ();
 FILLER_ASAP7_75t_R FILLER_185_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_462 ();
 DECAPx1_ASAP7_75t_R FILLER_185_488 ();
 DECAPx10_ASAP7_75t_R FILLER_185_498 ();
 DECAPx6_ASAP7_75t_R FILLER_185_520 ();
 DECAPx6_ASAP7_75t_R FILLER_185_547 ();
 FILLER_ASAP7_75t_R FILLER_185_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_563 ();
 DECAPx4_ASAP7_75t_R FILLER_185_576 ();
 FILLER_ASAP7_75t_R FILLER_185_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_588 ();
 FILLER_ASAP7_75t_R FILLER_185_621 ();
 DECAPx1_ASAP7_75t_R FILLER_185_655 ();
 DECAPx4_ASAP7_75t_R FILLER_185_679 ();
 FILLER_ASAP7_75t_R FILLER_185_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_691 ();
 DECAPx2_ASAP7_75t_R FILLER_185_713 ();
 DECAPx10_ASAP7_75t_R FILLER_185_727 ();
 DECAPx10_ASAP7_75t_R FILLER_185_749 ();
 DECAPx4_ASAP7_75t_R FILLER_185_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_781 ();
 DECAPx4_ASAP7_75t_R FILLER_185_788 ();
 FILLER_ASAP7_75t_R FILLER_185_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_800 ();
 DECAPx6_ASAP7_75t_R FILLER_185_815 ();
 DECAPx2_ASAP7_75t_R FILLER_185_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_835 ();
 FILLER_ASAP7_75t_R FILLER_185_839 ();
 DECAPx6_ASAP7_75t_R FILLER_185_844 ();
 DECAPx2_ASAP7_75t_R FILLER_185_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_893 ();
 DECAPx1_ASAP7_75t_R FILLER_185_920 ();
 FILLER_ASAP7_75t_R FILLER_185_926 ();
 DECAPx2_ASAP7_75t_R FILLER_185_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_942 ();
 FILLER_ASAP7_75t_R FILLER_185_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_955 ();
 DECAPx6_ASAP7_75t_R FILLER_185_986 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1064 ();
 FILLER_ASAP7_75t_R FILLER_185_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1191 ();
 FILLER_ASAP7_75t_R FILLER_185_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1267 ();
 FILLER_ASAP7_75t_R FILLER_185_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1331 ();
 FILLER_ASAP7_75t_R FILLER_185_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1399 ();
 DECAPx6_ASAP7_75t_R FILLER_186_2 ();
 DECAPx1_ASAP7_75t_R FILLER_186_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_58 ();
 DECAPx4_ASAP7_75t_R FILLER_186_65 ();
 FILLER_ASAP7_75t_R FILLER_186_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_77 ();
 DECAPx2_ASAP7_75t_R FILLER_186_81 ();
 FILLER_ASAP7_75t_R FILLER_186_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_89 ();
 FILLER_ASAP7_75t_R FILLER_186_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_95 ();
 FILLER_ASAP7_75t_R FILLER_186_120 ();
 FILLER_ASAP7_75t_R FILLER_186_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_157 ();
 DECAPx6_ASAP7_75t_R FILLER_186_164 ();
 DECAPx6_ASAP7_75t_R FILLER_186_192 ();
 DECAPx1_ASAP7_75t_R FILLER_186_220 ();
 FILLER_ASAP7_75t_R FILLER_186_230 ();
 DECAPx1_ASAP7_75t_R FILLER_186_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_244 ();
 DECAPx1_ASAP7_75t_R FILLER_186_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_255 ();
 DECAPx2_ASAP7_75t_R FILLER_186_278 ();
 FILLER_ASAP7_75t_R FILLER_186_284 ();
 DECAPx6_ASAP7_75t_R FILLER_186_292 ();
 DECAPx1_ASAP7_75t_R FILLER_186_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_310 ();
 DECAPx4_ASAP7_75t_R FILLER_186_317 ();
 FILLER_ASAP7_75t_R FILLER_186_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_329 ();
 DECAPx1_ASAP7_75t_R FILLER_186_336 ();
 DECAPx10_ASAP7_75t_R FILLER_186_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_371 ();
 DECAPx1_ASAP7_75t_R FILLER_186_378 ();
 DECAPx2_ASAP7_75t_R FILLER_186_388 ();
 FILLER_ASAP7_75t_R FILLER_186_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_406 ();
 DECAPx2_ASAP7_75t_R FILLER_186_419 ();
 FILLER_ASAP7_75t_R FILLER_186_425 ();
 DECAPx4_ASAP7_75t_R FILLER_186_433 ();
 FILLER_ASAP7_75t_R FILLER_186_443 ();
 DECAPx2_ASAP7_75t_R FILLER_186_453 ();
 FILLER_ASAP7_75t_R FILLER_186_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_461 ();
 FILLER_ASAP7_75t_R FILLER_186_487 ();
 DECAPx4_ASAP7_75t_R FILLER_186_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_528 ();
 DECAPx1_ASAP7_75t_R FILLER_186_587 ();
 DECAPx10_ASAP7_75t_R FILLER_186_647 ();
 DECAPx6_ASAP7_75t_R FILLER_186_669 ();
 FILLER_ASAP7_75t_R FILLER_186_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_685 ();
 DECAPx2_ASAP7_75t_R FILLER_186_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_700 ();
 FILLER_ASAP7_75t_R FILLER_186_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_722 ();
 DECAPx10_ASAP7_75t_R FILLER_186_728 ();
 DECAPx6_ASAP7_75t_R FILLER_186_750 ();
 DECAPx2_ASAP7_75t_R FILLER_186_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_791 ();
 DECAPx2_ASAP7_75t_R FILLER_186_803 ();
 FILLER_ASAP7_75t_R FILLER_186_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_811 ();
 DECAPx6_ASAP7_75t_R FILLER_186_822 ();
 DECAPx1_ASAP7_75t_R FILLER_186_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_840 ();
 DECAPx10_ASAP7_75t_R FILLER_186_847 ();
 DECAPx6_ASAP7_75t_R FILLER_186_869 ();
 DECAPx2_ASAP7_75t_R FILLER_186_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_889 ();
 DECAPx6_ASAP7_75t_R FILLER_186_893 ();
 FILLER_ASAP7_75t_R FILLER_186_907 ();
 DECAPx4_ASAP7_75t_R FILLER_186_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_922 ();
 DECAPx10_ASAP7_75t_R FILLER_186_931 ();
 DECAPx2_ASAP7_75t_R FILLER_186_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_959 ();
 DECAPx2_ASAP7_75t_R FILLER_186_981 ();
 FILLER_ASAP7_75t_R FILLER_186_987 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1077 ();
 FILLER_ASAP7_75t_R FILLER_186_1083 ();
 FILLER_ASAP7_75t_R FILLER_186_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1149 ();
 FILLER_ASAP7_75t_R FILLER_186_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1258 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1304 ();
 FILLER_ASAP7_75t_R FILLER_186_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1312 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1316 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1330 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1357 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1364 ();
 FILLER_ASAP7_75t_R FILLER_186_1378 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1380 ();
 FILLER_ASAP7_75t_R FILLER_186_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1388 ();
 FILLER_ASAP7_75t_R FILLER_186_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1404 ();
 FILLER_ASAP7_75t_R FILLER_187_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_4 ();
 DECAPx4_ASAP7_75t_R FILLER_187_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_41 ();
 FILLER_ASAP7_75t_R FILLER_187_45 ();
 FILLER_ASAP7_75t_R FILLER_187_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_75 ();
 FILLER_ASAP7_75t_R FILLER_187_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_81 ();
 FILLER_ASAP7_75t_R FILLER_187_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_169 ();
 DECAPx4_ASAP7_75t_R FILLER_187_173 ();
 FILLER_ASAP7_75t_R FILLER_187_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_185 ();
 DECAPx4_ASAP7_75t_R FILLER_187_189 ();
 FILLER_ASAP7_75t_R FILLER_187_199 ();
 DECAPx1_ASAP7_75t_R FILLER_187_208 ();
 DECAPx2_ASAP7_75t_R FILLER_187_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_224 ();
 DECAPx1_ASAP7_75t_R FILLER_187_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_239 ();
 DECAPx1_ASAP7_75t_R FILLER_187_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_280 ();
 DECAPx1_ASAP7_75t_R FILLER_187_299 ();
 DECAPx1_ASAP7_75t_R FILLER_187_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_315 ();
 DECAPx1_ASAP7_75t_R FILLER_187_330 ();
 DECAPx10_ASAP7_75t_R FILLER_187_342 ();
 DECAPx10_ASAP7_75t_R FILLER_187_364 ();
 DECAPx4_ASAP7_75t_R FILLER_187_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_396 ();
 DECAPx1_ASAP7_75t_R FILLER_187_435 ();
 DECAPx1_ASAP7_75t_R FILLER_187_458 ();
 FILLER_ASAP7_75t_R FILLER_187_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_480 ();
 DECAPx1_ASAP7_75t_R FILLER_187_487 ();
 DECAPx1_ASAP7_75t_R FILLER_187_497 ();
 DECAPx4_ASAP7_75t_R FILLER_187_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_536 ();
 DECAPx2_ASAP7_75t_R FILLER_187_543 ();
 DECAPx2_ASAP7_75t_R FILLER_187_552 ();
 DECAPx2_ASAP7_75t_R FILLER_187_567 ();
 FILLER_ASAP7_75t_R FILLER_187_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_578 ();
 DECAPx4_ASAP7_75t_R FILLER_187_624 ();
 FILLER_ASAP7_75t_R FILLER_187_634 ();
 DECAPx10_ASAP7_75t_R FILLER_187_639 ();
 DECAPx1_ASAP7_75t_R FILLER_187_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_665 ();
 DECAPx4_ASAP7_75t_R FILLER_187_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_686 ();
 DECAPx4_ASAP7_75t_R FILLER_187_699 ();
 FILLER_ASAP7_75t_R FILLER_187_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_711 ();
 DECAPx10_ASAP7_75t_R FILLER_187_732 ();
 DECAPx6_ASAP7_75t_R FILLER_187_760 ();
 FILLER_ASAP7_75t_R FILLER_187_774 ();
 DECAPx10_ASAP7_75t_R FILLER_187_792 ();
 DECAPx4_ASAP7_75t_R FILLER_187_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_824 ();
 DECAPx6_ASAP7_75t_R FILLER_187_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_846 ();
 DECAPx2_ASAP7_75t_R FILLER_187_859 ();
 FILLER_ASAP7_75t_R FILLER_187_865 ();
 FILLER_ASAP7_75t_R FILLER_187_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_882 ();
 DECAPx10_ASAP7_75t_R FILLER_187_898 ();
 DECAPx1_ASAP7_75t_R FILLER_187_920 ();
 FILLER_ASAP7_75t_R FILLER_187_926 ();
 DECAPx4_ASAP7_75t_R FILLER_187_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_944 ();
 DECAPx4_ASAP7_75t_R FILLER_187_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_961 ();
 DECAPx1_ASAP7_75t_R FILLER_187_965 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1025 ();
 FILLER_ASAP7_75t_R FILLER_187_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1095 ();
 FILLER_ASAP7_75t_R FILLER_187_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1201 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1236 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1243 ();
 FILLER_ASAP7_75t_R FILLER_187_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1293 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1368 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1382 ();
 DECAPx6_ASAP7_75t_R FILLER_188_2 ();
 FILLER_ASAP7_75t_R FILLER_188_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_18 ();
 FILLER_ASAP7_75t_R FILLER_188_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_50 ();
 DECAPx1_ASAP7_75t_R FILLER_188_94 ();
 FILLER_ASAP7_75t_R FILLER_188_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_103 ();
 DECAPx1_ASAP7_75t_R FILLER_188_136 ();
 DECAPx4_ASAP7_75t_R FILLER_188_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_156 ();
 FILLER_ASAP7_75t_R FILLER_188_167 ();
 DECAPx1_ASAP7_75t_R FILLER_188_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_176 ();
 DECAPx2_ASAP7_75t_R FILLER_188_183 ();
 FILLER_ASAP7_75t_R FILLER_188_189 ();
 DECAPx2_ASAP7_75t_R FILLER_188_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_225 ();
 FILLER_ASAP7_75t_R FILLER_188_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_254 ();
 DECAPx10_ASAP7_75t_R FILLER_188_261 ();
 FILLER_ASAP7_75t_R FILLER_188_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_300 ();
 DECAPx10_ASAP7_75t_R FILLER_188_307 ();
 DECAPx10_ASAP7_75t_R FILLER_188_329 ();
 DECAPx2_ASAP7_75t_R FILLER_188_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_357 ();
 FILLER_ASAP7_75t_R FILLER_188_378 ();
 DECAPx4_ASAP7_75t_R FILLER_188_386 ();
 FILLER_ASAP7_75t_R FILLER_188_396 ();
 FILLER_ASAP7_75t_R FILLER_188_416 ();
 FILLER_ASAP7_75t_R FILLER_188_450 ();
 DECAPx1_ASAP7_75t_R FILLER_188_458 ();
 DECAPx10_ASAP7_75t_R FILLER_188_477 ();
 DECAPx1_ASAP7_75t_R FILLER_188_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_503 ();
 DECAPx1_ASAP7_75t_R FILLER_188_507 ();
 DECAPx2_ASAP7_75t_R FILLER_188_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_537 ();
 DECAPx2_ASAP7_75t_R FILLER_188_544 ();
 FILLER_ASAP7_75t_R FILLER_188_550 ();
 DECAPx2_ASAP7_75t_R FILLER_188_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_584 ();
 DECAPx4_ASAP7_75t_R FILLER_188_614 ();
 FILLER_ASAP7_75t_R FILLER_188_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_649 ();
 DECAPx4_ASAP7_75t_R FILLER_188_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_670 ();
 DECAPx10_ASAP7_75t_R FILLER_188_677 ();
 DECAPx10_ASAP7_75t_R FILLER_188_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_721 ();
 DECAPx6_ASAP7_75t_R FILLER_188_769 ();
 DECAPx2_ASAP7_75t_R FILLER_188_783 ();
 DECAPx10_ASAP7_75t_R FILLER_188_796 ();
 FILLER_ASAP7_75t_R FILLER_188_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_820 ();
 DECAPx2_ASAP7_75t_R FILLER_188_859 ();
 FILLER_ASAP7_75t_R FILLER_188_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_893 ();
 DECAPx4_ASAP7_75t_R FILLER_188_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_957 ();
 DECAPx6_ASAP7_75t_R FILLER_188_973 ();
 DECAPx1_ASAP7_75t_R FILLER_188_987 ();
 FILLER_ASAP7_75t_R FILLER_188_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_996 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1005 ();
 FILLER_ASAP7_75t_R FILLER_188_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_188_1080 ();
 FILLER_ASAP7_75t_R FILLER_188_1090 ();
 FILLER_ASAP7_75t_R FILLER_188_1102 ();
 FILLER_ASAP7_75t_R FILLER_188_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1146 ();
 FILLER_ASAP7_75t_R FILLER_188_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_188_1248 ();
 FILLER_ASAP7_75t_R FILLER_188_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1284 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1318 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1339 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1354 ();
 FILLER_ASAP7_75t_R FILLER_188_1384 ();
 DECAPx4_ASAP7_75t_R FILLER_188_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1404 ();
 FILLER_ASAP7_75t_R FILLER_189_2 ();
 FILLER_ASAP7_75t_R FILLER_189_67 ();
 DECAPx2_ASAP7_75t_R FILLER_189_76 ();
 FILLER_ASAP7_75t_R FILLER_189_82 ();
 FILLER_ASAP7_75t_R FILLER_189_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_112 ();
 FILLER_ASAP7_75t_R FILLER_189_116 ();
 FILLER_ASAP7_75t_R FILLER_189_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_123 ();
 DECAPx1_ASAP7_75t_R FILLER_189_150 ();
 DECAPx1_ASAP7_75t_R FILLER_189_180 ();
 DECAPx1_ASAP7_75t_R FILLER_189_198 ();
 DECAPx2_ASAP7_75t_R FILLER_189_230 ();
 DECAPx10_ASAP7_75t_R FILLER_189_250 ();
 DECAPx10_ASAP7_75t_R FILLER_189_272 ();
 DECAPx10_ASAP7_75t_R FILLER_189_294 ();
 DECAPx6_ASAP7_75t_R FILLER_189_316 ();
 FILLER_ASAP7_75t_R FILLER_189_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_332 ();
 FILLER_ASAP7_75t_R FILLER_189_341 ();
 DECAPx6_ASAP7_75t_R FILLER_189_351 ();
 DECAPx2_ASAP7_75t_R FILLER_189_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_371 ();
 DECAPx10_ASAP7_75t_R FILLER_189_378 ();
 DECAPx10_ASAP7_75t_R FILLER_189_400 ();
 DECAPx4_ASAP7_75t_R FILLER_189_422 ();
 FILLER_ASAP7_75t_R FILLER_189_432 ();
 DECAPx10_ASAP7_75t_R FILLER_189_462 ();
 DECAPx10_ASAP7_75t_R FILLER_189_484 ();
 FILLER_ASAP7_75t_R FILLER_189_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_508 ();
 DECAPx1_ASAP7_75t_R FILLER_189_521 ();
 FILLER_ASAP7_75t_R FILLER_189_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_537 ();
 DECAPx2_ASAP7_75t_R FILLER_189_560 ();
 DECAPx1_ASAP7_75t_R FILLER_189_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_605 ();
 DECAPx6_ASAP7_75t_R FILLER_189_612 ();
 DECAPx2_ASAP7_75t_R FILLER_189_626 ();
 DECAPx2_ASAP7_75t_R FILLER_189_662 ();
 DECAPx10_ASAP7_75t_R FILLER_189_674 ();
 DECAPx2_ASAP7_75t_R FILLER_189_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_718 ();
 DECAPx10_ASAP7_75t_R FILLER_189_726 ();
 DECAPx4_ASAP7_75t_R FILLER_189_748 ();
 FILLER_ASAP7_75t_R FILLER_189_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_760 ();
 DECAPx10_ASAP7_75t_R FILLER_189_771 ();
 DECAPx10_ASAP7_75t_R FILLER_189_793 ();
 DECAPx4_ASAP7_75t_R FILLER_189_815 ();
 DECAPx4_ASAP7_75t_R FILLER_189_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_850 ();
 FILLER_ASAP7_75t_R FILLER_189_863 ();
 DECAPx1_ASAP7_75t_R FILLER_189_877 ();
 DECAPx2_ASAP7_75t_R FILLER_189_884 ();
 FILLER_ASAP7_75t_R FILLER_189_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_904 ();
 FILLER_ASAP7_75t_R FILLER_189_926 ();
 FILLER_ASAP7_75t_R FILLER_189_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_971 ();
 DECAPx6_ASAP7_75t_R FILLER_189_981 ();
 DECAPx1_ASAP7_75t_R FILLER_189_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_999 ();
 FILLER_ASAP7_75t_R FILLER_189_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1057 ();
 FILLER_ASAP7_75t_R FILLER_189_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1071 ();
 FILLER_ASAP7_75t_R FILLER_189_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1082 ();
 FILLER_ASAP7_75t_R FILLER_189_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1227 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1254 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1272 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1289 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1332 ();
 FILLER_ASAP7_75t_R FILLER_189_1338 ();
 FILLER_ASAP7_75t_R FILLER_189_1377 ();
 DECAPx6_ASAP7_75t_R FILLER_190_2 ();
 FILLER_ASAP7_75t_R FILLER_190_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_18 ();
 FILLER_ASAP7_75t_R FILLER_190_60 ();
 DECAPx2_ASAP7_75t_R FILLER_190_65 ();
 FILLER_ASAP7_75t_R FILLER_190_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_73 ();
 DECAPx4_ASAP7_75t_R FILLER_190_80 ();
 DECAPx4_ASAP7_75t_R FILLER_190_96 ();
 DECAPx6_ASAP7_75t_R FILLER_190_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_127 ();
 DECAPx1_ASAP7_75t_R FILLER_190_135 ();
 DECAPx10_ASAP7_75t_R FILLER_190_142 ();
 DECAPx1_ASAP7_75t_R FILLER_190_164 ();
 DECAPx4_ASAP7_75t_R FILLER_190_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_190 ();
 DECAPx2_ASAP7_75t_R FILLER_190_197 ();
 FILLER_ASAP7_75t_R FILLER_190_203 ();
 FILLER_ASAP7_75t_R FILLER_190_219 ();
 DECAPx1_ASAP7_75t_R FILLER_190_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_235 ();
 DECAPx10_ASAP7_75t_R FILLER_190_244 ();
 DECAPx10_ASAP7_75t_R FILLER_190_273 ();
 DECAPx4_ASAP7_75t_R FILLER_190_295 ();
 DECAPx2_ASAP7_75t_R FILLER_190_311 ();
 DECAPx4_ASAP7_75t_R FILLER_190_323 ();
 FILLER_ASAP7_75t_R FILLER_190_371 ();
 FILLER_ASAP7_75t_R FILLER_190_381 ();
 DECAPx4_ASAP7_75t_R FILLER_190_405 ();
 FILLER_ASAP7_75t_R FILLER_190_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_431 ();
 DECAPx6_ASAP7_75t_R FILLER_190_464 ();
 DECAPx2_ASAP7_75t_R FILLER_190_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_484 ();
 DECAPx10_ASAP7_75t_R FILLER_190_499 ();
 DECAPx6_ASAP7_75t_R FILLER_190_521 ();
 DECAPx1_ASAP7_75t_R FILLER_190_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_549 ();
 DECAPx4_ASAP7_75t_R FILLER_190_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_566 ();
 DECAPx2_ASAP7_75t_R FILLER_190_573 ();
 FILLER_ASAP7_75t_R FILLER_190_579 ();
 DECAPx4_ASAP7_75t_R FILLER_190_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_621 ();
 DECAPx10_ASAP7_75t_R FILLER_190_644 ();
 DECAPx2_ASAP7_75t_R FILLER_190_666 ();
 FILLER_ASAP7_75t_R FILLER_190_672 ();
 FILLER_ASAP7_75t_R FILLER_190_679 ();
 DECAPx2_ASAP7_75t_R FILLER_190_692 ();
 FILLER_ASAP7_75t_R FILLER_190_698 ();
 DECAPx10_ASAP7_75t_R FILLER_190_723 ();
 DECAPx6_ASAP7_75t_R FILLER_190_745 ();
 DECAPx1_ASAP7_75t_R FILLER_190_759 ();
 DECAPx10_ASAP7_75t_R FILLER_190_772 ();
 DECAPx2_ASAP7_75t_R FILLER_190_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_800 ();
 DECAPx6_ASAP7_75t_R FILLER_190_813 ();
 FILLER_ASAP7_75t_R FILLER_190_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_829 ();
 DECAPx10_ASAP7_75t_R FILLER_190_843 ();
 DECAPx4_ASAP7_75t_R FILLER_190_865 ();
 FILLER_ASAP7_75t_R FILLER_190_875 ();
 FILLER_ASAP7_75t_R FILLER_190_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_888 ();
 DECAPx4_ASAP7_75t_R FILLER_190_892 ();
 FILLER_ASAP7_75t_R FILLER_190_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_938 ();
 DECAPx2_ASAP7_75t_R FILLER_190_951 ();
 FILLER_ASAP7_75t_R FILLER_190_957 ();
 FILLER_ASAP7_75t_R FILLER_190_971 ();
 DECAPx6_ASAP7_75t_R FILLER_190_993 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1036 ();
 FILLER_ASAP7_75t_R FILLER_190_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1063 ();
 FILLER_ASAP7_75t_R FILLER_190_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1108 ();
 FILLER_ASAP7_75t_R FILLER_190_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1133 ();
 FILLER_ASAP7_75t_R FILLER_190_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1241 ();
 FILLER_ASAP7_75t_R FILLER_190_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1312 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1339 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1385 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1388 ();
 FILLER_ASAP7_75t_R FILLER_190_1394 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_191_2 ();
 DECAPx4_ASAP7_75t_R FILLER_191_24 ();
 FILLER_ASAP7_75t_R FILLER_191_34 ();
 DECAPx2_ASAP7_75t_R FILLER_191_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_48 ();
 FILLER_ASAP7_75t_R FILLER_191_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_60 ();
 DECAPx1_ASAP7_75t_R FILLER_191_64 ();
 DECAPx2_ASAP7_75t_R FILLER_191_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_80 ();
 DECAPx2_ASAP7_75t_R FILLER_191_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_132 ();
 FILLER_ASAP7_75t_R FILLER_191_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_148 ();
 DECAPx1_ASAP7_75t_R FILLER_191_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_159 ();
 DECAPx2_ASAP7_75t_R FILLER_191_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_169 ();
 DECAPx6_ASAP7_75t_R FILLER_191_176 ();
 DECAPx10_ASAP7_75t_R FILLER_191_196 ();
 DECAPx6_ASAP7_75t_R FILLER_191_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_232 ();
 DECAPx2_ASAP7_75t_R FILLER_191_239 ();
 FILLER_ASAP7_75t_R FILLER_191_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_247 ();
 FILLER_ASAP7_75t_R FILLER_191_256 ();
 DECAPx2_ASAP7_75t_R FILLER_191_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_271 ();
 DECAPx4_ASAP7_75t_R FILLER_191_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_288 ();
 DECAPx1_ASAP7_75t_R FILLER_191_295 ();
 DECAPx1_ASAP7_75t_R FILLER_191_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_323 ();
 DECAPx2_ASAP7_75t_R FILLER_191_332 ();
 FILLER_ASAP7_75t_R FILLER_191_338 ();
 DECAPx2_ASAP7_75t_R FILLER_191_370 ();
 DECAPx2_ASAP7_75t_R FILLER_191_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_402 ();
 FILLER_ASAP7_75t_R FILLER_191_410 ();
 FILLER_ASAP7_75t_R FILLER_191_431 ();
 FILLER_ASAP7_75t_R FILLER_191_455 ();
 DECAPx2_ASAP7_75t_R FILLER_191_472 ();
 FILLER_ASAP7_75t_R FILLER_191_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_480 ();
 FILLER_ASAP7_75t_R FILLER_191_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_507 ();
 DECAPx4_ASAP7_75t_R FILLER_191_514 ();
 DECAPx6_ASAP7_75t_R FILLER_191_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_541 ();
 DECAPx1_ASAP7_75t_R FILLER_191_558 ();
 DECAPx6_ASAP7_75t_R FILLER_191_588 ();
 DECAPx2_ASAP7_75t_R FILLER_191_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_608 ();
 DECAPx10_ASAP7_75t_R FILLER_191_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_634 ();
 DECAPx4_ASAP7_75t_R FILLER_191_640 ();
 FILLER_ASAP7_75t_R FILLER_191_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_652 ();
 DECAPx1_ASAP7_75t_R FILLER_191_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_667 ();
 DECAPx4_ASAP7_75t_R FILLER_191_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_703 ();
 DECAPx6_ASAP7_75t_R FILLER_191_712 ();
 DECAPx2_ASAP7_75t_R FILLER_191_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_732 ();
 DECAPx4_ASAP7_75t_R FILLER_191_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_749 ();
 DECAPx6_ASAP7_75t_R FILLER_191_756 ();
 DECAPx2_ASAP7_75t_R FILLER_191_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_776 ();
 DECAPx10_ASAP7_75t_R FILLER_191_784 ();
 DECAPx10_ASAP7_75t_R FILLER_191_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_854 ();
 FILLER_ASAP7_75t_R FILLER_191_864 ();
 DECAPx6_ASAP7_75t_R FILLER_191_905 ();
 DECAPx1_ASAP7_75t_R FILLER_191_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_923 ();
 DECAPx6_ASAP7_75t_R FILLER_191_926 ();
 DECAPx10_ASAP7_75t_R FILLER_191_946 ();
 DECAPx4_ASAP7_75t_R FILLER_191_968 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1124 ();
 FILLER_ASAP7_75t_R FILLER_191_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1148 ();
 FILLER_ASAP7_75t_R FILLER_191_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1161 ();
 FILLER_ASAP7_75t_R FILLER_191_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1204 ();
 FILLER_ASAP7_75t_R FILLER_191_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1246 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1267 ();
 FILLER_ASAP7_75t_R FILLER_191_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1293 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1301 ();
 FILLER_ASAP7_75t_R FILLER_191_1311 ();
 FILLER_ASAP7_75t_R FILLER_191_1326 ();
 FILLER_ASAP7_75t_R FILLER_191_1380 ();
 DECAPx4_ASAP7_75t_R FILLER_191_1388 ();
 FILLER_ASAP7_75t_R FILLER_191_1398 ();
 DECAPx4_ASAP7_75t_R FILLER_192_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_12 ();
 DECAPx6_ASAP7_75t_R FILLER_192_46 ();
 FILLER_ASAP7_75t_R FILLER_192_60 ();
 FILLER_ASAP7_75t_R FILLER_192_69 ();
 DECAPx6_ASAP7_75t_R FILLER_192_97 ();
 FILLER_ASAP7_75t_R FILLER_192_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_113 ();
 DECAPx2_ASAP7_75t_R FILLER_192_117 ();
 FILLER_ASAP7_75t_R FILLER_192_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_129 ();
 FILLER_ASAP7_75t_R FILLER_192_156 ();
 DECAPx2_ASAP7_75t_R FILLER_192_186 ();
 FILLER_ASAP7_75t_R FILLER_192_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_208 ();
 DECAPx1_ASAP7_75t_R FILLER_192_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_219 ();
 DECAPx4_ASAP7_75t_R FILLER_192_226 ();
 FILLER_ASAP7_75t_R FILLER_192_236 ();
 DECAPx4_ASAP7_75t_R FILLER_192_258 ();
 FILLER_ASAP7_75t_R FILLER_192_268 ();
 DECAPx2_ASAP7_75t_R FILLER_192_276 ();
 FILLER_ASAP7_75t_R FILLER_192_282 ();
 DECAPx6_ASAP7_75t_R FILLER_192_310 ();
 DECAPx1_ASAP7_75t_R FILLER_192_324 ();
 FILLER_ASAP7_75t_R FILLER_192_336 ();
 DECAPx4_ASAP7_75t_R FILLER_192_348 ();
 DECAPx4_ASAP7_75t_R FILLER_192_364 ();
 FILLER_ASAP7_75t_R FILLER_192_374 ();
 DECAPx1_ASAP7_75t_R FILLER_192_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_386 ();
 DECAPx6_ASAP7_75t_R FILLER_192_393 ();
 DECAPx1_ASAP7_75t_R FILLER_192_407 ();
 DECAPx6_ASAP7_75t_R FILLER_192_433 ();
 DECAPx2_ASAP7_75t_R FILLER_192_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_464 ();
 DECAPx10_ASAP7_75t_R FILLER_192_479 ();
 FILLER_ASAP7_75t_R FILLER_192_501 ();
 DECAPx2_ASAP7_75t_R FILLER_192_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_542 ();
 DECAPx4_ASAP7_75t_R FILLER_192_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_559 ();
 DECAPx1_ASAP7_75t_R FILLER_192_573 ();
 FILLER_ASAP7_75t_R FILLER_192_580 ();
 DECAPx1_ASAP7_75t_R FILLER_192_612 ();
 DECAPx4_ASAP7_75t_R FILLER_192_619 ();
 FILLER_ASAP7_75t_R FILLER_192_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_648 ();
 DECAPx10_ASAP7_75t_R FILLER_192_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_691 ();
 DECAPx6_ASAP7_75t_R FILLER_192_697 ();
 FILLER_ASAP7_75t_R FILLER_192_711 ();
 DECAPx6_ASAP7_75t_R FILLER_192_719 ();
 FILLER_ASAP7_75t_R FILLER_192_733 ();
 DECAPx4_ASAP7_75t_R FILLER_192_741 ();
 FILLER_ASAP7_75t_R FILLER_192_751 ();
 DECAPx10_ASAP7_75t_R FILLER_192_762 ();
 DECAPx6_ASAP7_75t_R FILLER_192_784 ();
 DECAPx1_ASAP7_75t_R FILLER_192_806 ();
 DECAPx6_ASAP7_75t_R FILLER_192_817 ();
 DECAPx2_ASAP7_75t_R FILLER_192_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_846 ();
 DECAPx2_ASAP7_75t_R FILLER_192_873 ();
 DECAPx6_ASAP7_75t_R FILLER_192_919 ();
 FILLER_ASAP7_75t_R FILLER_192_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_935 ();
 FILLER_ASAP7_75t_R FILLER_192_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_941 ();
 DECAPx1_ASAP7_75t_R FILLER_192_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_954 ();
 DECAPx2_ASAP7_75t_R FILLER_192_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_975 ();
 DECAPx4_ASAP7_75t_R FILLER_192_985 ();
 FILLER_ASAP7_75t_R FILLER_192_995 ();
 FILLER_ASAP7_75t_R FILLER_192_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1012 ();
 FILLER_ASAP7_75t_R FILLER_192_1022 ();
 FILLER_ASAP7_75t_R FILLER_192_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1036 ();
 FILLER_ASAP7_75t_R FILLER_192_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1118 ();
 FILLER_ASAP7_75t_R FILLER_192_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_192_1173 ();
 FILLER_ASAP7_75t_R FILLER_192_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_192_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_192_1227 ();
 FILLER_ASAP7_75t_R FILLER_192_1233 ();
 FILLER_ASAP7_75t_R FILLER_192_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1253 ();
 FILLER_ASAP7_75t_R FILLER_192_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1269 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1280 ();
 FILLER_ASAP7_75t_R FILLER_192_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1354 ();
 FILLER_ASAP7_75t_R FILLER_192_1384 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1395 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1399 ();
 DECAPx6_ASAP7_75t_R FILLER_193_2 ();
 DECAPx1_ASAP7_75t_R FILLER_193_16 ();
 DECAPx1_ASAP7_75t_R FILLER_193_23 ();
 DECAPx1_ASAP7_75t_R FILLER_193_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_76 ();
 FILLER_ASAP7_75t_R FILLER_193_80 ();
 DECAPx6_ASAP7_75t_R FILLER_193_111 ();
 DECAPx1_ASAP7_75t_R FILLER_193_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_136 ();
 DECAPx6_ASAP7_75t_R FILLER_193_140 ();
 FILLER_ASAP7_75t_R FILLER_193_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_156 ();
 DECAPx1_ASAP7_75t_R FILLER_193_169 ();
 DECAPx2_ASAP7_75t_R FILLER_193_186 ();
 FILLER_ASAP7_75t_R FILLER_193_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_194 ();
 DECAPx6_ASAP7_75t_R FILLER_193_201 ();
 DECAPx1_ASAP7_75t_R FILLER_193_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_219 ();
 DECAPx4_ASAP7_75t_R FILLER_193_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_245 ();
 DECAPx2_ASAP7_75t_R FILLER_193_252 ();
 FILLER_ASAP7_75t_R FILLER_193_258 ();
 DECAPx10_ASAP7_75t_R FILLER_193_282 ();
 DECAPx4_ASAP7_75t_R FILLER_193_304 ();
 DECAPx6_ASAP7_75t_R FILLER_193_320 ();
 DECAPx4_ASAP7_75t_R FILLER_193_340 ();
 DECAPx1_ASAP7_75t_R FILLER_193_372 ();
 FILLER_ASAP7_75t_R FILLER_193_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_386 ();
 DECAPx1_ASAP7_75t_R FILLER_193_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_399 ();
 DECAPx6_ASAP7_75t_R FILLER_193_412 ();
 FILLER_ASAP7_75t_R FILLER_193_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_428 ();
 DECAPx10_ASAP7_75t_R FILLER_193_435 ();
 DECAPx1_ASAP7_75t_R FILLER_193_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_461 ();
 DECAPx10_ASAP7_75t_R FILLER_193_474 ();
 DECAPx10_ASAP7_75t_R FILLER_193_496 ();
 DECAPx2_ASAP7_75t_R FILLER_193_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_524 ();
 DECAPx4_ASAP7_75t_R FILLER_193_535 ();
 FILLER_ASAP7_75t_R FILLER_193_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_547 ();
 DECAPx6_ASAP7_75t_R FILLER_193_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_578 ();
 FILLER_ASAP7_75t_R FILLER_193_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_594 ();
 DECAPx1_ASAP7_75t_R FILLER_193_627 ();
 DECAPx10_ASAP7_75t_R FILLER_193_641 ();
 DECAPx2_ASAP7_75t_R FILLER_193_663 ();
 FILLER_ASAP7_75t_R FILLER_193_669 ();
 DECAPx1_ASAP7_75t_R FILLER_193_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_690 ();
 FILLER_ASAP7_75t_R FILLER_193_697 ();
 FILLER_ASAP7_75t_R FILLER_193_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_719 ();
 DECAPx2_ASAP7_75t_R FILLER_193_728 ();
 DECAPx10_ASAP7_75t_R FILLER_193_746 ();
 DECAPx10_ASAP7_75t_R FILLER_193_768 ();
 DECAPx1_ASAP7_75t_R FILLER_193_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_794 ();
 DECAPx2_ASAP7_75t_R FILLER_193_805 ();
 DECAPx10_ASAP7_75t_R FILLER_193_826 ();
 FILLER_ASAP7_75t_R FILLER_193_848 ();
 DECAPx2_ASAP7_75t_R FILLER_193_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_863 ();
 FILLER_ASAP7_75t_R FILLER_193_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_869 ();
 FILLER_ASAP7_75t_R FILLER_193_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_897 ();
 FILLER_ASAP7_75t_R FILLER_193_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_962 ();
 DECAPx2_ASAP7_75t_R FILLER_193_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_983 ();
 DECAPx1_ASAP7_75t_R FILLER_193_991 ();
 FILLER_ASAP7_75t_R FILLER_193_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1080 ();
 FILLER_ASAP7_75t_R FILLER_193_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1232 ();
 DECAPx4_ASAP7_75t_R FILLER_193_1246 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1308 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1330 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1344 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1354 ();
 FILLER_ASAP7_75t_R FILLER_193_1376 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1378 ();
 FILLER_ASAP7_75t_R FILLER_194_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_4 ();
 FILLER_ASAP7_75t_R FILLER_194_31 ();
 DECAPx1_ASAP7_75t_R FILLER_194_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_63 ();
 DECAPx6_ASAP7_75t_R FILLER_194_67 ();
 DECAPx2_ASAP7_75t_R FILLER_194_81 ();
 DECAPx1_ASAP7_75t_R FILLER_194_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_107 ();
 FILLER_ASAP7_75t_R FILLER_194_121 ();
 DECAPx2_ASAP7_75t_R FILLER_194_155 ();
 FILLER_ASAP7_75t_R FILLER_194_161 ();
 DECAPx4_ASAP7_75t_R FILLER_194_185 ();
 FILLER_ASAP7_75t_R FILLER_194_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_197 ();
 DECAPx1_ASAP7_75t_R FILLER_194_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_216 ();
 DECAPx2_ASAP7_75t_R FILLER_194_223 ();
 FILLER_ASAP7_75t_R FILLER_194_229 ();
 DECAPx2_ASAP7_75t_R FILLER_194_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_261 ();
 DECAPx2_ASAP7_75t_R FILLER_194_281 ();
 FILLER_ASAP7_75t_R FILLER_194_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_289 ();
 FILLER_ASAP7_75t_R FILLER_194_300 ();
 DECAPx4_ASAP7_75t_R FILLER_194_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_336 ();
 FILLER_ASAP7_75t_R FILLER_194_347 ();
 DECAPx6_ASAP7_75t_R FILLER_194_362 ();
 FILLER_ASAP7_75t_R FILLER_194_376 ();
 DECAPx2_ASAP7_75t_R FILLER_194_386 ();
 FILLER_ASAP7_75t_R FILLER_194_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_394 ();
 DECAPx6_ASAP7_75t_R FILLER_194_409 ();
 FILLER_ASAP7_75t_R FILLER_194_423 ();
 DECAPx1_ASAP7_75t_R FILLER_194_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_437 ();
 DECAPx1_ASAP7_75t_R FILLER_194_445 ();
 DECAPx1_ASAP7_75t_R FILLER_194_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_461 ();
 DECAPx6_ASAP7_75t_R FILLER_194_464 ();
 DECAPx1_ASAP7_75t_R FILLER_194_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_500 ();
 DECAPx2_ASAP7_75t_R FILLER_194_508 ();
 FILLER_ASAP7_75t_R FILLER_194_514 ();
 DECAPx10_ASAP7_75t_R FILLER_194_522 ();
 DECAPx10_ASAP7_75t_R FILLER_194_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_566 ();
 DECAPx6_ASAP7_75t_R FILLER_194_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_595 ();
 DECAPx1_ASAP7_75t_R FILLER_194_599 ();
 DECAPx6_ASAP7_75t_R FILLER_194_611 ();
 DECAPx2_ASAP7_75t_R FILLER_194_625 ();
 DECAPx4_ASAP7_75t_R FILLER_194_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_672 ();
 DECAPx1_ASAP7_75t_R FILLER_194_683 ();
 DECAPx2_ASAP7_75t_R FILLER_194_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_703 ();
 DECAPx2_ASAP7_75t_R FILLER_194_707 ();
 DECAPx2_ASAP7_75t_R FILLER_194_733 ();
 FILLER_ASAP7_75t_R FILLER_194_739 ();
 DECAPx10_ASAP7_75t_R FILLER_194_745 ();
 DECAPx10_ASAP7_75t_R FILLER_194_767 ();
 DECAPx6_ASAP7_75t_R FILLER_194_789 ();
 FILLER_ASAP7_75t_R FILLER_194_803 ();
 DECAPx1_ASAP7_75t_R FILLER_194_813 ();
 DECAPx1_ASAP7_75t_R FILLER_194_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_827 ();
 DECAPx1_ASAP7_75t_R FILLER_194_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_851 ();
 DECAPx10_ASAP7_75t_R FILLER_194_858 ();
 FILLER_ASAP7_75t_R FILLER_194_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_882 ();
 FILLER_ASAP7_75t_R FILLER_194_886 ();
 DECAPx1_ASAP7_75t_R FILLER_194_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_902 ();
 DECAPx6_ASAP7_75t_R FILLER_194_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_923 ();
 FILLER_ASAP7_75t_R FILLER_194_938 ();
 DECAPx2_ASAP7_75t_R FILLER_194_947 ();
 FILLER_ASAP7_75t_R FILLER_194_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_955 ();
 FILLER_ASAP7_75t_R FILLER_194_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_964 ();
 FILLER_ASAP7_75t_R FILLER_194_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_977 ();
 FILLER_ASAP7_75t_R FILLER_194_993 ();
 DECAPx6_ASAP7_75t_R FILLER_194_1003 ();
 FILLER_ASAP7_75t_R FILLER_194_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1032 ();
 FILLER_ASAP7_75t_R FILLER_194_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1154 ();
 FILLER_ASAP7_75t_R FILLER_194_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_194_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1209 ();
 FILLER_ASAP7_75t_R FILLER_194_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_194_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1312 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_194_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1375 ();
 FILLER_ASAP7_75t_R FILLER_194_1384 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_195_2 ();
 DECAPx6_ASAP7_75t_R FILLER_195_30 ();
 FILLER_ASAP7_75t_R FILLER_195_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_46 ();
 DECAPx1_ASAP7_75t_R FILLER_195_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_60 ();
 FILLER_ASAP7_75t_R FILLER_195_71 ();
 DECAPx10_ASAP7_75t_R FILLER_195_79 ();
 DECAPx6_ASAP7_75t_R FILLER_195_127 ();
 DECAPx4_ASAP7_75t_R FILLER_195_155 ();
 DECAPx10_ASAP7_75t_R FILLER_195_193 ();
 DECAPx2_ASAP7_75t_R FILLER_195_239 ();
 DECAPx10_ASAP7_75t_R FILLER_195_257 ();
 FILLER_ASAP7_75t_R FILLER_195_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_281 ();
 FILLER_ASAP7_75t_R FILLER_195_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_290 ();
 DECAPx1_ASAP7_75t_R FILLER_195_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_305 ();
 DECAPx4_ASAP7_75t_R FILLER_195_314 ();
 FILLER_ASAP7_75t_R FILLER_195_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_326 ();
 DECAPx4_ASAP7_75t_R FILLER_195_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_345 ();
 DECAPx1_ASAP7_75t_R FILLER_195_352 ();
 DECAPx6_ASAP7_75t_R FILLER_195_362 ();
 DECAPx10_ASAP7_75t_R FILLER_195_382 ();
 DECAPx4_ASAP7_75t_R FILLER_195_404 ();
 DECAPx1_ASAP7_75t_R FILLER_195_422 ();
 DECAPx6_ASAP7_75t_R FILLER_195_432 ();
 FILLER_ASAP7_75t_R FILLER_195_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_454 ();
 DECAPx4_ASAP7_75t_R FILLER_195_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_480 ();
 FILLER_ASAP7_75t_R FILLER_195_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_501 ();
 DECAPx1_ASAP7_75t_R FILLER_195_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_541 ();
 FILLER_ASAP7_75t_R FILLER_195_548 ();
 DECAPx2_ASAP7_75t_R FILLER_195_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_566 ();
 DECAPx10_ASAP7_75t_R FILLER_195_577 ();
 DECAPx6_ASAP7_75t_R FILLER_195_599 ();
 DECAPx1_ASAP7_75t_R FILLER_195_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_617 ();
 DECAPx6_ASAP7_75t_R FILLER_195_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_644 ();
 DECAPx4_ASAP7_75t_R FILLER_195_692 ();
 FILLER_ASAP7_75t_R FILLER_195_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_744 ();
 FILLER_ASAP7_75t_R FILLER_195_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_757 ();
 FILLER_ASAP7_75t_R FILLER_195_764 ();
 DECAPx4_ASAP7_75t_R FILLER_195_786 ();
 DECAPx10_ASAP7_75t_R FILLER_195_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_839 ();
 FILLER_ASAP7_75t_R FILLER_195_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_887 ();
 FILLER_ASAP7_75t_R FILLER_195_891 ();
 FILLER_ASAP7_75t_R FILLER_195_896 ();
 DECAPx4_ASAP7_75t_R FILLER_195_949 ();
 FILLER_ASAP7_75t_R FILLER_195_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_961 ();
 DECAPx1_ASAP7_75t_R FILLER_195_968 ();
 DECAPx6_ASAP7_75t_R FILLER_195_975 ();
 FILLER_ASAP7_75t_R FILLER_195_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_991 ();
 DECAPx10_ASAP7_75t_R FILLER_195_998 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1058 ();
 FILLER_ASAP7_75t_R FILLER_195_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1091 ();
 FILLER_ASAP7_75t_R FILLER_195_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1163 ();
 FILLER_ASAP7_75t_R FILLER_195_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1234 ();
 FILLER_ASAP7_75t_R FILLER_195_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1259 ();
 FILLER_ASAP7_75t_R FILLER_195_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1278 ();
 FILLER_ASAP7_75t_R FILLER_195_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1325 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1355 ();
 FILLER_ASAP7_75t_R FILLER_195_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1404 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_2 ();
 DECAPx4_ASAP7_75t_R FILLER_196_41 ();
 FILLER_ASAP7_75t_R FILLER_196_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_53 ();
 FILLER_ASAP7_75t_R FILLER_196_80 ();
 FILLER_ASAP7_75t_R FILLER_196_88 ();
 DECAPx6_ASAP7_75t_R FILLER_196_97 ();
 DECAPx1_ASAP7_75t_R FILLER_196_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_115 ();
 DECAPx6_ASAP7_75t_R FILLER_196_126 ();
 DECAPx4_ASAP7_75t_R FILLER_196_156 ();
 FILLER_ASAP7_75t_R FILLER_196_178 ();
 DECAPx6_ASAP7_75t_R FILLER_196_188 ();
 DECAPx2_ASAP7_75t_R FILLER_196_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_208 ();
 FILLER_ASAP7_75t_R FILLER_196_215 ();
 DECAPx1_ASAP7_75t_R FILLER_196_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_238 ();
 DECAPx6_ASAP7_75t_R FILLER_196_253 ();
 DECAPx2_ASAP7_75t_R FILLER_196_267 ();
 DECAPx2_ASAP7_75t_R FILLER_196_285 ();
 FILLER_ASAP7_75t_R FILLER_196_291 ();
 FILLER_ASAP7_75t_R FILLER_196_299 ();
 DECAPx2_ASAP7_75t_R FILLER_196_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_319 ();
 DECAPx10_ASAP7_75t_R FILLER_196_332 ();
 DECAPx2_ASAP7_75t_R FILLER_196_368 ();
 FILLER_ASAP7_75t_R FILLER_196_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_376 ();
 DECAPx4_ASAP7_75t_R FILLER_196_383 ();
 FILLER_ASAP7_75t_R FILLER_196_393 ();
 DECAPx2_ASAP7_75t_R FILLER_196_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_407 ();
 DECAPx10_ASAP7_75t_R FILLER_196_424 ();
 DECAPx6_ASAP7_75t_R FILLER_196_446 ();
 FILLER_ASAP7_75t_R FILLER_196_460 ();
 DECAPx2_ASAP7_75t_R FILLER_196_474 ();
 FILLER_ASAP7_75t_R FILLER_196_480 ();
 DECAPx6_ASAP7_75t_R FILLER_196_488 ();
 DECAPx2_ASAP7_75t_R FILLER_196_508 ();
 DECAPx4_ASAP7_75t_R FILLER_196_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_539 ();
 FILLER_ASAP7_75t_R FILLER_196_566 ();
 DECAPx4_ASAP7_75t_R FILLER_196_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_585 ();
 FILLER_ASAP7_75t_R FILLER_196_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_614 ();
 DECAPx10_ASAP7_75t_R FILLER_196_641 ();
 DECAPx2_ASAP7_75t_R FILLER_196_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_669 ();
 DECAPx10_ASAP7_75t_R FILLER_196_677 ();
 DECAPx6_ASAP7_75t_R FILLER_196_699 ();
 DECAPx2_ASAP7_75t_R FILLER_196_713 ();
 FILLER_ASAP7_75t_R FILLER_196_727 ();
 DECAPx10_ASAP7_75t_R FILLER_196_750 ();
 DECAPx10_ASAP7_75t_R FILLER_196_772 ();
 DECAPx2_ASAP7_75t_R FILLER_196_803 ();
 FILLER_ASAP7_75t_R FILLER_196_809 ();
 DECAPx6_ASAP7_75t_R FILLER_196_819 ();
 DECAPx2_ASAP7_75t_R FILLER_196_833 ();
 DECAPx2_ASAP7_75t_R FILLER_196_845 ();
 FILLER_ASAP7_75t_R FILLER_196_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_857 ();
 FILLER_ASAP7_75t_R FILLER_196_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_872 ();
 FILLER_ASAP7_75t_R FILLER_196_899 ();
 DECAPx2_ASAP7_75t_R FILLER_196_908 ();
 FILLER_ASAP7_75t_R FILLER_196_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_916 ();
 DECAPx6_ASAP7_75t_R FILLER_196_920 ();
 FILLER_ASAP7_75t_R FILLER_196_934 ();
 FILLER_ASAP7_75t_R FILLER_196_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_960 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1003 ();
 FILLER_ASAP7_75t_R FILLER_196_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1094 ();
 FILLER_ASAP7_75t_R FILLER_196_1121 ();
 FILLER_ASAP7_75t_R FILLER_196_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1147 ();
 FILLER_ASAP7_75t_R FILLER_196_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1156 ();
 FILLER_ASAP7_75t_R FILLER_196_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1199 ();
 FILLER_ASAP7_75t_R FILLER_196_1228 ();
 FILLER_ASAP7_75t_R FILLER_196_1240 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1270 ();
 FILLER_ASAP7_75t_R FILLER_196_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1321 ();
 FILLER_ASAP7_75t_R FILLER_196_1327 ();
 FILLER_ASAP7_75t_R FILLER_196_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1382 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1388 ();
 FILLER_ASAP7_75t_R FILLER_196_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1404 ();
 DECAPx1_ASAP7_75t_R FILLER_197_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_43 ();
 FILLER_ASAP7_75t_R FILLER_197_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_111 ();
 FILLER_ASAP7_75t_R FILLER_197_138 ();
 DECAPx10_ASAP7_75t_R FILLER_197_166 ();
 DECAPx1_ASAP7_75t_R FILLER_197_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_221 ();
 DECAPx6_ASAP7_75t_R FILLER_197_229 ();
 DECAPx1_ASAP7_75t_R FILLER_197_243 ();
 FILLER_ASAP7_75t_R FILLER_197_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_264 ();
 DECAPx10_ASAP7_75t_R FILLER_197_287 ();
 DECAPx10_ASAP7_75t_R FILLER_197_309 ();
 DECAPx1_ASAP7_75t_R FILLER_197_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_350 ();
 DECAPx2_ASAP7_75t_R FILLER_197_359 ();
 FILLER_ASAP7_75t_R FILLER_197_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_367 ();
 DECAPx1_ASAP7_75t_R FILLER_197_384 ();
 DECAPx10_ASAP7_75t_R FILLER_197_410 ();
 DECAPx4_ASAP7_75t_R FILLER_197_450 ();
 FILLER_ASAP7_75t_R FILLER_197_460 ();
 DECAPx1_ASAP7_75t_R FILLER_197_470 ();
 DECAPx10_ASAP7_75t_R FILLER_197_486 ();
 DECAPx6_ASAP7_75t_R FILLER_197_508 ();
 DECAPx2_ASAP7_75t_R FILLER_197_522 ();
 FILLER_ASAP7_75t_R FILLER_197_548 ();
 FILLER_ASAP7_75t_R FILLER_197_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_562 ();
 DECAPx1_ASAP7_75t_R FILLER_197_595 ();
 FILLER_ASAP7_75t_R FILLER_197_625 ();
 DECAPx6_ASAP7_75t_R FILLER_197_658 ();
 FILLER_ASAP7_75t_R FILLER_197_672 ();
 FILLER_ASAP7_75t_R FILLER_197_681 ();
 FILLER_ASAP7_75t_R FILLER_197_701 ();
 FILLER_ASAP7_75t_R FILLER_197_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_719 ();
 DECAPx4_ASAP7_75t_R FILLER_197_726 ();
 FILLER_ASAP7_75t_R FILLER_197_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_738 ();
 DECAPx6_ASAP7_75t_R FILLER_197_747 ();
 FILLER_ASAP7_75t_R FILLER_197_761 ();
 DECAPx2_ASAP7_75t_R FILLER_197_767 ();
 FILLER_ASAP7_75t_R FILLER_197_773 ();
 DECAPx2_ASAP7_75t_R FILLER_197_785 ();
 FILLER_ASAP7_75t_R FILLER_197_791 ();
 DECAPx2_ASAP7_75t_R FILLER_197_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_819 ();
 DECAPx4_ASAP7_75t_R FILLER_197_833 ();
 DECAPx10_ASAP7_75t_R FILLER_197_855 ();
 DECAPx6_ASAP7_75t_R FILLER_197_877 ();
 DECAPx2_ASAP7_75t_R FILLER_197_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_897 ();
 DECAPx6_ASAP7_75t_R FILLER_197_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_940 ();
 DECAPx1_ASAP7_75t_R FILLER_197_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_957 ();
 DECAPx2_ASAP7_75t_R FILLER_197_967 ();
 FILLER_ASAP7_75t_R FILLER_197_973 ();
 DECAPx2_ASAP7_75t_R FILLER_197_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1008 ();
 FILLER_ASAP7_75t_R FILLER_197_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1109 ();
 FILLER_ASAP7_75t_R FILLER_197_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1166 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1185 ();
 FILLER_ASAP7_75t_R FILLER_197_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1210 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1241 ();
 FILLER_ASAP7_75t_R FILLER_197_1251 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1272 ();
 FILLER_ASAP7_75t_R FILLER_197_1282 ();
 FILLER_ASAP7_75t_R FILLER_197_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1292 ();
 FILLER_ASAP7_75t_R FILLER_197_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1324 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1335 ();
 FILLER_ASAP7_75t_R FILLER_197_1341 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1369 ();
 DECAPx6_ASAP7_75t_R FILLER_198_2 ();
 FILLER_ASAP7_75t_R FILLER_198_16 ();
 DECAPx1_ASAP7_75t_R FILLER_198_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_28 ();
 DECAPx1_ASAP7_75t_R FILLER_198_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_39 ();
 DECAPx4_ASAP7_75t_R FILLER_198_66 ();
 DECAPx2_ASAP7_75t_R FILLER_198_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_95 ();
 DECAPx4_ASAP7_75t_R FILLER_198_105 ();
 FILLER_ASAP7_75t_R FILLER_198_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_117 ();
 FILLER_ASAP7_75t_R FILLER_198_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_126 ();
 DECAPx2_ASAP7_75t_R FILLER_198_130 ();
 FILLER_ASAP7_75t_R FILLER_198_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_138 ();
 DECAPx2_ASAP7_75t_R FILLER_198_146 ();
 FILLER_ASAP7_75t_R FILLER_198_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_154 ();
 DECAPx6_ASAP7_75t_R FILLER_198_158 ();
 FILLER_ASAP7_75t_R FILLER_198_172 ();
 DECAPx10_ASAP7_75t_R FILLER_198_188 ();
 DECAPx10_ASAP7_75t_R FILLER_198_210 ();
 DECAPx10_ASAP7_75t_R FILLER_198_232 ();
 FILLER_ASAP7_75t_R FILLER_198_254 ();
 FILLER_ASAP7_75t_R FILLER_198_270 ();
 DECAPx10_ASAP7_75t_R FILLER_198_278 ();
 DECAPx2_ASAP7_75t_R FILLER_198_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_306 ();
 DECAPx4_ASAP7_75t_R FILLER_198_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_325 ();
 DECAPx4_ASAP7_75t_R FILLER_198_343 ();
 DECAPx2_ASAP7_75t_R FILLER_198_386 ();
 DECAPx6_ASAP7_75t_R FILLER_198_398 ();
 DECAPx1_ASAP7_75t_R FILLER_198_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_416 ();
 DECAPx1_ASAP7_75t_R FILLER_198_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_479 ();
 FILLER_ASAP7_75t_R FILLER_198_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_517 ();
 FILLER_ASAP7_75t_R FILLER_198_524 ();
 DECAPx6_ASAP7_75t_R FILLER_198_532 ();
 DECAPx1_ASAP7_75t_R FILLER_198_546 ();
 DECAPx2_ASAP7_75t_R FILLER_198_576 ();
 FILLER_ASAP7_75t_R FILLER_198_582 ();
 DECAPx1_ASAP7_75t_R FILLER_198_587 ();
 FILLER_ASAP7_75t_R FILLER_198_606 ();
 DECAPx1_ASAP7_75t_R FILLER_198_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_630 ();
 DECAPx6_ASAP7_75t_R FILLER_198_637 ();
 DECAPx1_ASAP7_75t_R FILLER_198_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_655 ();
 DECAPx2_ASAP7_75t_R FILLER_198_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_668 ();
 DECAPx1_ASAP7_75t_R FILLER_198_679 ();
 DECAPx4_ASAP7_75t_R FILLER_198_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_714 ();
 DECAPx1_ASAP7_75t_R FILLER_198_758 ();
 DECAPx10_ASAP7_75t_R FILLER_198_768 ();
 DECAPx4_ASAP7_75t_R FILLER_198_790 ();
 FILLER_ASAP7_75t_R FILLER_198_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_805 ();
 DECAPx10_ASAP7_75t_R FILLER_198_832 ();
 FILLER_ASAP7_75t_R FILLER_198_854 ();
 DECAPx1_ASAP7_75t_R FILLER_198_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_899 ();
 DECAPx4_ASAP7_75t_R FILLER_198_906 ();
 DECAPx10_ASAP7_75t_R FILLER_198_919 ();
 DECAPx2_ASAP7_75t_R FILLER_198_941 ();
 DECAPx6_ASAP7_75t_R FILLER_198_977 ();
 DECAPx1_ASAP7_75t_R FILLER_198_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_995 ();
 FILLER_ASAP7_75t_R FILLER_198_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1004 ();
 FILLER_ASAP7_75t_R FILLER_198_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1013 ();
 FILLER_ASAP7_75t_R FILLER_198_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1034 ();
 FILLER_ASAP7_75t_R FILLER_198_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1045 ();
 FILLER_ASAP7_75t_R FILLER_198_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1071 ();
 FILLER_ASAP7_75t_R FILLER_198_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1113 ();
 FILLER_ASAP7_75t_R FILLER_198_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1181 ();
 FILLER_ASAP7_75t_R FILLER_198_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1201 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1223 ();
 FILLER_ASAP7_75t_R FILLER_198_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1269 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1307 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1316 ();
 FILLER_ASAP7_75t_R FILLER_198_1326 ();
 FILLER_ASAP7_75t_R FILLER_198_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1360 ();
 FILLER_ASAP7_75t_R FILLER_198_1388 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1393 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_199_2 ();
 DECAPx2_ASAP7_75t_R FILLER_199_24 ();
 FILLER_ASAP7_75t_R FILLER_199_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_32 ();
 DECAPx4_ASAP7_75t_R FILLER_199_42 ();
 FILLER_ASAP7_75t_R FILLER_199_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_54 ();
 DECAPx10_ASAP7_75t_R FILLER_199_58 ();
 DECAPx10_ASAP7_75t_R FILLER_199_80 ();
 DECAPx2_ASAP7_75t_R FILLER_199_102 ();
 DECAPx4_ASAP7_75t_R FILLER_199_123 ();
 FILLER_ASAP7_75t_R FILLER_199_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_135 ();
 FILLER_ASAP7_75t_R FILLER_199_162 ();
 FILLER_ASAP7_75t_R FILLER_199_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_182 ();
 DECAPx1_ASAP7_75t_R FILLER_199_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_195 ();
 DECAPx6_ASAP7_75t_R FILLER_199_210 ();
 DECAPx2_ASAP7_75t_R FILLER_199_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_230 ();
 DECAPx6_ASAP7_75t_R FILLER_199_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_255 ();
 DECAPx1_ASAP7_75t_R FILLER_199_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_274 ();
 DECAPx1_ASAP7_75t_R FILLER_199_289 ();
 DECAPx4_ASAP7_75t_R FILLER_199_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_329 ();
 DECAPx6_ASAP7_75t_R FILLER_199_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_352 ();
 DECAPx2_ASAP7_75t_R FILLER_199_365 ();
 FILLER_ASAP7_75t_R FILLER_199_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_373 ();
 DECAPx4_ASAP7_75t_R FILLER_199_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_390 ();
 DECAPx6_ASAP7_75t_R FILLER_199_411 ();
 DECAPx1_ASAP7_75t_R FILLER_199_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_429 ();
 DECAPx2_ASAP7_75t_R FILLER_199_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_454 ();
 DECAPx2_ASAP7_75t_R FILLER_199_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_472 ();
 DECAPx2_ASAP7_75t_R FILLER_199_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_491 ();
 FILLER_ASAP7_75t_R FILLER_199_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_534 ();
 DECAPx2_ASAP7_75t_R FILLER_199_545 ();
 DECAPx2_ASAP7_75t_R FILLER_199_557 ();
 FILLER_ASAP7_75t_R FILLER_199_563 ();
 DECAPx10_ASAP7_75t_R FILLER_199_568 ();
 DECAPx10_ASAP7_75t_R FILLER_199_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_612 ();
 DECAPx4_ASAP7_75t_R FILLER_199_620 ();
 DECAPx1_ASAP7_75t_R FILLER_199_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_641 ();
 FILLER_ASAP7_75t_R FILLER_199_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_682 ();
 DECAPx4_ASAP7_75t_R FILLER_199_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_705 ();
 DECAPx10_ASAP7_75t_R FILLER_199_710 ();
 DECAPx10_ASAP7_75t_R FILLER_199_732 ();
 DECAPx6_ASAP7_75t_R FILLER_199_754 ();
 DECAPx1_ASAP7_75t_R FILLER_199_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_772 ();
 FILLER_ASAP7_75t_R FILLER_199_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_797 ();
 DECAPx4_ASAP7_75t_R FILLER_199_808 ();
 FILLER_ASAP7_75t_R FILLER_199_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_820 ();
 DECAPx1_ASAP7_75t_R FILLER_199_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_828 ();
 FILLER_ASAP7_75t_R FILLER_199_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_837 ();
 DECAPx2_ASAP7_75t_R FILLER_199_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_853 ();
 DECAPx2_ASAP7_75t_R FILLER_199_858 ();
 FILLER_ASAP7_75t_R FILLER_199_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_866 ();
 FILLER_ASAP7_75t_R FILLER_199_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_875 ();
 DECAPx2_ASAP7_75t_R FILLER_199_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_920 ();
 DECAPx2_ASAP7_75t_R FILLER_199_926 ();
 DECAPx2_ASAP7_75t_R FILLER_199_937 ();
 DECAPx4_ASAP7_75t_R FILLER_199_952 ();
 FILLER_ASAP7_75t_R FILLER_199_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_964 ();
 DECAPx6_ASAP7_75t_R FILLER_199_971 ();
 DECAPx1_ASAP7_75t_R FILLER_199_990 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1117 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1166 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1173 ();
 FILLER_ASAP7_75t_R FILLER_199_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1268 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1282 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1286 ();
 FILLER_ASAP7_75t_R FILLER_199_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1308 ();
 FILLER_ASAP7_75t_R FILLER_199_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1328 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1335 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1361 ();
 FILLER_ASAP7_75t_R FILLER_199_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1401 ();
 DECAPx4_ASAP7_75t_R FILLER_200_2 ();
 FILLER_ASAP7_75t_R FILLER_200_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_54 ();
 DECAPx4_ASAP7_75t_R FILLER_200_81 ();
 FILLER_ASAP7_75t_R FILLER_200_91 ();
 DECAPx1_ASAP7_75t_R FILLER_200_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_103 ();
 FILLER_ASAP7_75t_R FILLER_200_130 ();
 DECAPx2_ASAP7_75t_R FILLER_200_135 ();
 DECAPx1_ASAP7_75t_R FILLER_200_147 ();
 DECAPx1_ASAP7_75t_R FILLER_200_154 ();
 DECAPx2_ASAP7_75t_R FILLER_200_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_188 ();
 FILLER_ASAP7_75t_R FILLER_200_217 ();
 DECAPx2_ASAP7_75t_R FILLER_200_225 ();
 DECAPx2_ASAP7_75t_R FILLER_200_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_245 ();
 DECAPx10_ASAP7_75t_R FILLER_200_256 ();
 FILLER_ASAP7_75t_R FILLER_200_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_291 ();
 DECAPx1_ASAP7_75t_R FILLER_200_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_302 ();
 DECAPx10_ASAP7_75t_R FILLER_200_315 ();
 DECAPx10_ASAP7_75t_R FILLER_200_337 ();
 DECAPx6_ASAP7_75t_R FILLER_200_359 ();
 DECAPx2_ASAP7_75t_R FILLER_200_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_379 ();
 DECAPx2_ASAP7_75t_R FILLER_200_386 ();
 FILLER_ASAP7_75t_R FILLER_200_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_394 ();
 DECAPx1_ASAP7_75t_R FILLER_200_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_407 ();
 DECAPx10_ASAP7_75t_R FILLER_200_415 ();
 DECAPx10_ASAP7_75t_R FILLER_200_437 ();
 FILLER_ASAP7_75t_R FILLER_200_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_461 ();
 DECAPx10_ASAP7_75t_R FILLER_200_472 ();
 DECAPx1_ASAP7_75t_R FILLER_200_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_498 ();
 DECAPx2_ASAP7_75t_R FILLER_200_506 ();
 FILLER_ASAP7_75t_R FILLER_200_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_514 ();
 FILLER_ASAP7_75t_R FILLER_200_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_553 ();
 DECAPx4_ASAP7_75t_R FILLER_200_561 ();
 FILLER_ASAP7_75t_R FILLER_200_571 ();
 DECAPx4_ASAP7_75t_R FILLER_200_586 ();
 DECAPx10_ASAP7_75t_R FILLER_200_599 ();
 DECAPx2_ASAP7_75t_R FILLER_200_621 ();
 FILLER_ASAP7_75t_R FILLER_200_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_650 ();
 FILLER_ASAP7_75t_R FILLER_200_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_659 ();
 DECAPx6_ASAP7_75t_R FILLER_200_666 ();
 DECAPx2_ASAP7_75t_R FILLER_200_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_686 ();
 DECAPx1_ASAP7_75t_R FILLER_200_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_712 ();
 DECAPx4_ASAP7_75t_R FILLER_200_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_729 ();
 FILLER_ASAP7_75t_R FILLER_200_740 ();
 DECAPx4_ASAP7_75t_R FILLER_200_748 ();
 FILLER_ASAP7_75t_R FILLER_200_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_771 ();
 DECAPx1_ASAP7_75t_R FILLER_200_784 ();
 DECAPx6_ASAP7_75t_R FILLER_200_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_828 ();
 DECAPx10_ASAP7_75t_R FILLER_200_857 ();
 DECAPx1_ASAP7_75t_R FILLER_200_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_883 ();
 FILLER_ASAP7_75t_R FILLER_200_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_898 ();
 DECAPx6_ASAP7_75t_R FILLER_200_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_995 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1056 ();
 FILLER_ASAP7_75t_R FILLER_200_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1132 ();
 FILLER_ASAP7_75t_R FILLER_200_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1189 ();
 FILLER_ASAP7_75t_R FILLER_200_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1240 ();
 FILLER_ASAP7_75t_R FILLER_200_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1317 ();
 FILLER_ASAP7_75t_R FILLER_200_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1332 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1354 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1368 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1372 ();
 FILLER_ASAP7_75t_R FILLER_200_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1385 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1388 ();
 FILLER_ASAP7_75t_R FILLER_200_1398 ();
 DECAPx10_ASAP7_75t_R FILLER_201_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_24 ();
 DECAPx4_ASAP7_75t_R FILLER_201_109 ();
 DECAPx1_ASAP7_75t_R FILLER_201_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_126 ();
 DECAPx10_ASAP7_75t_R FILLER_201_133 ();
 DECAPx6_ASAP7_75t_R FILLER_201_155 ();
 DECAPx2_ASAP7_75t_R FILLER_201_169 ();
 DECAPx10_ASAP7_75t_R FILLER_201_181 ();
 DECAPx1_ASAP7_75t_R FILLER_201_203 ();
 FILLER_ASAP7_75t_R FILLER_201_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_215 ();
 FILLER_ASAP7_75t_R FILLER_201_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_233 ();
 FILLER_ASAP7_75t_R FILLER_201_250 ();
 DECAPx1_ASAP7_75t_R FILLER_201_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_264 ();
 DECAPx10_ASAP7_75t_R FILLER_201_271 ();
 DECAPx6_ASAP7_75t_R FILLER_201_293 ();
 DECAPx2_ASAP7_75t_R FILLER_201_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_313 ();
 DECAPx10_ASAP7_75t_R FILLER_201_320 ();
 DECAPx6_ASAP7_75t_R FILLER_201_342 ();
 DECAPx2_ASAP7_75t_R FILLER_201_356 ();
 DECAPx4_ASAP7_75t_R FILLER_201_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_379 ();
 DECAPx1_ASAP7_75t_R FILLER_201_388 ();
 FILLER_ASAP7_75t_R FILLER_201_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_408 ();
 DECAPx4_ASAP7_75t_R FILLER_201_426 ();
 FILLER_ASAP7_75t_R FILLER_201_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_438 ();
 DECAPx4_ASAP7_75t_R FILLER_201_445 ();
 FILLER_ASAP7_75t_R FILLER_201_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_457 ();
 DECAPx1_ASAP7_75t_R FILLER_201_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_468 ();
 FILLER_ASAP7_75t_R FILLER_201_483 ();
 DECAPx6_ASAP7_75t_R FILLER_201_491 ();
 DECAPx1_ASAP7_75t_R FILLER_201_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_509 ();
 FILLER_ASAP7_75t_R FILLER_201_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_522 ();
 DECAPx1_ASAP7_75t_R FILLER_201_549 ();
 FILLER_ASAP7_75t_R FILLER_201_579 ();
 DECAPx6_ASAP7_75t_R FILLER_201_607 ();
 FILLER_ASAP7_75t_R FILLER_201_621 ();
 DECAPx6_ASAP7_75t_R FILLER_201_631 ();
 DECAPx2_ASAP7_75t_R FILLER_201_645 ();
 DECAPx4_ASAP7_75t_R FILLER_201_665 ();
 DECAPx4_ASAP7_75t_R FILLER_201_681 ();
 FILLER_ASAP7_75t_R FILLER_201_703 ();
 FILLER_ASAP7_75t_R FILLER_201_717 ();
 DECAPx2_ASAP7_75t_R FILLER_201_725 ();
 FILLER_ASAP7_75t_R FILLER_201_731 ();
 FILLER_ASAP7_75t_R FILLER_201_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_743 ();
 DECAPx2_ASAP7_75t_R FILLER_201_770 ();
 FILLER_ASAP7_75t_R FILLER_201_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_778 ();
 DECAPx4_ASAP7_75t_R FILLER_201_792 ();
 DECAPx2_ASAP7_75t_R FILLER_201_805 ();
 FILLER_ASAP7_75t_R FILLER_201_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_813 ();
 DECAPx2_ASAP7_75t_R FILLER_201_817 ();
 DECAPx6_ASAP7_75t_R FILLER_201_833 ();
 DECAPx6_ASAP7_75t_R FILLER_201_871 ();
 DECAPx1_ASAP7_75t_R FILLER_201_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_889 ();
 DECAPx2_ASAP7_75t_R FILLER_201_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_902 ();
 DECAPx2_ASAP7_75t_R FILLER_201_915 ();
 FILLER_ASAP7_75t_R FILLER_201_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_923 ();
 DECAPx6_ASAP7_75t_R FILLER_201_926 ();
 DECAPx2_ASAP7_75t_R FILLER_201_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_946 ();
 DECAPx1_ASAP7_75t_R FILLER_201_954 ();
 DECAPx1_ASAP7_75t_R FILLER_201_980 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1020 ();
 FILLER_ASAP7_75t_R FILLER_201_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1247 ();
 FILLER_ASAP7_75t_R FILLER_201_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1268 ();
 FILLER_ASAP7_75t_R FILLER_201_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1284 ();
 FILLER_ASAP7_75t_R FILLER_201_1290 ();
 FILLER_ASAP7_75t_R FILLER_201_1344 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1378 ();
 DECAPx6_ASAP7_75t_R FILLER_202_2 ();
 DECAPx1_ASAP7_75t_R FILLER_202_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_20 ();
 FILLER_ASAP7_75t_R FILLER_202_27 ();
 DECAPx6_ASAP7_75t_R FILLER_202_32 ();
 FILLER_ASAP7_75t_R FILLER_202_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_48 ();
 DECAPx1_ASAP7_75t_R FILLER_202_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_56 ();
 FILLER_ASAP7_75t_R FILLER_202_63 ();
 FILLER_ASAP7_75t_R FILLER_202_86 ();
 DECAPx1_ASAP7_75t_R FILLER_202_94 ();
 DECAPx4_ASAP7_75t_R FILLER_202_101 ();
 FILLER_ASAP7_75t_R FILLER_202_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_119 ();
 FILLER_ASAP7_75t_R FILLER_202_123 ();
 DECAPx1_ASAP7_75t_R FILLER_202_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_170 ();
 DECAPx2_ASAP7_75t_R FILLER_202_187 ();
 FILLER_ASAP7_75t_R FILLER_202_193 ();
 DECAPx10_ASAP7_75t_R FILLER_202_209 ();
 FILLER_ASAP7_75t_R FILLER_202_231 ();
 DECAPx2_ASAP7_75t_R FILLER_202_239 ();
 FILLER_ASAP7_75t_R FILLER_202_245 ();
 DECAPx2_ASAP7_75t_R FILLER_202_267 ();
 FILLER_ASAP7_75t_R FILLER_202_273 ();
 DECAPx10_ASAP7_75t_R FILLER_202_301 ();
 DECAPx2_ASAP7_75t_R FILLER_202_331 ();
 DECAPx10_ASAP7_75t_R FILLER_202_392 ();
 FILLER_ASAP7_75t_R FILLER_202_414 ();
 DECAPx2_ASAP7_75t_R FILLER_202_422 ();
 FILLER_ASAP7_75t_R FILLER_202_428 ();
 DECAPx4_ASAP7_75t_R FILLER_202_450 ();
 FILLER_ASAP7_75t_R FILLER_202_460 ();
 DECAPx4_ASAP7_75t_R FILLER_202_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_474 ();
 DECAPx10_ASAP7_75t_R FILLER_202_498 ();
 DECAPx1_ASAP7_75t_R FILLER_202_520 ();
 FILLER_ASAP7_75t_R FILLER_202_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_538 ();
 DECAPx1_ASAP7_75t_R FILLER_202_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_555 ();
 DECAPx2_ASAP7_75t_R FILLER_202_562 ();
 DECAPx1_ASAP7_75t_R FILLER_202_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_575 ();
 DECAPx1_ASAP7_75t_R FILLER_202_583 ();
 DECAPx2_ASAP7_75t_R FILLER_202_613 ();
 FILLER_ASAP7_75t_R FILLER_202_619 ();
 DECAPx6_ASAP7_75t_R FILLER_202_635 ();
 DECAPx1_ASAP7_75t_R FILLER_202_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_653 ();
 FILLER_ASAP7_75t_R FILLER_202_665 ();
 FILLER_ASAP7_75t_R FILLER_202_673 ();
 DECAPx2_ASAP7_75t_R FILLER_202_690 ();
 FILLER_ASAP7_75t_R FILLER_202_704 ();
 FILLER_ASAP7_75t_R FILLER_202_740 ();
 DECAPx4_ASAP7_75t_R FILLER_202_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_762 ();
 DECAPx4_ASAP7_75t_R FILLER_202_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_799 ();
 FILLER_ASAP7_75t_R FILLER_202_810 ();
 DECAPx6_ASAP7_75t_R FILLER_202_838 ();
 FILLER_ASAP7_75t_R FILLER_202_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_866 ();
 DECAPx2_ASAP7_75t_R FILLER_202_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_893 ();
 DECAPx1_ASAP7_75t_R FILLER_202_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_914 ();
 DECAPx1_ASAP7_75t_R FILLER_202_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_945 ();
 DECAPx4_ASAP7_75t_R FILLER_202_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_962 ();
 DECAPx10_ASAP7_75t_R FILLER_202_969 ();
 DECAPx4_ASAP7_75t_R FILLER_202_991 ();
 FILLER_ASAP7_75t_R FILLER_202_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1029 ();
 FILLER_ASAP7_75t_R FILLER_202_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1077 ();
 FILLER_ASAP7_75t_R FILLER_202_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1116 ();
 FILLER_ASAP7_75t_R FILLER_202_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1135 ();
 FILLER_ASAP7_75t_R FILLER_202_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1155 ();
 FILLER_ASAP7_75t_R FILLER_202_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1177 ();
 FILLER_ASAP7_75t_R FILLER_202_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1209 ();
 FILLER_ASAP7_75t_R FILLER_202_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1309 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1323 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1330 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1344 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1395 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1399 ();
 FILLER_ASAP7_75t_R FILLER_203_2 ();
 DECAPx4_ASAP7_75t_R FILLER_203_36 ();
 FILLER_ASAP7_75t_R FILLER_203_46 ();
 DECAPx4_ASAP7_75t_R FILLER_203_57 ();
 FILLER_ASAP7_75t_R FILLER_203_67 ();
 DECAPx10_ASAP7_75t_R FILLER_203_72 ();
 FILLER_ASAP7_75t_R FILLER_203_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_96 ();
 FILLER_ASAP7_75t_R FILLER_203_103 ();
 DECAPx1_ASAP7_75t_R FILLER_203_137 ();
 DECAPx10_ASAP7_75t_R FILLER_203_177 ();
 DECAPx4_ASAP7_75t_R FILLER_203_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_209 ();
 DECAPx10_ASAP7_75t_R FILLER_203_226 ();
 DECAPx1_ASAP7_75t_R FILLER_203_248 ();
 DECAPx4_ASAP7_75t_R FILLER_203_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_273 ();
 DECAPx4_ASAP7_75t_R FILLER_203_280 ();
 FILLER_ASAP7_75t_R FILLER_203_290 ();
 DECAPx10_ASAP7_75t_R FILLER_203_308 ();
 DECAPx10_ASAP7_75t_R FILLER_203_330 ();
 DECAPx2_ASAP7_75t_R FILLER_203_352 ();
 FILLER_ASAP7_75t_R FILLER_203_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_375 ();
 DECAPx6_ASAP7_75t_R FILLER_203_382 ();
 DECAPx2_ASAP7_75t_R FILLER_203_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_402 ();
 DECAPx10_ASAP7_75t_R FILLER_203_410 ();
 DECAPx10_ASAP7_75t_R FILLER_203_432 ();
 DECAPx2_ASAP7_75t_R FILLER_203_454 ();
 DECAPx2_ASAP7_75t_R FILLER_203_475 ();
 FILLER_ASAP7_75t_R FILLER_203_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_483 ();
 DECAPx2_ASAP7_75t_R FILLER_203_490 ();
 FILLER_ASAP7_75t_R FILLER_203_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_498 ();
 DECAPx4_ASAP7_75t_R FILLER_203_535 ();
 FILLER_ASAP7_75t_R FILLER_203_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_547 ();
 DECAPx6_ASAP7_75t_R FILLER_203_560 ();
 FILLER_ASAP7_75t_R FILLER_203_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_576 ();
 DECAPx6_ASAP7_75t_R FILLER_203_583 ();
 DECAPx1_ASAP7_75t_R FILLER_203_597 ();
 DECAPx4_ASAP7_75t_R FILLER_203_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_625 ();
 FILLER_ASAP7_75t_R FILLER_203_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_644 ();
 DECAPx4_ASAP7_75t_R FILLER_203_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_675 ();
 DECAPx1_ASAP7_75t_R FILLER_203_682 ();
 DECAPx2_ASAP7_75t_R FILLER_203_696 ();
 DECAPx1_ASAP7_75t_R FILLER_203_708 ();
 DECAPx6_ASAP7_75t_R FILLER_203_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_740 ();
 DECAPx6_ASAP7_75t_R FILLER_203_759 ();
 DECAPx1_ASAP7_75t_R FILLER_203_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_777 ();
 FILLER_ASAP7_75t_R FILLER_203_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_783 ();
 DECAPx4_ASAP7_75t_R FILLER_203_787 ();
 FILLER_ASAP7_75t_R FILLER_203_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_799 ();
 DECAPx2_ASAP7_75t_R FILLER_203_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_816 ();
 DECAPx1_ASAP7_75t_R FILLER_203_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_837 ();
 DECAPx10_ASAP7_75t_R FILLER_203_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_872 ();
 DECAPx4_ASAP7_75t_R FILLER_203_885 ();
 FILLER_ASAP7_75t_R FILLER_203_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_897 ();
 DECAPx4_ASAP7_75t_R FILLER_203_926 ();
 FILLER_ASAP7_75t_R FILLER_203_944 ();
 DECAPx2_ASAP7_75t_R FILLER_203_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_986 ();
 DECAPx6_ASAP7_75t_R FILLER_203_993 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1029 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1040 ();
 FILLER_ASAP7_75t_R FILLER_203_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1088 ();
 FILLER_ASAP7_75t_R FILLER_203_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1116 ();
 FILLER_ASAP7_75t_R FILLER_203_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1137 ();
 FILLER_ASAP7_75t_R FILLER_203_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1233 ();
 FILLER_ASAP7_75t_R FILLER_203_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1252 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1290 ();
 FILLER_ASAP7_75t_R FILLER_203_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1317 ();
 FILLER_ASAP7_75t_R FILLER_203_1323 ();
 FILLER_ASAP7_75t_R FILLER_203_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1330 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1354 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1388 ();
 DECAPx6_ASAP7_75t_R FILLER_204_2 ();
 FILLER_ASAP7_75t_R FILLER_204_16 ();
 DECAPx1_ASAP7_75t_R FILLER_204_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_25 ();
 DECAPx2_ASAP7_75t_R FILLER_204_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_38 ();
 FILLER_ASAP7_75t_R FILLER_204_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_73 ();
 DECAPx1_ASAP7_75t_R FILLER_204_77 ();
 FILLER_ASAP7_75t_R FILLER_204_87 ();
 DECAPx4_ASAP7_75t_R FILLER_204_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_125 ();
 DECAPx2_ASAP7_75t_R FILLER_204_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_138 ();
 FILLER_ASAP7_75t_R FILLER_204_154 ();
 FILLER_ASAP7_75t_R FILLER_204_159 ();
 FILLER_ASAP7_75t_R FILLER_204_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_201 ();
 FILLER_ASAP7_75t_R FILLER_204_208 ();
 DECAPx1_ASAP7_75t_R FILLER_204_244 ();
 DECAPx1_ASAP7_75t_R FILLER_204_258 ();
 FILLER_ASAP7_75t_R FILLER_204_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_295 ();
 DECAPx1_ASAP7_75t_R FILLER_204_310 ();
 DECAPx4_ASAP7_75t_R FILLER_204_320 ();
 DECAPx6_ASAP7_75t_R FILLER_204_337 ();
 DECAPx2_ASAP7_75t_R FILLER_204_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_357 ();
 DECAPx2_ASAP7_75t_R FILLER_204_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_378 ();
 DECAPx6_ASAP7_75t_R FILLER_204_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_445 ();
 DECAPx1_ASAP7_75t_R FILLER_204_452 ();
 DECAPx1_ASAP7_75t_R FILLER_204_470 ();
 DECAPx10_ASAP7_75t_R FILLER_204_480 ();
 FILLER_ASAP7_75t_R FILLER_204_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_504 ();
 DECAPx4_ASAP7_75t_R FILLER_204_527 ();
 FILLER_ASAP7_75t_R FILLER_204_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_549 ();
 DECAPx1_ASAP7_75t_R FILLER_204_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_560 ();
 DECAPx4_ASAP7_75t_R FILLER_204_587 ();
 FILLER_ASAP7_75t_R FILLER_204_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_599 ();
 DECAPx4_ASAP7_75t_R FILLER_204_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_618 ();
 DECAPx1_ASAP7_75t_R FILLER_204_649 ();
 DECAPx1_ASAP7_75t_R FILLER_204_665 ();
 DECAPx10_ASAP7_75t_R FILLER_204_690 ();
 DECAPx10_ASAP7_75t_R FILLER_204_712 ();
 DECAPx4_ASAP7_75t_R FILLER_204_734 ();
 FILLER_ASAP7_75t_R FILLER_204_744 ();
 DECAPx1_ASAP7_75t_R FILLER_204_758 ();
 DECAPx6_ASAP7_75t_R FILLER_204_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_815 ();
 DECAPx6_ASAP7_75t_R FILLER_204_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_836 ();
 DECAPx2_ASAP7_75t_R FILLER_204_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_855 ();
 FILLER_ASAP7_75t_R FILLER_204_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_870 ();
 DECAPx10_ASAP7_75t_R FILLER_204_889 ();
 DECAPx1_ASAP7_75t_R FILLER_204_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_915 ();
 DECAPx4_ASAP7_75t_R FILLER_204_919 ();
 DECAPx4_ASAP7_75t_R FILLER_204_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_942 ();
 DECAPx4_ASAP7_75t_R FILLER_204_961 ();
 FILLER_ASAP7_75t_R FILLER_204_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_973 ();
 DECAPx6_ASAP7_75t_R FILLER_204_990 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1080 ();
 FILLER_ASAP7_75t_R FILLER_204_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1190 ();
 FILLER_ASAP7_75t_R FILLER_204_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1273 ();
 FILLER_ASAP7_75t_R FILLER_204_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1285 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1299 ();
 FILLER_ASAP7_75t_R FILLER_204_1303 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1372 ();
 FILLER_ASAP7_75t_R FILLER_204_1384 ();
 FILLER_ASAP7_75t_R FILLER_204_1388 ();
 DECAPx4_ASAP7_75t_R FILLER_205_2 ();
 FILLER_ASAP7_75t_R FILLER_205_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_102 ();
 DECAPx6_ASAP7_75t_R FILLER_205_106 ();
 FILLER_ASAP7_75t_R FILLER_205_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_122 ();
 DECAPx4_ASAP7_75t_R FILLER_205_130 ();
 FILLER_ASAP7_75t_R FILLER_205_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_142 ();
 DECAPx2_ASAP7_75t_R FILLER_205_149 ();
 FILLER_ASAP7_75t_R FILLER_205_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_157 ();
 DECAPx6_ASAP7_75t_R FILLER_205_161 ();
 DECAPx1_ASAP7_75t_R FILLER_205_205 ();
 DECAPx6_ASAP7_75t_R FILLER_205_217 ();
 DECAPx10_ASAP7_75t_R FILLER_205_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_274 ();
 DECAPx4_ASAP7_75t_R FILLER_205_281 ();
 DECAPx10_ASAP7_75t_R FILLER_205_303 ();
 DECAPx10_ASAP7_75t_R FILLER_205_325 ();
 DECAPx6_ASAP7_75t_R FILLER_205_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_361 ();
 DECAPx4_ASAP7_75t_R FILLER_205_370 ();
 DECAPx10_ASAP7_75t_R FILLER_205_394 ();
 DECAPx1_ASAP7_75t_R FILLER_205_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_420 ();
 DECAPx1_ASAP7_75t_R FILLER_205_437 ();
 DECAPx10_ASAP7_75t_R FILLER_205_455 ();
 DECAPx1_ASAP7_75t_R FILLER_205_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_481 ();
 DECAPx2_ASAP7_75t_R FILLER_205_490 ();
 FILLER_ASAP7_75t_R FILLER_205_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_507 ();
 DECAPx4_ASAP7_75t_R FILLER_205_518 ();
 FILLER_ASAP7_75t_R FILLER_205_528 ();
 DECAPx1_ASAP7_75t_R FILLER_205_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_545 ();
 FILLER_ASAP7_75t_R FILLER_205_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_601 ();
 DECAPx2_ASAP7_75t_R FILLER_205_623 ();
 FILLER_ASAP7_75t_R FILLER_205_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_631 ();
 DECAPx4_ASAP7_75t_R FILLER_205_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_649 ();
 FILLER_ASAP7_75t_R FILLER_205_656 ();
 DECAPx2_ASAP7_75t_R FILLER_205_664 ();
 FILLER_ASAP7_75t_R FILLER_205_670 ();
 DECAPx10_ASAP7_75t_R FILLER_205_679 ();
 FILLER_ASAP7_75t_R FILLER_205_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_703 ();
 FILLER_ASAP7_75t_R FILLER_205_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_767 ();
 FILLER_ASAP7_75t_R FILLER_205_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_778 ();
 DECAPx1_ASAP7_75t_R FILLER_205_800 ();
 DECAPx4_ASAP7_75t_R FILLER_205_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_840 ();
 FILLER_ASAP7_75t_R FILLER_205_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_855 ();
 DECAPx4_ASAP7_75t_R FILLER_205_882 ();
 DECAPx1_ASAP7_75t_R FILLER_205_907 ();
 DECAPx4_ASAP7_75t_R FILLER_205_914 ();
 DECAPx2_ASAP7_75t_R FILLER_205_926 ();
 DECAPx4_ASAP7_75t_R FILLER_205_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_948 ();
 DECAPx6_ASAP7_75t_R FILLER_205_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_966 ();
 DECAPx6_ASAP7_75t_R FILLER_205_974 ();
 FILLER_ASAP7_75t_R FILLER_205_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_990 ();
 FILLER_ASAP7_75t_R FILLER_205_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1047 ();
 FILLER_ASAP7_75t_R FILLER_205_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1170 ();
 FILLER_ASAP7_75t_R FILLER_205_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1190 ();
 FILLER_ASAP7_75t_R FILLER_205_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1225 ();
 FILLER_ASAP7_75t_R FILLER_205_1241 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1246 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1264 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1318 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1361 ();
 DECAPx6_ASAP7_75t_R FILLER_206_2 ();
 DECAPx2_ASAP7_75t_R FILLER_206_16 ();
 FILLER_ASAP7_75t_R FILLER_206_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_30 ();
 DECAPx1_ASAP7_75t_R FILLER_206_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_57 ();
 DECAPx6_ASAP7_75t_R FILLER_206_64 ();
 DECAPx2_ASAP7_75t_R FILLER_206_99 ();
 DECAPx1_ASAP7_75t_R FILLER_206_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_173 ();
 DECAPx1_ASAP7_75t_R FILLER_206_181 ();
 DECAPx2_ASAP7_75t_R FILLER_206_204 ();
 FILLER_ASAP7_75t_R FILLER_206_232 ();
 DECAPx10_ASAP7_75t_R FILLER_206_240 ();
 DECAPx2_ASAP7_75t_R FILLER_206_262 ();
 FILLER_ASAP7_75t_R FILLER_206_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_270 ();
 DECAPx10_ASAP7_75t_R FILLER_206_277 ();
 DECAPx6_ASAP7_75t_R FILLER_206_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_313 ();
 DECAPx10_ASAP7_75t_R FILLER_206_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_342 ();
 DECAPx2_ASAP7_75t_R FILLER_206_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_373 ();
 DECAPx10_ASAP7_75t_R FILLER_206_381 ();
 DECAPx6_ASAP7_75t_R FILLER_206_403 ();
 DECAPx2_ASAP7_75t_R FILLER_206_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_439 ();
 DECAPx1_ASAP7_75t_R FILLER_206_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_464 ();
 DECAPx2_ASAP7_75t_R FILLER_206_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_477 ();
 FILLER_ASAP7_75t_R FILLER_206_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_486 ();
 DECAPx6_ASAP7_75t_R FILLER_206_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_527 ();
 DECAPx2_ASAP7_75t_R FILLER_206_554 ();
 DECAPx1_ASAP7_75t_R FILLER_206_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_570 ();
 DECAPx2_ASAP7_75t_R FILLER_206_581 ();
 FILLER_ASAP7_75t_R FILLER_206_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_589 ();
 DECAPx4_ASAP7_75t_R FILLER_206_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_603 ();
 DECAPx1_ASAP7_75t_R FILLER_206_614 ();
 DECAPx10_ASAP7_75t_R FILLER_206_621 ();
 DECAPx4_ASAP7_75t_R FILLER_206_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_653 ();
 DECAPx6_ASAP7_75t_R FILLER_206_660 ();
 DECAPx2_ASAP7_75t_R FILLER_206_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_680 ();
 DECAPx10_ASAP7_75t_R FILLER_206_715 ();
 DECAPx2_ASAP7_75t_R FILLER_206_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_778 ();
 DECAPx2_ASAP7_75t_R FILLER_206_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_793 ();
 DECAPx4_ASAP7_75t_R FILLER_206_804 ();
 FILLER_ASAP7_75t_R FILLER_206_814 ();
 FILLER_ASAP7_75t_R FILLER_206_827 ();
 DECAPx6_ASAP7_75t_R FILLER_206_841 ();
 FILLER_ASAP7_75t_R FILLER_206_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_857 ();
 DECAPx6_ASAP7_75t_R FILLER_206_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_895 ();
 DECAPx4_ASAP7_75t_R FILLER_206_951 ();
 FILLER_ASAP7_75t_R FILLER_206_961 ();
 DECAPx1_ASAP7_75t_R FILLER_206_983 ();
 FILLER_ASAP7_75t_R FILLER_206_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1178 ();
 FILLER_ASAP7_75t_R FILLER_206_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1190 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1217 ();
 FILLER_ASAP7_75t_R FILLER_206_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1242 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1253 ();
 FILLER_ASAP7_75t_R FILLER_206_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1261 ();
 FILLER_ASAP7_75t_R FILLER_206_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1267 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1277 ();
 FILLER_ASAP7_75t_R FILLER_206_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1314 ();
 FILLER_ASAP7_75t_R FILLER_206_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1339 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1347 ();
 FILLER_ASAP7_75t_R FILLER_206_1357 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1394 ();
 DECAPx10_ASAP7_75t_R FILLER_207_2 ();
 DECAPx1_ASAP7_75t_R FILLER_207_24 ();
 DECAPx6_ASAP7_75t_R FILLER_207_106 ();
 FILLER_ASAP7_75t_R FILLER_207_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_122 ();
 DECAPx4_ASAP7_75t_R FILLER_207_126 ();
 FILLER_ASAP7_75t_R FILLER_207_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_138 ();
 DECAPx10_ASAP7_75t_R FILLER_207_152 ();
 DECAPx2_ASAP7_75t_R FILLER_207_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_180 ();
 DECAPx10_ASAP7_75t_R FILLER_207_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_209 ();
 DECAPx6_ASAP7_75t_R FILLER_207_216 ();
 DECAPx1_ASAP7_75t_R FILLER_207_230 ();
 DECAPx4_ASAP7_75t_R FILLER_207_240 ();
 DECAPx10_ASAP7_75t_R FILLER_207_272 ();
 DECAPx10_ASAP7_75t_R FILLER_207_294 ();
 DECAPx2_ASAP7_75t_R FILLER_207_316 ();
 DECAPx2_ASAP7_75t_R FILLER_207_330 ();
 DECAPx6_ASAP7_75t_R FILLER_207_344 ();
 FILLER_ASAP7_75t_R FILLER_207_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_360 ();
 DECAPx2_ASAP7_75t_R FILLER_207_365 ();
 FILLER_ASAP7_75t_R FILLER_207_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_373 ();
 DECAPx6_ASAP7_75t_R FILLER_207_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_402 ();
 FILLER_ASAP7_75t_R FILLER_207_409 ();
 DECAPx10_ASAP7_75t_R FILLER_207_417 ();
 DECAPx2_ASAP7_75t_R FILLER_207_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_445 ();
 DECAPx1_ASAP7_75t_R FILLER_207_452 ();
 DECAPx2_ASAP7_75t_R FILLER_207_472 ();
 DECAPx1_ASAP7_75t_R FILLER_207_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_496 ();
 DECAPx2_ASAP7_75t_R FILLER_207_513 ();
 FILLER_ASAP7_75t_R FILLER_207_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_521 ();
 DECAPx2_ASAP7_75t_R FILLER_207_535 ();
 FILLER_ASAP7_75t_R FILLER_207_541 ();
 DECAPx6_ASAP7_75t_R FILLER_207_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_560 ();
 DECAPx2_ASAP7_75t_R FILLER_207_567 ();
 DECAPx10_ASAP7_75t_R FILLER_207_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_602 ();
 DECAPx2_ASAP7_75t_R FILLER_207_629 ();
 FILLER_ASAP7_75t_R FILLER_207_635 ();
 DECAPx1_ASAP7_75t_R FILLER_207_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_683 ();
 FILLER_ASAP7_75t_R FILLER_207_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_694 ();
 FILLER_ASAP7_75t_R FILLER_207_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_703 ();
 DECAPx1_ASAP7_75t_R FILLER_207_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_714 ();
 DECAPx2_ASAP7_75t_R FILLER_207_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_739 ();
 FILLER_ASAP7_75t_R FILLER_207_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_754 ();
 FILLER_ASAP7_75t_R FILLER_207_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_786 ();
 DECAPx2_ASAP7_75t_R FILLER_207_796 ();
 FILLER_ASAP7_75t_R FILLER_207_802 ();
 FILLER_ASAP7_75t_R FILLER_207_826 ();
 DECAPx6_ASAP7_75t_R FILLER_207_848 ();
 FILLER_ASAP7_75t_R FILLER_207_862 ();
 DECAPx6_ASAP7_75t_R FILLER_207_867 ();
 DECAPx2_ASAP7_75t_R FILLER_207_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_887 ();
 DECAPx10_ASAP7_75t_R FILLER_207_894 ();
 DECAPx1_ASAP7_75t_R FILLER_207_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_923 ();
 DECAPx6_ASAP7_75t_R FILLER_207_926 ();
 DECAPx1_ASAP7_75t_R FILLER_207_940 ();
 DECAPx2_ASAP7_75t_R FILLER_207_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_963 ();
 DECAPx6_ASAP7_75t_R FILLER_207_973 ();
 DECAPx10_ASAP7_75t_R FILLER_207_991 ();
 FILLER_ASAP7_75t_R FILLER_207_1013 ();
 FILLER_ASAP7_75t_R FILLER_207_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1070 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1081 ();
 FILLER_ASAP7_75t_R FILLER_207_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1235 ();
 FILLER_ASAP7_75t_R FILLER_207_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1310 ();
 FILLER_ASAP7_75t_R FILLER_207_1318 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1372 ();
 DECAPx10_ASAP7_75t_R FILLER_208_2 ();
 DECAPx1_ASAP7_75t_R FILLER_208_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_28 ();
 FILLER_ASAP7_75t_R FILLER_208_35 ();
 DECAPx6_ASAP7_75t_R FILLER_208_52 ();
 DECAPx1_ASAP7_75t_R FILLER_208_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_70 ();
 DECAPx6_ASAP7_75t_R FILLER_208_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_88 ();
 FILLER_ASAP7_75t_R FILLER_208_115 ();
 FILLER_ASAP7_75t_R FILLER_208_120 ();
 FILLER_ASAP7_75t_R FILLER_208_125 ();
 DECAPx1_ASAP7_75t_R FILLER_208_133 ();
 DECAPx6_ASAP7_75t_R FILLER_208_163 ();
 DECAPx1_ASAP7_75t_R FILLER_208_177 ();
 DECAPx6_ASAP7_75t_R FILLER_208_187 ();
 FILLER_ASAP7_75t_R FILLER_208_201 ();
 DECAPx10_ASAP7_75t_R FILLER_208_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_239 ();
 DECAPx1_ASAP7_75t_R FILLER_208_246 ();
 DECAPx4_ASAP7_75t_R FILLER_208_258 ();
 FILLER_ASAP7_75t_R FILLER_208_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_270 ();
 DECAPx4_ASAP7_75t_R FILLER_208_279 ();
 FILLER_ASAP7_75t_R FILLER_208_289 ();
 DECAPx1_ASAP7_75t_R FILLER_208_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_303 ();
 DECAPx10_ASAP7_75t_R FILLER_208_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_332 ();
 DECAPx10_ASAP7_75t_R FILLER_208_341 ();
 DECAPx6_ASAP7_75t_R FILLER_208_363 ();
 DECAPx2_ASAP7_75t_R FILLER_208_377 ();
 FILLER_ASAP7_75t_R FILLER_208_391 ();
 DECAPx4_ASAP7_75t_R FILLER_208_413 ();
 FILLER_ASAP7_75t_R FILLER_208_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_425 ();
 DECAPx2_ASAP7_75t_R FILLER_208_432 ();
 FILLER_ASAP7_75t_R FILLER_208_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_470 ();
 DECAPx6_ASAP7_75t_R FILLER_208_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_497 ();
 DECAPx2_ASAP7_75t_R FILLER_208_516 ();
 DECAPx1_ASAP7_75t_R FILLER_208_564 ();
 FILLER_ASAP7_75t_R FILLER_208_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_602 ();
 DECAPx2_ASAP7_75t_R FILLER_208_666 ();
 FILLER_ASAP7_75t_R FILLER_208_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_696 ();
 DECAPx6_ASAP7_75t_R FILLER_208_703 ();
 FILLER_ASAP7_75t_R FILLER_208_717 ();
 DECAPx1_ASAP7_75t_R FILLER_208_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_729 ();
 DECAPx1_ASAP7_75t_R FILLER_208_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_737 ();
 DECAPx1_ASAP7_75t_R FILLER_208_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_789 ();
 DECAPx6_ASAP7_75t_R FILLER_208_812 ();
 DECAPx2_ASAP7_75t_R FILLER_208_826 ();
 DECAPx2_ASAP7_75t_R FILLER_208_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_883 ();
 DECAPx4_ASAP7_75t_R FILLER_208_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_907 ();
 DECAPx1_ASAP7_75t_R FILLER_208_934 ();
 DECAPx4_ASAP7_75t_R FILLER_208_969 ();
 FILLER_ASAP7_75t_R FILLER_208_979 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1004 ();
 FILLER_ASAP7_75t_R FILLER_208_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1060 ();
 FILLER_ASAP7_75t_R FILLER_208_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1078 ();
 FILLER_ASAP7_75t_R FILLER_208_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1090 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1143 ();
 FILLER_ASAP7_75t_R FILLER_208_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1177 ();
 FILLER_ASAP7_75t_R FILLER_208_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1228 ();
 FILLER_ASAP7_75t_R FILLER_208_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1255 ();
 FILLER_ASAP7_75t_R FILLER_208_1265 ();
 FILLER_ASAP7_75t_R FILLER_208_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1277 ();
 FILLER_ASAP7_75t_R FILLER_208_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1338 ();
 FILLER_ASAP7_75t_R FILLER_208_1345 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_209_2 ();
 FILLER_ASAP7_75t_R FILLER_209_24 ();
 DECAPx4_ASAP7_75t_R FILLER_209_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_66 ();
 DECAPx2_ASAP7_75t_R FILLER_209_79 ();
 FILLER_ASAP7_75t_R FILLER_209_85 ();
 DECAPx1_ASAP7_75t_R FILLER_209_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_106 ();
 FILLER_ASAP7_75t_R FILLER_209_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_135 ();
 DECAPx2_ASAP7_75t_R FILLER_209_142 ();
 FILLER_ASAP7_75t_R FILLER_209_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_150 ();
 DECAPx1_ASAP7_75t_R FILLER_209_154 ();
 FILLER_ASAP7_75t_R FILLER_209_173 ();
 DECAPx4_ASAP7_75t_R FILLER_209_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_220 ();
 DECAPx1_ASAP7_75t_R FILLER_209_237 ();
 DECAPx10_ASAP7_75t_R FILLER_209_247 ();
 DECAPx1_ASAP7_75t_R FILLER_209_269 ();
 DECAPx10_ASAP7_75t_R FILLER_209_287 ();
 DECAPx4_ASAP7_75t_R FILLER_209_309 ();
 FILLER_ASAP7_75t_R FILLER_209_326 ();
 DECAPx6_ASAP7_75t_R FILLER_209_331 ();
 DECAPx1_ASAP7_75t_R FILLER_209_345 ();
 DECAPx4_ASAP7_75t_R FILLER_209_355 ();
 FILLER_ASAP7_75t_R FILLER_209_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_367 ();
 FILLER_ASAP7_75t_R FILLER_209_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_384 ();
 DECAPx4_ASAP7_75t_R FILLER_209_391 ();
 DECAPx4_ASAP7_75t_R FILLER_209_409 ();
 FILLER_ASAP7_75t_R FILLER_209_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_421 ();
 DECAPx2_ASAP7_75t_R FILLER_209_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_442 ();
 DECAPx10_ASAP7_75t_R FILLER_209_449 ();
 DECAPx4_ASAP7_75t_R FILLER_209_471 ();
 FILLER_ASAP7_75t_R FILLER_209_481 ();
 DECAPx6_ASAP7_75t_R FILLER_209_489 ();
 DECAPx2_ASAP7_75t_R FILLER_209_503 ();
 DECAPx2_ASAP7_75t_R FILLER_209_521 ();
 FILLER_ASAP7_75t_R FILLER_209_527 ();
 DECAPx10_ASAP7_75t_R FILLER_209_535 ();
 DECAPx1_ASAP7_75t_R FILLER_209_557 ();
 FILLER_ASAP7_75t_R FILLER_209_587 ();
 DECAPx4_ASAP7_75t_R FILLER_209_621 ();
 FILLER_ASAP7_75t_R FILLER_209_631 ();
 FILLER_ASAP7_75t_R FILLER_209_640 ();
 FILLER_ASAP7_75t_R FILLER_209_675 ();
 DECAPx2_ASAP7_75t_R FILLER_209_690 ();
 FILLER_ASAP7_75t_R FILLER_209_696 ();
 FILLER_ASAP7_75t_R FILLER_209_753 ();
 DECAPx1_ASAP7_75t_R FILLER_209_789 ();
 DECAPx2_ASAP7_75t_R FILLER_209_819 ();
 FILLER_ASAP7_75t_R FILLER_209_825 ();
 DECAPx2_ASAP7_75t_R FILLER_209_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_845 ();
 DECAPx1_ASAP7_75t_R FILLER_209_872 ();
 DECAPx2_ASAP7_75t_R FILLER_209_933 ();
 FILLER_ASAP7_75t_R FILLER_209_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_941 ();
 DECAPx6_ASAP7_75t_R FILLER_209_949 ();
 FILLER_ASAP7_75t_R FILLER_209_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_965 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1016 ();
 FILLER_ASAP7_75t_R FILLER_209_1022 ();
 FILLER_ASAP7_75t_R FILLER_209_1034 ();
 FILLER_ASAP7_75t_R FILLER_209_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1089 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_209_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1219 ();
 FILLER_ASAP7_75t_R FILLER_209_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_209_1255 ();
 FILLER_ASAP7_75t_R FILLER_209_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1267 ();
 FILLER_ASAP7_75t_R FILLER_209_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1318 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1324 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1328 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_210_2 ();
 DECAPx2_ASAP7_75t_R FILLER_210_24 ();
 FILLER_ASAP7_75t_R FILLER_210_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_32 ();
 DECAPx2_ASAP7_75t_R FILLER_210_48 ();
 FILLER_ASAP7_75t_R FILLER_210_54 ();
 FILLER_ASAP7_75t_R FILLER_210_62 ();
 DECAPx6_ASAP7_75t_R FILLER_210_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_107 ();
 DECAPx1_ASAP7_75t_R FILLER_210_144 ();
 FILLER_ASAP7_75t_R FILLER_210_151 ();
 FILLER_ASAP7_75t_R FILLER_210_179 ();
 DECAPx1_ASAP7_75t_R FILLER_210_189 ();
 DECAPx4_ASAP7_75t_R FILLER_210_203 ();
 FILLER_ASAP7_75t_R FILLER_210_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_215 ();
 DECAPx2_ASAP7_75t_R FILLER_210_224 ();
 FILLER_ASAP7_75t_R FILLER_210_230 ();
 DECAPx4_ASAP7_75t_R FILLER_210_246 ();
 FILLER_ASAP7_75t_R FILLER_210_273 ();
 DECAPx1_ASAP7_75t_R FILLER_210_291 ();
 DECAPx4_ASAP7_75t_R FILLER_210_300 ();
 FILLER_ASAP7_75t_R FILLER_210_310 ();
 FILLER_ASAP7_75t_R FILLER_210_320 ();
 FILLER_ASAP7_75t_R FILLER_210_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_330 ();
 DECAPx1_ASAP7_75t_R FILLER_210_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_349 ();
 DECAPx4_ASAP7_75t_R FILLER_210_369 ();
 FILLER_ASAP7_75t_R FILLER_210_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_381 ();
 DECAPx1_ASAP7_75t_R FILLER_210_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_402 ();
 FILLER_ASAP7_75t_R FILLER_210_410 ();
 DECAPx1_ASAP7_75t_R FILLER_210_418 ();
 DECAPx1_ASAP7_75t_R FILLER_210_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_434 ();
 DECAPx2_ASAP7_75t_R FILLER_210_453 ();
 FILLER_ASAP7_75t_R FILLER_210_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_461 ();
 FILLER_ASAP7_75t_R FILLER_210_478 ();
 FILLER_ASAP7_75t_R FILLER_210_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_485 ();
 DECAPx2_ASAP7_75t_R FILLER_210_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_504 ();
 DECAPx1_ASAP7_75t_R FILLER_210_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_524 ();
 DECAPx4_ASAP7_75t_R FILLER_210_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_538 ();
 DECAPx1_ASAP7_75t_R FILLER_210_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_560 ();
 DECAPx2_ASAP7_75t_R FILLER_210_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_574 ();
 DECAPx2_ASAP7_75t_R FILLER_210_578 ();
 DECAPx4_ASAP7_75t_R FILLER_210_620 ();
 DECAPx2_ASAP7_75t_R FILLER_210_651 ();
 FILLER_ASAP7_75t_R FILLER_210_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_699 ();
 DECAPx4_ASAP7_75t_R FILLER_210_706 ();
 FILLER_ASAP7_75t_R FILLER_210_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_718 ();
 DECAPx6_ASAP7_75t_R FILLER_210_725 ();
 DECAPx2_ASAP7_75t_R FILLER_210_739 ();
 DECAPx1_ASAP7_75t_R FILLER_210_763 ();
 DECAPx6_ASAP7_75t_R FILLER_210_777 ();
 FILLER_ASAP7_75t_R FILLER_210_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_793 ();
 DECAPx2_ASAP7_75t_R FILLER_210_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_806 ();
 DECAPx10_ASAP7_75t_R FILLER_210_810 ();
 DECAPx10_ASAP7_75t_R FILLER_210_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_854 ();
 DECAPx2_ASAP7_75t_R FILLER_210_864 ();
 DECAPx2_ASAP7_75t_R FILLER_210_896 ();
 DECAPx6_ASAP7_75t_R FILLER_210_905 ();
 DECAPx1_ASAP7_75t_R FILLER_210_919 ();
 DECAPx1_ASAP7_75t_R FILLER_210_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_930 ();
 DECAPx6_ASAP7_75t_R FILLER_210_937 ();
 FILLER_ASAP7_75t_R FILLER_210_951 ();
 DECAPx2_ASAP7_75t_R FILLER_210_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_967 ();
 DECAPx10_ASAP7_75t_R FILLER_210_973 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1049 ();
 FILLER_ASAP7_75t_R FILLER_210_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1072 ();
 FILLER_ASAP7_75t_R FILLER_210_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1165 ();
 FILLER_ASAP7_75t_R FILLER_210_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1233 ();
 FILLER_ASAP7_75t_R FILLER_210_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_210_1273 ();
 FILLER_ASAP7_75t_R FILLER_210_1283 ();
 FILLER_ASAP7_75t_R FILLER_210_1298 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1326 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1340 ();
 FILLER_ASAP7_75t_R FILLER_210_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_211_2 ();
 DECAPx2_ASAP7_75t_R FILLER_211_24 ();
 FILLER_ASAP7_75t_R FILLER_211_30 ();
 DECAPx1_ASAP7_75t_R FILLER_211_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_71 ();
 FILLER_ASAP7_75t_R FILLER_211_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_77 ();
 DECAPx2_ASAP7_75t_R FILLER_211_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_102 ();
 DECAPx1_ASAP7_75t_R FILLER_211_106 ();
 DECAPx2_ASAP7_75t_R FILLER_211_125 ();
 FILLER_ASAP7_75t_R FILLER_211_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_133 ();
 FILLER_ASAP7_75t_R FILLER_211_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_162 ();
 DECAPx6_ASAP7_75t_R FILLER_211_202 ();
 DECAPx1_ASAP7_75t_R FILLER_211_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_220 ();
 DECAPx1_ASAP7_75t_R FILLER_211_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_285 ();
 DECAPx1_ASAP7_75t_R FILLER_211_307 ();
 DECAPx4_ASAP7_75t_R FILLER_211_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_343 ();
 DECAPx6_ASAP7_75t_R FILLER_211_350 ();
 DECAPx1_ASAP7_75t_R FILLER_211_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_368 ();
 FILLER_ASAP7_75t_R FILLER_211_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_384 ();
 DECAPx2_ASAP7_75t_R FILLER_211_391 ();
 FILLER_ASAP7_75t_R FILLER_211_397 ();
 DECAPx2_ASAP7_75t_R FILLER_211_411 ();
 FILLER_ASAP7_75t_R FILLER_211_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_419 ();
 FILLER_ASAP7_75t_R FILLER_211_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_443 ();
 FILLER_ASAP7_75t_R FILLER_211_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_452 ();
 DECAPx4_ASAP7_75t_R FILLER_211_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_466 ();
 DECAPx2_ASAP7_75t_R FILLER_211_476 ();
 FILLER_ASAP7_75t_R FILLER_211_482 ();
 DECAPx2_ASAP7_75t_R FILLER_211_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_568 ();
 FILLER_ASAP7_75t_R FILLER_211_579 ();
 DECAPx4_ASAP7_75t_R FILLER_211_619 ();
 FILLER_ASAP7_75t_R FILLER_211_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_631 ();
 DECAPx2_ASAP7_75t_R FILLER_211_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_645 ();
 DECAPx2_ASAP7_75t_R FILLER_211_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_707 ();
 FILLER_ASAP7_75t_R FILLER_211_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_716 ();
 DECAPx6_ASAP7_75t_R FILLER_211_725 ();
 DECAPx2_ASAP7_75t_R FILLER_211_746 ();
 FILLER_ASAP7_75t_R FILLER_211_752 ();
 DECAPx10_ASAP7_75t_R FILLER_211_780 ();
 DECAPx2_ASAP7_75t_R FILLER_211_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_808 ();
 DECAPx2_ASAP7_75t_R FILLER_211_833 ();
 FILLER_ASAP7_75t_R FILLER_211_839 ();
 DECAPx10_ASAP7_75t_R FILLER_211_849 ();
 DECAPx6_ASAP7_75t_R FILLER_211_871 ();
 DECAPx10_ASAP7_75t_R FILLER_211_888 ();
 DECAPx6_ASAP7_75t_R FILLER_211_910 ();
 DECAPx2_ASAP7_75t_R FILLER_211_926 ();
 FILLER_ASAP7_75t_R FILLER_211_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_945 ();
 DECAPx6_ASAP7_75t_R FILLER_211_991 ();
 FILLER_ASAP7_75t_R FILLER_211_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_211_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1137 ();
 FILLER_ASAP7_75t_R FILLER_211_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1243 ();
 FILLER_ASAP7_75t_R FILLER_211_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_212_2 ();
 DECAPx4_ASAP7_75t_R FILLER_212_24 ();
 DECAPx1_ASAP7_75t_R FILLER_212_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_44 ();
 FILLER_ASAP7_75t_R FILLER_212_74 ();
 FILLER_ASAP7_75t_R FILLER_212_102 ();
 DECAPx2_ASAP7_75t_R FILLER_212_134 ();
 FILLER_ASAP7_75t_R FILLER_212_140 ();
 DECAPx1_ASAP7_75t_R FILLER_212_150 ();
 DECAPx2_ASAP7_75t_R FILLER_212_160 ();
 FILLER_ASAP7_75t_R FILLER_212_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_168 ();
 DECAPx4_ASAP7_75t_R FILLER_212_172 ();
 FILLER_ASAP7_75t_R FILLER_212_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_191 ();
 DECAPx1_ASAP7_75t_R FILLER_212_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_212 ();
 DECAPx2_ASAP7_75t_R FILLER_212_223 ();
 FILLER_ASAP7_75t_R FILLER_212_229 ();
 DECAPx2_ASAP7_75t_R FILLER_212_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_243 ();
 DECAPx2_ASAP7_75t_R FILLER_212_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_272 ();
 FILLER_ASAP7_75t_R FILLER_212_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_294 ();
 DECAPx1_ASAP7_75t_R FILLER_212_307 ();
 DECAPx6_ASAP7_75t_R FILLER_212_324 ();
 DECAPx1_ASAP7_75t_R FILLER_212_338 ();
 DECAPx6_ASAP7_75t_R FILLER_212_350 ();
 DECAPx1_ASAP7_75t_R FILLER_212_364 ();
 DECAPx2_ASAP7_75t_R FILLER_212_374 ();
 FILLER_ASAP7_75t_R FILLER_212_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_382 ();
 DECAPx6_ASAP7_75t_R FILLER_212_393 ();
 DECAPx1_ASAP7_75t_R FILLER_212_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_417 ();
 DECAPx6_ASAP7_75t_R FILLER_212_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_435 ();
 FILLER_ASAP7_75t_R FILLER_212_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_466 ();
 DECAPx2_ASAP7_75t_R FILLER_212_493 ();
 FILLER_ASAP7_75t_R FILLER_212_499 ();
 DECAPx1_ASAP7_75t_R FILLER_212_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_508 ();
 DECAPx1_ASAP7_75t_R FILLER_212_515 ();
 DECAPx4_ASAP7_75t_R FILLER_212_525 ();
 FILLER_ASAP7_75t_R FILLER_212_535 ();
 DECAPx2_ASAP7_75t_R FILLER_212_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_549 ();
 DECAPx4_ASAP7_75t_R FILLER_212_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_563 ();
 DECAPx1_ASAP7_75t_R FILLER_212_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_594 ();
 DECAPx6_ASAP7_75t_R FILLER_212_607 ();
 FILLER_ASAP7_75t_R FILLER_212_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_623 ();
 DECAPx10_ASAP7_75t_R FILLER_212_631 ();
 FILLER_ASAP7_75t_R FILLER_212_653 ();
 DECAPx2_ASAP7_75t_R FILLER_212_662 ();
 FILLER_ASAP7_75t_R FILLER_212_668 ();
 FILLER_ASAP7_75t_R FILLER_212_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_743 ();
 DECAPx2_ASAP7_75t_R FILLER_212_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_758 ();
 DECAPx2_ASAP7_75t_R FILLER_212_765 ();
 FILLER_ASAP7_75t_R FILLER_212_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_773 ();
 DECAPx1_ASAP7_75t_R FILLER_212_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_785 ();
 DECAPx2_ASAP7_75t_R FILLER_212_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_812 ();
 DECAPx2_ASAP7_75t_R FILLER_212_821 ();
 FILLER_ASAP7_75t_R FILLER_212_835 ();
 FILLER_ASAP7_75t_R FILLER_212_843 ();
 DECAPx2_ASAP7_75t_R FILLER_212_858 ();
 FILLER_ASAP7_75t_R FILLER_212_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_866 ();
 DECAPx10_ASAP7_75t_R FILLER_212_875 ();
 DECAPx4_ASAP7_75t_R FILLER_212_897 ();
 FILLER_ASAP7_75t_R FILLER_212_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_919 ();
 DECAPx6_ASAP7_75t_R FILLER_212_923 ();
 FILLER_ASAP7_75t_R FILLER_212_937 ();
 DECAPx6_ASAP7_75t_R FILLER_212_977 ();
 DECAPx2_ASAP7_75t_R FILLER_212_991 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1063 ();
 FILLER_ASAP7_75t_R FILLER_212_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1132 ();
 FILLER_ASAP7_75t_R FILLER_212_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1224 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1260 ();
 FILLER_ASAP7_75t_R FILLER_212_1267 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1297 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1335 ();
 FILLER_ASAP7_75t_R FILLER_212_1345 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1357 ();
 FILLER_ASAP7_75t_R FILLER_212_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_213_2 ();
 DECAPx10_ASAP7_75t_R FILLER_213_24 ();
 DECAPx6_ASAP7_75t_R FILLER_213_46 ();
 FILLER_ASAP7_75t_R FILLER_213_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_62 ();
 DECAPx10_ASAP7_75t_R FILLER_213_66 ();
 DECAPx1_ASAP7_75t_R FILLER_213_88 ();
 DECAPx4_ASAP7_75t_R FILLER_213_95 ();
 FILLER_ASAP7_75t_R FILLER_213_105 ();
 DECAPx6_ASAP7_75t_R FILLER_213_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_133 ();
 DECAPx1_ASAP7_75t_R FILLER_213_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_141 ();
 DECAPx6_ASAP7_75t_R FILLER_213_168 ();
 DECAPx2_ASAP7_75t_R FILLER_213_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_188 ();
 DECAPx2_ASAP7_75t_R FILLER_213_200 ();
 FILLER_ASAP7_75t_R FILLER_213_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_208 ();
 FILLER_ASAP7_75t_R FILLER_213_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_227 ();
 DECAPx4_ASAP7_75t_R FILLER_213_236 ();
 DECAPx6_ASAP7_75t_R FILLER_213_254 ();
 FILLER_ASAP7_75t_R FILLER_213_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_270 ();
 DECAPx2_ASAP7_75t_R FILLER_213_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_287 ();
 DECAPx10_ASAP7_75t_R FILLER_213_298 ();
 DECAPx1_ASAP7_75t_R FILLER_213_320 ();
 DECAPx4_ASAP7_75t_R FILLER_213_327 ();
 FILLER_ASAP7_75t_R FILLER_213_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_339 ();
 FILLER_ASAP7_75t_R FILLER_213_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_348 ();
 DECAPx10_ASAP7_75t_R FILLER_213_355 ();
 DECAPx10_ASAP7_75t_R FILLER_213_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_399 ();
 DECAPx4_ASAP7_75t_R FILLER_213_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_439 ();
 DECAPx2_ASAP7_75t_R FILLER_213_446 ();
 DECAPx4_ASAP7_75t_R FILLER_213_455 ();
 FILLER_ASAP7_75t_R FILLER_213_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_467 ();
 DECAPx2_ASAP7_75t_R FILLER_213_474 ();
 FILLER_ASAP7_75t_R FILLER_213_480 ();
 DECAPx1_ASAP7_75t_R FILLER_213_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_489 ();
 DECAPx6_ASAP7_75t_R FILLER_213_496 ();
 DECAPx6_ASAP7_75t_R FILLER_213_550 ();
 DECAPx2_ASAP7_75t_R FILLER_213_564 ();
 DECAPx2_ASAP7_75t_R FILLER_213_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_596 ();
 DECAPx6_ASAP7_75t_R FILLER_213_648 ();
 DECAPx10_ASAP7_75t_R FILLER_213_689 ();
 DECAPx10_ASAP7_75t_R FILLER_213_711 ();
 DECAPx4_ASAP7_75t_R FILLER_213_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_743 ();
 DECAPx2_ASAP7_75t_R FILLER_213_750 ();
 FILLER_ASAP7_75t_R FILLER_213_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_758 ();
 DECAPx4_ASAP7_75t_R FILLER_213_766 ();
 DECAPx10_ASAP7_75t_R FILLER_213_810 ();
 FILLER_ASAP7_75t_R FILLER_213_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_834 ();
 DECAPx4_ASAP7_75t_R FILLER_213_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_899 ();
 FILLER_ASAP7_75t_R FILLER_213_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_923 ();
 DECAPx2_ASAP7_75t_R FILLER_213_934 ();
 DECAPx1_ASAP7_75t_R FILLER_213_955 ();
 DECAPx2_ASAP7_75t_R FILLER_213_999 ();
 FILLER_ASAP7_75t_R FILLER_213_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1023 ();
 FILLER_ASAP7_75t_R FILLER_213_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1031 ();
 FILLER_ASAP7_75t_R FILLER_213_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1219 ();
 FILLER_ASAP7_75t_R FILLER_213_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1243 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1262 ();
 FILLER_ASAP7_75t_R FILLER_213_1305 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1339 ();
 FILLER_ASAP7_75t_R FILLER_213_1351 ();
 DECAPx10_ASAP7_75t_R FILLER_214_2 ();
 DECAPx10_ASAP7_75t_R FILLER_214_24 ();
 DECAPx10_ASAP7_75t_R FILLER_214_46 ();
 DECAPx1_ASAP7_75t_R FILLER_214_68 ();
 DECAPx6_ASAP7_75t_R FILLER_214_93 ();
 DECAPx1_ASAP7_75t_R FILLER_214_107 ();
 DECAPx4_ASAP7_75t_R FILLER_214_137 ();
 FILLER_ASAP7_75t_R FILLER_214_154 ();
 DECAPx4_ASAP7_75t_R FILLER_214_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_169 ();
 DECAPx4_ASAP7_75t_R FILLER_214_180 ();
 DECAPx6_ASAP7_75t_R FILLER_214_196 ();
 FILLER_ASAP7_75t_R FILLER_214_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_218 ();
 FILLER_ASAP7_75t_R FILLER_214_225 ();
 DECAPx2_ASAP7_75t_R FILLER_214_233 ();
 FILLER_ASAP7_75t_R FILLER_214_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_247 ();
 DECAPx2_ASAP7_75t_R FILLER_214_266 ();
 FILLER_ASAP7_75t_R FILLER_214_272 ();
 DECAPx4_ASAP7_75t_R FILLER_214_284 ();
 FILLER_ASAP7_75t_R FILLER_214_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_296 ();
 DECAPx10_ASAP7_75t_R FILLER_214_307 ();
 FILLER_ASAP7_75t_R FILLER_214_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_346 ();
 FILLER_ASAP7_75t_R FILLER_214_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_355 ();
 DECAPx1_ASAP7_75t_R FILLER_214_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_374 ();
 DECAPx6_ASAP7_75t_R FILLER_214_387 ();
 FILLER_ASAP7_75t_R FILLER_214_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_403 ();
 DECAPx6_ASAP7_75t_R FILLER_214_410 ();
 DECAPx1_ASAP7_75t_R FILLER_214_424 ();
 DECAPx6_ASAP7_75t_R FILLER_214_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_450 ();
 FILLER_ASAP7_75t_R FILLER_214_460 ();
 DECAPx6_ASAP7_75t_R FILLER_214_464 ();
 DECAPx1_ASAP7_75t_R FILLER_214_478 ();
 DECAPx6_ASAP7_75t_R FILLER_214_511 ();
 DECAPx2_ASAP7_75t_R FILLER_214_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_531 ();
 DECAPx1_ASAP7_75t_R FILLER_214_543 ();
 DECAPx10_ASAP7_75t_R FILLER_214_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_599 ();
 DECAPx2_ASAP7_75t_R FILLER_214_606 ();
 DECAPx4_ASAP7_75t_R FILLER_214_615 ();
 FILLER_ASAP7_75t_R FILLER_214_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_627 ();
 DECAPx2_ASAP7_75t_R FILLER_214_634 ();
 FILLER_ASAP7_75t_R FILLER_214_640 ();
 DECAPx1_ASAP7_75t_R FILLER_214_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_667 ();
 DECAPx2_ASAP7_75t_R FILLER_214_698 ();
 FILLER_ASAP7_75t_R FILLER_214_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_706 ();
 DECAPx4_ASAP7_75t_R FILLER_214_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_737 ();
 DECAPx4_ASAP7_75t_R FILLER_214_773 ();
 FILLER_ASAP7_75t_R FILLER_214_783 ();
 DECAPx2_ASAP7_75t_R FILLER_214_791 ();
 FILLER_ASAP7_75t_R FILLER_214_797 ();
 FILLER_ASAP7_75t_R FILLER_214_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_811 ();
 DECAPx2_ASAP7_75t_R FILLER_214_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_825 ();
 FILLER_ASAP7_75t_R FILLER_214_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_844 ();
 DECAPx4_ASAP7_75t_R FILLER_214_853 ();
 FILLER_ASAP7_75t_R FILLER_214_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_905 ();
 DECAPx1_ASAP7_75t_R FILLER_214_924 ();
 FILLER_ASAP7_75t_R FILLER_214_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_950 ();
 DECAPx4_ASAP7_75t_R FILLER_214_988 ();
 FILLER_ASAP7_75t_R FILLER_214_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1000 ();
 FILLER_ASAP7_75t_R FILLER_214_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1097 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1101 ();
 FILLER_ASAP7_75t_R FILLER_214_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1182 ();
 FILLER_ASAP7_75t_R FILLER_214_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1201 ();
 FILLER_ASAP7_75t_R FILLER_214_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1220 ();
 FILLER_ASAP7_75t_R FILLER_214_1242 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1270 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1279 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1296 ();
 FILLER_ASAP7_75t_R FILLER_214_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1320 ();
 FILLER_ASAP7_75t_R FILLER_214_1326 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1331 ();
 FILLER_ASAP7_75t_R FILLER_214_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1339 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1376 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1394 ();
 DECAPx10_ASAP7_75t_R FILLER_215_2 ();
 DECAPx10_ASAP7_75t_R FILLER_215_24 ();
 DECAPx6_ASAP7_75t_R FILLER_215_46 ();
 DECAPx1_ASAP7_75t_R FILLER_215_60 ();
 DECAPx1_ASAP7_75t_R FILLER_215_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_112 ();
 DECAPx2_ASAP7_75t_R FILLER_215_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_125 ();
 DECAPx2_ASAP7_75t_R FILLER_215_135 ();
 FILLER_ASAP7_75t_R FILLER_215_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_143 ();
 DECAPx2_ASAP7_75t_R FILLER_215_157 ();
 FILLER_ASAP7_75t_R FILLER_215_206 ();
 DECAPx2_ASAP7_75t_R FILLER_215_224 ();
 FILLER_ASAP7_75t_R FILLER_215_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_249 ();
 DECAPx6_ASAP7_75t_R FILLER_215_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_270 ();
 DECAPx10_ASAP7_75t_R FILLER_215_281 ();
 DECAPx4_ASAP7_75t_R FILLER_215_303 ();
 FILLER_ASAP7_75t_R FILLER_215_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_315 ();
 DECAPx10_ASAP7_75t_R FILLER_215_336 ();
 DECAPx4_ASAP7_75t_R FILLER_215_358 ();
 DECAPx1_ASAP7_75t_R FILLER_215_376 ();
 DECAPx1_ASAP7_75t_R FILLER_215_389 ();
 DECAPx4_ASAP7_75t_R FILLER_215_399 ();
 DECAPx1_ASAP7_75t_R FILLER_215_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_425 ();
 DECAPx4_ASAP7_75t_R FILLER_215_432 ();
 DECAPx2_ASAP7_75t_R FILLER_215_448 ();
 DECAPx4_ASAP7_75t_R FILLER_215_476 ();
 FILLER_ASAP7_75t_R FILLER_215_486 ();
 DECAPx1_ASAP7_75t_R FILLER_215_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_498 ();
 FILLER_ASAP7_75t_R FILLER_215_502 ();
 FILLER_ASAP7_75t_R FILLER_215_510 ();
 DECAPx4_ASAP7_75t_R FILLER_215_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_534 ();
 DECAPx1_ASAP7_75t_R FILLER_215_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_549 ();
 DECAPx2_ASAP7_75t_R FILLER_215_569 ();
 FILLER_ASAP7_75t_R FILLER_215_575 ();
 DECAPx10_ASAP7_75t_R FILLER_215_606 ();
 DECAPx6_ASAP7_75t_R FILLER_215_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_664 ();
 FILLER_ASAP7_75t_R FILLER_215_692 ();
 DECAPx1_ASAP7_75t_R FILLER_215_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_719 ();
 DECAPx4_ASAP7_75t_R FILLER_215_746 ();
 FILLER_ASAP7_75t_R FILLER_215_756 ();
 DECAPx2_ASAP7_75t_R FILLER_215_761 ();
 FILLER_ASAP7_75t_R FILLER_215_767 ();
 DECAPx10_ASAP7_75t_R FILLER_215_779 ();
 DECAPx6_ASAP7_75t_R FILLER_215_809 ();
 DECAPx1_ASAP7_75t_R FILLER_215_823 ();
 FILLER_ASAP7_75t_R FILLER_215_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_837 ();
 DECAPx10_ASAP7_75t_R FILLER_215_844 ();
 DECAPx4_ASAP7_75t_R FILLER_215_874 ();
 FILLER_ASAP7_75t_R FILLER_215_884 ();
 DECAPx6_ASAP7_75t_R FILLER_215_898 ();
 DECAPx2_ASAP7_75t_R FILLER_215_912 ();
 DECAPx6_ASAP7_75t_R FILLER_215_938 ();
 DECAPx2_ASAP7_75t_R FILLER_215_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_958 ();
 DECAPx2_ASAP7_75t_R FILLER_215_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_973 ();
 DECAPx2_ASAP7_75t_R FILLER_215_977 ();
 FILLER_ASAP7_75t_R FILLER_215_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_985 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1012 ();
 FILLER_ASAP7_75t_R FILLER_215_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1077 ();
 FILLER_ASAP7_75t_R FILLER_215_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1107 ();
 FILLER_ASAP7_75t_R FILLER_215_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1142 ();
 FILLER_ASAP7_75t_R FILLER_215_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1221 ();
 FILLER_ASAP7_75t_R FILLER_215_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1331 ();
 FILLER_ASAP7_75t_R FILLER_215_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1362 ();
 FILLER_ASAP7_75t_R FILLER_215_1389 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1391 ();
 DECAPx10_ASAP7_75t_R FILLER_216_2 ();
 DECAPx10_ASAP7_75t_R FILLER_216_24 ();
 DECAPx10_ASAP7_75t_R FILLER_216_46 ();
 DECAPx1_ASAP7_75t_R FILLER_216_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_72 ();
 DECAPx2_ASAP7_75t_R FILLER_216_125 ();
 FILLER_ASAP7_75t_R FILLER_216_131 ();
 DECAPx4_ASAP7_75t_R FILLER_216_159 ();
 DECAPx1_ASAP7_75t_R FILLER_216_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_180 ();
 DECAPx2_ASAP7_75t_R FILLER_216_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_193 ();
 FILLER_ASAP7_75t_R FILLER_216_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_210 ();
 DECAPx2_ASAP7_75t_R FILLER_216_217 ();
 FILLER_ASAP7_75t_R FILLER_216_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_225 ();
 DECAPx2_ASAP7_75t_R FILLER_216_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_238 ();
 DECAPx10_ASAP7_75t_R FILLER_216_245 ();
 DECAPx2_ASAP7_75t_R FILLER_216_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_273 ();
 FILLER_ASAP7_75t_R FILLER_216_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_282 ();
 DECAPx2_ASAP7_75t_R FILLER_216_289 ();
 FILLER_ASAP7_75t_R FILLER_216_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_313 ();
 DECAPx10_ASAP7_75t_R FILLER_216_334 ();
 DECAPx2_ASAP7_75t_R FILLER_216_356 ();
 FILLER_ASAP7_75t_R FILLER_216_362 ();
 FILLER_ASAP7_75t_R FILLER_216_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_396 ();
 DECAPx1_ASAP7_75t_R FILLER_216_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_432 ();
 DECAPx4_ASAP7_75t_R FILLER_216_439 ();
 FILLER_ASAP7_75t_R FILLER_216_449 ();
 FILLER_ASAP7_75t_R FILLER_216_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_461 ();
 DECAPx1_ASAP7_75t_R FILLER_216_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_468 ();
 DECAPx2_ASAP7_75t_R FILLER_216_489 ();
 FILLER_ASAP7_75t_R FILLER_216_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_497 ();
 DECAPx6_ASAP7_75t_R FILLER_216_530 ();
 DECAPx1_ASAP7_75t_R FILLER_216_544 ();
 DECAPx6_ASAP7_75t_R FILLER_216_574 ();
 DECAPx2_ASAP7_75t_R FILLER_216_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_594 ();
 DECAPx6_ASAP7_75t_R FILLER_216_598 ();
 DECAPx1_ASAP7_75t_R FILLER_216_612 ();
 DECAPx2_ASAP7_75t_R FILLER_216_639 ();
 DECAPx1_ASAP7_75t_R FILLER_216_665 ();
 DECAPx1_ASAP7_75t_R FILLER_216_697 ();
 DECAPx6_ASAP7_75t_R FILLER_216_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_742 ();
 FILLER_ASAP7_75t_R FILLER_216_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_753 ();
 FILLER_ASAP7_75t_R FILLER_216_760 ();
 DECAPx4_ASAP7_75t_R FILLER_216_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_780 ();
 DECAPx6_ASAP7_75t_R FILLER_216_787 ();
 DECAPx2_ASAP7_75t_R FILLER_216_801 ();
 DECAPx4_ASAP7_75t_R FILLER_216_826 ();
 FILLER_ASAP7_75t_R FILLER_216_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_844 ();
 FILLER_ASAP7_75t_R FILLER_216_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_858 ();
 DECAPx4_ASAP7_75t_R FILLER_216_875 ();
 FILLER_ASAP7_75t_R FILLER_216_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_887 ();
 DECAPx2_ASAP7_75t_R FILLER_216_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_905 ();
 DECAPx4_ASAP7_75t_R FILLER_216_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_922 ();
 FILLER_ASAP7_75t_R FILLER_216_938 ();
 DECAPx10_ASAP7_75t_R FILLER_216_952 ();
 DECAPx2_ASAP7_75t_R FILLER_216_974 ();
 FILLER_ASAP7_75t_R FILLER_216_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_982 ();
 DECAPx6_ASAP7_75t_R FILLER_216_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1006 ();
 FILLER_ASAP7_75t_R FILLER_216_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1058 ();
 FILLER_ASAP7_75t_R FILLER_216_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1074 ();
 FILLER_ASAP7_75t_R FILLER_216_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1117 ();
 FILLER_ASAP7_75t_R FILLER_216_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1129 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1166 ();
 FILLER_ASAP7_75t_R FILLER_216_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1181 ();
 FILLER_ASAP7_75t_R FILLER_216_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1243 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1247 ();
 FILLER_ASAP7_75t_R FILLER_216_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1280 ();
 FILLER_ASAP7_75t_R FILLER_216_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1298 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1334 ();
 FILLER_ASAP7_75t_R FILLER_216_1377 ();
 FILLER_ASAP7_75t_R FILLER_216_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_217_2 ();
 DECAPx10_ASAP7_75t_R FILLER_217_24 ();
 DECAPx10_ASAP7_75t_R FILLER_217_46 ();
 DECAPx10_ASAP7_75t_R FILLER_217_68 ();
 FILLER_ASAP7_75t_R FILLER_217_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_92 ();
 DECAPx4_ASAP7_75t_R FILLER_217_96 ();
 DECAPx10_ASAP7_75t_R FILLER_217_109 ();
 DECAPx2_ASAP7_75t_R FILLER_217_139 ();
 FILLER_ASAP7_75t_R FILLER_217_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_147 ();
 DECAPx2_ASAP7_75t_R FILLER_217_187 ();
 FILLER_ASAP7_75t_R FILLER_217_193 ();
 DECAPx4_ASAP7_75t_R FILLER_217_201 ();
 DECAPx2_ASAP7_75t_R FILLER_217_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_223 ();
 DECAPx4_ASAP7_75t_R FILLER_217_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_252 ();
 DECAPx1_ASAP7_75t_R FILLER_217_272 ();
 DECAPx1_ASAP7_75t_R FILLER_217_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_288 ();
 DECAPx2_ASAP7_75t_R FILLER_217_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_301 ();
 DECAPx1_ASAP7_75t_R FILLER_217_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_312 ();
 DECAPx4_ASAP7_75t_R FILLER_217_327 ();
 FILLER_ASAP7_75t_R FILLER_217_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_347 ();
 FILLER_ASAP7_75t_R FILLER_217_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_357 ();
 DECAPx4_ASAP7_75t_R FILLER_217_374 ();
 FILLER_ASAP7_75t_R FILLER_217_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_398 ();
 DECAPx6_ASAP7_75t_R FILLER_217_411 ();
 FILLER_ASAP7_75t_R FILLER_217_425 ();
 DECAPx1_ASAP7_75t_R FILLER_217_447 ();
 DECAPx1_ASAP7_75t_R FILLER_217_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_461 ();
 DECAPx10_ASAP7_75t_R FILLER_217_468 ();
 FILLER_ASAP7_75t_R FILLER_217_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_492 ();
 DECAPx2_ASAP7_75t_R FILLER_217_501 ();
 FILLER_ASAP7_75t_R FILLER_217_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_509 ();
 DECAPx2_ASAP7_75t_R FILLER_217_539 ();
 FILLER_ASAP7_75t_R FILLER_217_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_547 ();
 DECAPx2_ASAP7_75t_R FILLER_217_554 ();
 DECAPx1_ASAP7_75t_R FILLER_217_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_590 ();
 DECAPx2_ASAP7_75t_R FILLER_217_597 ();
 FILLER_ASAP7_75t_R FILLER_217_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_605 ();
 DECAPx10_ASAP7_75t_R FILLER_217_644 ();
 DECAPx4_ASAP7_75t_R FILLER_217_666 ();
 FILLER_ASAP7_75t_R FILLER_217_683 ();
 FILLER_ASAP7_75t_R FILLER_217_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_693 ();
 DECAPx4_ASAP7_75t_R FILLER_217_708 ();
 FILLER_ASAP7_75t_R FILLER_217_718 ();
 DECAPx2_ASAP7_75t_R FILLER_217_727 ();
 FILLER_ASAP7_75t_R FILLER_217_733 ();
 DECAPx1_ASAP7_75t_R FILLER_217_789 ();
 FILLER_ASAP7_75t_R FILLER_217_808 ();
 FILLER_ASAP7_75t_R FILLER_217_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_844 ();
 DECAPx1_ASAP7_75t_R FILLER_217_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_923 ();
 FILLER_ASAP7_75t_R FILLER_217_926 ();
 DECAPx6_ASAP7_75t_R FILLER_217_940 ();
 FILLER_ASAP7_75t_R FILLER_217_954 ();
 FILLER_ASAP7_75t_R FILLER_217_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_973 ();
 DECAPx2_ASAP7_75t_R FILLER_217_985 ();
 FILLER_ASAP7_75t_R FILLER_217_991 ();
 DECAPx4_ASAP7_75t_R FILLER_217_996 ();
 FILLER_ASAP7_75t_R FILLER_217_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1046 ();
 FILLER_ASAP7_75t_R FILLER_217_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1054 ();
 FILLER_ASAP7_75t_R FILLER_217_1081 ();
 FILLER_ASAP7_75t_R FILLER_217_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1109 ();
 FILLER_ASAP7_75t_R FILLER_217_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1129 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1142 ();
 FILLER_ASAP7_75t_R FILLER_217_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1195 ();
 FILLER_ASAP7_75t_R FILLER_217_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1203 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1207 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1234 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1260 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_217_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1314 ();
 FILLER_ASAP7_75t_R FILLER_217_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1325 ();
 FILLER_ASAP7_75t_R FILLER_217_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1351 ();
 FILLER_ASAP7_75t_R FILLER_217_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_218_2 ();
 DECAPx10_ASAP7_75t_R FILLER_218_24 ();
 DECAPx10_ASAP7_75t_R FILLER_218_46 ();
 DECAPx6_ASAP7_75t_R FILLER_218_68 ();
 DECAPx2_ASAP7_75t_R FILLER_218_82 ();
 DECAPx4_ASAP7_75t_R FILLER_218_100 ();
 FILLER_ASAP7_75t_R FILLER_218_110 ();
 FILLER_ASAP7_75t_R FILLER_218_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_123 ();
 FILLER_ASAP7_75t_R FILLER_218_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_141 ();
 DECAPx2_ASAP7_75t_R FILLER_218_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_155 ();
 DECAPx1_ASAP7_75t_R FILLER_218_159 ();
 DECAPx2_ASAP7_75t_R FILLER_218_169 ();
 DECAPx10_ASAP7_75t_R FILLER_218_178 ();
 DECAPx1_ASAP7_75t_R FILLER_218_200 ();
 DECAPx1_ASAP7_75t_R FILLER_218_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_248 ();
 DECAPx2_ASAP7_75t_R FILLER_218_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_271 ();
 DECAPx6_ASAP7_75t_R FILLER_218_292 ();
 DECAPx1_ASAP7_75t_R FILLER_218_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_310 ();
 DECAPx1_ASAP7_75t_R FILLER_218_325 ();
 DECAPx10_ASAP7_75t_R FILLER_218_359 ();
 DECAPx6_ASAP7_75t_R FILLER_218_381 ();
 DECAPx1_ASAP7_75t_R FILLER_218_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_399 ();
 DECAPx6_ASAP7_75t_R FILLER_218_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_422 ();
 FILLER_ASAP7_75t_R FILLER_218_442 ();
 DECAPx2_ASAP7_75t_R FILLER_218_456 ();
 DECAPx1_ASAP7_75t_R FILLER_218_464 ();
 DECAPx10_ASAP7_75t_R FILLER_218_474 ();
 DECAPx1_ASAP7_75t_R FILLER_218_496 ();
 DECAPx2_ASAP7_75t_R FILLER_218_518 ();
 FILLER_ASAP7_75t_R FILLER_218_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_526 ();
 DECAPx2_ASAP7_75t_R FILLER_218_530 ();
 DECAPx2_ASAP7_75t_R FILLER_218_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_551 ();
 DECAPx10_ASAP7_75t_R FILLER_218_556 ();
 DECAPx4_ASAP7_75t_R FILLER_218_578 ();
 FILLER_ASAP7_75t_R FILLER_218_588 ();
 FILLER_ASAP7_75t_R FILLER_218_596 ();
 DECAPx1_ASAP7_75t_R FILLER_218_610 ();
 DECAPx2_ASAP7_75t_R FILLER_218_617 ();
 FILLER_ASAP7_75t_R FILLER_218_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_625 ();
 FILLER_ASAP7_75t_R FILLER_218_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_647 ();
 DECAPx1_ASAP7_75t_R FILLER_218_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_660 ();
 DECAPx6_ASAP7_75t_R FILLER_218_667 ();
 FILLER_ASAP7_75t_R FILLER_218_681 ();
 DECAPx10_ASAP7_75t_R FILLER_218_696 ();
 DECAPx6_ASAP7_75t_R FILLER_218_718 ();
 DECAPx1_ASAP7_75t_R FILLER_218_732 ();
 DECAPx10_ASAP7_75t_R FILLER_218_744 ();
 DECAPx1_ASAP7_75t_R FILLER_218_766 ();
 FILLER_ASAP7_75t_R FILLER_218_777 ();
 DECAPx6_ASAP7_75t_R FILLER_218_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_827 ();
 DECAPx4_ASAP7_75t_R FILLER_218_854 ();
 FILLER_ASAP7_75t_R FILLER_218_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_866 ();
 DECAPx1_ASAP7_75t_R FILLER_218_875 ();
 DECAPx6_ASAP7_75t_R FILLER_218_905 ();
 FILLER_ASAP7_75t_R FILLER_218_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_921 ();
 DECAPx2_ASAP7_75t_R FILLER_218_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_939 ();
 FILLER_ASAP7_75t_R FILLER_218_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_977 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1086 ();
 FILLER_ASAP7_75t_R FILLER_218_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1214 ();
 FILLER_ASAP7_75t_R FILLER_218_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1244 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1306 ();
 FILLER_ASAP7_75t_R FILLER_218_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1320 ();
 FILLER_ASAP7_75t_R FILLER_218_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_219_2 ();
 DECAPx10_ASAP7_75t_R FILLER_219_24 ();
 DECAPx10_ASAP7_75t_R FILLER_219_46 ();
 DECAPx2_ASAP7_75t_R FILLER_219_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_74 ();
 FILLER_ASAP7_75t_R FILLER_219_139 ();
 DECAPx2_ASAP7_75t_R FILLER_219_170 ();
 FILLER_ASAP7_75t_R FILLER_219_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_186 ();
 DECAPx4_ASAP7_75t_R FILLER_219_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_222 ();
 FILLER_ASAP7_75t_R FILLER_219_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_233 ();
 DECAPx1_ASAP7_75t_R FILLER_219_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_244 ();
 DECAPx6_ASAP7_75t_R FILLER_219_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_275 ();
 DECAPx2_ASAP7_75t_R FILLER_219_292 ();
 DECAPx10_ASAP7_75t_R FILLER_219_308 ();
 DECAPx2_ASAP7_75t_R FILLER_219_330 ();
 FILLER_ASAP7_75t_R FILLER_219_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_338 ();
 DECAPx10_ASAP7_75t_R FILLER_219_357 ();
 DECAPx2_ASAP7_75t_R FILLER_219_379 ();
 FILLER_ASAP7_75t_R FILLER_219_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_395 ();
 DECAPx2_ASAP7_75t_R FILLER_219_412 ();
 DECAPx4_ASAP7_75t_R FILLER_219_426 ();
 FILLER_ASAP7_75t_R FILLER_219_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_438 ();
 DECAPx2_ASAP7_75t_R FILLER_219_457 ();
 FILLER_ASAP7_75t_R FILLER_219_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_465 ();
 DECAPx2_ASAP7_75t_R FILLER_219_480 ();
 FILLER_ASAP7_75t_R FILLER_219_486 ();
 DECAPx10_ASAP7_75t_R FILLER_219_502 ();
 DECAPx4_ASAP7_75t_R FILLER_219_524 ();
 DECAPx4_ASAP7_75t_R FILLER_219_560 ();
 DECAPx4_ASAP7_75t_R FILLER_219_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_597 ();
 DECAPx6_ASAP7_75t_R FILLER_219_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_621 ();
 FILLER_ASAP7_75t_R FILLER_219_639 ();
 DECAPx1_ASAP7_75t_R FILLER_219_658 ();
 DECAPx2_ASAP7_75t_R FILLER_219_674 ();
 FILLER_ASAP7_75t_R FILLER_219_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_682 ();
 DECAPx4_ASAP7_75t_R FILLER_219_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_714 ();
 DECAPx2_ASAP7_75t_R FILLER_219_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_729 ();
 DECAPx6_ASAP7_75t_R FILLER_219_741 ();
 FILLER_ASAP7_75t_R FILLER_219_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_757 ();
 DECAPx6_ASAP7_75t_R FILLER_219_765 ();
 FILLER_ASAP7_75t_R FILLER_219_779 ();
 DECAPx1_ASAP7_75t_R FILLER_219_789 ();
 DECAPx2_ASAP7_75t_R FILLER_219_796 ();
 FILLER_ASAP7_75t_R FILLER_219_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_804 ();
 DECAPx10_ASAP7_75t_R FILLER_219_811 ();
 DECAPx10_ASAP7_75t_R FILLER_219_833 ();
 DECAPx4_ASAP7_75t_R FILLER_219_855 ();
 DECAPx4_ASAP7_75t_R FILLER_219_872 ();
 DECAPx10_ASAP7_75t_R FILLER_219_886 ();
 DECAPx2_ASAP7_75t_R FILLER_219_908 ();
 FILLER_ASAP7_75t_R FILLER_219_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_916 ();
 DECAPx2_ASAP7_75t_R FILLER_219_929 ();
 FILLER_ASAP7_75t_R FILLER_219_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_950 ();
 DECAPx6_ASAP7_75t_R FILLER_219_963 ();
 FILLER_ASAP7_75t_R FILLER_219_977 ();
 DECAPx1_ASAP7_75t_R FILLER_219_987 ();
 DECAPx4_ASAP7_75t_R FILLER_219_994 ();
 FILLER_ASAP7_75t_R FILLER_219_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_219_1016 ();
 FILLER_ASAP7_75t_R FILLER_219_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1144 ();
 FILLER_ASAP7_75t_R FILLER_219_1157 ();
 FILLER_ASAP7_75t_R FILLER_219_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1216 ();
 FILLER_ASAP7_75t_R FILLER_219_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1304 ();
 FILLER_ASAP7_75t_R FILLER_219_1326 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1338 ();
 FILLER_ASAP7_75t_R FILLER_219_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_220_2 ();
 DECAPx10_ASAP7_75t_R FILLER_220_24 ();
 DECAPx10_ASAP7_75t_R FILLER_220_46 ();
 DECAPx6_ASAP7_75t_R FILLER_220_68 ();
 DECAPx1_ASAP7_75t_R FILLER_220_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_86 ();
 FILLER_ASAP7_75t_R FILLER_220_119 ();
 DECAPx1_ASAP7_75t_R FILLER_220_124 ();
 DECAPx6_ASAP7_75t_R FILLER_220_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_168 ();
 FILLER_ASAP7_75t_R FILLER_220_188 ();
 DECAPx1_ASAP7_75t_R FILLER_220_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_200 ();
 DECAPx1_ASAP7_75t_R FILLER_220_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_225 ();
 DECAPx1_ASAP7_75t_R FILLER_220_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_236 ();
 FILLER_ASAP7_75t_R FILLER_220_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_261 ();
 DECAPx4_ASAP7_75t_R FILLER_220_278 ();
 FILLER_ASAP7_75t_R FILLER_220_288 ();
 FILLER_ASAP7_75t_R FILLER_220_300 ();
 DECAPx4_ASAP7_75t_R FILLER_220_320 ();
 FILLER_ASAP7_75t_R FILLER_220_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_338 ();
 FILLER_ASAP7_75t_R FILLER_220_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_344 ();
 DECAPx6_ASAP7_75t_R FILLER_220_351 ();
 FILLER_ASAP7_75t_R FILLER_220_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_395 ();
 DECAPx1_ASAP7_75t_R FILLER_220_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_412 ();
 DECAPx6_ASAP7_75t_R FILLER_220_422 ();
 FILLER_ASAP7_75t_R FILLER_220_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_438 ();
 FILLER_ASAP7_75t_R FILLER_220_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_455 ();
 DECAPx1_ASAP7_75t_R FILLER_220_464 ();
 FILLER_ASAP7_75t_R FILLER_220_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_507 ();
 DECAPx1_ASAP7_75t_R FILLER_220_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_535 ();
 FILLER_ASAP7_75t_R FILLER_220_542 ();
 DECAPx1_ASAP7_75t_R FILLER_220_558 ();
 DECAPx1_ASAP7_75t_R FILLER_220_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_581 ();
 DECAPx6_ASAP7_75t_R FILLER_220_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_606 ();
 DECAPx2_ASAP7_75t_R FILLER_220_621 ();
 DECAPx1_ASAP7_75t_R FILLER_220_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_637 ();
 DECAPx4_ASAP7_75t_R FILLER_220_644 ();
 FILLER_ASAP7_75t_R FILLER_220_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_656 ();
 FILLER_ASAP7_75t_R FILLER_220_671 ();
 DECAPx10_ASAP7_75t_R FILLER_220_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_739 ();
 FILLER_ASAP7_75t_R FILLER_220_756 ();
 DECAPx2_ASAP7_75t_R FILLER_220_774 ();
 FILLER_ASAP7_75t_R FILLER_220_780 ();
 DECAPx2_ASAP7_75t_R FILLER_220_790 ();
 DECAPx4_ASAP7_75t_R FILLER_220_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_838 ();
 DECAPx4_ASAP7_75t_R FILLER_220_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_864 ();
 DECAPx2_ASAP7_75t_R FILLER_220_886 ();
 FILLER_ASAP7_75t_R FILLER_220_892 ();
 FILLER_ASAP7_75t_R FILLER_220_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_912 ();
 DECAPx10_ASAP7_75t_R FILLER_220_934 ();
 DECAPx4_ASAP7_75t_R FILLER_220_956 ();
 FILLER_ASAP7_75t_R FILLER_220_966 ();
 FILLER_ASAP7_75t_R FILLER_220_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1018 ();
 FILLER_ASAP7_75t_R FILLER_220_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1182 ();
 FILLER_ASAP7_75t_R FILLER_220_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1190 ();
 FILLER_ASAP7_75t_R FILLER_220_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1232 ();
 FILLER_ASAP7_75t_R FILLER_220_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1240 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1269 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1283 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1308 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1385 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1394 ();
 DECAPx10_ASAP7_75t_R FILLER_221_2 ();
 DECAPx10_ASAP7_75t_R FILLER_221_24 ();
 DECAPx10_ASAP7_75t_R FILLER_221_46 ();
 DECAPx10_ASAP7_75t_R FILLER_221_68 ();
 DECAPx2_ASAP7_75t_R FILLER_221_90 ();
 FILLER_ASAP7_75t_R FILLER_221_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_101 ();
 DECAPx10_ASAP7_75t_R FILLER_221_105 ();
 DECAPx2_ASAP7_75t_R FILLER_221_127 ();
 FILLER_ASAP7_75t_R FILLER_221_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_141 ();
 DECAPx6_ASAP7_75t_R FILLER_221_145 ();
 DECAPx2_ASAP7_75t_R FILLER_221_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_191 ();
 DECAPx2_ASAP7_75t_R FILLER_221_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_209 ();
 DECAPx1_ASAP7_75t_R FILLER_221_222 ();
 DECAPx4_ASAP7_75t_R FILLER_221_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_242 ();
 DECAPx4_ASAP7_75t_R FILLER_221_249 ();
 FILLER_ASAP7_75t_R FILLER_221_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_261 ();
 DECAPx4_ASAP7_75t_R FILLER_221_268 ();
 FILLER_ASAP7_75t_R FILLER_221_278 ();
 DECAPx1_ASAP7_75t_R FILLER_221_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_312 ();
 FILLER_ASAP7_75t_R FILLER_221_345 ();
 DECAPx6_ASAP7_75t_R FILLER_221_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_380 ();
 DECAPx6_ASAP7_75t_R FILLER_221_387 ();
 DECAPx2_ASAP7_75t_R FILLER_221_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_407 ();
 DECAPx4_ASAP7_75t_R FILLER_221_417 ();
 FILLER_ASAP7_75t_R FILLER_221_427 ();
 DECAPx4_ASAP7_75t_R FILLER_221_435 ();
 FILLER_ASAP7_75t_R FILLER_221_445 ();
 DECAPx4_ASAP7_75t_R FILLER_221_453 ();
 FILLER_ASAP7_75t_R FILLER_221_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_465 ();
 DECAPx2_ASAP7_75t_R FILLER_221_480 ();
 FILLER_ASAP7_75t_R FILLER_221_486 ();
 DECAPx2_ASAP7_75t_R FILLER_221_562 ();
 DECAPx2_ASAP7_75t_R FILLER_221_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_589 ();
 DECAPx6_ASAP7_75t_R FILLER_221_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_622 ();
 DECAPx10_ASAP7_75t_R FILLER_221_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_653 ();
 FILLER_ASAP7_75t_R FILLER_221_660 ();
 DECAPx4_ASAP7_75t_R FILLER_221_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_685 ();
 DECAPx6_ASAP7_75t_R FILLER_221_694 ();
 DECAPx2_ASAP7_75t_R FILLER_221_708 ();
 DECAPx1_ASAP7_75t_R FILLER_221_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_745 ();
 DECAPx1_ASAP7_75t_R FILLER_221_754 ();
 DECAPx6_ASAP7_75t_R FILLER_221_770 ();
 FILLER_ASAP7_75t_R FILLER_221_784 ();
 DECAPx6_ASAP7_75t_R FILLER_221_792 ();
 FILLER_ASAP7_75t_R FILLER_221_812 ();
 FILLER_ASAP7_75t_R FILLER_221_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_837 ();
 DECAPx1_ASAP7_75t_R FILLER_221_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_917 ();
 FILLER_ASAP7_75t_R FILLER_221_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_947 ();
 FILLER_ASAP7_75t_R FILLER_221_952 ();
 FILLER_ASAP7_75t_R FILLER_221_963 ();
 DECAPx2_ASAP7_75t_R FILLER_221_985 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1005 ();
 FILLER_ASAP7_75t_R FILLER_221_1012 ();
 FILLER_ASAP7_75t_R FILLER_221_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1116 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1146 ();
 FILLER_ASAP7_75t_R FILLER_221_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1157 ();
 FILLER_ASAP7_75t_R FILLER_221_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1181 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1213 ();
 FILLER_ASAP7_75t_R FILLER_221_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1286 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1313 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1331 ();
 FILLER_ASAP7_75t_R FILLER_221_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_222_2 ();
 DECAPx10_ASAP7_75t_R FILLER_222_24 ();
 DECAPx10_ASAP7_75t_R FILLER_222_46 ();
 DECAPx10_ASAP7_75t_R FILLER_222_68 ();
 DECAPx10_ASAP7_75t_R FILLER_222_90 ();
 DECAPx1_ASAP7_75t_R FILLER_222_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_116 ();
 DECAPx2_ASAP7_75t_R FILLER_222_143 ();
 DECAPx4_ASAP7_75t_R FILLER_222_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_172 ();
 FILLER_ASAP7_75t_R FILLER_222_176 ();
 DECAPx10_ASAP7_75t_R FILLER_222_210 ();
 DECAPx10_ASAP7_75t_R FILLER_222_232 ();
 DECAPx6_ASAP7_75t_R FILLER_222_254 ();
 FILLER_ASAP7_75t_R FILLER_222_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_270 ();
 DECAPx2_ASAP7_75t_R FILLER_222_292 ();
 DECAPx4_ASAP7_75t_R FILLER_222_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_318 ();
 FILLER_ASAP7_75t_R FILLER_222_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_330 ();
 DECAPx2_ASAP7_75t_R FILLER_222_389 ();
 DECAPx6_ASAP7_75t_R FILLER_222_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_461 ();
 DECAPx6_ASAP7_75t_R FILLER_222_464 ();
 DECAPx1_ASAP7_75t_R FILLER_222_478 ();
 DECAPx10_ASAP7_75t_R FILLER_222_488 ();
 DECAPx10_ASAP7_75t_R FILLER_222_510 ();
 DECAPx10_ASAP7_75t_R FILLER_222_532 ();
 FILLER_ASAP7_75t_R FILLER_222_560 ();
 DECAPx10_ASAP7_75t_R FILLER_222_568 ();
 DECAPx10_ASAP7_75t_R FILLER_222_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_625 ();
 FILLER_ASAP7_75t_R FILLER_222_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_642 ();
 DECAPx1_ASAP7_75t_R FILLER_222_659 ();
 FILLER_ASAP7_75t_R FILLER_222_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_673 ();
 DECAPx2_ASAP7_75t_R FILLER_222_718 ();
 FILLER_ASAP7_75t_R FILLER_222_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_726 ();
 DECAPx10_ASAP7_75t_R FILLER_222_735 ();
 DECAPx1_ASAP7_75t_R FILLER_222_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_761 ();
 DECAPx4_ASAP7_75t_R FILLER_222_770 ();
 FILLER_ASAP7_75t_R FILLER_222_780 ();
 DECAPx6_ASAP7_75t_R FILLER_222_804 ();
 DECAPx6_ASAP7_75t_R FILLER_222_824 ();
 DECAPx2_ASAP7_75t_R FILLER_222_838 ();
 DECAPx2_ASAP7_75t_R FILLER_222_873 ();
 DECAPx4_ASAP7_75t_R FILLER_222_912 ();
 FILLER_ASAP7_75t_R FILLER_222_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_924 ();
 FILLER_ASAP7_75t_R FILLER_222_938 ();
 FILLER_ASAP7_75t_R FILLER_222_980 ();
 DECAPx1_ASAP7_75t_R FILLER_222_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_999 ();
 FILLER_ASAP7_75t_R FILLER_222_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1040 ();
 FILLER_ASAP7_75t_R FILLER_222_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_222_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_222_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1181 ();
 FILLER_ASAP7_75t_R FILLER_222_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1234 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1277 ();
 FILLER_ASAP7_75t_R FILLER_222_1285 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1293 ();
 FILLER_ASAP7_75t_R FILLER_222_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1352 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1356 ();
 FILLER_ASAP7_75t_R FILLER_222_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1385 ();
 FILLER_ASAP7_75t_R FILLER_222_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_223_2 ();
 DECAPx10_ASAP7_75t_R FILLER_223_24 ();
 DECAPx10_ASAP7_75t_R FILLER_223_46 ();
 DECAPx10_ASAP7_75t_R FILLER_223_68 ();
 DECAPx10_ASAP7_75t_R FILLER_223_90 ();
 DECAPx6_ASAP7_75t_R FILLER_223_112 ();
 FILLER_ASAP7_75t_R FILLER_223_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_128 ();
 DECAPx2_ASAP7_75t_R FILLER_223_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_145 ();
 DECAPx6_ASAP7_75t_R FILLER_223_172 ();
 DECAPx2_ASAP7_75t_R FILLER_223_186 ();
 DECAPx4_ASAP7_75t_R FILLER_223_201 ();
 FILLER_ASAP7_75t_R FILLER_223_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_239 ();
 FILLER_ASAP7_75t_R FILLER_223_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_249 ();
 DECAPx1_ASAP7_75t_R FILLER_223_253 ();
 DECAPx10_ASAP7_75t_R FILLER_223_270 ();
 DECAPx10_ASAP7_75t_R FILLER_223_292 ();
 DECAPx6_ASAP7_75t_R FILLER_223_314 ();
 DECAPx2_ASAP7_75t_R FILLER_223_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_334 ();
 DECAPx1_ASAP7_75t_R FILLER_223_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_348 ();
 FILLER_ASAP7_75t_R FILLER_223_375 ();
 DECAPx2_ASAP7_75t_R FILLER_223_380 ();
 FILLER_ASAP7_75t_R FILLER_223_386 ();
 DECAPx4_ASAP7_75t_R FILLER_223_395 ();
 DECAPx6_ASAP7_75t_R FILLER_223_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_425 ();
 DECAPx1_ASAP7_75t_R FILLER_223_432 ();
 DECAPx1_ASAP7_75t_R FILLER_223_439 ();
 DECAPx4_ASAP7_75t_R FILLER_223_469 ();
 FILLER_ASAP7_75t_R FILLER_223_479 ();
 FILLER_ASAP7_75t_R FILLER_223_488 ();
 DECAPx6_ASAP7_75t_R FILLER_223_499 ();
 FILLER_ASAP7_75t_R FILLER_223_513 ();
 DECAPx10_ASAP7_75t_R FILLER_223_522 ();
 DECAPx2_ASAP7_75t_R FILLER_223_544 ();
 FILLER_ASAP7_75t_R FILLER_223_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_552 ();
 FILLER_ASAP7_75t_R FILLER_223_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_569 ();
 DECAPx4_ASAP7_75t_R FILLER_223_590 ();
 DECAPx6_ASAP7_75t_R FILLER_223_607 ();
 DECAPx2_ASAP7_75t_R FILLER_223_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_639 ();
 DECAPx4_ASAP7_75t_R FILLER_223_649 ();
 FILLER_ASAP7_75t_R FILLER_223_666 ();
 DECAPx10_ASAP7_75t_R FILLER_223_674 ();
 DECAPx10_ASAP7_75t_R FILLER_223_696 ();
 FILLER_ASAP7_75t_R FILLER_223_724 ();
 DECAPx6_ASAP7_75t_R FILLER_223_744 ();
 FILLER_ASAP7_75t_R FILLER_223_758 ();
 FILLER_ASAP7_75t_R FILLER_223_774 ();
 DECAPx2_ASAP7_75t_R FILLER_223_799 ();
 FILLER_ASAP7_75t_R FILLER_223_805 ();
 DECAPx6_ASAP7_75t_R FILLER_223_821 ();
 FILLER_ASAP7_75t_R FILLER_223_835 ();
 DECAPx10_ASAP7_75t_R FILLER_223_843 ();
 DECAPx6_ASAP7_75t_R FILLER_223_865 ();
 DECAPx1_ASAP7_75t_R FILLER_223_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_883 ();
 DECAPx6_ASAP7_75t_R FILLER_223_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_904 ();
 FILLER_ASAP7_75t_R FILLER_223_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_914 ();
 DECAPx1_ASAP7_75t_R FILLER_223_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_923 ();
 DECAPx6_ASAP7_75t_R FILLER_223_926 ();
 FILLER_ASAP7_75t_R FILLER_223_940 ();
 DECAPx2_ASAP7_75t_R FILLER_223_948 ();
 DECAPx1_ASAP7_75t_R FILLER_223_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_964 ();
 DECAPx4_ASAP7_75t_R FILLER_223_985 ();
 FILLER_ASAP7_75t_R FILLER_223_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_997 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_223_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1063 ();
 FILLER_ASAP7_75t_R FILLER_223_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1071 ();
 FILLER_ASAP7_75t_R FILLER_223_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1181 ();
 FILLER_ASAP7_75t_R FILLER_223_1187 ();
 FILLER_ASAP7_75t_R FILLER_223_1219 ();
 FILLER_ASAP7_75t_R FILLER_223_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1270 ();
 DECAPx4_ASAP7_75t_R FILLER_223_1300 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1349 ();
 DECAPx10_ASAP7_75t_R FILLER_224_2 ();
 DECAPx10_ASAP7_75t_R FILLER_224_24 ();
 DECAPx10_ASAP7_75t_R FILLER_224_46 ();
 DECAPx10_ASAP7_75t_R FILLER_224_68 ();
 DECAPx10_ASAP7_75t_R FILLER_224_90 ();
 DECAPx10_ASAP7_75t_R FILLER_224_112 ();
 DECAPx4_ASAP7_75t_R FILLER_224_134 ();
 FILLER_ASAP7_75t_R FILLER_224_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_159 ();
 DECAPx2_ASAP7_75t_R FILLER_224_163 ();
 FILLER_ASAP7_75t_R FILLER_224_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_171 ();
 FILLER_ASAP7_75t_R FILLER_224_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_184 ();
 FILLER_ASAP7_75t_R FILLER_224_188 ();
 FILLER_ASAP7_75t_R FILLER_224_223 ();
 DECAPx6_ASAP7_75t_R FILLER_224_283 ();
 DECAPx2_ASAP7_75t_R FILLER_224_304 ();
 FILLER_ASAP7_75t_R FILLER_224_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_312 ();
 DECAPx2_ASAP7_75t_R FILLER_224_345 ();
 FILLER_ASAP7_75t_R FILLER_224_351 ();
 DECAPx1_ASAP7_75t_R FILLER_224_359 ();
 DECAPx6_ASAP7_75t_R FILLER_224_366 ();
 FILLER_ASAP7_75t_R FILLER_224_380 ();
 DECAPx2_ASAP7_75t_R FILLER_224_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_420 ();
 DECAPx4_ASAP7_75t_R FILLER_224_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_470 ();
 FILLER_ASAP7_75t_R FILLER_224_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_479 ();
 DECAPx2_ASAP7_75t_R FILLER_224_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_512 ();
 DECAPx2_ASAP7_75t_R FILLER_224_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_545 ();
 DECAPx6_ASAP7_75t_R FILLER_224_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_572 ();
 DECAPx2_ASAP7_75t_R FILLER_224_583 ();
 FILLER_ASAP7_75t_R FILLER_224_607 ();
 DECAPx2_ASAP7_75t_R FILLER_224_628 ();
 FILLER_ASAP7_75t_R FILLER_224_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_636 ();
 DECAPx1_ASAP7_75t_R FILLER_224_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_655 ();
 DECAPx1_ASAP7_75t_R FILLER_224_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_689 ();
 DECAPx2_ASAP7_75t_R FILLER_224_696 ();
 FILLER_ASAP7_75t_R FILLER_224_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_704 ();
 FILLER_ASAP7_75t_R FILLER_224_717 ();
 DECAPx1_ASAP7_75t_R FILLER_224_727 ();
 DECAPx4_ASAP7_75t_R FILLER_224_743 ();
 DECAPx6_ASAP7_75t_R FILLER_224_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_806 ();
 FILLER_ASAP7_75t_R FILLER_224_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_824 ();
 DECAPx1_ASAP7_75t_R FILLER_224_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_836 ();
 DECAPx2_ASAP7_75t_R FILLER_224_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_850 ();
 DECAPx2_ASAP7_75t_R FILLER_224_858 ();
 DECAPx6_ASAP7_75t_R FILLER_224_883 ();
 FILLER_ASAP7_75t_R FILLER_224_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_904 ();
 FILLER_ASAP7_75t_R FILLER_224_932 ();
 DECAPx6_ASAP7_75t_R FILLER_224_937 ();
 DECAPx2_ASAP7_75t_R FILLER_224_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_957 ();
 DECAPx4_ASAP7_75t_R FILLER_224_961 ();
 FILLER_ASAP7_75t_R FILLER_224_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_977 ();
 DECAPx2_ASAP7_75t_R FILLER_224_986 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1028 ();
 FILLER_ASAP7_75t_R FILLER_224_1034 ();
 FILLER_ASAP7_75t_R FILLER_224_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1145 ();
 FILLER_ASAP7_75t_R FILLER_224_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1246 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1265 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1276 ();
 FILLER_ASAP7_75t_R FILLER_224_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1314 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1328 ();
 FILLER_ASAP7_75t_R FILLER_224_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1380 ();
 FILLER_ASAP7_75t_R FILLER_224_1398 ();
 DECAPx10_ASAP7_75t_R FILLER_225_2 ();
 DECAPx10_ASAP7_75t_R FILLER_225_24 ();
 DECAPx10_ASAP7_75t_R FILLER_225_46 ();
 DECAPx10_ASAP7_75t_R FILLER_225_68 ();
 DECAPx10_ASAP7_75t_R FILLER_225_90 ();
 DECAPx10_ASAP7_75t_R FILLER_225_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_134 ();
 FILLER_ASAP7_75t_R FILLER_225_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_170 ();
 DECAPx1_ASAP7_75t_R FILLER_225_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_207 ();
 FILLER_ASAP7_75t_R FILLER_225_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_230 ();
 DECAPx6_ASAP7_75t_R FILLER_225_238 ();
 DECAPx2_ASAP7_75t_R FILLER_225_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_258 ();
 FILLER_ASAP7_75t_R FILLER_225_265 ();
 DECAPx1_ASAP7_75t_R FILLER_225_285 ();
 DECAPx2_ASAP7_75t_R FILLER_225_321 ();
 DECAPx10_ASAP7_75t_R FILLER_225_330 ();
 DECAPx2_ASAP7_75t_R FILLER_225_352 ();
 FILLER_ASAP7_75t_R FILLER_225_374 ();
 DECAPx1_ASAP7_75t_R FILLER_225_382 ();
 DECAPx6_ASAP7_75t_R FILLER_225_444 ();
 FILLER_ASAP7_75t_R FILLER_225_458 ();
 DECAPx1_ASAP7_75t_R FILLER_225_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_516 ();
 DECAPx1_ASAP7_75t_R FILLER_225_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_527 ();
 DECAPx10_ASAP7_75t_R FILLER_225_531 ();
 DECAPx10_ASAP7_75t_R FILLER_225_553 ();
 DECAPx10_ASAP7_75t_R FILLER_225_575 ();
 DECAPx10_ASAP7_75t_R FILLER_225_597 ();
 DECAPx4_ASAP7_75t_R FILLER_225_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_645 ();
 DECAPx10_ASAP7_75t_R FILLER_225_652 ();
 DECAPx2_ASAP7_75t_R FILLER_225_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_680 ();
 DECAPx1_ASAP7_75t_R FILLER_225_702 ();
 FILLER_ASAP7_75t_R FILLER_225_728 ();
 DECAPx2_ASAP7_75t_R FILLER_225_744 ();
 FILLER_ASAP7_75t_R FILLER_225_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_752 ();
 FILLER_ASAP7_75t_R FILLER_225_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_767 ();
 DECAPx1_ASAP7_75t_R FILLER_225_782 ();
 DECAPx2_ASAP7_75t_R FILLER_225_792 ();
 FILLER_ASAP7_75t_R FILLER_225_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_904 ();
 DECAPx4_ASAP7_75t_R FILLER_225_911 ();
 FILLER_ASAP7_75t_R FILLER_225_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_929 ();
 FILLER_ASAP7_75t_R FILLER_225_936 ();
 FILLER_ASAP7_75t_R FILLER_225_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_962 ();
 DECAPx4_ASAP7_75t_R FILLER_225_970 ();
 FILLER_ASAP7_75t_R FILLER_225_980 ();
 FILLER_ASAP7_75t_R FILLER_225_1021 ();
 FILLER_ASAP7_75t_R FILLER_225_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1065 ();
 FILLER_ASAP7_75t_R FILLER_225_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1085 ();
 FILLER_ASAP7_75t_R FILLER_225_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1178 ();
 FILLER_ASAP7_75t_R FILLER_225_1206 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1218 ();
 FILLER_ASAP7_75t_R FILLER_225_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1259 ();
 FILLER_ASAP7_75t_R FILLER_225_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1283 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1290 ();
 FILLER_ASAP7_75t_R FILLER_225_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1298 ();
 FILLER_ASAP7_75t_R FILLER_225_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_226_2 ();
 DECAPx10_ASAP7_75t_R FILLER_226_24 ();
 DECAPx10_ASAP7_75t_R FILLER_226_46 ();
 DECAPx10_ASAP7_75t_R FILLER_226_68 ();
 DECAPx10_ASAP7_75t_R FILLER_226_90 ();
 DECAPx10_ASAP7_75t_R FILLER_226_112 ();
 DECAPx2_ASAP7_75t_R FILLER_226_134 ();
 FILLER_ASAP7_75t_R FILLER_226_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_142 ();
 DECAPx1_ASAP7_75t_R FILLER_226_169 ();
 DECAPx6_ASAP7_75t_R FILLER_226_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_223 ();
 DECAPx1_ASAP7_75t_R FILLER_226_227 ();
 DECAPx4_ASAP7_75t_R FILLER_226_238 ();
 DECAPx4_ASAP7_75t_R FILLER_226_274 ();
 FILLER_ASAP7_75t_R FILLER_226_284 ();
 DECAPx1_ASAP7_75t_R FILLER_226_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_308 ();
 DECAPx4_ASAP7_75t_R FILLER_226_312 ();
 DECAPx2_ASAP7_75t_R FILLER_226_329 ();
 DECAPx2_ASAP7_75t_R FILLER_226_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_354 ();
 DECAPx1_ASAP7_75t_R FILLER_226_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_392 ();
 FILLER_ASAP7_75t_R FILLER_226_400 ();
 DECAPx1_ASAP7_75t_R FILLER_226_405 ();
 DECAPx10_ASAP7_75t_R FILLER_226_412 ();
 DECAPx2_ASAP7_75t_R FILLER_226_434 ();
 FILLER_ASAP7_75t_R FILLER_226_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_442 ();
 FILLER_ASAP7_75t_R FILLER_226_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_458 ();
 DECAPx4_ASAP7_75t_R FILLER_226_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_474 ();
 DECAPx4_ASAP7_75t_R FILLER_226_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_488 ();
 DECAPx2_ASAP7_75t_R FILLER_226_496 ();
 FILLER_ASAP7_75t_R FILLER_226_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_504 ();
 DECAPx10_ASAP7_75t_R FILLER_226_508 ();
 DECAPx4_ASAP7_75t_R FILLER_226_530 ();
 FILLER_ASAP7_75t_R FILLER_226_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_542 ();
 DECAPx4_ASAP7_75t_R FILLER_226_549 ();
 FILLER_ASAP7_75t_R FILLER_226_559 ();
 DECAPx6_ASAP7_75t_R FILLER_226_567 ();
 DECAPx1_ASAP7_75t_R FILLER_226_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_585 ();
 DECAPx2_ASAP7_75t_R FILLER_226_589 ();
 FILLER_ASAP7_75t_R FILLER_226_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_597 ();
 DECAPx1_ASAP7_75t_R FILLER_226_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_617 ();
 DECAPx2_ASAP7_75t_R FILLER_226_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_638 ();
 DECAPx1_ASAP7_75t_R FILLER_226_659 ();
 DECAPx10_ASAP7_75t_R FILLER_226_676 ();
 DECAPx6_ASAP7_75t_R FILLER_226_698 ();
 DECAPx1_ASAP7_75t_R FILLER_226_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_716 ();
 FILLER_ASAP7_75t_R FILLER_226_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_731 ();
 DECAPx10_ASAP7_75t_R FILLER_226_738 ();
 DECAPx2_ASAP7_75t_R FILLER_226_775 ();
 FILLER_ASAP7_75t_R FILLER_226_781 ();
 DECAPx2_ASAP7_75t_R FILLER_226_797 ();
 FILLER_ASAP7_75t_R FILLER_226_803 ();
 DECAPx10_ASAP7_75t_R FILLER_226_826 ();
 DECAPx1_ASAP7_75t_R FILLER_226_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_852 ();
 DECAPx2_ASAP7_75t_R FILLER_226_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_865 ();
 FILLER_ASAP7_75t_R FILLER_226_883 ();
 DECAPx10_ASAP7_75t_R FILLER_226_895 ();
 DECAPx4_ASAP7_75t_R FILLER_226_917 ();
 FILLER_ASAP7_75t_R FILLER_226_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_929 ();
 FILLER_ASAP7_75t_R FILLER_226_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_940 ();
 FILLER_ASAP7_75t_R FILLER_226_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_964 ();
 DECAPx6_ASAP7_75t_R FILLER_226_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1000 ();
 FILLER_ASAP7_75t_R FILLER_226_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1053 ();
 FILLER_ASAP7_75t_R FILLER_226_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1069 ();
 FILLER_ASAP7_75t_R FILLER_226_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1158 ();
 FILLER_ASAP7_75t_R FILLER_226_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1176 ();
 FILLER_ASAP7_75t_R FILLER_226_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1272 ();
 FILLER_ASAP7_75t_R FILLER_226_1281 ();
 FILLER_ASAP7_75t_R FILLER_226_1290 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1356 ();
 FILLER_ASAP7_75t_R FILLER_226_1365 ();
 FILLER_ASAP7_75t_R FILLER_226_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_227_2 ();
 DECAPx10_ASAP7_75t_R FILLER_227_24 ();
 DECAPx10_ASAP7_75t_R FILLER_227_46 ();
 DECAPx10_ASAP7_75t_R FILLER_227_68 ();
 DECAPx10_ASAP7_75t_R FILLER_227_90 ();
 DECAPx10_ASAP7_75t_R FILLER_227_112 ();
 DECAPx4_ASAP7_75t_R FILLER_227_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_144 ();
 DECAPx2_ASAP7_75t_R FILLER_227_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_157 ();
 FILLER_ASAP7_75t_R FILLER_227_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_166 ();
 DECAPx2_ASAP7_75t_R FILLER_227_199 ();
 FILLER_ASAP7_75t_R FILLER_227_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_207 ();
 DECAPx1_ASAP7_75t_R FILLER_227_222 ();
 DECAPx4_ASAP7_75t_R FILLER_227_252 ();
 DECAPx6_ASAP7_75t_R FILLER_227_265 ();
 DECAPx1_ASAP7_75t_R FILLER_227_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_283 ();
 DECAPx1_ASAP7_75t_R FILLER_227_310 ();
 DECAPx1_ASAP7_75t_R FILLER_227_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_370 ();
 DECAPx6_ASAP7_75t_R FILLER_227_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_411 ();
 DECAPx2_ASAP7_75t_R FILLER_227_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_426 ();
 DECAPx1_ASAP7_75t_R FILLER_227_430 ();
 DECAPx2_ASAP7_75t_R FILLER_227_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_443 ();
 DECAPx6_ASAP7_75t_R FILLER_227_470 ();
 DECAPx1_ASAP7_75t_R FILLER_227_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_488 ();
 DECAPx10_ASAP7_75t_R FILLER_227_495 ();
 DECAPx10_ASAP7_75t_R FILLER_227_517 ();
 FILLER_ASAP7_75t_R FILLER_227_539 ();
 FILLER_ASAP7_75t_R FILLER_227_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_550 ();
 FILLER_ASAP7_75t_R FILLER_227_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_567 ();
 FILLER_ASAP7_75t_R FILLER_227_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_618 ();
 DECAPx6_ASAP7_75t_R FILLER_227_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_646 ();
 FILLER_ASAP7_75t_R FILLER_227_653 ();
 DECAPx6_ASAP7_75t_R FILLER_227_687 ();
 FILLER_ASAP7_75t_R FILLER_227_701 ();
 DECAPx2_ASAP7_75t_R FILLER_227_717 ();
 FILLER_ASAP7_75t_R FILLER_227_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_725 ();
 DECAPx2_ASAP7_75t_R FILLER_227_740 ();
 FILLER_ASAP7_75t_R FILLER_227_746 ();
 DECAPx10_ASAP7_75t_R FILLER_227_756 ();
 DECAPx1_ASAP7_75t_R FILLER_227_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_782 ();
 DECAPx6_ASAP7_75t_R FILLER_227_792 ();
 FILLER_ASAP7_75t_R FILLER_227_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_815 ();
 DECAPx10_ASAP7_75t_R FILLER_227_822 ();
 DECAPx10_ASAP7_75t_R FILLER_227_844 ();
 DECAPx10_ASAP7_75t_R FILLER_227_866 ();
 FILLER_ASAP7_75t_R FILLER_227_888 ();
 FILLER_ASAP7_75t_R FILLER_227_904 ();
 DECAPx2_ASAP7_75t_R FILLER_227_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_923 ();
 FILLER_ASAP7_75t_R FILLER_227_938 ();
 DECAPx4_ASAP7_75t_R FILLER_227_947 ();
 FILLER_ASAP7_75t_R FILLER_227_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_963 ();
 DECAPx2_ASAP7_75t_R FILLER_227_977 ();
 DECAPx2_ASAP7_75t_R FILLER_227_995 ();
 FILLER_ASAP7_75t_R FILLER_227_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1037 ();
 FILLER_ASAP7_75t_R FILLER_227_1043 ();
 FILLER_ASAP7_75t_R FILLER_227_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_227_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_227_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1179 ();
 FILLER_ASAP7_75t_R FILLER_227_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_227_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1268 ();
 FILLER_ASAP7_75t_R FILLER_227_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1308 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_228_2 ();
 DECAPx10_ASAP7_75t_R FILLER_228_24 ();
 DECAPx10_ASAP7_75t_R FILLER_228_46 ();
 DECAPx10_ASAP7_75t_R FILLER_228_68 ();
 DECAPx10_ASAP7_75t_R FILLER_228_90 ();
 DECAPx10_ASAP7_75t_R FILLER_228_112 ();
 DECAPx10_ASAP7_75t_R FILLER_228_134 ();
 DECAPx6_ASAP7_75t_R FILLER_228_156 ();
 FILLER_ASAP7_75t_R FILLER_228_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_172 ();
 FILLER_ASAP7_75t_R FILLER_228_178 ();
 DECAPx4_ASAP7_75t_R FILLER_228_186 ();
 DECAPx6_ASAP7_75t_R FILLER_228_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_236 ();
 DECAPx10_ASAP7_75t_R FILLER_228_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_280 ();
 DECAPx1_ASAP7_75t_R FILLER_228_287 ();
 DECAPx1_ASAP7_75t_R FILLER_228_329 ();
 DECAPx2_ASAP7_75t_R FILLER_228_336 ();
 FILLER_ASAP7_75t_R FILLER_228_342 ();
 DECAPx1_ASAP7_75t_R FILLER_228_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_354 ();
 DECAPx10_ASAP7_75t_R FILLER_228_358 ();
 DECAPx1_ASAP7_75t_R FILLER_228_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_384 ();
 DECAPx4_ASAP7_75t_R FILLER_228_388 ();
 FILLER_ASAP7_75t_R FILLER_228_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_411 ();
 DECAPx2_ASAP7_75t_R FILLER_228_438 ();
 FILLER_ASAP7_75t_R FILLER_228_444 ();
 DECAPx4_ASAP7_75t_R FILLER_228_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_522 ();
 DECAPx4_ASAP7_75t_R FILLER_228_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_542 ();
 DECAPx10_ASAP7_75t_R FILLER_228_555 ();
 DECAPx2_ASAP7_75t_R FILLER_228_577 ();
 DECAPx10_ASAP7_75t_R FILLER_228_589 ();
 DECAPx10_ASAP7_75t_R FILLER_228_611 ();
 DECAPx1_ASAP7_75t_R FILLER_228_633 ();
 DECAPx2_ASAP7_75t_R FILLER_228_649 ();
 FILLER_ASAP7_75t_R FILLER_228_655 ();
 DECAPx1_ASAP7_75t_R FILLER_228_664 ();
 DECAPx4_ASAP7_75t_R FILLER_228_674 ();
 FILLER_ASAP7_75t_R FILLER_228_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_686 ();
 FILLER_ASAP7_75t_R FILLER_228_695 ();
 DECAPx1_ASAP7_75t_R FILLER_228_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_766 ();
 DECAPx2_ASAP7_75t_R FILLER_228_774 ();
 FILLER_ASAP7_75t_R FILLER_228_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_782 ();
 DECAPx1_ASAP7_75t_R FILLER_228_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_801 ();
 FILLER_ASAP7_75t_R FILLER_228_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_817 ();
 DECAPx2_ASAP7_75t_R FILLER_228_828 ();
 DECAPx10_ASAP7_75t_R FILLER_228_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_872 ();
 DECAPx6_ASAP7_75t_R FILLER_228_885 ();
 DECAPx1_ASAP7_75t_R FILLER_228_907 ();
 DECAPx6_ASAP7_75t_R FILLER_228_947 ();
 FILLER_ASAP7_75t_R FILLER_228_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_963 ();
 DECAPx1_ASAP7_75t_R FILLER_228_985 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1001 ();
 FILLER_ASAP7_75t_R FILLER_228_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1078 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_228_1122 ();
 FILLER_ASAP7_75t_R FILLER_228_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1153 ();
 FILLER_ASAP7_75t_R FILLER_228_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1203 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1239 ();
 FILLER_ASAP7_75t_R FILLER_228_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1300 ();
 FILLER_ASAP7_75t_R FILLER_228_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1331 ();
 FILLER_ASAP7_75t_R FILLER_228_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1385 ();
 FILLER_ASAP7_75t_R FILLER_228_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_229_2 ();
 DECAPx10_ASAP7_75t_R FILLER_229_24 ();
 DECAPx10_ASAP7_75t_R FILLER_229_46 ();
 DECAPx10_ASAP7_75t_R FILLER_229_68 ();
 DECAPx10_ASAP7_75t_R FILLER_229_90 ();
 DECAPx10_ASAP7_75t_R FILLER_229_112 ();
 DECAPx10_ASAP7_75t_R FILLER_229_134 ();
 FILLER_ASAP7_75t_R FILLER_229_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_158 ();
 DECAPx2_ASAP7_75t_R FILLER_229_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_171 ();
 DECAPx1_ASAP7_75t_R FILLER_229_179 ();
 DECAPx4_ASAP7_75t_R FILLER_229_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_228 ();
 FILLER_ASAP7_75t_R FILLER_229_255 ();
 DECAPx1_ASAP7_75t_R FILLER_229_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_294 ();
 DECAPx1_ASAP7_75t_R FILLER_229_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_309 ();
 DECAPx4_ASAP7_75t_R FILLER_229_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_346 ();
 DECAPx2_ASAP7_75t_R FILLER_229_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_360 ();
 DECAPx2_ASAP7_75t_R FILLER_229_370 ();
 FILLER_ASAP7_75t_R FILLER_229_441 ();
 DECAPx1_ASAP7_75t_R FILLER_229_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_507 ();
 DECAPx10_ASAP7_75t_R FILLER_229_534 ();
 DECAPx10_ASAP7_75t_R FILLER_229_556 ();
 DECAPx10_ASAP7_75t_R FILLER_229_578 ();
 FILLER_ASAP7_75t_R FILLER_229_600 ();
 DECAPx2_ASAP7_75t_R FILLER_229_616 ();
 FILLER_ASAP7_75t_R FILLER_229_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_624 ();
 DECAPx2_ASAP7_75t_R FILLER_229_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_637 ();
 DECAPx1_ASAP7_75t_R FILLER_229_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_649 ();
 DECAPx4_ASAP7_75t_R FILLER_229_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_674 ();
 DECAPx6_ASAP7_75t_R FILLER_229_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_697 ();
 FILLER_ASAP7_75t_R FILLER_229_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_730 ();
 DECAPx4_ASAP7_75t_R FILLER_229_740 ();
 FILLER_ASAP7_75t_R FILLER_229_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_752 ();
 FILLER_ASAP7_75t_R FILLER_229_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_809 ();
 DECAPx2_ASAP7_75t_R FILLER_229_826 ();
 FILLER_ASAP7_75t_R FILLER_229_832 ();
 DECAPx1_ASAP7_75t_R FILLER_229_855 ();
 DECAPx4_ASAP7_75t_R FILLER_229_880 ();
 DECAPx4_ASAP7_75t_R FILLER_229_914 ();
 DECAPx10_ASAP7_75t_R FILLER_229_940 ();
 DECAPx2_ASAP7_75t_R FILLER_229_962 ();
 FILLER_ASAP7_75t_R FILLER_229_968 ();
 DECAPx6_ASAP7_75t_R FILLER_229_976 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1064 ();
 FILLER_ASAP7_75t_R FILLER_229_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1080 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1182 ();
 FILLER_ASAP7_75t_R FILLER_229_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1204 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1301 ();
 FILLER_ASAP7_75t_R FILLER_229_1321 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1349 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1363 ();
 DECAPx10_ASAP7_75t_R FILLER_230_2 ();
 DECAPx10_ASAP7_75t_R FILLER_230_24 ();
 DECAPx10_ASAP7_75t_R FILLER_230_46 ();
 DECAPx10_ASAP7_75t_R FILLER_230_68 ();
 DECAPx10_ASAP7_75t_R FILLER_230_90 ();
 DECAPx10_ASAP7_75t_R FILLER_230_112 ();
 DECAPx6_ASAP7_75t_R FILLER_230_134 ();
 DECAPx2_ASAP7_75t_R FILLER_230_148 ();
 DECAPx1_ASAP7_75t_R FILLER_230_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_165 ();
 DECAPx1_ASAP7_75t_R FILLER_230_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_196 ();
 DECAPx6_ASAP7_75t_R FILLER_230_200 ();
 DECAPx1_ASAP7_75t_R FILLER_230_214 ();
 FILLER_ASAP7_75t_R FILLER_230_244 ();
 DECAPx10_ASAP7_75t_R FILLER_230_282 ();
 DECAPx4_ASAP7_75t_R FILLER_230_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_314 ();
 FILLER_ASAP7_75t_R FILLER_230_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_324 ();
 FILLER_ASAP7_75t_R FILLER_230_340 ();
 FILLER_ASAP7_75t_R FILLER_230_368 ();
 FILLER_ASAP7_75t_R FILLER_230_396 ();
 FILLER_ASAP7_75t_R FILLER_230_404 ();
 DECAPx2_ASAP7_75t_R FILLER_230_409 ();
 FILLER_ASAP7_75t_R FILLER_230_415 ();
 DECAPx4_ASAP7_75t_R FILLER_230_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_456 ();
 FILLER_ASAP7_75t_R FILLER_230_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_470 ();
 DECAPx6_ASAP7_75t_R FILLER_230_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_495 ();
 DECAPx2_ASAP7_75t_R FILLER_230_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_505 ();
 DECAPx6_ASAP7_75t_R FILLER_230_522 ();
 FILLER_ASAP7_75t_R FILLER_230_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_538 ();
 DECAPx6_ASAP7_75t_R FILLER_230_545 ();
 FILLER_ASAP7_75t_R FILLER_230_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_561 ();
 DECAPx2_ASAP7_75t_R FILLER_230_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_581 ();
 FILLER_ASAP7_75t_R FILLER_230_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_598 ();
 DECAPx6_ASAP7_75t_R FILLER_230_606 ();
 DECAPx1_ASAP7_75t_R FILLER_230_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_624 ();
 DECAPx2_ASAP7_75t_R FILLER_230_643 ();
 FILLER_ASAP7_75t_R FILLER_230_649 ();
 DECAPx1_ASAP7_75t_R FILLER_230_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_671 ();
 DECAPx6_ASAP7_75t_R FILLER_230_675 ();
 DECAPx2_ASAP7_75t_R FILLER_230_689 ();
 DECAPx2_ASAP7_75t_R FILLER_230_715 ();
 FILLER_ASAP7_75t_R FILLER_230_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_723 ();
 DECAPx1_ASAP7_75t_R FILLER_230_744 ();
 DECAPx4_ASAP7_75t_R FILLER_230_770 ();
 FILLER_ASAP7_75t_R FILLER_230_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_782 ();
 DECAPx1_ASAP7_75t_R FILLER_230_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_797 ();
 DECAPx1_ASAP7_75t_R FILLER_230_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_851 ();
 DECAPx1_ASAP7_75t_R FILLER_230_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_900 ();
 DECAPx6_ASAP7_75t_R FILLER_230_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_921 ();
 DECAPx2_ASAP7_75t_R FILLER_230_936 ();
 DECAPx4_ASAP7_75t_R FILLER_230_970 ();
 FILLER_ASAP7_75t_R FILLER_230_980 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1073 ();
 FILLER_ASAP7_75t_R FILLER_230_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_230_1150 ();
 FILLER_ASAP7_75t_R FILLER_230_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1199 ();
 FILLER_ASAP7_75t_R FILLER_230_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1336 ();
 FILLER_ASAP7_75t_R FILLER_230_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_231_2 ();
 DECAPx10_ASAP7_75t_R FILLER_231_24 ();
 DECAPx10_ASAP7_75t_R FILLER_231_46 ();
 DECAPx10_ASAP7_75t_R FILLER_231_68 ();
 DECAPx10_ASAP7_75t_R FILLER_231_90 ();
 DECAPx10_ASAP7_75t_R FILLER_231_112 ();
 DECAPx6_ASAP7_75t_R FILLER_231_134 ();
 DECAPx1_ASAP7_75t_R FILLER_231_148 ();
 FILLER_ASAP7_75t_R FILLER_231_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_180 ();
 DECAPx2_ASAP7_75t_R FILLER_231_184 ();
 FILLER_ASAP7_75t_R FILLER_231_190 ();
 DECAPx1_ASAP7_75t_R FILLER_231_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_212 ();
 DECAPx1_ASAP7_75t_R FILLER_231_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_243 ();
 DECAPx4_ASAP7_75t_R FILLER_231_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_267 ();
 FILLER_ASAP7_75t_R FILLER_231_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_273 ();
 DECAPx10_ASAP7_75t_R FILLER_231_280 ();
 DECAPx6_ASAP7_75t_R FILLER_231_302 ();
 DECAPx1_ASAP7_75t_R FILLER_231_316 ();
 FILLER_ASAP7_75t_R FILLER_231_346 ();
 FILLER_ASAP7_75t_R FILLER_231_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_362 ();
 FILLER_ASAP7_75t_R FILLER_231_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_368 ();
 DECAPx4_ASAP7_75t_R FILLER_231_414 ();
 FILLER_ASAP7_75t_R FILLER_231_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_426 ();
 DECAPx2_ASAP7_75t_R FILLER_231_492 ();
 FILLER_ASAP7_75t_R FILLER_231_498 ();
 DECAPx2_ASAP7_75t_R FILLER_231_513 ();
 FILLER_ASAP7_75t_R FILLER_231_519 ();
 DECAPx4_ASAP7_75t_R FILLER_231_524 ();
 FILLER_ASAP7_75t_R FILLER_231_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_556 ();
 DECAPx6_ASAP7_75t_R FILLER_231_578 ();
 DECAPx1_ASAP7_75t_R FILLER_231_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_603 ();
 DECAPx6_ASAP7_75t_R FILLER_231_610 ();
 FILLER_ASAP7_75t_R FILLER_231_624 ();
 FILLER_ASAP7_75t_R FILLER_231_635 ();
 DECAPx1_ASAP7_75t_R FILLER_231_652 ();
 FILLER_ASAP7_75t_R FILLER_231_662 ();
 DECAPx1_ASAP7_75t_R FILLER_231_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_678 ();
 DECAPx4_ASAP7_75t_R FILLER_231_695 ();
 DECAPx4_ASAP7_75t_R FILLER_231_717 ();
 FILLER_ASAP7_75t_R FILLER_231_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_754 ();
 FILLER_ASAP7_75t_R FILLER_231_758 ();
 DECAPx6_ASAP7_75t_R FILLER_231_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_780 ();
 DECAPx2_ASAP7_75t_R FILLER_231_789 ();
 FILLER_ASAP7_75t_R FILLER_231_795 ();
 FILLER_ASAP7_75t_R FILLER_231_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_812 ();
 DECAPx6_ASAP7_75t_R FILLER_231_819 ();
 FILLER_ASAP7_75t_R FILLER_231_833 ();
 DECAPx2_ASAP7_75t_R FILLER_231_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_862 ();
 FILLER_ASAP7_75t_R FILLER_231_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_880 ();
 DECAPx6_ASAP7_75t_R FILLER_231_901 ();
 FILLER_ASAP7_75t_R FILLER_231_915 ();
 DECAPx1_ASAP7_75t_R FILLER_231_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_938 ();
 FILLER_ASAP7_75t_R FILLER_231_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_970 ();
 FILLER_ASAP7_75t_R FILLER_231_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_991 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1030 ();
 FILLER_ASAP7_75t_R FILLER_231_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1065 ();
 FILLER_ASAP7_75t_R FILLER_231_1071 ();
 FILLER_ASAP7_75t_R FILLER_231_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1097 ();
 FILLER_ASAP7_75t_R FILLER_231_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1149 ();
 FILLER_ASAP7_75t_R FILLER_231_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1278 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1300 ();
 FILLER_ASAP7_75t_R FILLER_231_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1365 ();
 DECAPx10_ASAP7_75t_R FILLER_232_2 ();
 DECAPx10_ASAP7_75t_R FILLER_232_24 ();
 DECAPx10_ASAP7_75t_R FILLER_232_46 ();
 DECAPx10_ASAP7_75t_R FILLER_232_68 ();
 DECAPx10_ASAP7_75t_R FILLER_232_90 ();
 DECAPx10_ASAP7_75t_R FILLER_232_112 ();
 DECAPx10_ASAP7_75t_R FILLER_232_134 ();
 DECAPx4_ASAP7_75t_R FILLER_232_156 ();
 DECAPx1_ASAP7_75t_R FILLER_232_169 ();
 DECAPx1_ASAP7_75t_R FILLER_232_180 ();
 DECAPx2_ASAP7_75t_R FILLER_232_219 ();
 FILLER_ASAP7_75t_R FILLER_232_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_227 ();
 DECAPx6_ASAP7_75t_R FILLER_232_231 ();
 DECAPx1_ASAP7_75t_R FILLER_232_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_301 ();
 DECAPx2_ASAP7_75t_R FILLER_232_305 ();
 DECAPx2_ASAP7_75t_R FILLER_232_326 ();
 FILLER_ASAP7_75t_R FILLER_232_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_334 ();
 DECAPx1_ASAP7_75t_R FILLER_232_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_342 ();
 FILLER_ASAP7_75t_R FILLER_232_375 ();
 DECAPx4_ASAP7_75t_R FILLER_232_423 ();
 FILLER_ASAP7_75t_R FILLER_232_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_435 ();
 DECAPx1_ASAP7_75t_R FILLER_232_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_495 ();
 DECAPx10_ASAP7_75t_R FILLER_232_532 ();
 DECAPx2_ASAP7_75t_R FILLER_232_554 ();
 FILLER_ASAP7_75t_R FILLER_232_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_562 ();
 DECAPx2_ASAP7_75t_R FILLER_232_573 ();
 FILLER_ASAP7_75t_R FILLER_232_579 ();
 DECAPx6_ASAP7_75t_R FILLER_232_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_601 ();
 DECAPx1_ASAP7_75t_R FILLER_232_626 ();
 DECAPx4_ASAP7_75t_R FILLER_232_637 ();
 FILLER_ASAP7_75t_R FILLER_232_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_674 ();
 DECAPx4_ASAP7_75t_R FILLER_232_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_707 ();
 DECAPx6_ASAP7_75t_R FILLER_232_718 ();
 FILLER_ASAP7_75t_R FILLER_232_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_772 ();
 FILLER_ASAP7_75t_R FILLER_232_779 ();
 DECAPx4_ASAP7_75t_R FILLER_232_791 ();
 FILLER_ASAP7_75t_R FILLER_232_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_803 ();
 DECAPx10_ASAP7_75t_R FILLER_232_820 ();
 DECAPx10_ASAP7_75t_R FILLER_232_842 ();
 DECAPx2_ASAP7_75t_R FILLER_232_864 ();
 DECAPx1_ASAP7_75t_R FILLER_232_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_878 ();
 FILLER_ASAP7_75t_R FILLER_232_903 ();
 DECAPx4_ASAP7_75t_R FILLER_232_911 ();
 FILLER_ASAP7_75t_R FILLER_232_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_923 ();
 FILLER_ASAP7_75t_R FILLER_232_936 ();
 DECAPx6_ASAP7_75t_R FILLER_232_964 ();
 DECAPx2_ASAP7_75t_R FILLER_232_978 ();
 DECAPx6_ASAP7_75t_R FILLER_232_990 ();
 FILLER_ASAP7_75t_R FILLER_232_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1023 ();
 FILLER_ASAP7_75t_R FILLER_232_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1098 ();
 FILLER_ASAP7_75t_R FILLER_232_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1171 ();
 FILLER_ASAP7_75t_R FILLER_232_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1252 ();
 FILLER_ASAP7_75t_R FILLER_232_1258 ();
 FILLER_ASAP7_75t_R FILLER_232_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1265 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1284 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1305 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1336 ();
 FILLER_ASAP7_75t_R FILLER_232_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1365 ();
 FILLER_ASAP7_75t_R FILLER_232_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1385 ();
 FILLER_ASAP7_75t_R FILLER_232_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_233_2 ();
 DECAPx10_ASAP7_75t_R FILLER_233_24 ();
 DECAPx10_ASAP7_75t_R FILLER_233_46 ();
 DECAPx10_ASAP7_75t_R FILLER_233_68 ();
 DECAPx10_ASAP7_75t_R FILLER_233_90 ();
 DECAPx10_ASAP7_75t_R FILLER_233_112 ();
 DECAPx10_ASAP7_75t_R FILLER_233_134 ();
 DECAPx4_ASAP7_75t_R FILLER_233_156 ();
 FILLER_ASAP7_75t_R FILLER_233_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_168 ();
 DECAPx2_ASAP7_75t_R FILLER_233_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_201 ();
 DECAPx2_ASAP7_75t_R FILLER_233_205 ();
 FILLER_ASAP7_75t_R FILLER_233_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_213 ();
 DECAPx2_ASAP7_75t_R FILLER_233_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_227 ();
 DECAPx4_ASAP7_75t_R FILLER_233_267 ();
 DECAPx1_ASAP7_75t_R FILLER_233_284 ();
 FILLER_ASAP7_75t_R FILLER_233_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_316 ();
 DECAPx6_ASAP7_75t_R FILLER_233_332 ();
 DECAPx1_ASAP7_75t_R FILLER_233_346 ();
 DECAPx1_ASAP7_75t_R FILLER_233_357 ();
 DECAPx2_ASAP7_75t_R FILLER_233_364 ();
 FILLER_ASAP7_75t_R FILLER_233_370 ();
 DECAPx6_ASAP7_75t_R FILLER_233_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_453 ();
 FILLER_ASAP7_75t_R FILLER_233_480 ();
 DECAPx1_ASAP7_75t_R FILLER_233_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_495 ();
 DECAPx2_ASAP7_75t_R FILLER_233_532 ();
 FILLER_ASAP7_75t_R FILLER_233_538 ();
 DECAPx6_ASAP7_75t_R FILLER_233_549 ();
 FILLER_ASAP7_75t_R FILLER_233_577 ();
 FILLER_ASAP7_75t_R FILLER_233_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_589 ();
 DECAPx10_ASAP7_75t_R FILLER_233_596 ();
 DECAPx6_ASAP7_75t_R FILLER_233_618 ();
 DECAPx4_ASAP7_75t_R FILLER_233_638 ();
 FILLER_ASAP7_75t_R FILLER_233_648 ();
 DECAPx1_ASAP7_75t_R FILLER_233_668 ();
 DECAPx10_ASAP7_75t_R FILLER_233_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_700 ();
 FILLER_ASAP7_75t_R FILLER_233_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_732 ();
 FILLER_ASAP7_75t_R FILLER_233_763 ();
 DECAPx1_ASAP7_75t_R FILLER_233_777 ();
 DECAPx4_ASAP7_75t_R FILLER_233_791 ();
 FILLER_ASAP7_75t_R FILLER_233_801 ();
 DECAPx4_ASAP7_75t_R FILLER_233_821 ();
 DECAPx4_ASAP7_75t_R FILLER_233_839 ();
 FILLER_ASAP7_75t_R FILLER_233_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_851 ();
 DECAPx4_ASAP7_75t_R FILLER_233_855 ();
 FILLER_ASAP7_75t_R FILLER_233_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_867 ();
 FILLER_ASAP7_75t_R FILLER_233_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_892 ();
 DECAPx10_ASAP7_75t_R FILLER_233_926 ();
 DECAPx1_ASAP7_75t_R FILLER_233_948 ();
 FILLER_ASAP7_75t_R FILLER_233_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_957 ();
 DECAPx1_ASAP7_75t_R FILLER_233_986 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1043 ();
 FILLER_ASAP7_75t_R FILLER_233_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1072 ();
 FILLER_ASAP7_75t_R FILLER_233_1078 ();
 FILLER_ASAP7_75t_R FILLER_233_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1169 ();
 FILLER_ASAP7_75t_R FILLER_233_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1187 ();
 FILLER_ASAP7_75t_R FILLER_233_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1234 ();
 FILLER_ASAP7_75t_R FILLER_233_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1248 ();
 FILLER_ASAP7_75t_R FILLER_233_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1325 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1347 ();
 FILLER_ASAP7_75t_R FILLER_233_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1363 ();
 DECAPx10_ASAP7_75t_R FILLER_234_2 ();
 DECAPx10_ASAP7_75t_R FILLER_234_24 ();
 DECAPx10_ASAP7_75t_R FILLER_234_46 ();
 DECAPx10_ASAP7_75t_R FILLER_234_68 ();
 DECAPx10_ASAP7_75t_R FILLER_234_90 ();
 DECAPx10_ASAP7_75t_R FILLER_234_112 ();
 DECAPx10_ASAP7_75t_R FILLER_234_134 ();
 DECAPx10_ASAP7_75t_R FILLER_234_156 ();
 DECAPx4_ASAP7_75t_R FILLER_234_178 ();
 FILLER_ASAP7_75t_R FILLER_234_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_203 ();
 DECAPx2_ASAP7_75t_R FILLER_234_207 ();
 DECAPx6_ASAP7_75t_R FILLER_234_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_280 ();
 FILLER_ASAP7_75t_R FILLER_234_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_289 ();
 DECAPx4_ASAP7_75t_R FILLER_234_293 ();
 FILLER_ASAP7_75t_R FILLER_234_303 ();
 DECAPx2_ASAP7_75t_R FILLER_234_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_337 ();
 FILLER_ASAP7_75t_R FILLER_234_344 ();
 DECAPx2_ASAP7_75t_R FILLER_234_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_407 ();
 DECAPx1_ASAP7_75t_R FILLER_234_411 ();
 DECAPx2_ASAP7_75t_R FILLER_234_421 ();
 FILLER_ASAP7_75t_R FILLER_234_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_429 ();
 DECAPx4_ASAP7_75t_R FILLER_234_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_443 ();
 DECAPx1_ASAP7_75t_R FILLER_234_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_461 ();
 DECAPx2_ASAP7_75t_R FILLER_234_473 ();
 FILLER_ASAP7_75t_R FILLER_234_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_481 ();
 DECAPx1_ASAP7_75t_R FILLER_234_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_538 ();
 DECAPx1_ASAP7_75t_R FILLER_234_559 ();
 DECAPx6_ASAP7_75t_R FILLER_234_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_587 ();
 DECAPx6_ASAP7_75t_R FILLER_234_596 ();
 DECAPx1_ASAP7_75t_R FILLER_234_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_614 ();
 DECAPx6_ASAP7_75t_R FILLER_234_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_636 ();
 DECAPx10_ASAP7_75t_R FILLER_234_643 ();
 DECAPx2_ASAP7_75t_R FILLER_234_665 ();
 FILLER_ASAP7_75t_R FILLER_234_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_673 ();
 FILLER_ASAP7_75t_R FILLER_234_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_682 ();
 DECAPx6_ASAP7_75t_R FILLER_234_691 ();
 FILLER_ASAP7_75t_R FILLER_234_705 ();
 FILLER_ASAP7_75t_R FILLER_234_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_724 ();
 DECAPx1_ASAP7_75t_R FILLER_234_737 ();
 DECAPx2_ASAP7_75t_R FILLER_234_773 ();
 FILLER_ASAP7_75t_R FILLER_234_779 ();
 DECAPx2_ASAP7_75t_R FILLER_234_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_805 ();
 DECAPx4_ASAP7_75t_R FILLER_234_818 ();
 DECAPx1_ASAP7_75t_R FILLER_234_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_846 ();
 FILLER_ASAP7_75t_R FILLER_234_898 ();
 DECAPx4_ASAP7_75t_R FILLER_234_907 ();
 DECAPx10_ASAP7_75t_R FILLER_234_921 ();
 DECAPx6_ASAP7_75t_R FILLER_234_943 ();
 DECAPx1_ASAP7_75t_R FILLER_234_957 ();
 DECAPx4_ASAP7_75t_R FILLER_234_967 ();
 FILLER_ASAP7_75t_R FILLER_234_977 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1031 ();
 FILLER_ASAP7_75t_R FILLER_234_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1087 ();
 FILLER_ASAP7_75t_R FILLER_234_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1108 ();
 FILLER_ASAP7_75t_R FILLER_234_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1342 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1380 ();
 FILLER_ASAP7_75t_R FILLER_234_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_235_2 ();
 DECAPx10_ASAP7_75t_R FILLER_235_24 ();
 DECAPx10_ASAP7_75t_R FILLER_235_46 ();
 DECAPx10_ASAP7_75t_R FILLER_235_68 ();
 DECAPx10_ASAP7_75t_R FILLER_235_90 ();
 DECAPx10_ASAP7_75t_R FILLER_235_112 ();
 DECAPx10_ASAP7_75t_R FILLER_235_134 ();
 DECAPx10_ASAP7_75t_R FILLER_235_156 ();
 DECAPx4_ASAP7_75t_R FILLER_235_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_215 ();
 FILLER_ASAP7_75t_R FILLER_235_222 ();
 DECAPx4_ASAP7_75t_R FILLER_235_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_263 ();
 DECAPx6_ASAP7_75t_R FILLER_235_303 ();
 FILLER_ASAP7_75t_R FILLER_235_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_319 ();
 FILLER_ASAP7_75t_R FILLER_235_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_325 ();
 FILLER_ASAP7_75t_R FILLER_235_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_345 ();
 FILLER_ASAP7_75t_R FILLER_235_383 ();
 FILLER_ASAP7_75t_R FILLER_235_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_399 ();
 DECAPx6_ASAP7_75t_R FILLER_235_407 ();
 DECAPx6_ASAP7_75t_R FILLER_235_434 ();
 FILLER_ASAP7_75t_R FILLER_235_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_450 ();
 DECAPx10_ASAP7_75t_R FILLER_235_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_494 ();
 DECAPx2_ASAP7_75t_R FILLER_235_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_510 ();
 DECAPx1_ASAP7_75t_R FILLER_235_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_521 ();
 DECAPx10_ASAP7_75t_R FILLER_235_525 ();
 DECAPx6_ASAP7_75t_R FILLER_235_547 ();
 DECAPx2_ASAP7_75t_R FILLER_235_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_567 ();
 DECAPx1_ASAP7_75t_R FILLER_235_574 ();
 DECAPx2_ASAP7_75t_R FILLER_235_594 ();
 FILLER_ASAP7_75t_R FILLER_235_600 ();
 DECAPx6_ASAP7_75t_R FILLER_235_610 ();
 DECAPx1_ASAP7_75t_R FILLER_235_624 ();
 DECAPx1_ASAP7_75t_R FILLER_235_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_647 ();
 DECAPx1_ASAP7_75t_R FILLER_235_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_705 ();
 DECAPx10_ASAP7_75t_R FILLER_235_736 ();
 DECAPx2_ASAP7_75t_R FILLER_235_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_764 ();
 DECAPx4_ASAP7_75t_R FILLER_235_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_785 ();
 DECAPx2_ASAP7_75t_R FILLER_235_795 ();
 DECAPx4_ASAP7_75t_R FILLER_235_821 ();
 FILLER_ASAP7_75t_R FILLER_235_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_844 ();
 FILLER_ASAP7_75t_R FILLER_235_889 ();
 DECAPx1_ASAP7_75t_R FILLER_235_897 ();
 FILLER_ASAP7_75t_R FILLER_235_922 ();
 FILLER_ASAP7_75t_R FILLER_235_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_928 ();
 DECAPx4_ASAP7_75t_R FILLER_235_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_945 ();
 FILLER_ASAP7_75t_R FILLER_235_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_956 ();
 DECAPx4_ASAP7_75t_R FILLER_235_967 ();
 FILLER_ASAP7_75t_R FILLER_235_977 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1013 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1050 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1141 ();
 FILLER_ASAP7_75t_R FILLER_235_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1189 ();
 FILLER_ASAP7_75t_R FILLER_235_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1224 ();
 FILLER_ASAP7_75t_R FILLER_235_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1304 ();
 FILLER_ASAP7_75t_R FILLER_235_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_236_2 ();
 DECAPx10_ASAP7_75t_R FILLER_236_24 ();
 DECAPx10_ASAP7_75t_R FILLER_236_46 ();
 DECAPx10_ASAP7_75t_R FILLER_236_68 ();
 DECAPx10_ASAP7_75t_R FILLER_236_90 ();
 DECAPx10_ASAP7_75t_R FILLER_236_112 ();
 DECAPx10_ASAP7_75t_R FILLER_236_134 ();
 DECAPx10_ASAP7_75t_R FILLER_236_156 ();
 DECAPx10_ASAP7_75t_R FILLER_236_178 ();
 DECAPx10_ASAP7_75t_R FILLER_236_200 ();
 DECAPx6_ASAP7_75t_R FILLER_236_222 ();
 DECAPx1_ASAP7_75t_R FILLER_236_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_240 ();
 FILLER_ASAP7_75t_R FILLER_236_276 ();
 DECAPx4_ASAP7_75t_R FILLER_236_310 ();
 DECAPx1_ASAP7_75t_R FILLER_236_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_461 ();
 FILLER_ASAP7_75t_R FILLER_236_464 ();
 FILLER_ASAP7_75t_R FILLER_236_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_471 ();
 DECAPx2_ASAP7_75t_R FILLER_236_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_481 ();
 DECAPx10_ASAP7_75t_R FILLER_236_514 ();
 DECAPx1_ASAP7_75t_R FILLER_236_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_540 ();
 DECAPx1_ASAP7_75t_R FILLER_236_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_559 ();
 DECAPx6_ASAP7_75t_R FILLER_236_567 ();
 DECAPx2_ASAP7_75t_R FILLER_236_581 ();
 DECAPx10_ASAP7_75t_R FILLER_236_597 ();
 DECAPx4_ASAP7_75t_R FILLER_236_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_629 ();
 DECAPx4_ASAP7_75t_R FILLER_236_636 ();
 FILLER_ASAP7_75t_R FILLER_236_652 ();
 DECAPx1_ASAP7_75t_R FILLER_236_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_672 ();
 DECAPx10_ASAP7_75t_R FILLER_236_685 ();
 DECAPx10_ASAP7_75t_R FILLER_236_707 ();
 DECAPx1_ASAP7_75t_R FILLER_236_729 ();
 FILLER_ASAP7_75t_R FILLER_236_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_738 ();
 DECAPx1_ASAP7_75t_R FILLER_236_749 ();
 DECAPx10_ASAP7_75t_R FILLER_236_756 ();
 FILLER_ASAP7_75t_R FILLER_236_778 ();
 DECAPx1_ASAP7_75t_R FILLER_236_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_790 ();
 DECAPx4_ASAP7_75t_R FILLER_236_799 ();
 FILLER_ASAP7_75t_R FILLER_236_809 ();
 DECAPx4_ASAP7_75t_R FILLER_236_814 ();
 FILLER_ASAP7_75t_R FILLER_236_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_826 ();
 DECAPx1_ASAP7_75t_R FILLER_236_830 ();
 DECAPx2_ASAP7_75t_R FILLER_236_842 ();
 FILLER_ASAP7_75t_R FILLER_236_848 ();
 DECAPx4_ASAP7_75t_R FILLER_236_863 ();
 FILLER_ASAP7_75t_R FILLER_236_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1002 ();
 FILLER_ASAP7_75t_R FILLER_236_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1063 ();
 FILLER_ASAP7_75t_R FILLER_236_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_236_1104 ();
 FILLER_ASAP7_75t_R FILLER_236_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1167 ();
 FILLER_ASAP7_75t_R FILLER_236_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_236_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1205 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1269 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1305 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1326 ();
 FILLER_ASAP7_75t_R FILLER_236_1330 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1338 ();
 FILLER_ASAP7_75t_R FILLER_236_1352 ();
 FILLER_ASAP7_75t_R FILLER_236_1364 ();
 FILLER_ASAP7_75t_R FILLER_236_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_237_2 ();
 DECAPx10_ASAP7_75t_R FILLER_237_24 ();
 DECAPx10_ASAP7_75t_R FILLER_237_46 ();
 DECAPx10_ASAP7_75t_R FILLER_237_68 ();
 DECAPx10_ASAP7_75t_R FILLER_237_90 ();
 DECAPx10_ASAP7_75t_R FILLER_237_112 ();
 DECAPx10_ASAP7_75t_R FILLER_237_134 ();
 DECAPx10_ASAP7_75t_R FILLER_237_156 ();
 DECAPx10_ASAP7_75t_R FILLER_237_178 ();
 DECAPx10_ASAP7_75t_R FILLER_237_200 ();
 DECAPx10_ASAP7_75t_R FILLER_237_222 ();
 DECAPx4_ASAP7_75t_R FILLER_237_244 ();
 FILLER_ASAP7_75t_R FILLER_237_254 ();
 DECAPx2_ASAP7_75t_R FILLER_237_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_265 ();
 DECAPx2_ASAP7_75t_R FILLER_237_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_288 ();
 DECAPx10_ASAP7_75t_R FILLER_237_347 ();
 DECAPx1_ASAP7_75t_R FILLER_237_369 ();
 DECAPx2_ASAP7_75t_R FILLER_237_376 ();
 DECAPx2_ASAP7_75t_R FILLER_237_408 ();
 DECAPx4_ASAP7_75t_R FILLER_237_417 ();
 FILLER_ASAP7_75t_R FILLER_237_433 ();
 DECAPx6_ASAP7_75t_R FILLER_237_531 ();
 FILLER_ASAP7_75t_R FILLER_237_545 ();
 DECAPx6_ASAP7_75t_R FILLER_237_556 ();
 FILLER_ASAP7_75t_R FILLER_237_570 ();
 DECAPx4_ASAP7_75t_R FILLER_237_595 ();
 DECAPx10_ASAP7_75t_R FILLER_237_621 ();
 DECAPx10_ASAP7_75t_R FILLER_237_651 ();
 FILLER_ASAP7_75t_R FILLER_237_673 ();
 DECAPx2_ASAP7_75t_R FILLER_237_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_691 ();
 DECAPx2_ASAP7_75t_R FILLER_237_721 ();
 FILLER_ASAP7_75t_R FILLER_237_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_763 ();
 FILLER_ASAP7_75t_R FILLER_237_774 ();
 FILLER_ASAP7_75t_R FILLER_237_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_804 ();
 DECAPx6_ASAP7_75t_R FILLER_237_838 ();
 DECAPx6_ASAP7_75t_R FILLER_237_858 ();
 DECAPx1_ASAP7_75t_R FILLER_237_872 ();
 FILLER_ASAP7_75t_R FILLER_237_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_884 ();
 DECAPx6_ASAP7_75t_R FILLER_237_891 ();
 FILLER_ASAP7_75t_R FILLER_237_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_907 ();
 DECAPx4_ASAP7_75t_R FILLER_237_914 ();
 FILLER_ASAP7_75t_R FILLER_237_926 ();
 FILLER_ASAP7_75t_R FILLER_237_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_944 ();
 FILLER_ASAP7_75t_R FILLER_237_956 ();
 DECAPx1_ASAP7_75t_R FILLER_237_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_990 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1144 ();
 FILLER_ASAP7_75t_R FILLER_237_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1152 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1229 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1251 ();
 FILLER_ASAP7_75t_R FILLER_237_1261 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1304 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1344 ();
 FILLER_ASAP7_75t_R FILLER_237_1361 ();
 DECAPx10_ASAP7_75t_R FILLER_238_2 ();
 DECAPx10_ASAP7_75t_R FILLER_238_24 ();
 DECAPx10_ASAP7_75t_R FILLER_238_46 ();
 DECAPx10_ASAP7_75t_R FILLER_238_68 ();
 DECAPx10_ASAP7_75t_R FILLER_238_90 ();
 DECAPx10_ASAP7_75t_R FILLER_238_112 ();
 DECAPx10_ASAP7_75t_R FILLER_238_134 ();
 DECAPx10_ASAP7_75t_R FILLER_238_156 ();
 DECAPx10_ASAP7_75t_R FILLER_238_178 ();
 DECAPx10_ASAP7_75t_R FILLER_238_200 ();
 DECAPx10_ASAP7_75t_R FILLER_238_222 ();
 FILLER_ASAP7_75t_R FILLER_238_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_246 ();
 DECAPx6_ASAP7_75t_R FILLER_238_285 ();
 FILLER_ASAP7_75t_R FILLER_238_299 ();
 DECAPx10_ASAP7_75t_R FILLER_238_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_335 ();
 DECAPx2_ASAP7_75t_R FILLER_238_339 ();
 DECAPx2_ASAP7_75t_R FILLER_238_351 ();
 DECAPx4_ASAP7_75t_R FILLER_238_360 ();
 DECAPx1_ASAP7_75t_R FILLER_238_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_377 ();
 DECAPx2_ASAP7_75t_R FILLER_238_390 ();
 FILLER_ASAP7_75t_R FILLER_238_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_401 ();
 DECAPx6_ASAP7_75t_R FILLER_238_405 ();
 DECAPx2_ASAP7_75t_R FILLER_238_419 ();
 DECAPx4_ASAP7_75t_R FILLER_238_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_506 ();
 DECAPx2_ASAP7_75t_R FILLER_238_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_519 ();
 DECAPx2_ASAP7_75t_R FILLER_238_523 ();
 FILLER_ASAP7_75t_R FILLER_238_529 ();
 FILLER_ASAP7_75t_R FILLER_238_539 ();
 DECAPx1_ASAP7_75t_R FILLER_238_548 ();
 DECAPx2_ASAP7_75t_R FILLER_238_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_567 ();
 DECAPx6_ASAP7_75t_R FILLER_238_584 ();
 DECAPx1_ASAP7_75t_R FILLER_238_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_602 ();
 DECAPx6_ASAP7_75t_R FILLER_238_611 ();
 DECAPx2_ASAP7_75t_R FILLER_238_625 ();
 DECAPx2_ASAP7_75t_R FILLER_238_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_657 ();
 DECAPx2_ASAP7_75t_R FILLER_238_670 ();
 DECAPx4_ASAP7_75t_R FILLER_238_692 ();
 FILLER_ASAP7_75t_R FILLER_238_702 ();
 DECAPx1_ASAP7_75t_R FILLER_238_730 ();
 DECAPx4_ASAP7_75t_R FILLER_238_740 ();
 FILLER_ASAP7_75t_R FILLER_238_750 ();
 DECAPx4_ASAP7_75t_R FILLER_238_762 ();
 FILLER_ASAP7_75t_R FILLER_238_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_774 ();
 FILLER_ASAP7_75t_R FILLER_238_794 ();
 DECAPx1_ASAP7_75t_R FILLER_238_832 ();
 DECAPx1_ASAP7_75t_R FILLER_238_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_843 ();
 DECAPx6_ASAP7_75t_R FILLER_238_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_874 ();
 DECAPx4_ASAP7_75t_R FILLER_238_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_890 ();
 DECAPx2_ASAP7_75t_R FILLER_238_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_901 ();
 DECAPx4_ASAP7_75t_R FILLER_238_909 ();
 DECAPx2_ASAP7_75t_R FILLER_238_922 ();
 FILLER_ASAP7_75t_R FILLER_238_928 ();
 DECAPx2_ASAP7_75t_R FILLER_238_936 ();
 DECAPx6_ASAP7_75t_R FILLER_238_949 ();
 DECAPx1_ASAP7_75t_R FILLER_238_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_967 ();
 FILLER_ASAP7_75t_R FILLER_238_980 ();
 DECAPx10_ASAP7_75t_R FILLER_238_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1130 ();
 FILLER_ASAP7_75t_R FILLER_238_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1174 ();
 FILLER_ASAP7_75t_R FILLER_238_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1182 ();
 FILLER_ASAP7_75t_R FILLER_238_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1206 ();
 FILLER_ASAP7_75t_R FILLER_238_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1230 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1281 ();
 FILLER_ASAP7_75t_R FILLER_238_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1314 ();
 FILLER_ASAP7_75t_R FILLER_238_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1326 ();
 FILLER_ASAP7_75t_R FILLER_238_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1371 ();
 DECAPx10_ASAP7_75t_R FILLER_239_2 ();
 DECAPx10_ASAP7_75t_R FILLER_239_24 ();
 DECAPx10_ASAP7_75t_R FILLER_239_46 ();
 DECAPx10_ASAP7_75t_R FILLER_239_68 ();
 DECAPx10_ASAP7_75t_R FILLER_239_90 ();
 DECAPx10_ASAP7_75t_R FILLER_239_112 ();
 DECAPx10_ASAP7_75t_R FILLER_239_134 ();
 DECAPx10_ASAP7_75t_R FILLER_239_156 ();
 DECAPx10_ASAP7_75t_R FILLER_239_178 ();
 DECAPx10_ASAP7_75t_R FILLER_239_200 ();
 DECAPx10_ASAP7_75t_R FILLER_239_222 ();
 DECAPx2_ASAP7_75t_R FILLER_239_244 ();
 FILLER_ASAP7_75t_R FILLER_239_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_252 ();
 DECAPx4_ASAP7_75t_R FILLER_239_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_302 ();
 DECAPx10_ASAP7_75t_R FILLER_239_309 ();
 DECAPx4_ASAP7_75t_R FILLER_239_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_341 ();
 FILLER_ASAP7_75t_R FILLER_239_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_370 ();
 DECAPx2_ASAP7_75t_R FILLER_239_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_403 ();
 DECAPx2_ASAP7_75t_R FILLER_239_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_425 ();
 DECAPx2_ASAP7_75t_R FILLER_239_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_438 ();
 DECAPx10_ASAP7_75t_R FILLER_239_442 ();
 DECAPx6_ASAP7_75t_R FILLER_239_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_478 ();
 DECAPx4_ASAP7_75t_R FILLER_239_482 ();
 FILLER_ASAP7_75t_R FILLER_239_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_494 ();
 DECAPx10_ASAP7_75t_R FILLER_239_498 ();
 DECAPx10_ASAP7_75t_R FILLER_239_520 ();
 DECAPx2_ASAP7_75t_R FILLER_239_554 ();
 FILLER_ASAP7_75t_R FILLER_239_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_570 ();
 DECAPx1_ASAP7_75t_R FILLER_239_585 ();
 DECAPx10_ASAP7_75t_R FILLER_239_595 ();
 DECAPx1_ASAP7_75t_R FILLER_239_617 ();
 DECAPx2_ASAP7_75t_R FILLER_239_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_659 ();
 FILLER_ASAP7_75t_R FILLER_239_677 ();
 DECAPx10_ASAP7_75t_R FILLER_239_695 ();
 DECAPx1_ASAP7_75t_R FILLER_239_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_721 ();
 DECAPx6_ASAP7_75t_R FILLER_239_732 ();
 FILLER_ASAP7_75t_R FILLER_239_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_748 ();
 DECAPx2_ASAP7_75t_R FILLER_239_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_771 ();
 DECAPx4_ASAP7_75t_R FILLER_239_778 ();
 DECAPx4_ASAP7_75t_R FILLER_239_794 ();
 DECAPx2_ASAP7_75t_R FILLER_239_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_816 ();
 DECAPx2_ASAP7_75t_R FILLER_239_820 ();
 FILLER_ASAP7_75t_R FILLER_239_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_828 ();
 FILLER_ASAP7_75t_R FILLER_239_842 ();
 DECAPx4_ASAP7_75t_R FILLER_239_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_882 ();
 FILLER_ASAP7_75t_R FILLER_239_895 ();
 DECAPx6_ASAP7_75t_R FILLER_239_932 ();
 FILLER_ASAP7_75t_R FILLER_239_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_948 ();
 DECAPx2_ASAP7_75t_R FILLER_239_961 ();
 DECAPx4_ASAP7_75t_R FILLER_239_973 ();
 FILLER_ASAP7_75t_R FILLER_239_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_985 ();
 FILLER_ASAP7_75t_R FILLER_239_993 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1001 ();
 FILLER_ASAP7_75t_R FILLER_239_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_239_1050 ();
 FILLER_ASAP7_75t_R FILLER_239_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1077 ();
 DECAPx6_ASAP7_75t_R FILLER_239_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1127 ();
 FILLER_ASAP7_75t_R FILLER_239_1133 ();
 FILLER_ASAP7_75t_R FILLER_239_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1182 ();
 FILLER_ASAP7_75t_R FILLER_239_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1190 ();
 FILLER_ASAP7_75t_R FILLER_239_1255 ();
 FILLER_ASAP7_75t_R FILLER_239_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1311 ();
 FILLER_ASAP7_75t_R FILLER_239_1319 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1321 ();
 DECAPx4_ASAP7_75t_R FILLER_239_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1365 ();
 FILLER_ASAP7_75t_R FILLER_239_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1371 ();
 FILLER_ASAP7_75t_R FILLER_239_1377 ();
 DECAPx10_ASAP7_75t_R FILLER_240_2 ();
 DECAPx10_ASAP7_75t_R FILLER_240_24 ();
 DECAPx10_ASAP7_75t_R FILLER_240_46 ();
 DECAPx10_ASAP7_75t_R FILLER_240_68 ();
 DECAPx10_ASAP7_75t_R FILLER_240_90 ();
 DECAPx10_ASAP7_75t_R FILLER_240_112 ();
 DECAPx10_ASAP7_75t_R FILLER_240_134 ();
 DECAPx10_ASAP7_75t_R FILLER_240_156 ();
 DECAPx10_ASAP7_75t_R FILLER_240_178 ();
 DECAPx10_ASAP7_75t_R FILLER_240_200 ();
 DECAPx10_ASAP7_75t_R FILLER_240_222 ();
 DECAPx6_ASAP7_75t_R FILLER_240_244 ();
 FILLER_ASAP7_75t_R FILLER_240_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_260 ();
 FILLER_ASAP7_75t_R FILLER_240_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_270 ();
 DECAPx4_ASAP7_75t_R FILLER_240_277 ();
 FILLER_ASAP7_75t_R FILLER_240_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_289 ();
 DECAPx2_ASAP7_75t_R FILLER_240_316 ();
 DECAPx2_ASAP7_75t_R FILLER_240_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_344 ();
 DECAPx1_ASAP7_75t_R FILLER_240_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_361 ();
 DECAPx6_ASAP7_75t_R FILLER_240_366 ();
 DECAPx1_ASAP7_75t_R FILLER_240_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_384 ();
 DECAPx4_ASAP7_75t_R FILLER_240_388 ();
 DECAPx6_ASAP7_75t_R FILLER_240_427 ();
 FILLER_ASAP7_75t_R FILLER_240_441 ();
 DECAPx1_ASAP7_75t_R FILLER_240_458 ();
 DECAPx10_ASAP7_75t_R FILLER_240_470 ();
 DECAPx10_ASAP7_75t_R FILLER_240_492 ();
 DECAPx6_ASAP7_75t_R FILLER_240_514 ();
 DECAPx1_ASAP7_75t_R FILLER_240_528 ();
 FILLER_ASAP7_75t_R FILLER_240_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_542 ();
 DECAPx4_ASAP7_75t_R FILLER_240_561 ();
 DECAPx1_ASAP7_75t_R FILLER_240_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_582 ();
 DECAPx4_ASAP7_75t_R FILLER_240_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_615 ();
 DECAPx4_ASAP7_75t_R FILLER_240_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_632 ();
 DECAPx1_ASAP7_75t_R FILLER_240_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_643 ();
 FILLER_ASAP7_75t_R FILLER_240_656 ();
 DECAPx2_ASAP7_75t_R FILLER_240_670 ();
 DECAPx6_ASAP7_75t_R FILLER_240_686 ();
 DECAPx2_ASAP7_75t_R FILLER_240_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_716 ();
 DECAPx10_ASAP7_75t_R FILLER_240_767 ();
 DECAPx4_ASAP7_75t_R FILLER_240_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_799 ();
 DECAPx6_ASAP7_75t_R FILLER_240_813 ();
 DECAPx1_ASAP7_75t_R FILLER_240_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_852 ();
 DECAPx2_ASAP7_75t_R FILLER_240_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_905 ();
 DECAPx4_ASAP7_75t_R FILLER_240_919 ();
 DECAPx1_ASAP7_75t_R FILLER_240_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_946 ();
 DECAPx4_ASAP7_75t_R FILLER_240_957 ();
 FILLER_ASAP7_75t_R FILLER_240_967 ();
 DECAPx1_ASAP7_75t_R FILLER_240_982 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1007 ();
 FILLER_ASAP7_75t_R FILLER_240_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1078 ();
 FILLER_ASAP7_75t_R FILLER_240_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1120 ();
 FILLER_ASAP7_75t_R FILLER_240_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1175 ();
 FILLER_ASAP7_75t_R FILLER_240_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1229 ();
 FILLER_ASAP7_75t_R FILLER_240_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1279 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1301 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1337 ();
 FILLER_ASAP7_75t_R FILLER_240_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_241_2 ();
 DECAPx10_ASAP7_75t_R FILLER_241_24 ();
 DECAPx10_ASAP7_75t_R FILLER_241_46 ();
 DECAPx10_ASAP7_75t_R FILLER_241_68 ();
 DECAPx10_ASAP7_75t_R FILLER_241_90 ();
 DECAPx10_ASAP7_75t_R FILLER_241_112 ();
 DECAPx10_ASAP7_75t_R FILLER_241_134 ();
 DECAPx10_ASAP7_75t_R FILLER_241_156 ();
 DECAPx10_ASAP7_75t_R FILLER_241_178 ();
 DECAPx10_ASAP7_75t_R FILLER_241_200 ();
 DECAPx10_ASAP7_75t_R FILLER_241_222 ();
 DECAPx6_ASAP7_75t_R FILLER_241_244 ();
 DECAPx2_ASAP7_75t_R FILLER_241_258 ();
 FILLER_ASAP7_75t_R FILLER_241_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_269 ();
 DECAPx2_ASAP7_75t_R FILLER_241_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_292 ();
 FILLER_ASAP7_75t_R FILLER_241_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_304 ();
 DECAPx2_ASAP7_75t_R FILLER_241_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_366 ();
 FILLER_ASAP7_75t_R FILLER_241_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_384 ();
 FILLER_ASAP7_75t_R FILLER_241_388 ();
 DECAPx4_ASAP7_75t_R FILLER_241_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_404 ();
 FILLER_ASAP7_75t_R FILLER_241_437 ();
 FILLER_ASAP7_75t_R FILLER_241_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_477 ();
 DECAPx10_ASAP7_75t_R FILLER_241_482 ();
 DECAPx10_ASAP7_75t_R FILLER_241_504 ();
 DECAPx2_ASAP7_75t_R FILLER_241_526 ();
 DECAPx1_ASAP7_75t_R FILLER_241_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_560 ();
 DECAPx2_ASAP7_75t_R FILLER_241_569 ();
 DECAPx10_ASAP7_75t_R FILLER_241_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_603 ();
 FILLER_ASAP7_75t_R FILLER_241_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_614 ();
 FILLER_ASAP7_75t_R FILLER_241_623 ();
 FILLER_ASAP7_75t_R FILLER_241_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_639 ();
 DECAPx6_ASAP7_75t_R FILLER_241_656 ();
 DECAPx1_ASAP7_75t_R FILLER_241_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_674 ();
 DECAPx6_ASAP7_75t_R FILLER_241_685 ();
 DECAPx1_ASAP7_75t_R FILLER_241_725 ();
 DECAPx2_ASAP7_75t_R FILLER_241_739 ();
 FILLER_ASAP7_75t_R FILLER_241_745 ();
 DECAPx1_ASAP7_75t_R FILLER_241_760 ();
 DECAPx1_ASAP7_75t_R FILLER_241_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_778 ();
 DECAPx1_ASAP7_75t_R FILLER_241_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_821 ();
 DECAPx10_ASAP7_75t_R FILLER_241_825 ();
 FILLER_ASAP7_75t_R FILLER_241_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_849 ();
 DECAPx10_ASAP7_75t_R FILLER_241_856 ();
 FILLER_ASAP7_75t_R FILLER_241_884 ();
 DECAPx6_ASAP7_75t_R FILLER_241_907 ();
 FILLER_ASAP7_75t_R FILLER_241_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_926 ();
 FILLER_ASAP7_75t_R FILLER_241_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_952 ();
 DECAPx4_ASAP7_75t_R FILLER_241_967 ();
 FILLER_ASAP7_75t_R FILLER_241_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_979 ();
 FILLER_ASAP7_75t_R FILLER_241_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1095 ();
 FILLER_ASAP7_75t_R FILLER_241_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1130 ();
 FILLER_ASAP7_75t_R FILLER_241_1144 ();
 FILLER_ASAP7_75t_R FILLER_241_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_241_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_241_1221 ();
 FILLER_ASAP7_75t_R FILLER_241_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1248 ();
 FILLER_ASAP7_75t_R FILLER_241_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1264 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1285 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1292 ();
 FILLER_ASAP7_75t_R FILLER_241_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1300 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1319 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1328 ();
 FILLER_ASAP7_75t_R FILLER_241_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1370 ();
 FILLER_ASAP7_75t_R FILLER_241_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_242_2 ();
 DECAPx10_ASAP7_75t_R FILLER_242_24 ();
 DECAPx10_ASAP7_75t_R FILLER_242_46 ();
 DECAPx10_ASAP7_75t_R FILLER_242_68 ();
 DECAPx10_ASAP7_75t_R FILLER_242_90 ();
 DECAPx10_ASAP7_75t_R FILLER_242_112 ();
 DECAPx10_ASAP7_75t_R FILLER_242_134 ();
 DECAPx10_ASAP7_75t_R FILLER_242_156 ();
 DECAPx10_ASAP7_75t_R FILLER_242_178 ();
 DECAPx10_ASAP7_75t_R FILLER_242_200 ();
 DECAPx10_ASAP7_75t_R FILLER_242_222 ();
 FILLER_ASAP7_75t_R FILLER_242_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_246 ();
 DECAPx1_ASAP7_75t_R FILLER_242_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_312 ();
 DECAPx4_ASAP7_75t_R FILLER_242_319 ();
 DECAPx6_ASAP7_75t_R FILLER_242_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_346 ();
 FILLER_ASAP7_75t_R FILLER_242_353 ();
 DECAPx2_ASAP7_75t_R FILLER_242_358 ();
 FILLER_ASAP7_75t_R FILLER_242_364 ();
 DECAPx6_ASAP7_75t_R FILLER_242_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_415 ();
 FILLER_ASAP7_75t_R FILLER_242_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_427 ();
 DECAPx6_ASAP7_75t_R FILLER_242_434 ();
 DECAPx1_ASAP7_75t_R FILLER_242_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_452 ();
 DECAPx2_ASAP7_75t_R FILLER_242_456 ();
 DECAPx10_ASAP7_75t_R FILLER_242_490 ();
 DECAPx10_ASAP7_75t_R FILLER_242_512 ();
 DECAPx4_ASAP7_75t_R FILLER_242_534 ();
 DECAPx2_ASAP7_75t_R FILLER_242_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_568 ();
 DECAPx1_ASAP7_75t_R FILLER_242_583 ();
 DECAPx10_ASAP7_75t_R FILLER_242_593 ();
 DECAPx1_ASAP7_75t_R FILLER_242_623 ();
 DECAPx10_ASAP7_75t_R FILLER_242_635 ();
 DECAPx4_ASAP7_75t_R FILLER_242_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_667 ();
 DECAPx2_ASAP7_75t_R FILLER_242_682 ();
 FILLER_ASAP7_75t_R FILLER_242_688 ();
 DECAPx2_ASAP7_75t_R FILLER_242_722 ();
 FILLER_ASAP7_75t_R FILLER_242_734 ();
 DECAPx10_ASAP7_75t_R FILLER_242_739 ();
 DECAPx2_ASAP7_75t_R FILLER_242_761 ();
 FILLER_ASAP7_75t_R FILLER_242_767 ();
 FILLER_ASAP7_75t_R FILLER_242_795 ();
 FILLER_ASAP7_75t_R FILLER_242_803 ();
 FILLER_ASAP7_75t_R FILLER_242_834 ();
 DECAPx2_ASAP7_75t_R FILLER_242_857 ();
 DECAPx2_ASAP7_75t_R FILLER_242_869 ();
 DECAPx4_ASAP7_75t_R FILLER_242_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_904 ();
 DECAPx2_ASAP7_75t_R FILLER_242_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_917 ();
 DECAPx6_ASAP7_75t_R FILLER_242_924 ();
 DECAPx2_ASAP7_75t_R FILLER_242_938 ();
 DECAPx1_ASAP7_75t_R FILLER_242_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_962 ();
 DECAPx10_ASAP7_75t_R FILLER_242_970 ();
 DECAPx6_ASAP7_75t_R FILLER_242_992 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_242_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_242_1158 ();
 FILLER_ASAP7_75t_R FILLER_242_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1174 ();
 FILLER_ASAP7_75t_R FILLER_242_1180 ();
 DECAPx6_ASAP7_75t_R FILLER_242_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1209 ();
 DECAPx6_ASAP7_75t_R FILLER_242_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1254 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1303 ();
 FILLER_ASAP7_75t_R FILLER_242_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1352 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1361 ();
 FILLER_ASAP7_75t_R FILLER_242_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_242_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_243_2 ();
 DECAPx10_ASAP7_75t_R FILLER_243_24 ();
 DECAPx10_ASAP7_75t_R FILLER_243_46 ();
 DECAPx10_ASAP7_75t_R FILLER_243_68 ();
 DECAPx10_ASAP7_75t_R FILLER_243_90 ();
 DECAPx10_ASAP7_75t_R FILLER_243_112 ();
 DECAPx10_ASAP7_75t_R FILLER_243_134 ();
 DECAPx10_ASAP7_75t_R FILLER_243_156 ();
 DECAPx10_ASAP7_75t_R FILLER_243_178 ();
 DECAPx10_ASAP7_75t_R FILLER_243_200 ();
 DECAPx10_ASAP7_75t_R FILLER_243_222 ();
 DECAPx10_ASAP7_75t_R FILLER_243_244 ();
 DECAPx10_ASAP7_75t_R FILLER_243_266 ();
 DECAPx1_ASAP7_75t_R FILLER_243_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_307 ();
 DECAPx4_ASAP7_75t_R FILLER_243_337 ();
 DECAPx1_ASAP7_75t_R FILLER_243_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_357 ();
 DECAPx1_ASAP7_75t_R FILLER_243_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_365 ();
 DECAPx2_ASAP7_75t_R FILLER_243_370 ();
 DECAPx4_ASAP7_75t_R FILLER_243_414 ();
 DECAPx10_ASAP7_75t_R FILLER_243_456 ();
 DECAPx10_ASAP7_75t_R FILLER_243_478 ();
 DECAPx10_ASAP7_75t_R FILLER_243_500 ();
 DECAPx4_ASAP7_75t_R FILLER_243_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_541 ();
 DECAPx6_ASAP7_75t_R FILLER_243_548 ();
 DECAPx1_ASAP7_75t_R FILLER_243_562 ();
 FILLER_ASAP7_75t_R FILLER_243_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_592 ();
 DECAPx2_ASAP7_75t_R FILLER_243_614 ();
 FILLER_ASAP7_75t_R FILLER_243_620 ();
 DECAPx4_ASAP7_75t_R FILLER_243_628 ();
 FILLER_ASAP7_75t_R FILLER_243_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_640 ();
 DECAPx2_ASAP7_75t_R FILLER_243_651 ();
 FILLER_ASAP7_75t_R FILLER_243_657 ();
 DECAPx1_ASAP7_75t_R FILLER_243_673 ();
 DECAPx6_ASAP7_75t_R FILLER_243_690 ();
 DECAPx4_ASAP7_75t_R FILLER_243_707 ();
 FILLER_ASAP7_75t_R FILLER_243_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_725 ();
 DECAPx2_ASAP7_75t_R FILLER_243_733 ();
 FILLER_ASAP7_75t_R FILLER_243_739 ();
 DECAPx6_ASAP7_75t_R FILLER_243_769 ();
 DECAPx2_ASAP7_75t_R FILLER_243_786 ();
 FILLER_ASAP7_75t_R FILLER_243_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_794 ();
 FILLER_ASAP7_75t_R FILLER_243_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_804 ();
 DECAPx10_ASAP7_75t_R FILLER_243_812 ();
 DECAPx2_ASAP7_75t_R FILLER_243_841 ();
 FILLER_ASAP7_75t_R FILLER_243_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_849 ();
 FILLER_ASAP7_75t_R FILLER_243_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_858 ();
 DECAPx2_ASAP7_75t_R FILLER_243_886 ();
 DECAPx1_ASAP7_75t_R FILLER_243_920 ();
 DECAPx1_ASAP7_75t_R FILLER_243_934 ();
 DECAPx1_ASAP7_75t_R FILLER_243_944 ();
 DECAPx2_ASAP7_75t_R FILLER_243_951 ();
 DECAPx2_ASAP7_75t_R FILLER_243_963 ();
 DECAPx4_ASAP7_75t_R FILLER_243_990 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1006 ();
 FILLER_ASAP7_75t_R FILLER_243_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1044 ();
 FILLER_ASAP7_75t_R FILLER_243_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_243_1115 ();
 FILLER_ASAP7_75t_R FILLER_243_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_243_1173 ();
 FILLER_ASAP7_75t_R FILLER_243_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_243_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1262 ();
 FILLER_ASAP7_75t_R FILLER_243_1272 ();
 FILLER_ASAP7_75t_R FILLER_243_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1327 ();
 FILLER_ASAP7_75t_R FILLER_243_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_243_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_244_2 ();
 DECAPx10_ASAP7_75t_R FILLER_244_24 ();
 DECAPx10_ASAP7_75t_R FILLER_244_46 ();
 DECAPx10_ASAP7_75t_R FILLER_244_68 ();
 DECAPx10_ASAP7_75t_R FILLER_244_90 ();
 DECAPx10_ASAP7_75t_R FILLER_244_112 ();
 DECAPx10_ASAP7_75t_R FILLER_244_134 ();
 DECAPx10_ASAP7_75t_R FILLER_244_156 ();
 DECAPx10_ASAP7_75t_R FILLER_244_178 ();
 DECAPx10_ASAP7_75t_R FILLER_244_200 ();
 DECAPx10_ASAP7_75t_R FILLER_244_222 ();
 DECAPx10_ASAP7_75t_R FILLER_244_244 ();
 DECAPx6_ASAP7_75t_R FILLER_244_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_306 ();
 DECAPx6_ASAP7_75t_R FILLER_244_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_342 ();
 DECAPx6_ASAP7_75t_R FILLER_244_369 ();
 FILLER_ASAP7_75t_R FILLER_244_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_385 ();
 FILLER_ASAP7_75t_R FILLER_244_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_435 ();
 DECAPx10_ASAP7_75t_R FILLER_244_467 ();
 DECAPx6_ASAP7_75t_R FILLER_244_489 ();
 DECAPx2_ASAP7_75t_R FILLER_244_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_509 ();
 DECAPx2_ASAP7_75t_R FILLER_244_531 ();
 DECAPx2_ASAP7_75t_R FILLER_244_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_567 ();
 DECAPx1_ASAP7_75t_R FILLER_244_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_580 ();
 DECAPx2_ASAP7_75t_R FILLER_244_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_598 ();
 DECAPx6_ASAP7_75t_R FILLER_244_605 ();
 DECAPx1_ASAP7_75t_R FILLER_244_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_623 ();
 DECAPx6_ASAP7_75t_R FILLER_244_636 ();
 DECAPx1_ASAP7_75t_R FILLER_244_650 ();
 DECAPx1_ASAP7_75t_R FILLER_244_661 ();
 DECAPx4_ASAP7_75t_R FILLER_244_696 ();
 FILLER_ASAP7_75t_R FILLER_244_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_718 ();
 FILLER_ASAP7_75t_R FILLER_244_732 ();
 DECAPx2_ASAP7_75t_R FILLER_244_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_798 ();
 DECAPx2_ASAP7_75t_R FILLER_244_834 ();
 DECAPx1_ASAP7_75t_R FILLER_244_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_847 ();
 FILLER_ASAP7_75t_R FILLER_244_851 ();
 DECAPx1_ASAP7_75t_R FILLER_244_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_866 ();
 DECAPx10_ASAP7_75t_R FILLER_244_873 ();
 DECAPx10_ASAP7_75t_R FILLER_244_895 ();
 DECAPx2_ASAP7_75t_R FILLER_244_917 ();
 DECAPx4_ASAP7_75t_R FILLER_244_987 ();
 FILLER_ASAP7_75t_R FILLER_244_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_999 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1128 ();
 FILLER_ASAP7_75t_R FILLER_244_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_244_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1255 ();
 FILLER_ASAP7_75t_R FILLER_244_1283 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1306 ();
 FILLER_ASAP7_75t_R FILLER_244_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1323 ();
 FILLER_ASAP7_75t_R FILLER_244_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1385 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1401 ();
 DECAPx10_ASAP7_75t_R FILLER_245_2 ();
 DECAPx10_ASAP7_75t_R FILLER_245_24 ();
 DECAPx10_ASAP7_75t_R FILLER_245_46 ();
 DECAPx10_ASAP7_75t_R FILLER_245_68 ();
 DECAPx10_ASAP7_75t_R FILLER_245_90 ();
 DECAPx10_ASAP7_75t_R FILLER_245_112 ();
 DECAPx10_ASAP7_75t_R FILLER_245_134 ();
 DECAPx10_ASAP7_75t_R FILLER_245_156 ();
 DECAPx10_ASAP7_75t_R FILLER_245_178 ();
 DECAPx10_ASAP7_75t_R FILLER_245_200 ();
 DECAPx10_ASAP7_75t_R FILLER_245_222 ();
 DECAPx10_ASAP7_75t_R FILLER_245_244 ();
 DECAPx10_ASAP7_75t_R FILLER_245_266 ();
 DECAPx2_ASAP7_75t_R FILLER_245_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_294 ();
 DECAPx4_ASAP7_75t_R FILLER_245_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_308 ();
 DECAPx2_ASAP7_75t_R FILLER_245_339 ();
 DECAPx1_ASAP7_75t_R FILLER_245_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_371 ();
 DECAPx2_ASAP7_75t_R FILLER_245_384 ();
 FILLER_ASAP7_75t_R FILLER_245_390 ();
 DECAPx2_ASAP7_75t_R FILLER_245_398 ();
 FILLER_ASAP7_75t_R FILLER_245_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_406 ();
 DECAPx2_ASAP7_75t_R FILLER_245_433 ();
 FILLER_ASAP7_75t_R FILLER_245_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_444 ();
 FILLER_ASAP7_75t_R FILLER_245_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_453 ();
 DECAPx10_ASAP7_75t_R FILLER_245_457 ();
 DECAPx10_ASAP7_75t_R FILLER_245_479 ();
 DECAPx4_ASAP7_75t_R FILLER_245_501 ();
 FILLER_ASAP7_75t_R FILLER_245_511 ();
 DECAPx1_ASAP7_75t_R FILLER_245_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_538 ();
 DECAPx2_ASAP7_75t_R FILLER_245_545 ();
 FILLER_ASAP7_75t_R FILLER_245_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_561 ();
 DECAPx10_ASAP7_75t_R FILLER_245_576 ();
 DECAPx6_ASAP7_75t_R FILLER_245_598 ();
 DECAPx1_ASAP7_75t_R FILLER_245_612 ();
 DECAPx1_ASAP7_75t_R FILLER_245_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_626 ();
 DECAPx6_ASAP7_75t_R FILLER_245_654 ();
 DECAPx2_ASAP7_75t_R FILLER_245_668 ();
 DECAPx1_ASAP7_75t_R FILLER_245_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_747 ();
 FILLER_ASAP7_75t_R FILLER_245_778 ();
 FILLER_ASAP7_75t_R FILLER_245_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_819 ();
 DECAPx4_ASAP7_75t_R FILLER_245_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_833 ();
 DECAPx1_ASAP7_75t_R FILLER_245_851 ();
 DECAPx10_ASAP7_75t_R FILLER_245_865 ();
 DECAPx6_ASAP7_75t_R FILLER_245_907 ();
 FILLER_ASAP7_75t_R FILLER_245_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_923 ();
 FILLER_ASAP7_75t_R FILLER_245_926 ();
 DECAPx10_ASAP7_75t_R FILLER_245_934 ();
 DECAPx1_ASAP7_75t_R FILLER_245_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_960 ();
 FILLER_ASAP7_75t_R FILLER_245_967 ();
 FILLER_ASAP7_75t_R FILLER_245_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1049 ();
 FILLER_ASAP7_75t_R FILLER_245_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1125 ();
 FILLER_ASAP7_75t_R FILLER_245_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_245_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1193 ();
 FILLER_ASAP7_75t_R FILLER_245_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1235 ();
 FILLER_ASAP7_75t_R FILLER_245_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1259 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1272 ();
 FILLER_ASAP7_75t_R FILLER_245_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1321 ();
 FILLER_ASAP7_75t_R FILLER_245_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1329 ();
 FILLER_ASAP7_75t_R FILLER_245_1339 ();
 FILLER_ASAP7_75t_R FILLER_245_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1349 ();
 FILLER_ASAP7_75t_R FILLER_245_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_245_1401 ();
 DECAPx10_ASAP7_75t_R FILLER_246_2 ();
 DECAPx10_ASAP7_75t_R FILLER_246_24 ();
 DECAPx10_ASAP7_75t_R FILLER_246_46 ();
 DECAPx10_ASAP7_75t_R FILLER_246_68 ();
 DECAPx10_ASAP7_75t_R FILLER_246_90 ();
 DECAPx10_ASAP7_75t_R FILLER_246_112 ();
 DECAPx10_ASAP7_75t_R FILLER_246_134 ();
 DECAPx10_ASAP7_75t_R FILLER_246_156 ();
 DECAPx10_ASAP7_75t_R FILLER_246_178 ();
 DECAPx10_ASAP7_75t_R FILLER_246_200 ();
 DECAPx10_ASAP7_75t_R FILLER_246_222 ();
 DECAPx10_ASAP7_75t_R FILLER_246_244 ();
 DECAPx10_ASAP7_75t_R FILLER_246_266 ();
 DECAPx10_ASAP7_75t_R FILLER_246_288 ();
 DECAPx4_ASAP7_75t_R FILLER_246_310 ();
 FILLER_ASAP7_75t_R FILLER_246_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_322 ();
 DECAPx6_ASAP7_75t_R FILLER_246_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_340 ();
 DECAPx2_ASAP7_75t_R FILLER_246_397 ();
 FILLER_ASAP7_75t_R FILLER_246_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_405 ();
 DECAPx2_ASAP7_75t_R FILLER_246_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_420 ();
 DECAPx6_ASAP7_75t_R FILLER_246_424 ();
 DECAPx1_ASAP7_75t_R FILLER_246_438 ();
 DECAPx6_ASAP7_75t_R FILLER_246_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_464 ();
 DECAPx10_ASAP7_75t_R FILLER_246_486 ();
 DECAPx10_ASAP7_75t_R FILLER_246_508 ();
 DECAPx4_ASAP7_75t_R FILLER_246_530 ();
 FILLER_ASAP7_75t_R FILLER_246_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_542 ();
 DECAPx2_ASAP7_75t_R FILLER_246_555 ();
 DECAPx2_ASAP7_75t_R FILLER_246_577 ();
 DECAPx1_ASAP7_75t_R FILLER_246_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_595 ();
 DECAPx1_ASAP7_75t_R FILLER_246_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_615 ();
 FILLER_ASAP7_75t_R FILLER_246_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_625 ();
 FILLER_ASAP7_75t_R FILLER_246_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_646 ();
 DECAPx4_ASAP7_75t_R FILLER_246_670 ();
 FILLER_ASAP7_75t_R FILLER_246_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_682 ();
 DECAPx1_ASAP7_75t_R FILLER_246_691 ();
 DECAPx6_ASAP7_75t_R FILLER_246_721 ();
 DECAPx4_ASAP7_75t_R FILLER_246_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_748 ();
 DECAPx1_ASAP7_75t_R FILLER_246_778 ();
 DECAPx2_ASAP7_75t_R FILLER_246_798 ();
 FILLER_ASAP7_75t_R FILLER_246_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_806 ();
 DECAPx10_ASAP7_75t_R FILLER_246_810 ();
 DECAPx2_ASAP7_75t_R FILLER_246_853 ();
 DECAPx1_ASAP7_75t_R FILLER_246_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_866 ();
 DECAPx10_ASAP7_75t_R FILLER_246_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_899 ();
 DECAPx6_ASAP7_75t_R FILLER_246_938 ();
 DECAPx1_ASAP7_75t_R FILLER_246_952 ();
 DECAPx10_ASAP7_75t_R FILLER_246_962 ();
 DECAPx6_ASAP7_75t_R FILLER_246_984 ();
 DECAPx1_ASAP7_75t_R FILLER_246_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_246_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_246_1081 ();
 FILLER_ASAP7_75t_R FILLER_246_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1132 ();
 FILLER_ASAP7_75t_R FILLER_246_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1150 ();
 FILLER_ASAP7_75t_R FILLER_246_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_246_1211 ();
 FILLER_ASAP7_75t_R FILLER_246_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_246_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1257 ();
 FILLER_ASAP7_75t_R FILLER_246_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1265 ();
 DECAPx6_ASAP7_75t_R FILLER_246_1272 ();
 FILLER_ASAP7_75t_R FILLER_246_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1316 ();
 FILLER_ASAP7_75t_R FILLER_246_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1340 ();
 DECAPx4_ASAP7_75t_R FILLER_246_1348 ();
 FILLER_ASAP7_75t_R FILLER_246_1358 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1396 ();
 FILLER_ASAP7_75t_R FILLER_246_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_247_2 ();
 DECAPx10_ASAP7_75t_R FILLER_247_24 ();
 DECAPx10_ASAP7_75t_R FILLER_247_46 ();
 DECAPx10_ASAP7_75t_R FILLER_247_68 ();
 DECAPx10_ASAP7_75t_R FILLER_247_90 ();
 DECAPx10_ASAP7_75t_R FILLER_247_112 ();
 DECAPx10_ASAP7_75t_R FILLER_247_134 ();
 DECAPx10_ASAP7_75t_R FILLER_247_156 ();
 DECAPx10_ASAP7_75t_R FILLER_247_178 ();
 DECAPx10_ASAP7_75t_R FILLER_247_200 ();
 DECAPx10_ASAP7_75t_R FILLER_247_222 ();
 DECAPx10_ASAP7_75t_R FILLER_247_244 ();
 DECAPx10_ASAP7_75t_R FILLER_247_266 ();
 DECAPx10_ASAP7_75t_R FILLER_247_288 ();
 DECAPx10_ASAP7_75t_R FILLER_247_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_332 ();
 DECAPx1_ASAP7_75t_R FILLER_247_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_359 ();
 DECAPx6_ASAP7_75t_R FILLER_247_363 ();
 DECAPx1_ASAP7_75t_R FILLER_247_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_381 ();
 DECAPx10_ASAP7_75t_R FILLER_247_385 ();
 DECAPx6_ASAP7_75t_R FILLER_247_407 ();
 DECAPx1_ASAP7_75t_R FILLER_247_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_425 ();
 DECAPx10_ASAP7_75t_R FILLER_247_453 ();
 DECAPx6_ASAP7_75t_R FILLER_247_475 ();
 FILLER_ASAP7_75t_R FILLER_247_489 ();
 DECAPx2_ASAP7_75t_R FILLER_247_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_518 ();
 DECAPx6_ASAP7_75t_R FILLER_247_527 ();
 FILLER_ASAP7_75t_R FILLER_247_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_543 ();
 DECAPx10_ASAP7_75t_R FILLER_247_552 ();
 DECAPx2_ASAP7_75t_R FILLER_247_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_580 ();
 FILLER_ASAP7_75t_R FILLER_247_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_607 ();
 DECAPx10_ASAP7_75t_R FILLER_247_623 ();
 DECAPx2_ASAP7_75t_R FILLER_247_645 ();
 FILLER_ASAP7_75t_R FILLER_247_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_669 ();
 DECAPx10_ASAP7_75t_R FILLER_247_678 ();
 DECAPx1_ASAP7_75t_R FILLER_247_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_708 ();
 DECAPx4_ASAP7_75t_R FILLER_247_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_722 ();
 DECAPx6_ASAP7_75t_R FILLER_247_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_750 ();
 DECAPx2_ASAP7_75t_R FILLER_247_754 ();
 DECAPx1_ASAP7_75t_R FILLER_247_770 ();
 DECAPx1_ASAP7_75t_R FILLER_247_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_781 ();
 FILLER_ASAP7_75t_R FILLER_247_798 ();
 DECAPx1_ASAP7_75t_R FILLER_247_807 ();
 DECAPx2_ASAP7_75t_R FILLER_247_814 ();
 FILLER_ASAP7_75t_R FILLER_247_820 ();
 DECAPx6_ASAP7_75t_R FILLER_247_832 ();
 FILLER_ASAP7_75t_R FILLER_247_846 ();
 DECAPx1_ASAP7_75t_R FILLER_247_855 ();
 DECAPx1_ASAP7_75t_R FILLER_247_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_892 ();
 DECAPx1_ASAP7_75t_R FILLER_247_920 ();
 FILLER_ASAP7_75t_R FILLER_247_926 ();
 FILLER_ASAP7_75t_R FILLER_247_972 ();
 FILLER_ASAP7_75t_R FILLER_247_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_984 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_247_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_247_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_247_1060 ();
 FILLER_ASAP7_75t_R FILLER_247_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_247_1097 ();
 FILLER_ASAP7_75t_R FILLER_247_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_247_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_247_1177 ();
 FILLER_ASAP7_75t_R FILLER_247_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_247_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_247_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1217 ();
 FILLER_ASAP7_75t_R FILLER_247_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_247_1284 ();
 FILLER_ASAP7_75t_R FILLER_247_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_247_1326 ();
 DECAPx6_ASAP7_75t_R FILLER_247_1390 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_248_2 ();
 DECAPx10_ASAP7_75t_R FILLER_248_24 ();
 DECAPx10_ASAP7_75t_R FILLER_248_46 ();
 DECAPx10_ASAP7_75t_R FILLER_248_68 ();
 DECAPx10_ASAP7_75t_R FILLER_248_90 ();
 DECAPx10_ASAP7_75t_R FILLER_248_112 ();
 DECAPx10_ASAP7_75t_R FILLER_248_134 ();
 DECAPx10_ASAP7_75t_R FILLER_248_156 ();
 DECAPx10_ASAP7_75t_R FILLER_248_178 ();
 DECAPx10_ASAP7_75t_R FILLER_248_200 ();
 DECAPx10_ASAP7_75t_R FILLER_248_222 ();
 DECAPx10_ASAP7_75t_R FILLER_248_244 ();
 DECAPx10_ASAP7_75t_R FILLER_248_266 ();
 DECAPx10_ASAP7_75t_R FILLER_248_288 ();
 DECAPx10_ASAP7_75t_R FILLER_248_310 ();
 DECAPx10_ASAP7_75t_R FILLER_248_332 ();
 DECAPx10_ASAP7_75t_R FILLER_248_354 ();
 DECAPx10_ASAP7_75t_R FILLER_248_376 ();
 DECAPx10_ASAP7_75t_R FILLER_248_398 ();
 DECAPx2_ASAP7_75t_R FILLER_248_420 ();
 FILLER_ASAP7_75t_R FILLER_248_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_520 ();
 DECAPx4_ASAP7_75t_R FILLER_248_535 ();
 FILLER_ASAP7_75t_R FILLER_248_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_547 ();
 DECAPx1_ASAP7_75t_R FILLER_248_566 ();
 DECAPx2_ASAP7_75t_R FILLER_248_578 ();
 DECAPx4_ASAP7_75t_R FILLER_248_599 ();
 FILLER_ASAP7_75t_R FILLER_248_609 ();
 DECAPx10_ASAP7_75t_R FILLER_248_627 ();
 DECAPx4_ASAP7_75t_R FILLER_248_649 ();
 DECAPx4_ASAP7_75t_R FILLER_248_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_676 ();
 DECAPx10_ASAP7_75t_R FILLER_248_687 ();
 DECAPx1_ASAP7_75t_R FILLER_248_709 ();
 DECAPx1_ASAP7_75t_R FILLER_248_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_757 ();
 DECAPx4_ASAP7_75t_R FILLER_248_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_794 ();
 DECAPx4_ASAP7_75t_R FILLER_248_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_831 ();
 FILLER_ASAP7_75t_R FILLER_248_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_837 ();
 DECAPx2_ASAP7_75t_R FILLER_248_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_850 ();
 DECAPx2_ASAP7_75t_R FILLER_248_857 ();
 FILLER_ASAP7_75t_R FILLER_248_863 ();
 FILLER_ASAP7_75t_R FILLER_248_874 ();
 DECAPx4_ASAP7_75t_R FILLER_248_883 ();
 FILLER_ASAP7_75t_R FILLER_248_893 ();
 DECAPx2_ASAP7_75t_R FILLER_248_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_927 ();
 FILLER_ASAP7_75t_R FILLER_248_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_937 ();
 DECAPx2_ASAP7_75t_R FILLER_248_965 ();
 FILLER_ASAP7_75t_R FILLER_248_971 ();
 FILLER_ASAP7_75t_R FILLER_248_988 ();
 FILLER_ASAP7_75t_R FILLER_248_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1003 ();
 FILLER_ASAP7_75t_R FILLER_248_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_248_1027 ();
 FILLER_ASAP7_75t_R FILLER_248_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_248_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_248_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_248_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_248_1168 ();
 FILLER_ASAP7_75t_R FILLER_248_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1299 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1320 ();
 FILLER_ASAP7_75t_R FILLER_248_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1329 ();
 FILLER_ASAP7_75t_R FILLER_248_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1348 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1355 ();
 DECAPx4_ASAP7_75t_R FILLER_248_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_248_1388 ();
 FILLER_ASAP7_75t_R FILLER_248_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_249_2 ();
 DECAPx10_ASAP7_75t_R FILLER_249_24 ();
 DECAPx10_ASAP7_75t_R FILLER_249_46 ();
 DECAPx10_ASAP7_75t_R FILLER_249_68 ();
 DECAPx10_ASAP7_75t_R FILLER_249_90 ();
 DECAPx10_ASAP7_75t_R FILLER_249_112 ();
 DECAPx10_ASAP7_75t_R FILLER_249_134 ();
 DECAPx10_ASAP7_75t_R FILLER_249_156 ();
 DECAPx10_ASAP7_75t_R FILLER_249_178 ();
 DECAPx10_ASAP7_75t_R FILLER_249_200 ();
 DECAPx10_ASAP7_75t_R FILLER_249_222 ();
 DECAPx10_ASAP7_75t_R FILLER_249_244 ();
 DECAPx10_ASAP7_75t_R FILLER_249_266 ();
 DECAPx10_ASAP7_75t_R FILLER_249_288 ();
 DECAPx10_ASAP7_75t_R FILLER_249_310 ();
 DECAPx10_ASAP7_75t_R FILLER_249_332 ();
 DECAPx10_ASAP7_75t_R FILLER_249_354 ();
 DECAPx10_ASAP7_75t_R FILLER_249_376 ();
 DECAPx10_ASAP7_75t_R FILLER_249_398 ();
 DECAPx4_ASAP7_75t_R FILLER_249_420 ();
 FILLER_ASAP7_75t_R FILLER_249_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_432 ();
 FILLER_ASAP7_75t_R FILLER_249_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_485 ();
 DECAPx1_ASAP7_75t_R FILLER_249_493 ();
 DECAPx1_ASAP7_75t_R FILLER_249_519 ();
 DECAPx4_ASAP7_75t_R FILLER_249_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_547 ();
 FILLER_ASAP7_75t_R FILLER_249_554 ();
 DECAPx1_ASAP7_75t_R FILLER_249_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_578 ();
 FILLER_ASAP7_75t_R FILLER_249_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_599 ();
 DECAPx2_ASAP7_75t_R FILLER_249_606 ();
 FILLER_ASAP7_75t_R FILLER_249_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_614 ();
 DECAPx2_ASAP7_75t_R FILLER_249_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_675 ();
 DECAPx2_ASAP7_75t_R FILLER_249_683 ();
 FILLER_ASAP7_75t_R FILLER_249_689 ();
 FILLER_ASAP7_75t_R FILLER_249_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_722 ();
 DECAPx4_ASAP7_75t_R FILLER_249_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_743 ();
 DECAPx2_ASAP7_75t_R FILLER_249_753 ();
 DECAPx1_ASAP7_75t_R FILLER_249_768 ();
 DECAPx1_ASAP7_75t_R FILLER_249_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_786 ();
 FILLER_ASAP7_75t_R FILLER_249_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_808 ();
 FILLER_ASAP7_75t_R FILLER_249_812 ();
 DECAPx1_ASAP7_75t_R FILLER_249_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_853 ();
 DECAPx4_ASAP7_75t_R FILLER_249_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_870 ();
 DECAPx6_ASAP7_75t_R FILLER_249_888 ();
 DECAPx1_ASAP7_75t_R FILLER_249_920 ();
 DECAPx4_ASAP7_75t_R FILLER_249_926 ();
 DECAPx4_ASAP7_75t_R FILLER_249_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_953 ();
 DECAPx2_ASAP7_75t_R FILLER_249_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_972 ();
 DECAPx2_ASAP7_75t_R FILLER_249_998 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_249_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_249_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1108 ();
 DECAPx1_ASAP7_75t_R FILLER_249_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1171 ();
 FILLER_ASAP7_75t_R FILLER_249_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1233 ();
 FILLER_ASAP7_75t_R FILLER_249_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1268 ();
 FILLER_ASAP7_75t_R FILLER_249_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_249_1283 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1290 ();
 FILLER_ASAP7_75t_R FILLER_249_1296 ();
 DECAPx4_ASAP7_75t_R FILLER_249_1331 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1347 ();
 FILLER_ASAP7_75t_R FILLER_249_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1355 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1389 ();
 FILLER_ASAP7_75t_R FILLER_249_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_250_2 ();
 DECAPx10_ASAP7_75t_R FILLER_250_24 ();
 DECAPx10_ASAP7_75t_R FILLER_250_46 ();
 DECAPx10_ASAP7_75t_R FILLER_250_68 ();
 DECAPx10_ASAP7_75t_R FILLER_250_90 ();
 DECAPx10_ASAP7_75t_R FILLER_250_112 ();
 DECAPx10_ASAP7_75t_R FILLER_250_134 ();
 DECAPx10_ASAP7_75t_R FILLER_250_156 ();
 DECAPx10_ASAP7_75t_R FILLER_250_178 ();
 DECAPx10_ASAP7_75t_R FILLER_250_200 ();
 DECAPx10_ASAP7_75t_R FILLER_250_222 ();
 DECAPx10_ASAP7_75t_R FILLER_250_244 ();
 DECAPx10_ASAP7_75t_R FILLER_250_266 ();
 DECAPx10_ASAP7_75t_R FILLER_250_288 ();
 DECAPx10_ASAP7_75t_R FILLER_250_310 ();
 DECAPx10_ASAP7_75t_R FILLER_250_332 ();
 DECAPx10_ASAP7_75t_R FILLER_250_354 ();
 DECAPx10_ASAP7_75t_R FILLER_250_376 ();
 DECAPx6_ASAP7_75t_R FILLER_250_398 ();
 DECAPx2_ASAP7_75t_R FILLER_250_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_418 ();
 DECAPx10_ASAP7_75t_R FILLER_250_425 ();
 DECAPx6_ASAP7_75t_R FILLER_250_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_461 ();
 DECAPx1_ASAP7_75t_R FILLER_250_464 ();
 FILLER_ASAP7_75t_R FILLER_250_474 ();
 FILLER_ASAP7_75t_R FILLER_250_482 ();
 DECAPx4_ASAP7_75t_R FILLER_250_497 ();
 FILLER_ASAP7_75t_R FILLER_250_507 ();
 FILLER_ASAP7_75t_R FILLER_250_517 ();
 DECAPx10_ASAP7_75t_R FILLER_250_554 ();
 DECAPx6_ASAP7_75t_R FILLER_250_576 ();
 DECAPx2_ASAP7_75t_R FILLER_250_590 ();
 FILLER_ASAP7_75t_R FILLER_250_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_613 ();
 FILLER_ASAP7_75t_R FILLER_250_623 ();
 DECAPx2_ASAP7_75t_R FILLER_250_638 ();
 FILLER_ASAP7_75t_R FILLER_250_644 ();
 DECAPx10_ASAP7_75t_R FILLER_250_662 ();
 DECAPx6_ASAP7_75t_R FILLER_250_684 ();
 DECAPx2_ASAP7_75t_R FILLER_250_724 ();
 DECAPx6_ASAP7_75t_R FILLER_250_743 ();
 DECAPx2_ASAP7_75t_R FILLER_250_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_776 ();
 FILLER_ASAP7_75t_R FILLER_250_784 ();
 DECAPx6_ASAP7_75t_R FILLER_250_815 ();
 FILLER_ASAP7_75t_R FILLER_250_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_831 ();
 DECAPx1_ASAP7_75t_R FILLER_250_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_839 ();
 FILLER_ASAP7_75t_R FILLER_250_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_855 ();
 DECAPx10_ASAP7_75t_R FILLER_250_866 ();
 DECAPx1_ASAP7_75t_R FILLER_250_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_892 ();
 DECAPx2_ASAP7_75t_R FILLER_250_899 ();
 FILLER_ASAP7_75t_R FILLER_250_905 ();
 DECAPx1_ASAP7_75t_R FILLER_250_936 ();
 DECAPx10_ASAP7_75t_R FILLER_250_949 ();
 DECAPx2_ASAP7_75t_R FILLER_250_971 ();
 DECAPx10_ASAP7_75t_R FILLER_250_983 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_250_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1052 ();
 FILLER_ASAP7_75t_R FILLER_250_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_250_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_250_1157 ();
 FILLER_ASAP7_75t_R FILLER_250_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_250_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1223 ();
 DECAPx4_ASAP7_75t_R FILLER_250_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1272 ();
 DECAPx6_ASAP7_75t_R FILLER_250_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1312 ();
 DECAPx6_ASAP7_75t_R FILLER_250_1323 ();
 FILLER_ASAP7_75t_R FILLER_250_1337 ();
 FILLER_ASAP7_75t_R FILLER_250_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1361 ();
 FILLER_ASAP7_75t_R FILLER_250_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1377 ();
 DECAPx1_ASAP7_75t_R FILLER_250_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_250_1388 ();
 FILLER_ASAP7_75t_R FILLER_250_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_251_2 ();
 DECAPx10_ASAP7_75t_R FILLER_251_24 ();
 DECAPx10_ASAP7_75t_R FILLER_251_46 ();
 DECAPx10_ASAP7_75t_R FILLER_251_68 ();
 DECAPx10_ASAP7_75t_R FILLER_251_90 ();
 DECAPx10_ASAP7_75t_R FILLER_251_112 ();
 DECAPx10_ASAP7_75t_R FILLER_251_134 ();
 DECAPx10_ASAP7_75t_R FILLER_251_156 ();
 DECAPx10_ASAP7_75t_R FILLER_251_178 ();
 DECAPx10_ASAP7_75t_R FILLER_251_200 ();
 DECAPx10_ASAP7_75t_R FILLER_251_222 ();
 DECAPx10_ASAP7_75t_R FILLER_251_244 ();
 DECAPx10_ASAP7_75t_R FILLER_251_266 ();
 DECAPx10_ASAP7_75t_R FILLER_251_288 ();
 DECAPx10_ASAP7_75t_R FILLER_251_310 ();
 DECAPx10_ASAP7_75t_R FILLER_251_332 ();
 DECAPx10_ASAP7_75t_R FILLER_251_354 ();
 DECAPx10_ASAP7_75t_R FILLER_251_376 ();
 DECAPx2_ASAP7_75t_R FILLER_251_398 ();
 DECAPx4_ASAP7_75t_R FILLER_251_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_441 ();
 DECAPx1_ASAP7_75t_R FILLER_251_452 ();
 DECAPx6_ASAP7_75t_R FILLER_251_462 ();
 DECAPx2_ASAP7_75t_R FILLER_251_476 ();
 DECAPx2_ASAP7_75t_R FILLER_251_494 ();
 DECAPx1_ASAP7_75t_R FILLER_251_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_537 ();
 DECAPx2_ASAP7_75t_R FILLER_251_546 ();
 FILLER_ASAP7_75t_R FILLER_251_552 ();
 DECAPx1_ASAP7_75t_R FILLER_251_562 ();
 DECAPx1_ASAP7_75t_R FILLER_251_572 ();
 DECAPx10_ASAP7_75t_R FILLER_251_582 ();
 DECAPx6_ASAP7_75t_R FILLER_251_604 ();
 DECAPx6_ASAP7_75t_R FILLER_251_626 ();
 DECAPx1_ASAP7_75t_R FILLER_251_640 ();
 DECAPx10_ASAP7_75t_R FILLER_251_656 ();
 DECAPx10_ASAP7_75t_R FILLER_251_678 ();
 DECAPx2_ASAP7_75t_R FILLER_251_700 ();
 DECAPx1_ASAP7_75t_R FILLER_251_709 ();
 DECAPx1_ASAP7_75t_R FILLER_251_716 ();
 FILLER_ASAP7_75t_R FILLER_251_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_800 ();
 DECAPx10_ASAP7_75t_R FILLER_251_804 ();
 DECAPx6_ASAP7_75t_R FILLER_251_826 ();
 FILLER_ASAP7_75t_R FILLER_251_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_848 ();
 DECAPx2_ASAP7_75t_R FILLER_251_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_883 ();
 FILLER_ASAP7_75t_R FILLER_251_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_906 ();
 FILLER_ASAP7_75t_R FILLER_251_913 ();
 FILLER_ASAP7_75t_R FILLER_251_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_923 ();
 DECAPx2_ASAP7_75t_R FILLER_251_926 ();
 FILLER_ASAP7_75t_R FILLER_251_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_934 ();
 DECAPx2_ASAP7_75t_R FILLER_251_957 ();
 FILLER_ASAP7_75t_R FILLER_251_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_996 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_251_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1050 ();
 FILLER_ASAP7_75t_R FILLER_251_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1093 ();
 FILLER_ASAP7_75t_R FILLER_251_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1109 ();
 FILLER_ASAP7_75t_R FILLER_251_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_251_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_251_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_251_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_251_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1293 ();
 FILLER_ASAP7_75t_R FILLER_251_1299 ();
 DECAPx4_ASAP7_75t_R FILLER_251_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1335 ();
 FILLER_ASAP7_75t_R FILLER_251_1362 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1390 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_252_2 ();
 DECAPx10_ASAP7_75t_R FILLER_252_24 ();
 DECAPx10_ASAP7_75t_R FILLER_252_46 ();
 DECAPx10_ASAP7_75t_R FILLER_252_68 ();
 DECAPx10_ASAP7_75t_R FILLER_252_90 ();
 DECAPx10_ASAP7_75t_R FILLER_252_112 ();
 DECAPx10_ASAP7_75t_R FILLER_252_134 ();
 DECAPx10_ASAP7_75t_R FILLER_252_156 ();
 DECAPx10_ASAP7_75t_R FILLER_252_178 ();
 DECAPx10_ASAP7_75t_R FILLER_252_200 ();
 DECAPx10_ASAP7_75t_R FILLER_252_222 ();
 DECAPx10_ASAP7_75t_R FILLER_252_244 ();
 DECAPx10_ASAP7_75t_R FILLER_252_266 ();
 DECAPx10_ASAP7_75t_R FILLER_252_288 ();
 DECAPx10_ASAP7_75t_R FILLER_252_310 ();
 DECAPx10_ASAP7_75t_R FILLER_252_332 ();
 DECAPx10_ASAP7_75t_R FILLER_252_354 ();
 DECAPx10_ASAP7_75t_R FILLER_252_376 ();
 DECAPx6_ASAP7_75t_R FILLER_252_398 ();
 DECAPx1_ASAP7_75t_R FILLER_252_412 ();
 DECAPx1_ASAP7_75t_R FILLER_252_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_427 ();
 DECAPx1_ASAP7_75t_R FILLER_252_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_440 ();
 DECAPx1_ASAP7_75t_R FILLER_252_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_468 ();
 FILLER_ASAP7_75t_R FILLER_252_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_484 ();
 DECAPx2_ASAP7_75t_R FILLER_252_522 ();
 FILLER_ASAP7_75t_R FILLER_252_528 ();
 DECAPx4_ASAP7_75t_R FILLER_252_544 ();
 FILLER_ASAP7_75t_R FILLER_252_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_556 ();
 FILLER_ASAP7_75t_R FILLER_252_564 ();
 DECAPx2_ASAP7_75t_R FILLER_252_586 ();
 DECAPx10_ASAP7_75t_R FILLER_252_606 ();
 FILLER_ASAP7_75t_R FILLER_252_628 ();
 DECAPx2_ASAP7_75t_R FILLER_252_637 ();
 FILLER_ASAP7_75t_R FILLER_252_643 ();
 DECAPx6_ASAP7_75t_R FILLER_252_655 ();
 DECAPx1_ASAP7_75t_R FILLER_252_669 ();
 DECAPx1_ASAP7_75t_R FILLER_252_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_687 ();
 FILLER_ASAP7_75t_R FILLER_252_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_693 ();
 DECAPx4_ASAP7_75t_R FILLER_252_701 ();
 DECAPx6_ASAP7_75t_R FILLER_252_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_733 ();
 DECAPx6_ASAP7_75t_R FILLER_252_737 ();
 DECAPx2_ASAP7_75t_R FILLER_252_751 ();
 DECAPx4_ASAP7_75t_R FILLER_252_766 ();
 FILLER_ASAP7_75t_R FILLER_252_776 ();
 DECAPx10_ASAP7_75t_R FILLER_252_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_831 ();
 DECAPx1_ASAP7_75t_R FILLER_252_853 ();
 DECAPx6_ASAP7_75t_R FILLER_252_865 ();
 FILLER_ASAP7_75t_R FILLER_252_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_911 ();
 DECAPx6_ASAP7_75t_R FILLER_252_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_953 ();
 FILLER_ASAP7_75t_R FILLER_252_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_972 ();
 FILLER_ASAP7_75t_R FILLER_252_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_996 ();
 DECAPx6_ASAP7_75t_R FILLER_252_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_252_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_252_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_252_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_252_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_252_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1245 ();
 FILLER_ASAP7_75t_R FILLER_252_1261 ();
 DECAPx1_ASAP7_75t_R FILLER_252_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_252_1307 ();
 FILLER_ASAP7_75t_R FILLER_252_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1319 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_252_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_252_1388 ();
 FILLER_ASAP7_75t_R FILLER_252_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_253_2 ();
 DECAPx10_ASAP7_75t_R FILLER_253_24 ();
 DECAPx10_ASAP7_75t_R FILLER_253_46 ();
 DECAPx10_ASAP7_75t_R FILLER_253_68 ();
 DECAPx10_ASAP7_75t_R FILLER_253_90 ();
 DECAPx10_ASAP7_75t_R FILLER_253_112 ();
 DECAPx10_ASAP7_75t_R FILLER_253_134 ();
 DECAPx10_ASAP7_75t_R FILLER_253_156 ();
 DECAPx10_ASAP7_75t_R FILLER_253_178 ();
 DECAPx10_ASAP7_75t_R FILLER_253_200 ();
 DECAPx10_ASAP7_75t_R FILLER_253_222 ();
 DECAPx10_ASAP7_75t_R FILLER_253_244 ();
 DECAPx10_ASAP7_75t_R FILLER_253_266 ();
 DECAPx10_ASAP7_75t_R FILLER_253_288 ();
 DECAPx10_ASAP7_75t_R FILLER_253_310 ();
 DECAPx10_ASAP7_75t_R FILLER_253_332 ();
 DECAPx10_ASAP7_75t_R FILLER_253_354 ();
 DECAPx10_ASAP7_75t_R FILLER_253_376 ();
 DECAPx2_ASAP7_75t_R FILLER_253_461 ();
 FILLER_ASAP7_75t_R FILLER_253_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_491 ();
 FILLER_ASAP7_75t_R FILLER_253_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_524 ();
 DECAPx1_ASAP7_75t_R FILLER_253_533 ();
 FILLER_ASAP7_75t_R FILLER_253_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_565 ();
 DECAPx1_ASAP7_75t_R FILLER_253_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_584 ();
 FILLER_ASAP7_75t_R FILLER_253_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_597 ();
 DECAPx4_ASAP7_75t_R FILLER_253_620 ();
 FILLER_ASAP7_75t_R FILLER_253_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_632 ();
 DECAPx6_ASAP7_75t_R FILLER_253_653 ();
 DECAPx2_ASAP7_75t_R FILLER_253_667 ();
 FILLER_ASAP7_75t_R FILLER_253_688 ();
 FILLER_ASAP7_75t_R FILLER_253_705 ();
 DECAPx4_ASAP7_75t_R FILLER_253_727 ();
 DECAPx6_ASAP7_75t_R FILLER_253_764 ();
 DECAPx1_ASAP7_75t_R FILLER_253_778 ();
 DECAPx6_ASAP7_75t_R FILLER_253_788 ();
 FILLER_ASAP7_75t_R FILLER_253_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_804 ();
 DECAPx10_ASAP7_75t_R FILLER_253_811 ();
 FILLER_ASAP7_75t_R FILLER_253_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_835 ();
 DECAPx1_ASAP7_75t_R FILLER_253_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_854 ();
 DECAPx1_ASAP7_75t_R FILLER_253_861 ();
 DECAPx6_ASAP7_75t_R FILLER_253_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_923 ();
 DECAPx6_ASAP7_75t_R FILLER_253_926 ();
 DECAPx1_ASAP7_75t_R FILLER_253_940 ();
 FILLER_ASAP7_75t_R FILLER_253_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_952 ();
 DECAPx4_ASAP7_75t_R FILLER_253_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_973 ();
 DECAPx2_ASAP7_75t_R FILLER_253_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_994 ();
 DECAPx1_ASAP7_75t_R FILLER_253_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1005 ();
 FILLER_ASAP7_75t_R FILLER_253_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_253_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1139 ();
 FILLER_ASAP7_75t_R FILLER_253_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_253_1168 ();
 FILLER_ASAP7_75t_R FILLER_253_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1190 ();
 FILLER_ASAP7_75t_R FILLER_253_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_253_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1288 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1353 ();
 FILLER_ASAP7_75t_R FILLER_253_1359 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_253_1386 ();
 DECAPx1_ASAP7_75t_R FILLER_253_1400 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_254_2 ();
 DECAPx10_ASAP7_75t_R FILLER_254_24 ();
 DECAPx10_ASAP7_75t_R FILLER_254_46 ();
 DECAPx10_ASAP7_75t_R FILLER_254_68 ();
 DECAPx10_ASAP7_75t_R FILLER_254_90 ();
 DECAPx10_ASAP7_75t_R FILLER_254_112 ();
 DECAPx10_ASAP7_75t_R FILLER_254_134 ();
 DECAPx10_ASAP7_75t_R FILLER_254_156 ();
 DECAPx10_ASAP7_75t_R FILLER_254_178 ();
 DECAPx10_ASAP7_75t_R FILLER_254_200 ();
 DECAPx10_ASAP7_75t_R FILLER_254_222 ();
 DECAPx10_ASAP7_75t_R FILLER_254_244 ();
 DECAPx10_ASAP7_75t_R FILLER_254_266 ();
 DECAPx10_ASAP7_75t_R FILLER_254_288 ();
 DECAPx10_ASAP7_75t_R FILLER_254_310 ();
 DECAPx10_ASAP7_75t_R FILLER_254_332 ();
 DECAPx10_ASAP7_75t_R FILLER_254_354 ();
 DECAPx10_ASAP7_75t_R FILLER_254_376 ();
 DECAPx6_ASAP7_75t_R FILLER_254_398 ();
 FILLER_ASAP7_75t_R FILLER_254_412 ();
 DECAPx2_ASAP7_75t_R FILLER_254_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_432 ();
 DECAPx4_ASAP7_75t_R FILLER_254_443 ();
 FILLER_ASAP7_75t_R FILLER_254_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_455 ();
 DECAPx1_ASAP7_75t_R FILLER_254_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_468 ();
 FILLER_ASAP7_75t_R FILLER_254_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_487 ();
 DECAPx1_ASAP7_75t_R FILLER_254_549 ();
 DECAPx1_ASAP7_75t_R FILLER_254_569 ();
 DECAPx2_ASAP7_75t_R FILLER_254_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_587 ();
 DECAPx1_ASAP7_75t_R FILLER_254_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_612 ();
 DECAPx2_ASAP7_75t_R FILLER_254_620 ();
 FILLER_ASAP7_75t_R FILLER_254_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_628 ();
 DECAPx6_ASAP7_75t_R FILLER_254_649 ();
 DECAPx1_ASAP7_75t_R FILLER_254_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_683 ();
 FILLER_ASAP7_75t_R FILLER_254_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_708 ();
 DECAPx4_ASAP7_75t_R FILLER_254_715 ();
 DECAPx2_ASAP7_75t_R FILLER_254_733 ();
 FILLER_ASAP7_75t_R FILLER_254_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_741 ();
 FILLER_ASAP7_75t_R FILLER_254_758 ();
 DECAPx2_ASAP7_75t_R FILLER_254_774 ();
 FILLER_ASAP7_75t_R FILLER_254_780 ();
 FILLER_ASAP7_75t_R FILLER_254_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_840 ();
 DECAPx1_ASAP7_75t_R FILLER_254_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_858 ();
 DECAPx6_ASAP7_75t_R FILLER_254_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_896 ();
 DECAPx10_ASAP7_75t_R FILLER_254_948 ();
 DECAPx10_ASAP7_75t_R FILLER_254_970 ();
 DECAPx10_ASAP7_75t_R FILLER_254_992 ();
 DECAPx2_ASAP7_75t_R FILLER_254_1014 ();
 FILLER_ASAP7_75t_R FILLER_254_1020 ();
 FILLER_ASAP7_75t_R FILLER_254_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1037 ();
 FILLER_ASAP7_75t_R FILLER_254_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_254_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_254_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1150 ();
 FILLER_ASAP7_75t_R FILLER_254_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_254_1220 ();
 FILLER_ASAP7_75t_R FILLER_254_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1228 ();
 FILLER_ASAP7_75t_R FILLER_254_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1257 ();
 DECAPx1_ASAP7_75t_R FILLER_254_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1280 ();
 FILLER_ASAP7_75t_R FILLER_254_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1303 ();
 FILLER_ASAP7_75t_R FILLER_254_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1340 ();
 FILLER_ASAP7_75t_R FILLER_254_1362 ();
 DECAPx6_ASAP7_75t_R FILLER_254_1388 ();
 FILLER_ASAP7_75t_R FILLER_254_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_255_2 ();
 DECAPx10_ASAP7_75t_R FILLER_255_24 ();
 DECAPx10_ASAP7_75t_R FILLER_255_46 ();
 DECAPx10_ASAP7_75t_R FILLER_255_68 ();
 DECAPx10_ASAP7_75t_R FILLER_255_90 ();
 DECAPx10_ASAP7_75t_R FILLER_255_112 ();
 DECAPx10_ASAP7_75t_R FILLER_255_134 ();
 DECAPx10_ASAP7_75t_R FILLER_255_156 ();
 DECAPx10_ASAP7_75t_R FILLER_255_178 ();
 DECAPx10_ASAP7_75t_R FILLER_255_200 ();
 DECAPx10_ASAP7_75t_R FILLER_255_222 ();
 DECAPx10_ASAP7_75t_R FILLER_255_244 ();
 DECAPx10_ASAP7_75t_R FILLER_255_266 ();
 DECAPx10_ASAP7_75t_R FILLER_255_288 ();
 DECAPx10_ASAP7_75t_R FILLER_255_310 ();
 DECAPx10_ASAP7_75t_R FILLER_255_332 ();
 DECAPx10_ASAP7_75t_R FILLER_255_354 ();
 DECAPx10_ASAP7_75t_R FILLER_255_376 ();
 DECAPx6_ASAP7_75t_R FILLER_255_398 ();
 DECAPx1_ASAP7_75t_R FILLER_255_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_416 ();
 DECAPx10_ASAP7_75t_R FILLER_255_423 ();
 FILLER_ASAP7_75t_R FILLER_255_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_447 ();
 DECAPx1_ASAP7_75t_R FILLER_255_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_459 ();
 DECAPx10_ASAP7_75t_R FILLER_255_468 ();
 DECAPx6_ASAP7_75t_R FILLER_255_490 ();
 FILLER_ASAP7_75t_R FILLER_255_504 ();
 FILLER_ASAP7_75t_R FILLER_255_527 ();
 DECAPx6_ASAP7_75t_R FILLER_255_535 ();
 DECAPx2_ASAP7_75t_R FILLER_255_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_555 ();
 DECAPx4_ASAP7_75t_R FILLER_255_562 ();
 FILLER_ASAP7_75t_R FILLER_255_572 ();
 DECAPx10_ASAP7_75t_R FILLER_255_580 ();
 DECAPx2_ASAP7_75t_R FILLER_255_602 ();
 FILLER_ASAP7_75t_R FILLER_255_608 ();
 DECAPx6_ASAP7_75t_R FILLER_255_632 ();
 FILLER_ASAP7_75t_R FILLER_255_646 ();
 DECAPx1_ASAP7_75t_R FILLER_255_656 ();
 DECAPx1_ASAP7_75t_R FILLER_255_668 ();
 DECAPx10_ASAP7_75t_R FILLER_255_706 ();
 DECAPx4_ASAP7_75t_R FILLER_255_728 ();
 FILLER_ASAP7_75t_R FILLER_255_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_740 ();
 DECAPx1_ASAP7_75t_R FILLER_255_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_804 ();
 DECAPx4_ASAP7_75t_R FILLER_255_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_831 ();
 FILLER_ASAP7_75t_R FILLER_255_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_852 ();
 DECAPx4_ASAP7_75t_R FILLER_255_859 ();
 FILLER_ASAP7_75t_R FILLER_255_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_887 ();
 DECAPx6_ASAP7_75t_R FILLER_255_934 ();
 DECAPx6_ASAP7_75t_R FILLER_255_959 ();
 DECAPx2_ASAP7_75t_R FILLER_255_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_979 ();
 FILLER_ASAP7_75t_R FILLER_255_995 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1026 ();
 FILLER_ASAP7_75t_R FILLER_255_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1050 ();
 DECAPx4_ASAP7_75t_R FILLER_255_1077 ();
 FILLER_ASAP7_75t_R FILLER_255_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_255_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_255_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_255_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_255_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1201 ();
 FILLER_ASAP7_75t_R FILLER_255_1228 ();
 DECAPx6_ASAP7_75t_R FILLER_255_1256 ();
 DECAPx2_ASAP7_75t_R FILLER_255_1270 ();
 DECAPx1_ASAP7_75t_R FILLER_255_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_255_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_255_1305 ();
 FILLER_ASAP7_75t_R FILLER_255_1345 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1350 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1372 ();
 DECAPx4_ASAP7_75t_R FILLER_255_1394 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_256_2 ();
 DECAPx10_ASAP7_75t_R FILLER_256_24 ();
 DECAPx10_ASAP7_75t_R FILLER_256_46 ();
 DECAPx10_ASAP7_75t_R FILLER_256_68 ();
 DECAPx10_ASAP7_75t_R FILLER_256_90 ();
 DECAPx10_ASAP7_75t_R FILLER_256_112 ();
 DECAPx10_ASAP7_75t_R FILLER_256_134 ();
 DECAPx10_ASAP7_75t_R FILLER_256_156 ();
 DECAPx10_ASAP7_75t_R FILLER_256_178 ();
 DECAPx10_ASAP7_75t_R FILLER_256_200 ();
 DECAPx10_ASAP7_75t_R FILLER_256_222 ();
 DECAPx10_ASAP7_75t_R FILLER_256_244 ();
 DECAPx10_ASAP7_75t_R FILLER_256_266 ();
 DECAPx10_ASAP7_75t_R FILLER_256_288 ();
 DECAPx10_ASAP7_75t_R FILLER_256_310 ();
 DECAPx10_ASAP7_75t_R FILLER_256_332 ();
 DECAPx10_ASAP7_75t_R FILLER_256_354 ();
 DECAPx10_ASAP7_75t_R FILLER_256_376 ();
 FILLER_ASAP7_75t_R FILLER_256_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_400 ();
 FILLER_ASAP7_75t_R FILLER_256_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_430 ();
 DECAPx4_ASAP7_75t_R FILLER_256_464 ();
 FILLER_ASAP7_75t_R FILLER_256_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_486 ();
 DECAPx6_ASAP7_75t_R FILLER_256_495 ();
 DECAPx2_ASAP7_75t_R FILLER_256_509 ();
 DECAPx4_ASAP7_75t_R FILLER_256_529 ();
 FILLER_ASAP7_75t_R FILLER_256_539 ();
 DECAPx4_ASAP7_75t_R FILLER_256_544 ();
 DECAPx6_ASAP7_75t_R FILLER_256_557 ();
 FILLER_ASAP7_75t_R FILLER_256_571 ();
 FILLER_ASAP7_75t_R FILLER_256_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_578 ();
 FILLER_ASAP7_75t_R FILLER_256_587 ();
 DECAPx4_ASAP7_75t_R FILLER_256_605 ();
 FILLER_ASAP7_75t_R FILLER_256_615 ();
 DECAPx1_ASAP7_75t_R FILLER_256_620 ();
 DECAPx4_ASAP7_75t_R FILLER_256_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_659 ();
 FILLER_ASAP7_75t_R FILLER_256_668 ();
 DECAPx6_ASAP7_75t_R FILLER_256_687 ();
 FILLER_ASAP7_75t_R FILLER_256_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_703 ();
 DECAPx6_ASAP7_75t_R FILLER_256_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_724 ();
 DECAPx6_ASAP7_75t_R FILLER_256_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_801 ();
 DECAPx10_ASAP7_75t_R FILLER_256_810 ();
 DECAPx1_ASAP7_75t_R FILLER_256_832 ();
 DECAPx1_ASAP7_75t_R FILLER_256_846 ();
 FILLER_ASAP7_75t_R FILLER_256_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_867 ();
 FILLER_ASAP7_75t_R FILLER_256_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_899 ();
 DECAPx6_ASAP7_75t_R FILLER_256_915 ();
 FILLER_ASAP7_75t_R FILLER_256_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_256_1032 ();
 FILLER_ASAP7_75t_R FILLER_256_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_256_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1069 ();
 FILLER_ASAP7_75t_R FILLER_256_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1105 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1124 ();
 FILLER_ASAP7_75t_R FILLER_256_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1197 ();
 FILLER_ASAP7_75t_R FILLER_256_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1205 ();
 FILLER_ASAP7_75t_R FILLER_256_1212 ();
 FILLER_ASAP7_75t_R FILLER_256_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1260 ();
 FILLER_ASAP7_75t_R FILLER_256_1266 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1312 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1388 ();
 FILLER_ASAP7_75t_R FILLER_256_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_257_2 ();
 DECAPx10_ASAP7_75t_R FILLER_257_24 ();
 DECAPx10_ASAP7_75t_R FILLER_257_46 ();
 DECAPx10_ASAP7_75t_R FILLER_257_68 ();
 DECAPx10_ASAP7_75t_R FILLER_257_90 ();
 DECAPx10_ASAP7_75t_R FILLER_257_112 ();
 DECAPx10_ASAP7_75t_R FILLER_257_134 ();
 DECAPx10_ASAP7_75t_R FILLER_257_156 ();
 DECAPx10_ASAP7_75t_R FILLER_257_178 ();
 DECAPx10_ASAP7_75t_R FILLER_257_200 ();
 DECAPx10_ASAP7_75t_R FILLER_257_222 ();
 DECAPx10_ASAP7_75t_R FILLER_257_244 ();
 DECAPx10_ASAP7_75t_R FILLER_257_266 ();
 DECAPx10_ASAP7_75t_R FILLER_257_288 ();
 DECAPx10_ASAP7_75t_R FILLER_257_310 ();
 DECAPx10_ASAP7_75t_R FILLER_257_332 ();
 DECAPx10_ASAP7_75t_R FILLER_257_354 ();
 DECAPx10_ASAP7_75t_R FILLER_257_376 ();
 DECAPx6_ASAP7_75t_R FILLER_257_398 ();
 FILLER_ASAP7_75t_R FILLER_257_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_414 ();
 DECAPx1_ASAP7_75t_R FILLER_257_422 ();
 FILLER_ASAP7_75t_R FILLER_257_447 ();
 DECAPx6_ASAP7_75t_R FILLER_257_455 ();
 DECAPx2_ASAP7_75t_R FILLER_257_520 ();
 DECAPx2_ASAP7_75t_R FILLER_257_532 ();
 DECAPx1_ASAP7_75t_R FILLER_257_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_571 ();
 DECAPx4_ASAP7_75t_R FILLER_257_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_597 ();
 FILLER_ASAP7_75t_R FILLER_257_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_606 ();
 FILLER_ASAP7_75t_R FILLER_257_613 ();
 FILLER_ASAP7_75t_R FILLER_257_621 ();
 DECAPx4_ASAP7_75t_R FILLER_257_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_646 ();
 DECAPx4_ASAP7_75t_R FILLER_257_659 ();
 FILLER_ASAP7_75t_R FILLER_257_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_671 ();
 DECAPx2_ASAP7_75t_R FILLER_257_684 ();
 DECAPx6_ASAP7_75t_R FILLER_257_696 ();
 DECAPx1_ASAP7_75t_R FILLER_257_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_714 ();
 DECAPx2_ASAP7_75t_R FILLER_257_743 ();
 DECAPx1_ASAP7_75t_R FILLER_257_759 ();
 DECAPx1_ASAP7_75t_R FILLER_257_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_773 ();
 DECAPx6_ASAP7_75t_R FILLER_257_796 ();
 DECAPx1_ASAP7_75t_R FILLER_257_810 ();
 DECAPx2_ASAP7_75t_R FILLER_257_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_841 ();
 DECAPx4_ASAP7_75t_R FILLER_257_869 ();
 DECAPx1_ASAP7_75t_R FILLER_257_885 ();
 FILLER_ASAP7_75t_R FILLER_257_896 ();
 DECAPx6_ASAP7_75t_R FILLER_257_904 ();
 DECAPx2_ASAP7_75t_R FILLER_257_918 ();
 DECAPx1_ASAP7_75t_R FILLER_257_926 ();
 FILLER_ASAP7_75t_R FILLER_257_946 ();
 DECAPx4_ASAP7_75t_R FILLER_257_959 ();
 DECAPx2_ASAP7_75t_R FILLER_257_976 ();
 FILLER_ASAP7_75t_R FILLER_257_982 ();
 DECAPx2_ASAP7_75t_R FILLER_257_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_257_1043 ();
 FILLER_ASAP7_75t_R FILLER_257_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_257_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_257_1134 ();
 FILLER_ASAP7_75t_R FILLER_257_1148 ();
 DECAPx6_ASAP7_75t_R FILLER_257_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_257_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_257_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_257_1219 ();
 FILLER_ASAP7_75t_R FILLER_257_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1227 ();
 DECAPx6_ASAP7_75t_R FILLER_257_1231 ();
 FILLER_ASAP7_75t_R FILLER_257_1245 ();
 FILLER_ASAP7_75t_R FILLER_257_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_257_1288 ();
 FILLER_ASAP7_75t_R FILLER_257_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1296 ();
 FILLER_ASAP7_75t_R FILLER_257_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1339 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1361 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1383 ();
 DECAPx10_ASAP7_75t_R FILLER_258_2 ();
 DECAPx10_ASAP7_75t_R FILLER_258_24 ();
 DECAPx10_ASAP7_75t_R FILLER_258_46 ();
 DECAPx10_ASAP7_75t_R FILLER_258_68 ();
 DECAPx10_ASAP7_75t_R FILLER_258_90 ();
 DECAPx10_ASAP7_75t_R FILLER_258_112 ();
 DECAPx10_ASAP7_75t_R FILLER_258_134 ();
 DECAPx10_ASAP7_75t_R FILLER_258_156 ();
 DECAPx10_ASAP7_75t_R FILLER_258_178 ();
 DECAPx10_ASAP7_75t_R FILLER_258_200 ();
 DECAPx10_ASAP7_75t_R FILLER_258_222 ();
 DECAPx10_ASAP7_75t_R FILLER_258_244 ();
 DECAPx10_ASAP7_75t_R FILLER_258_266 ();
 DECAPx10_ASAP7_75t_R FILLER_258_288 ();
 DECAPx10_ASAP7_75t_R FILLER_258_310 ();
 DECAPx10_ASAP7_75t_R FILLER_258_332 ();
 DECAPx10_ASAP7_75t_R FILLER_258_354 ();
 DECAPx10_ASAP7_75t_R FILLER_258_376 ();
 FILLER_ASAP7_75t_R FILLER_258_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_406 ();
 DECAPx4_ASAP7_75t_R FILLER_258_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_423 ();
 FILLER_ASAP7_75t_R FILLER_258_432 ();
 DECAPx10_ASAP7_75t_R FILLER_258_440 ();
 DECAPx1_ASAP7_75t_R FILLER_258_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_495 ();
 DECAPx1_ASAP7_75t_R FILLER_258_549 ();
 DECAPx4_ASAP7_75t_R FILLER_258_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_620 ();
 DECAPx1_ASAP7_75t_R FILLER_258_637 ();
 DECAPx4_ASAP7_75t_R FILLER_258_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_657 ();
 DECAPx2_ASAP7_75t_R FILLER_258_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_670 ();
 DECAPx1_ASAP7_75t_R FILLER_258_678 ();
 DECAPx4_ASAP7_75t_R FILLER_258_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_706 ();
 DECAPx10_ASAP7_75t_R FILLER_258_740 ();
 DECAPx2_ASAP7_75t_R FILLER_258_762 ();
 FILLER_ASAP7_75t_R FILLER_258_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_770 ();
 DECAPx10_ASAP7_75t_R FILLER_258_783 ();
 DECAPx2_ASAP7_75t_R FILLER_258_805 ();
 FILLER_ASAP7_75t_R FILLER_258_811 ();
 DECAPx1_ASAP7_75t_R FILLER_258_848 ();
 DECAPx4_ASAP7_75t_R FILLER_258_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_883 ();
 DECAPx2_ASAP7_75t_R FILLER_258_920 ();
 FILLER_ASAP7_75t_R FILLER_258_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_979 ();
 DECAPx6_ASAP7_75t_R FILLER_258_987 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1023 ();
 FILLER_ASAP7_75t_R FILLER_258_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1031 ();
 FILLER_ASAP7_75t_R FILLER_258_1040 ();
 FILLER_ASAP7_75t_R FILLER_258_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1058 ();
 FILLER_ASAP7_75t_R FILLER_258_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1069 ();
 FILLER_ASAP7_75t_R FILLER_258_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_258_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_258_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_258_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1135 ();
 FILLER_ASAP7_75t_R FILLER_258_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1216 ();
 DECAPx6_ASAP7_75t_R FILLER_258_1225 ();
 FILLER_ASAP7_75t_R FILLER_258_1239 ();
 DECAPx4_ASAP7_75t_R FILLER_258_1244 ();
 FILLER_ASAP7_75t_R FILLER_258_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_258_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1352 ();
 DECAPx4_ASAP7_75t_R FILLER_258_1374 ();
 FILLER_ASAP7_75t_R FILLER_258_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_258_1388 ();
 FILLER_ASAP7_75t_R FILLER_258_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_259_2 ();
 DECAPx10_ASAP7_75t_R FILLER_259_24 ();
 DECAPx10_ASAP7_75t_R FILLER_259_46 ();
 DECAPx10_ASAP7_75t_R FILLER_259_68 ();
 DECAPx10_ASAP7_75t_R FILLER_259_90 ();
 DECAPx10_ASAP7_75t_R FILLER_259_112 ();
 DECAPx10_ASAP7_75t_R FILLER_259_134 ();
 DECAPx10_ASAP7_75t_R FILLER_259_156 ();
 DECAPx10_ASAP7_75t_R FILLER_259_178 ();
 DECAPx10_ASAP7_75t_R FILLER_259_200 ();
 DECAPx10_ASAP7_75t_R FILLER_259_222 ();
 DECAPx10_ASAP7_75t_R FILLER_259_244 ();
 DECAPx10_ASAP7_75t_R FILLER_259_266 ();
 DECAPx10_ASAP7_75t_R FILLER_259_288 ();
 DECAPx10_ASAP7_75t_R FILLER_259_310 ();
 DECAPx10_ASAP7_75t_R FILLER_259_332 ();
 DECAPx10_ASAP7_75t_R FILLER_259_354 ();
 DECAPx2_ASAP7_75t_R FILLER_259_376 ();
 FILLER_ASAP7_75t_R FILLER_259_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_384 ();
 DECAPx1_ASAP7_75t_R FILLER_259_406 ();
 DECAPx4_ASAP7_75t_R FILLER_259_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_428 ();
 DECAPx10_ASAP7_75t_R FILLER_259_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_461 ();
 DECAPx1_ASAP7_75t_R FILLER_259_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_472 ();
 DECAPx2_ASAP7_75t_R FILLER_259_479 ();
 FILLER_ASAP7_75t_R FILLER_259_485 ();
 DECAPx4_ASAP7_75t_R FILLER_259_493 ();
 FILLER_ASAP7_75t_R FILLER_259_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_505 ();
 DECAPx2_ASAP7_75t_R FILLER_259_520 ();
 FILLER_ASAP7_75t_R FILLER_259_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_528 ();
 DECAPx4_ASAP7_75t_R FILLER_259_534 ();
 FILLER_ASAP7_75t_R FILLER_259_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_546 ();
 FILLER_ASAP7_75t_R FILLER_259_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_562 ();
 DECAPx2_ASAP7_75t_R FILLER_259_592 ();
 DECAPx6_ASAP7_75t_R FILLER_259_604 ();
 DECAPx2_ASAP7_75t_R FILLER_259_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_624 ();
 FILLER_ASAP7_75t_R FILLER_259_631 ();
 FILLER_ASAP7_75t_R FILLER_259_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_647 ();
 DECAPx2_ASAP7_75t_R FILLER_259_656 ();
 FILLER_ASAP7_75t_R FILLER_259_662 ();
 DECAPx2_ASAP7_75t_R FILLER_259_753 ();
 FILLER_ASAP7_75t_R FILLER_259_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_764 ();
 DECAPx10_ASAP7_75t_R FILLER_259_814 ();
 DECAPx10_ASAP7_75t_R FILLER_259_836 ();
 DECAPx2_ASAP7_75t_R FILLER_259_858 ();
 FILLER_ASAP7_75t_R FILLER_259_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_866 ();
 FILLER_ASAP7_75t_R FILLER_259_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_875 ();
 DECAPx2_ASAP7_75t_R FILLER_259_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_892 ();
 DECAPx10_ASAP7_75t_R FILLER_259_896 ();
 DECAPx2_ASAP7_75t_R FILLER_259_918 ();
 DECAPx10_ASAP7_75t_R FILLER_259_934 ();
 FILLER_ASAP7_75t_R FILLER_259_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_958 ();
 DECAPx1_ASAP7_75t_R FILLER_259_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_984 ();
 DECAPx10_ASAP7_75t_R FILLER_259_999 ();
 DECAPx4_ASAP7_75t_R FILLER_259_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_259_1058 ();
 FILLER_ASAP7_75t_R FILLER_259_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_259_1079 ();
 FILLER_ASAP7_75t_R FILLER_259_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_259_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_259_1161 ();
 FILLER_ASAP7_75t_R FILLER_259_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1184 ();
 FILLER_ASAP7_75t_R FILLER_259_1195 ();
 DECAPx6_ASAP7_75t_R FILLER_259_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_259_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1377 ();
 DECAPx2_ASAP7_75t_R FILLER_259_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_260_2 ();
 DECAPx10_ASAP7_75t_R FILLER_260_24 ();
 DECAPx10_ASAP7_75t_R FILLER_260_46 ();
 DECAPx10_ASAP7_75t_R FILLER_260_68 ();
 DECAPx10_ASAP7_75t_R FILLER_260_90 ();
 DECAPx10_ASAP7_75t_R FILLER_260_112 ();
 DECAPx10_ASAP7_75t_R FILLER_260_134 ();
 DECAPx10_ASAP7_75t_R FILLER_260_156 ();
 DECAPx10_ASAP7_75t_R FILLER_260_178 ();
 DECAPx10_ASAP7_75t_R FILLER_260_200 ();
 DECAPx10_ASAP7_75t_R FILLER_260_222 ();
 DECAPx10_ASAP7_75t_R FILLER_260_244 ();
 DECAPx10_ASAP7_75t_R FILLER_260_266 ();
 DECAPx10_ASAP7_75t_R FILLER_260_288 ();
 DECAPx10_ASAP7_75t_R FILLER_260_310 ();
 DECAPx10_ASAP7_75t_R FILLER_260_332 ();
 DECAPx10_ASAP7_75t_R FILLER_260_354 ();
 DECAPx10_ASAP7_75t_R FILLER_260_376 ();
 FILLER_ASAP7_75t_R FILLER_260_405 ();
 DECAPx1_ASAP7_75t_R FILLER_260_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_453 ();
 DECAPx1_ASAP7_75t_R FILLER_260_487 ();
 DECAPx10_ASAP7_75t_R FILLER_260_498 ();
 DECAPx2_ASAP7_75t_R FILLER_260_520 ();
 DECAPx1_ASAP7_75t_R FILLER_260_534 ();
 FILLER_ASAP7_75t_R FILLER_260_550 ();
 DECAPx6_ASAP7_75t_R FILLER_260_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_574 ();
 DECAPx10_ASAP7_75t_R FILLER_260_583 ();
 DECAPx1_ASAP7_75t_R FILLER_260_605 ();
 DECAPx6_ASAP7_75t_R FILLER_260_622 ();
 DECAPx2_ASAP7_75t_R FILLER_260_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_642 ();
 DECAPx2_ASAP7_75t_R FILLER_260_670 ();
 FILLER_ASAP7_75t_R FILLER_260_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_678 ();
 DECAPx6_ASAP7_75t_R FILLER_260_691 ();
 FILLER_ASAP7_75t_R FILLER_260_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_719 ();
 DECAPx4_ASAP7_75t_R FILLER_260_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_774 ();
 DECAPx1_ASAP7_75t_R FILLER_260_786 ();
 DECAPx4_ASAP7_75t_R FILLER_260_824 ();
 DECAPx10_ASAP7_75t_R FILLER_260_840 ();
 DECAPx4_ASAP7_75t_R FILLER_260_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_890 ();
 DECAPx10_ASAP7_75t_R FILLER_260_908 ();
 DECAPx10_ASAP7_75t_R FILLER_260_930 ();
 DECAPx2_ASAP7_75t_R FILLER_260_952 ();
 FILLER_ASAP7_75t_R FILLER_260_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_960 ();
 DECAPx1_ASAP7_75t_R FILLER_260_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_986 ();
 DECAPx2_ASAP7_75t_R FILLER_260_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_260_1027 ();
 FILLER_ASAP7_75t_R FILLER_260_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1043 ();
 FILLER_ASAP7_75t_R FILLER_260_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_260_1141 ();
 FILLER_ASAP7_75t_R FILLER_260_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_260_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_260_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_260_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_260_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_260_1239 ();
 FILLER_ASAP7_75t_R FILLER_260_1253 ();
 DECAPx4_ASAP7_75t_R FILLER_260_1281 ();
 DECAPx2_ASAP7_75t_R FILLER_260_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_260_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_260_1381 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_260_1388 ();
 FILLER_ASAP7_75t_R FILLER_260_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_261_2 ();
 DECAPx10_ASAP7_75t_R FILLER_261_24 ();
 DECAPx10_ASAP7_75t_R FILLER_261_46 ();
 DECAPx10_ASAP7_75t_R FILLER_261_68 ();
 DECAPx10_ASAP7_75t_R FILLER_261_90 ();
 DECAPx10_ASAP7_75t_R FILLER_261_112 ();
 DECAPx10_ASAP7_75t_R FILLER_261_134 ();
 DECAPx10_ASAP7_75t_R FILLER_261_156 ();
 DECAPx10_ASAP7_75t_R FILLER_261_178 ();
 DECAPx10_ASAP7_75t_R FILLER_261_200 ();
 DECAPx10_ASAP7_75t_R FILLER_261_222 ();
 DECAPx10_ASAP7_75t_R FILLER_261_244 ();
 DECAPx10_ASAP7_75t_R FILLER_261_266 ();
 DECAPx10_ASAP7_75t_R FILLER_261_288 ();
 DECAPx10_ASAP7_75t_R FILLER_261_310 ();
 DECAPx10_ASAP7_75t_R FILLER_261_332 ();
 DECAPx10_ASAP7_75t_R FILLER_261_354 ();
 DECAPx6_ASAP7_75t_R FILLER_261_376 ();
 DECAPx2_ASAP7_75t_R FILLER_261_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_396 ();
 FILLER_ASAP7_75t_R FILLER_261_404 ();
 FILLER_ASAP7_75t_R FILLER_261_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_424 ();
 FILLER_ASAP7_75t_R FILLER_261_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_439 ();
 DECAPx10_ASAP7_75t_R FILLER_261_468 ();
 DECAPx10_ASAP7_75t_R FILLER_261_490 ();
 FILLER_ASAP7_75t_R FILLER_261_512 ();
 DECAPx2_ASAP7_75t_R FILLER_261_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_550 ();
 DECAPx6_ASAP7_75t_R FILLER_261_557 ();
 DECAPx4_ASAP7_75t_R FILLER_261_579 ();
 FILLER_ASAP7_75t_R FILLER_261_589 ();
 DECAPx2_ASAP7_75t_R FILLER_261_597 ();
 FILLER_ASAP7_75t_R FILLER_261_603 ();
 DECAPx2_ASAP7_75t_R FILLER_261_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_635 ();
 FILLER_ASAP7_75t_R FILLER_261_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_644 ();
 FILLER_ASAP7_75t_R FILLER_261_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_660 ();
 DECAPx6_ASAP7_75t_R FILLER_261_680 ();
 FILLER_ASAP7_75t_R FILLER_261_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_696 ();
 DECAPx6_ASAP7_75t_R FILLER_261_703 ();
 DECAPx2_ASAP7_75t_R FILLER_261_717 ();
 DECAPx4_ASAP7_75t_R FILLER_261_729 ();
 FILLER_ASAP7_75t_R FILLER_261_739 ();
 FILLER_ASAP7_75t_R FILLER_261_744 ();
 DECAPx4_ASAP7_75t_R FILLER_261_754 ();
 FILLER_ASAP7_75t_R FILLER_261_764 ();
 DECAPx2_ASAP7_75t_R FILLER_261_799 ();
 DECAPx1_ASAP7_75t_R FILLER_261_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_812 ();
 FILLER_ASAP7_75t_R FILLER_261_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_844 ();
 FILLER_ASAP7_75t_R FILLER_261_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_857 ();
 DECAPx2_ASAP7_75t_R FILLER_261_868 ();
 FILLER_ASAP7_75t_R FILLER_261_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_876 ();
 DECAPx1_ASAP7_75t_R FILLER_261_929 ();
 FILLER_ASAP7_75t_R FILLER_261_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_955 ();
 DECAPx6_ASAP7_75t_R FILLER_261_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_980 ();
 DECAPx6_ASAP7_75t_R FILLER_261_991 ();
 FILLER_ASAP7_75t_R FILLER_261_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_261_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1046 ();
 FILLER_ASAP7_75t_R FILLER_261_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_261_1073 ();
 FILLER_ASAP7_75t_R FILLER_261_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_261_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_261_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_261_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_261_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1252 ();
 FILLER_ASAP7_75t_R FILLER_261_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1359 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1381 ();
 FILLER_ASAP7_75t_R FILLER_261_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_262_2 ();
 DECAPx10_ASAP7_75t_R FILLER_262_24 ();
 DECAPx10_ASAP7_75t_R FILLER_262_46 ();
 DECAPx10_ASAP7_75t_R FILLER_262_68 ();
 DECAPx10_ASAP7_75t_R FILLER_262_90 ();
 DECAPx10_ASAP7_75t_R FILLER_262_112 ();
 DECAPx10_ASAP7_75t_R FILLER_262_134 ();
 DECAPx10_ASAP7_75t_R FILLER_262_156 ();
 DECAPx10_ASAP7_75t_R FILLER_262_178 ();
 DECAPx10_ASAP7_75t_R FILLER_262_200 ();
 DECAPx10_ASAP7_75t_R FILLER_262_222 ();
 DECAPx10_ASAP7_75t_R FILLER_262_244 ();
 DECAPx10_ASAP7_75t_R FILLER_262_266 ();
 DECAPx10_ASAP7_75t_R FILLER_262_288 ();
 DECAPx10_ASAP7_75t_R FILLER_262_310 ();
 DECAPx10_ASAP7_75t_R FILLER_262_332 ();
 DECAPx10_ASAP7_75t_R FILLER_262_354 ();
 DECAPx2_ASAP7_75t_R FILLER_262_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_382 ();
 DECAPx10_ASAP7_75t_R FILLER_262_418 ();
 DECAPx6_ASAP7_75t_R FILLER_262_440 ();
 FILLER_ASAP7_75t_R FILLER_262_454 ();
 DECAPx2_ASAP7_75t_R FILLER_262_470 ();
 FILLER_ASAP7_75t_R FILLER_262_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_500 ();
 DECAPx6_ASAP7_75t_R FILLER_262_507 ();
 FILLER_ASAP7_75t_R FILLER_262_521 ();
 DECAPx2_ASAP7_75t_R FILLER_262_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_541 ();
 DECAPx6_ASAP7_75t_R FILLER_262_550 ();
 FILLER_ASAP7_75t_R FILLER_262_564 ();
 FILLER_ASAP7_75t_R FILLER_262_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_589 ();
 FILLER_ASAP7_75t_R FILLER_262_598 ();
 DECAPx1_ASAP7_75t_R FILLER_262_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_611 ();
 DECAPx2_ASAP7_75t_R FILLER_262_624 ();
 DECAPx6_ASAP7_75t_R FILLER_262_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_665 ();
 DECAPx6_ASAP7_75t_R FILLER_262_674 ();
 DECAPx2_ASAP7_75t_R FILLER_262_688 ();
 DECAPx4_ASAP7_75t_R FILLER_262_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_720 ();
 DECAPx10_ASAP7_75t_R FILLER_262_736 ();
 DECAPx6_ASAP7_75t_R FILLER_262_758 ();
 DECAPx1_ASAP7_75t_R FILLER_262_778 ();
 DECAPx2_ASAP7_75t_R FILLER_262_790 ();
 FILLER_ASAP7_75t_R FILLER_262_796 ();
 DECAPx10_ASAP7_75t_R FILLER_262_801 ();
 DECAPx6_ASAP7_75t_R FILLER_262_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_849 ();
 DECAPx4_ASAP7_75t_R FILLER_262_856 ();
 DECAPx2_ASAP7_75t_R FILLER_262_874 ();
 FILLER_ASAP7_75t_R FILLER_262_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_882 ();
 DECAPx2_ASAP7_75t_R FILLER_262_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_920 ();
 DECAPx4_ASAP7_75t_R FILLER_262_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_938 ();
 DECAPx10_ASAP7_75t_R FILLER_262_960 ();
 DECAPx2_ASAP7_75t_R FILLER_262_982 ();
 FILLER_ASAP7_75t_R FILLER_262_988 ();
 DECAPx4_ASAP7_75t_R FILLER_262_998 ();
 FILLER_ASAP7_75t_R FILLER_262_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_262_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_262_1058 ();
 FILLER_ASAP7_75t_R FILLER_262_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_262_1109 ();
 FILLER_ASAP7_75t_R FILLER_262_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1125 ();
 DECAPx4_ASAP7_75t_R FILLER_262_1139 ();
 FILLER_ASAP7_75t_R FILLER_262_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_262_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_262_1194 ();
 FILLER_ASAP7_75t_R FILLER_262_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_262_1246 ();
 FILLER_ASAP7_75t_R FILLER_262_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_262_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1299 ();
 DECAPx6_ASAP7_75t_R FILLER_262_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_262_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1347 ();
 DECAPx6_ASAP7_75t_R FILLER_262_1369 ();
 FILLER_ASAP7_75t_R FILLER_262_1383 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_262_1388 ();
 FILLER_ASAP7_75t_R FILLER_262_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_263_2 ();
 DECAPx10_ASAP7_75t_R FILLER_263_24 ();
 DECAPx10_ASAP7_75t_R FILLER_263_46 ();
 DECAPx10_ASAP7_75t_R FILLER_263_68 ();
 DECAPx10_ASAP7_75t_R FILLER_263_90 ();
 DECAPx10_ASAP7_75t_R FILLER_263_112 ();
 DECAPx10_ASAP7_75t_R FILLER_263_134 ();
 DECAPx10_ASAP7_75t_R FILLER_263_156 ();
 DECAPx10_ASAP7_75t_R FILLER_263_178 ();
 DECAPx10_ASAP7_75t_R FILLER_263_200 ();
 DECAPx10_ASAP7_75t_R FILLER_263_222 ();
 DECAPx10_ASAP7_75t_R FILLER_263_244 ();
 DECAPx10_ASAP7_75t_R FILLER_263_266 ();
 DECAPx10_ASAP7_75t_R FILLER_263_288 ();
 DECAPx10_ASAP7_75t_R FILLER_263_310 ();
 DECAPx10_ASAP7_75t_R FILLER_263_332 ();
 DECAPx10_ASAP7_75t_R FILLER_263_354 ();
 DECAPx10_ASAP7_75t_R FILLER_263_376 ();
 DECAPx1_ASAP7_75t_R FILLER_263_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_402 ();
 DECAPx6_ASAP7_75t_R FILLER_263_422 ();
 FILLER_ASAP7_75t_R FILLER_263_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_438 ();
 DECAPx4_ASAP7_75t_R FILLER_263_449 ();
 FILLER_ASAP7_75t_R FILLER_263_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_474 ();
 DECAPx2_ASAP7_75t_R FILLER_263_491 ();
 FILLER_ASAP7_75t_R FILLER_263_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_499 ();
 DECAPx2_ASAP7_75t_R FILLER_263_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_522 ();
 DECAPx1_ASAP7_75t_R FILLER_263_529 ();
 FILLER_ASAP7_75t_R FILLER_263_560 ();
 FILLER_ASAP7_75t_R FILLER_263_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_585 ();
 DECAPx1_ASAP7_75t_R FILLER_263_592 ();
 DECAPx6_ASAP7_75t_R FILLER_263_604 ();
 DECAPx1_ASAP7_75t_R FILLER_263_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_622 ();
 DECAPx2_ASAP7_75t_R FILLER_263_626 ();
 FILLER_ASAP7_75t_R FILLER_263_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_634 ();
 DECAPx10_ASAP7_75t_R FILLER_263_643 ();
 DECAPx2_ASAP7_75t_R FILLER_263_665 ();
 DECAPx2_ASAP7_75t_R FILLER_263_679 ();
 DECAPx1_ASAP7_75t_R FILLER_263_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_695 ();
 DECAPx2_ASAP7_75t_R FILLER_263_702 ();
 FILLER_ASAP7_75t_R FILLER_263_708 ();
 DECAPx2_ASAP7_75t_R FILLER_263_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_753 ();
 DECAPx6_ASAP7_75t_R FILLER_263_757 ();
 DECAPx1_ASAP7_75t_R FILLER_263_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_775 ();
 DECAPx2_ASAP7_75t_R FILLER_263_810 ();
 FILLER_ASAP7_75t_R FILLER_263_816 ();
 DECAPx1_ASAP7_75t_R FILLER_263_830 ();
 DECAPx4_ASAP7_75t_R FILLER_263_864 ();
 FILLER_ASAP7_75t_R FILLER_263_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_876 ();
 DECAPx6_ASAP7_75t_R FILLER_263_895 ();
 DECAPx1_ASAP7_75t_R FILLER_263_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_913 ();
 DECAPx1_ASAP7_75t_R FILLER_263_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_934 ();
 DECAPx4_ASAP7_75t_R FILLER_263_947 ();
 FILLER_ASAP7_75t_R FILLER_263_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_959 ();
 DECAPx1_ASAP7_75t_R FILLER_263_970 ();
 DECAPx4_ASAP7_75t_R FILLER_263_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_990 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_263_1028 ();
 FILLER_ASAP7_75t_R FILLER_263_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_263_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_263_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1089 ();
 FILLER_ASAP7_75t_R FILLER_263_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1106 ();
 FILLER_ASAP7_75t_R FILLER_263_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1135 ();
 FILLER_ASAP7_75t_R FILLER_263_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1194 ();
 FILLER_ASAP7_75t_R FILLER_263_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1217 ();
 FILLER_ASAP7_75t_R FILLER_263_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1349 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1371 ();
 DECAPx4_ASAP7_75t_R FILLER_263_1393 ();
 FILLER_ASAP7_75t_R FILLER_263_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_264_2 ();
 DECAPx10_ASAP7_75t_R FILLER_264_24 ();
 DECAPx10_ASAP7_75t_R FILLER_264_46 ();
 DECAPx10_ASAP7_75t_R FILLER_264_68 ();
 DECAPx10_ASAP7_75t_R FILLER_264_90 ();
 DECAPx10_ASAP7_75t_R FILLER_264_112 ();
 DECAPx10_ASAP7_75t_R FILLER_264_134 ();
 DECAPx10_ASAP7_75t_R FILLER_264_156 ();
 DECAPx10_ASAP7_75t_R FILLER_264_178 ();
 DECAPx10_ASAP7_75t_R FILLER_264_200 ();
 DECAPx10_ASAP7_75t_R FILLER_264_222 ();
 DECAPx10_ASAP7_75t_R FILLER_264_244 ();
 DECAPx10_ASAP7_75t_R FILLER_264_266 ();
 DECAPx10_ASAP7_75t_R FILLER_264_288 ();
 DECAPx10_ASAP7_75t_R FILLER_264_310 ();
 DECAPx10_ASAP7_75t_R FILLER_264_332 ();
 DECAPx10_ASAP7_75t_R FILLER_264_354 ();
 DECAPx4_ASAP7_75t_R FILLER_264_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_386 ();
 FILLER_ASAP7_75t_R FILLER_264_408 ();
 FILLER_ASAP7_75t_R FILLER_264_420 ();
 DECAPx1_ASAP7_75t_R FILLER_264_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_432 ();
 DECAPx1_ASAP7_75t_R FILLER_264_464 ();
 FILLER_ASAP7_75t_R FILLER_264_488 ();
 FILLER_ASAP7_75t_R FILLER_264_520 ();
 DECAPx2_ASAP7_75t_R FILLER_264_540 ();
 DECAPx2_ASAP7_75t_R FILLER_264_552 ();
 DECAPx1_ASAP7_75t_R FILLER_264_564 ();
 FILLER_ASAP7_75t_R FILLER_264_580 ();
 DECAPx6_ASAP7_75t_R FILLER_264_610 ();
 DECAPx4_ASAP7_75t_R FILLER_264_635 ();
 FILLER_ASAP7_75t_R FILLER_264_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_647 ();
 DECAPx1_ASAP7_75t_R FILLER_264_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_660 ();
 DECAPx10_ASAP7_75t_R FILLER_264_683 ();
 FILLER_ASAP7_75t_R FILLER_264_705 ();
 DECAPx1_ASAP7_75t_R FILLER_264_719 ();
 FILLER_ASAP7_75t_R FILLER_264_737 ();
 DECAPx1_ASAP7_75t_R FILLER_264_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_779 ();
 DECAPx2_ASAP7_75t_R FILLER_264_786 ();
 FILLER_ASAP7_75t_R FILLER_264_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_794 ();
 DECAPx2_ASAP7_75t_R FILLER_264_842 ();
 FILLER_ASAP7_75t_R FILLER_264_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_850 ();
 DECAPx1_ASAP7_75t_R FILLER_264_854 ();
 DECAPx10_ASAP7_75t_R FILLER_264_864 ();
 DECAPx4_ASAP7_75t_R FILLER_264_886 ();
 DECAPx1_ASAP7_75t_R FILLER_264_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_907 ();
 DECAPx10_ASAP7_75t_R FILLER_264_924 ();
 DECAPx1_ASAP7_75t_R FILLER_264_946 ();
 FILLER_ASAP7_75t_R FILLER_264_977 ();
 FILLER_ASAP7_75t_R FILLER_264_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_989 ();
 DECAPx2_ASAP7_75t_R FILLER_264_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1003 ();
 FILLER_ASAP7_75t_R FILLER_264_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_264_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_264_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_264_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_264_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_264_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1189 ();
 FILLER_ASAP7_75t_R FILLER_264_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_264_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_264_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_264_1388 ();
 FILLER_ASAP7_75t_R FILLER_264_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_265_2 ();
 DECAPx10_ASAP7_75t_R FILLER_265_24 ();
 DECAPx10_ASAP7_75t_R FILLER_265_46 ();
 DECAPx10_ASAP7_75t_R FILLER_265_68 ();
 DECAPx10_ASAP7_75t_R FILLER_265_90 ();
 DECAPx10_ASAP7_75t_R FILLER_265_112 ();
 DECAPx10_ASAP7_75t_R FILLER_265_134 ();
 DECAPx10_ASAP7_75t_R FILLER_265_156 ();
 DECAPx10_ASAP7_75t_R FILLER_265_178 ();
 DECAPx10_ASAP7_75t_R FILLER_265_200 ();
 DECAPx10_ASAP7_75t_R FILLER_265_222 ();
 DECAPx10_ASAP7_75t_R FILLER_265_244 ();
 DECAPx10_ASAP7_75t_R FILLER_265_266 ();
 DECAPx10_ASAP7_75t_R FILLER_265_288 ();
 DECAPx10_ASAP7_75t_R FILLER_265_310 ();
 DECAPx10_ASAP7_75t_R FILLER_265_332 ();
 DECAPx10_ASAP7_75t_R FILLER_265_354 ();
 DECAPx10_ASAP7_75t_R FILLER_265_376 ();
 DECAPx2_ASAP7_75t_R FILLER_265_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_404 ();
 DECAPx1_ASAP7_75t_R FILLER_265_426 ();
 DECAPx1_ASAP7_75t_R FILLER_265_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_462 ();
 DECAPx10_ASAP7_75t_R FILLER_265_482 ();
 DECAPx2_ASAP7_75t_R FILLER_265_516 ();
 DECAPx2_ASAP7_75t_R FILLER_265_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_534 ();
 DECAPx2_ASAP7_75t_R FILLER_265_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_544 ();
 DECAPx1_ASAP7_75t_R FILLER_265_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_573 ();
 DECAPx2_ASAP7_75t_R FILLER_265_580 ();
 FILLER_ASAP7_75t_R FILLER_265_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_595 ();
 DECAPx2_ASAP7_75t_R FILLER_265_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_608 ();
 FILLER_ASAP7_75t_R FILLER_265_617 ();
 DECAPx2_ASAP7_75t_R FILLER_265_640 ();
 FILLER_ASAP7_75t_R FILLER_265_646 ();
 DECAPx2_ASAP7_75t_R FILLER_265_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_683 ();
 FILLER_ASAP7_75t_R FILLER_265_695 ();
 FILLER_ASAP7_75t_R FILLER_265_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_707 ();
 FILLER_ASAP7_75t_R FILLER_265_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_727 ();
 DECAPx10_ASAP7_75t_R FILLER_265_734 ();
 DECAPx2_ASAP7_75t_R FILLER_265_788 ();
 FILLER_ASAP7_75t_R FILLER_265_822 ();
 DECAPx1_ASAP7_75t_R FILLER_265_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_847 ();
 DECAPx1_ASAP7_75t_R FILLER_265_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_902 ();
 DECAPx1_ASAP7_75t_R FILLER_265_932 ();
 DECAPx2_ASAP7_75t_R FILLER_265_943 ();
 FILLER_ASAP7_75t_R FILLER_265_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_963 ();
 FILLER_ASAP7_75t_R FILLER_265_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1043 ();
 FILLER_ASAP7_75t_R FILLER_265_1050 ();
 FILLER_ASAP7_75t_R FILLER_265_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1088 ();
 DECAPx6_ASAP7_75t_R FILLER_265_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_265_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_265_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_265_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_265_1397 ();
 FILLER_ASAP7_75t_R FILLER_265_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_266_2 ();
 DECAPx10_ASAP7_75t_R FILLER_266_24 ();
 DECAPx10_ASAP7_75t_R FILLER_266_46 ();
 DECAPx10_ASAP7_75t_R FILLER_266_68 ();
 DECAPx10_ASAP7_75t_R FILLER_266_90 ();
 DECAPx10_ASAP7_75t_R FILLER_266_112 ();
 DECAPx10_ASAP7_75t_R FILLER_266_134 ();
 DECAPx10_ASAP7_75t_R FILLER_266_156 ();
 DECAPx10_ASAP7_75t_R FILLER_266_178 ();
 DECAPx10_ASAP7_75t_R FILLER_266_200 ();
 DECAPx10_ASAP7_75t_R FILLER_266_222 ();
 DECAPx10_ASAP7_75t_R FILLER_266_244 ();
 DECAPx10_ASAP7_75t_R FILLER_266_266 ();
 DECAPx10_ASAP7_75t_R FILLER_266_288 ();
 DECAPx10_ASAP7_75t_R FILLER_266_310 ();
 DECAPx10_ASAP7_75t_R FILLER_266_332 ();
 DECAPx10_ASAP7_75t_R FILLER_266_354 ();
 DECAPx10_ASAP7_75t_R FILLER_266_376 ();
 DECAPx6_ASAP7_75t_R FILLER_266_404 ();
 FILLER_ASAP7_75t_R FILLER_266_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_420 ();
 FILLER_ASAP7_75t_R FILLER_266_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_461 ();
 DECAPx10_ASAP7_75t_R FILLER_266_464 ();
 DECAPx6_ASAP7_75t_R FILLER_266_486 ();
 FILLER_ASAP7_75t_R FILLER_266_500 ();
 DECAPx1_ASAP7_75t_R FILLER_266_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_576 ();
 FILLER_ASAP7_75t_R FILLER_266_583 ();
 DECAPx1_ASAP7_75t_R FILLER_266_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_611 ();
 DECAPx1_ASAP7_75t_R FILLER_266_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_627 ();
 DECAPx4_ASAP7_75t_R FILLER_266_634 ();
 DECAPx2_ASAP7_75t_R FILLER_266_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_659 ();
 DECAPx1_ASAP7_75t_R FILLER_266_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_685 ();
 DECAPx6_ASAP7_75t_R FILLER_266_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_727 ();
 FILLER_ASAP7_75t_R FILLER_266_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_773 ();
 DECAPx10_ASAP7_75t_R FILLER_266_783 ();
 DECAPx2_ASAP7_75t_R FILLER_266_818 ();
 FILLER_ASAP7_75t_R FILLER_266_824 ();
 DECAPx2_ASAP7_75t_R FILLER_266_833 ();
 FILLER_ASAP7_75t_R FILLER_266_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_841 ();
 DECAPx4_ASAP7_75t_R FILLER_266_848 ();
 FILLER_ASAP7_75t_R FILLER_266_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_860 ();
 DECAPx1_ASAP7_75t_R FILLER_266_883 ();
 DECAPx2_ASAP7_75t_R FILLER_266_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_920 ();
 DECAPx2_ASAP7_75t_R FILLER_266_929 ();
 FILLER_ASAP7_75t_R FILLER_266_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_949 ();
 DECAPx1_ASAP7_75t_R FILLER_266_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_971 ();
 DECAPx2_ASAP7_75t_R FILLER_266_985 ();
 FILLER_ASAP7_75t_R FILLER_266_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_993 ();
 DECAPx2_ASAP7_75t_R FILLER_266_1000 ();
 FILLER_ASAP7_75t_R FILLER_266_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_266_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1037 ();
 FILLER_ASAP7_75t_R FILLER_266_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1050 ();
 DECAPx4_ASAP7_75t_R FILLER_266_1058 ();
 FILLER_ASAP7_75t_R FILLER_266_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_266_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_266_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_266_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1119 ();
 FILLER_ASAP7_75t_R FILLER_266_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1143 ();
 FILLER_ASAP7_75t_R FILLER_266_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_266_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_266_1209 ();
 FILLER_ASAP7_75t_R FILLER_266_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1362 ();
 FILLER_ASAP7_75t_R FILLER_266_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_266_1388 ();
 FILLER_ASAP7_75t_R FILLER_266_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_267_2 ();
 DECAPx10_ASAP7_75t_R FILLER_267_24 ();
 DECAPx10_ASAP7_75t_R FILLER_267_46 ();
 DECAPx10_ASAP7_75t_R FILLER_267_68 ();
 DECAPx10_ASAP7_75t_R FILLER_267_90 ();
 DECAPx10_ASAP7_75t_R FILLER_267_112 ();
 DECAPx10_ASAP7_75t_R FILLER_267_134 ();
 DECAPx10_ASAP7_75t_R FILLER_267_156 ();
 DECAPx10_ASAP7_75t_R FILLER_267_178 ();
 DECAPx10_ASAP7_75t_R FILLER_267_200 ();
 DECAPx10_ASAP7_75t_R FILLER_267_222 ();
 DECAPx10_ASAP7_75t_R FILLER_267_244 ();
 DECAPx10_ASAP7_75t_R FILLER_267_266 ();
 DECAPx10_ASAP7_75t_R FILLER_267_288 ();
 DECAPx10_ASAP7_75t_R FILLER_267_310 ();
 DECAPx10_ASAP7_75t_R FILLER_267_332 ();
 DECAPx10_ASAP7_75t_R FILLER_267_354 ();
 DECAPx6_ASAP7_75t_R FILLER_267_376 ();
 DECAPx2_ASAP7_75t_R FILLER_267_390 ();
 FILLER_ASAP7_75t_R FILLER_267_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_405 ();
 DECAPx4_ASAP7_75t_R FILLER_267_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_447 ();
 DECAPx2_ASAP7_75t_R FILLER_267_469 ();
 FILLER_ASAP7_75t_R FILLER_267_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_499 ();
 FILLER_ASAP7_75t_R FILLER_267_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_515 ();
 FILLER_ASAP7_75t_R FILLER_267_537 ();
 DECAPx4_ASAP7_75t_R FILLER_267_547 ();
 DECAPx4_ASAP7_75t_R FILLER_267_565 ();
 FILLER_ASAP7_75t_R FILLER_267_575 ();
 DECAPx1_ASAP7_75t_R FILLER_267_591 ();
 DECAPx10_ASAP7_75t_R FILLER_267_601 ();
 FILLER_ASAP7_75t_R FILLER_267_623 ();
 DECAPx1_ASAP7_75t_R FILLER_267_631 ();
 DECAPx4_ASAP7_75t_R FILLER_267_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_669 ();
 FILLER_ASAP7_75t_R FILLER_267_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_698 ();
 DECAPx6_ASAP7_75t_R FILLER_267_707 ();
 FILLER_ASAP7_75t_R FILLER_267_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_747 ();
 DECAPx2_ASAP7_75t_R FILLER_267_761 ();
 FILLER_ASAP7_75t_R FILLER_267_767 ();
 FILLER_ASAP7_75t_R FILLER_267_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_803 ();
 FILLER_ASAP7_75t_R FILLER_267_834 ();
 DECAPx4_ASAP7_75t_R FILLER_267_856 ();
 FILLER_ASAP7_75t_R FILLER_267_866 ();
 DECAPx4_ASAP7_75t_R FILLER_267_882 ();
 DECAPx2_ASAP7_75t_R FILLER_267_898 ();
 FILLER_ASAP7_75t_R FILLER_267_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_906 ();
 DECAPx4_ASAP7_75t_R FILLER_267_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_923 ();
 DECAPx2_ASAP7_75t_R FILLER_267_926 ();
 FILLER_ASAP7_75t_R FILLER_267_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_934 ();
 FILLER_ASAP7_75t_R FILLER_267_942 ();
 FILLER_ASAP7_75t_R FILLER_267_950 ();
 DECAPx10_ASAP7_75t_R FILLER_267_964 ();
 DECAPx10_ASAP7_75t_R FILLER_267_986 ();
 FILLER_ASAP7_75t_R FILLER_267_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_267_1039 ();
 FILLER_ASAP7_75t_R FILLER_267_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_267_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1073 ();
 FILLER_ASAP7_75t_R FILLER_267_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_267_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_267_1162 ();
 FILLER_ASAP7_75t_R FILLER_267_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1358 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1380 ();
 FILLER_ASAP7_75t_R FILLER_267_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_268_2 ();
 DECAPx10_ASAP7_75t_R FILLER_268_24 ();
 DECAPx10_ASAP7_75t_R FILLER_268_46 ();
 DECAPx10_ASAP7_75t_R FILLER_268_68 ();
 DECAPx10_ASAP7_75t_R FILLER_268_90 ();
 DECAPx10_ASAP7_75t_R FILLER_268_112 ();
 DECAPx10_ASAP7_75t_R FILLER_268_134 ();
 DECAPx10_ASAP7_75t_R FILLER_268_156 ();
 DECAPx10_ASAP7_75t_R FILLER_268_178 ();
 DECAPx10_ASAP7_75t_R FILLER_268_200 ();
 DECAPx10_ASAP7_75t_R FILLER_268_222 ();
 DECAPx10_ASAP7_75t_R FILLER_268_244 ();
 DECAPx10_ASAP7_75t_R FILLER_268_266 ();
 DECAPx10_ASAP7_75t_R FILLER_268_288 ();
 DECAPx10_ASAP7_75t_R FILLER_268_310 ();
 DECAPx10_ASAP7_75t_R FILLER_268_332 ();
 DECAPx10_ASAP7_75t_R FILLER_268_354 ();
 DECAPx2_ASAP7_75t_R FILLER_268_376 ();
 FILLER_ASAP7_75t_R FILLER_268_437 ();
 FILLER_ASAP7_75t_R FILLER_268_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_461 ();
 FILLER_ASAP7_75t_R FILLER_268_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_466 ();
 DECAPx1_ASAP7_75t_R FILLER_268_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_606 ();
 DECAPx2_ASAP7_75t_R FILLER_268_636 ();
 DECAPx2_ASAP7_75t_R FILLER_268_650 ();
 DECAPx6_ASAP7_75t_R FILLER_268_664 ();
 FILLER_ASAP7_75t_R FILLER_268_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_721 ();
 DECAPx10_ASAP7_75t_R FILLER_268_738 ();
 DECAPx6_ASAP7_75t_R FILLER_268_760 ();
 DECAPx1_ASAP7_75t_R FILLER_268_774 ();
 FILLER_ASAP7_75t_R FILLER_268_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_808 ();
 DECAPx1_ASAP7_75t_R FILLER_268_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_841 ();
 DECAPx2_ASAP7_75t_R FILLER_268_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_863 ();
 DECAPx2_ASAP7_75t_R FILLER_268_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_882 ();
 FILLER_ASAP7_75t_R FILLER_268_896 ();
 DECAPx6_ASAP7_75t_R FILLER_268_906 ();
 DECAPx4_ASAP7_75t_R FILLER_268_926 ();
 FILLER_ASAP7_75t_R FILLER_268_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_957 ();
 DECAPx1_ASAP7_75t_R FILLER_268_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_970 ();
 DECAPx4_ASAP7_75t_R FILLER_268_981 ();
 DECAPx2_ASAP7_75t_R FILLER_268_997 ();
 FILLER_ASAP7_75t_R FILLER_268_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_268_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_268_1039 ();
 FILLER_ASAP7_75t_R FILLER_268_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_268_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_268_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_268_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_268_1161 ();
 FILLER_ASAP7_75t_R FILLER_268_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1178 ();
 FILLER_ASAP7_75t_R FILLER_268_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_268_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_268_1378 ();
 FILLER_ASAP7_75t_R FILLER_268_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_268_1388 ();
 FILLER_ASAP7_75t_R FILLER_268_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_269_2 ();
 DECAPx10_ASAP7_75t_R FILLER_269_24 ();
 DECAPx10_ASAP7_75t_R FILLER_269_46 ();
 DECAPx10_ASAP7_75t_R FILLER_269_68 ();
 DECAPx10_ASAP7_75t_R FILLER_269_90 ();
 DECAPx10_ASAP7_75t_R FILLER_269_112 ();
 DECAPx10_ASAP7_75t_R FILLER_269_134 ();
 DECAPx10_ASAP7_75t_R FILLER_269_156 ();
 DECAPx10_ASAP7_75t_R FILLER_269_178 ();
 DECAPx10_ASAP7_75t_R FILLER_269_200 ();
 DECAPx10_ASAP7_75t_R FILLER_269_222 ();
 DECAPx10_ASAP7_75t_R FILLER_269_244 ();
 DECAPx10_ASAP7_75t_R FILLER_269_266 ();
 DECAPx10_ASAP7_75t_R FILLER_269_288 ();
 DECAPx10_ASAP7_75t_R FILLER_269_310 ();
 DECAPx10_ASAP7_75t_R FILLER_269_332 ();
 DECAPx10_ASAP7_75t_R FILLER_269_354 ();
 DECAPx10_ASAP7_75t_R FILLER_269_376 ();
 DECAPx1_ASAP7_75t_R FILLER_269_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_431 ();
 DECAPx1_ASAP7_75t_R FILLER_269_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_452 ();
 DECAPx2_ASAP7_75t_R FILLER_269_469 ();
 FILLER_ASAP7_75t_R FILLER_269_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_477 ();
 DECAPx1_ASAP7_75t_R FILLER_269_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_496 ();
 DECAPx6_ASAP7_75t_R FILLER_269_515 ();
 DECAPx1_ASAP7_75t_R FILLER_269_529 ();
 DECAPx6_ASAP7_75t_R FILLER_269_547 ();
 DECAPx2_ASAP7_75t_R FILLER_269_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_594 ();
 DECAPx6_ASAP7_75t_R FILLER_269_601 ();
 FILLER_ASAP7_75t_R FILLER_269_615 ();
 DECAPx1_ASAP7_75t_R FILLER_269_644 ();
 DECAPx2_ASAP7_75t_R FILLER_269_669 ();
 DECAPx10_ASAP7_75t_R FILLER_269_696 ();
 DECAPx4_ASAP7_75t_R FILLER_269_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_728 ();
 DECAPx2_ASAP7_75t_R FILLER_269_737 ();
 FILLER_ASAP7_75t_R FILLER_269_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_745 ();
 DECAPx1_ASAP7_75t_R FILLER_269_786 ();
 DECAPx4_ASAP7_75t_R FILLER_269_798 ();
 FILLER_ASAP7_75t_R FILLER_269_808 ();
 DECAPx1_ASAP7_75t_R FILLER_269_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_826 ();
 FILLER_ASAP7_75t_R FILLER_269_848 ();
 DECAPx2_ASAP7_75t_R FILLER_269_866 ();
 FILLER_ASAP7_75t_R FILLER_269_901 ();
 FILLER_ASAP7_75t_R FILLER_269_912 ();
 FILLER_ASAP7_75t_R FILLER_269_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_944 ();
 DECAPx1_ASAP7_75t_R FILLER_269_951 ();
 DECAPx2_ASAP7_75t_R FILLER_269_976 ();
 FILLER_ASAP7_75t_R FILLER_269_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1002 ();
 FILLER_ASAP7_75t_R FILLER_269_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_269_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_269_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_269_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_269_1136 ();
 FILLER_ASAP7_75t_R FILLER_269_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1152 ();
 FILLER_ASAP7_75t_R FILLER_269_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1169 ();
 FILLER_ASAP7_75t_R FILLER_269_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1200 ();
 DECAPx4_ASAP7_75t_R FILLER_269_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1366 ();
 DECAPx6_ASAP7_75t_R FILLER_269_1388 ();
 FILLER_ASAP7_75t_R FILLER_269_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_270_2 ();
 DECAPx10_ASAP7_75t_R FILLER_270_24 ();
 DECAPx10_ASAP7_75t_R FILLER_270_46 ();
 DECAPx10_ASAP7_75t_R FILLER_270_68 ();
 DECAPx10_ASAP7_75t_R FILLER_270_90 ();
 DECAPx10_ASAP7_75t_R FILLER_270_112 ();
 DECAPx10_ASAP7_75t_R FILLER_270_134 ();
 DECAPx10_ASAP7_75t_R FILLER_270_156 ();
 DECAPx10_ASAP7_75t_R FILLER_270_178 ();
 DECAPx10_ASAP7_75t_R FILLER_270_200 ();
 DECAPx10_ASAP7_75t_R FILLER_270_222 ();
 DECAPx10_ASAP7_75t_R FILLER_270_244 ();
 DECAPx10_ASAP7_75t_R FILLER_270_266 ();
 DECAPx10_ASAP7_75t_R FILLER_270_288 ();
 DECAPx10_ASAP7_75t_R FILLER_270_310 ();
 DECAPx10_ASAP7_75t_R FILLER_270_332 ();
 DECAPx10_ASAP7_75t_R FILLER_270_354 ();
 DECAPx10_ASAP7_75t_R FILLER_270_376 ();
 DECAPx4_ASAP7_75t_R FILLER_270_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_408 ();
 DECAPx1_ASAP7_75t_R FILLER_270_419 ();
 DECAPx2_ASAP7_75t_R FILLER_270_456 ();
 DECAPx10_ASAP7_75t_R FILLER_270_464 ();
 DECAPx6_ASAP7_75t_R FILLER_270_486 ();
 DECAPx1_ASAP7_75t_R FILLER_270_500 ();
 DECAPx10_ASAP7_75t_R FILLER_270_511 ();
 FILLER_ASAP7_75t_R FILLER_270_533 ();
 DECAPx10_ASAP7_75t_R FILLER_270_542 ();
 DECAPx10_ASAP7_75t_R FILLER_270_564 ();
 DECAPx10_ASAP7_75t_R FILLER_270_586 ();
 DECAPx6_ASAP7_75t_R FILLER_270_608 ();
 DECAPx1_ASAP7_75t_R FILLER_270_622 ();
 DECAPx10_ASAP7_75t_R FILLER_270_634 ();
 DECAPx10_ASAP7_75t_R FILLER_270_669 ();
 DECAPx1_ASAP7_75t_R FILLER_270_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_695 ();
 DECAPx2_ASAP7_75t_R FILLER_270_710 ();
 FILLER_ASAP7_75t_R FILLER_270_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_718 ();
 FILLER_ASAP7_75t_R FILLER_270_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_729 ();
 DECAPx1_ASAP7_75t_R FILLER_270_760 ();
 DECAPx6_ASAP7_75t_R FILLER_270_783 ();
 FILLER_ASAP7_75t_R FILLER_270_797 ();
 DECAPx10_ASAP7_75t_R FILLER_270_805 ();
 DECAPx10_ASAP7_75t_R FILLER_270_827 ();
 DECAPx2_ASAP7_75t_R FILLER_270_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_855 ();
 DECAPx2_ASAP7_75t_R FILLER_270_862 ();
 FILLER_ASAP7_75t_R FILLER_270_868 ();
 FILLER_ASAP7_75t_R FILLER_270_879 ();
 DECAPx6_ASAP7_75t_R FILLER_270_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_911 ();
 DECAPx1_ASAP7_75t_R FILLER_270_933 ();
 DECAPx2_ASAP7_75t_R FILLER_270_945 ();
 FILLER_ASAP7_75t_R FILLER_270_951 ();
 FILLER_ASAP7_75t_R FILLER_270_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_965 ();
 DECAPx1_ASAP7_75t_R FILLER_270_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_988 ();
 DECAPx2_ASAP7_75t_R FILLER_270_1010 ();
 FILLER_ASAP7_75t_R FILLER_270_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_270_1064 ();
 FILLER_ASAP7_75t_R FILLER_270_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_270_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_270_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_270_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_270_1163 ();
 FILLER_ASAP7_75t_R FILLER_270_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_270_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_270_1382 ();
 DECAPx6_ASAP7_75t_R FILLER_270_1388 ();
 FILLER_ASAP7_75t_R FILLER_270_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_271_2 ();
 DECAPx10_ASAP7_75t_R FILLER_271_24 ();
 DECAPx10_ASAP7_75t_R FILLER_271_46 ();
 DECAPx10_ASAP7_75t_R FILLER_271_68 ();
 DECAPx10_ASAP7_75t_R FILLER_271_90 ();
 DECAPx10_ASAP7_75t_R FILLER_271_112 ();
 DECAPx10_ASAP7_75t_R FILLER_271_134 ();
 DECAPx10_ASAP7_75t_R FILLER_271_156 ();
 DECAPx10_ASAP7_75t_R FILLER_271_178 ();
 DECAPx10_ASAP7_75t_R FILLER_271_200 ();
 DECAPx10_ASAP7_75t_R FILLER_271_222 ();
 DECAPx10_ASAP7_75t_R FILLER_271_244 ();
 DECAPx10_ASAP7_75t_R FILLER_271_266 ();
 DECAPx10_ASAP7_75t_R FILLER_271_288 ();
 DECAPx10_ASAP7_75t_R FILLER_271_310 ();
 DECAPx10_ASAP7_75t_R FILLER_271_332 ();
 DECAPx10_ASAP7_75t_R FILLER_271_354 ();
 DECAPx10_ASAP7_75t_R FILLER_271_376 ();
 DECAPx10_ASAP7_75t_R FILLER_271_398 ();
 DECAPx10_ASAP7_75t_R FILLER_271_420 ();
 DECAPx6_ASAP7_75t_R FILLER_271_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_456 ();
 DECAPx1_ASAP7_75t_R FILLER_271_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_475 ();
 DECAPx2_ASAP7_75t_R FILLER_271_496 ();
 FILLER_ASAP7_75t_R FILLER_271_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_504 ();
 DECAPx6_ASAP7_75t_R FILLER_271_519 ();
 DECAPx1_ASAP7_75t_R FILLER_271_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_537 ();
 DECAPx4_ASAP7_75t_R FILLER_271_545 ();
 DECAPx4_ASAP7_75t_R FILLER_271_562 ();
 FILLER_ASAP7_75t_R FILLER_271_572 ();
 DECAPx6_ASAP7_75t_R FILLER_271_581 ();
 FILLER_ASAP7_75t_R FILLER_271_598 ();
 DECAPx4_ASAP7_75t_R FILLER_271_614 ();
 DECAPx4_ASAP7_75t_R FILLER_271_631 ();
 DECAPx1_ASAP7_75t_R FILLER_271_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_652 ();
 DECAPx4_ASAP7_75t_R FILLER_271_656 ();
 DECAPx4_ASAP7_75t_R FILLER_271_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_707 ();
 DECAPx2_ASAP7_75t_R FILLER_271_714 ();
 FILLER_ASAP7_75t_R FILLER_271_720 ();
 DECAPx1_ASAP7_75t_R FILLER_271_738 ();
 DECAPx6_ASAP7_75t_R FILLER_271_777 ();
 DECAPx2_ASAP7_75t_R FILLER_271_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_797 ();
 DECAPx1_ASAP7_75t_R FILLER_271_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_814 ();
 DECAPx2_ASAP7_75t_R FILLER_271_827 ();
 FILLER_ASAP7_75t_R FILLER_271_833 ();
 DECAPx4_ASAP7_75t_R FILLER_271_841 ();
 FILLER_ASAP7_75t_R FILLER_271_871 ();
 FILLER_ASAP7_75t_R FILLER_271_879 ();
 DECAPx4_ASAP7_75t_R FILLER_271_887 ();
 FILLER_ASAP7_75t_R FILLER_271_897 ();
 DECAPx1_ASAP7_75t_R FILLER_271_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_923 ();
 DECAPx1_ASAP7_75t_R FILLER_271_940 ();
 DECAPx10_ASAP7_75t_R FILLER_271_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_984 ();
 DECAPx4_ASAP7_75t_R FILLER_271_1003 ();
 FILLER_ASAP7_75t_R FILLER_271_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_271_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_271_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1101 ();
 FILLER_ASAP7_75t_R FILLER_271_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1185 ();
 FILLER_ASAP7_75t_R FILLER_271_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_271_1397 ();
 FILLER_ASAP7_75t_R FILLER_271_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_272_2 ();
 DECAPx10_ASAP7_75t_R FILLER_272_24 ();
 DECAPx10_ASAP7_75t_R FILLER_272_46 ();
 DECAPx10_ASAP7_75t_R FILLER_272_68 ();
 DECAPx10_ASAP7_75t_R FILLER_272_90 ();
 DECAPx10_ASAP7_75t_R FILLER_272_112 ();
 DECAPx10_ASAP7_75t_R FILLER_272_134 ();
 DECAPx10_ASAP7_75t_R FILLER_272_156 ();
 DECAPx10_ASAP7_75t_R FILLER_272_178 ();
 DECAPx10_ASAP7_75t_R FILLER_272_200 ();
 DECAPx10_ASAP7_75t_R FILLER_272_222 ();
 DECAPx10_ASAP7_75t_R FILLER_272_244 ();
 DECAPx10_ASAP7_75t_R FILLER_272_266 ();
 DECAPx10_ASAP7_75t_R FILLER_272_288 ();
 DECAPx10_ASAP7_75t_R FILLER_272_310 ();
 DECAPx10_ASAP7_75t_R FILLER_272_332 ();
 DECAPx10_ASAP7_75t_R FILLER_272_354 ();
 DECAPx10_ASAP7_75t_R FILLER_272_376 ();
 DECAPx2_ASAP7_75t_R FILLER_272_408 ();
 DECAPx6_ASAP7_75t_R FILLER_272_420 ();
 DECAPx2_ASAP7_75t_R FILLER_272_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_440 ();
 DECAPx4_ASAP7_75t_R FILLER_272_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_481 ();
 DECAPx4_ASAP7_75t_R FILLER_272_490 ();
 DECAPx1_ASAP7_75t_R FILLER_272_518 ();
 DECAPx6_ASAP7_75t_R FILLER_272_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_561 ();
 DECAPx1_ASAP7_75t_R FILLER_272_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_572 ();
 DECAPx2_ASAP7_75t_R FILLER_272_610 ();
 FILLER_ASAP7_75t_R FILLER_272_616 ();
 DECAPx1_ASAP7_75t_R FILLER_272_621 ();
 DECAPx4_ASAP7_75t_R FILLER_272_631 ();
 FILLER_ASAP7_75t_R FILLER_272_641 ();
 DECAPx2_ASAP7_75t_R FILLER_272_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_658 ();
 DECAPx2_ASAP7_75t_R FILLER_272_665 ();
 FILLER_ASAP7_75t_R FILLER_272_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_721 ();
 DECAPx10_ASAP7_75t_R FILLER_272_743 ();
 DECAPx6_ASAP7_75t_R FILLER_272_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_779 ();
 DECAPx4_ASAP7_75t_R FILLER_272_786 ();
 DECAPx1_ASAP7_75t_R FILLER_272_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_816 ();
 DECAPx1_ASAP7_75t_R FILLER_272_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_837 ();
 DECAPx4_ASAP7_75t_R FILLER_272_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_868 ();
 DECAPx10_ASAP7_75t_R FILLER_272_875 ();
 DECAPx6_ASAP7_75t_R FILLER_272_897 ();
 FILLER_ASAP7_75t_R FILLER_272_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_913 ();
 FILLER_ASAP7_75t_R FILLER_272_920 ();
 DECAPx2_ASAP7_75t_R FILLER_272_970 ();
 FILLER_ASAP7_75t_R FILLER_272_976 ();
 DECAPx4_ASAP7_75t_R FILLER_272_984 ();
 DECAPx6_ASAP7_75t_R FILLER_272_1002 ();
 FILLER_ASAP7_75t_R FILLER_272_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_272_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1052 ();
 FILLER_ASAP7_75t_R FILLER_272_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_272_1107 ();
 FILLER_ASAP7_75t_R FILLER_272_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_272_1119 ();
 FILLER_ASAP7_75t_R FILLER_272_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_272_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1174 ();
 DECAPx4_ASAP7_75t_R FILLER_272_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1342 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1364 ();
 DECAPx6_ASAP7_75t_R FILLER_272_1388 ();
 FILLER_ASAP7_75t_R FILLER_272_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_273_2 ();
 DECAPx10_ASAP7_75t_R FILLER_273_24 ();
 DECAPx10_ASAP7_75t_R FILLER_273_46 ();
 DECAPx10_ASAP7_75t_R FILLER_273_68 ();
 DECAPx10_ASAP7_75t_R FILLER_273_90 ();
 DECAPx10_ASAP7_75t_R FILLER_273_112 ();
 DECAPx10_ASAP7_75t_R FILLER_273_134 ();
 DECAPx10_ASAP7_75t_R FILLER_273_156 ();
 DECAPx10_ASAP7_75t_R FILLER_273_178 ();
 DECAPx10_ASAP7_75t_R FILLER_273_200 ();
 DECAPx10_ASAP7_75t_R FILLER_273_222 ();
 DECAPx10_ASAP7_75t_R FILLER_273_244 ();
 DECAPx10_ASAP7_75t_R FILLER_273_266 ();
 DECAPx10_ASAP7_75t_R FILLER_273_288 ();
 DECAPx10_ASAP7_75t_R FILLER_273_310 ();
 DECAPx10_ASAP7_75t_R FILLER_273_332 ();
 DECAPx10_ASAP7_75t_R FILLER_273_354 ();
 DECAPx10_ASAP7_75t_R FILLER_273_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_398 ();
 DECAPx2_ASAP7_75t_R FILLER_273_407 ();
 DECAPx2_ASAP7_75t_R FILLER_273_428 ();
 DECAPx4_ASAP7_75t_R FILLER_273_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_458 ();
 DECAPx1_ASAP7_75t_R FILLER_273_465 ();
 DECAPx2_ASAP7_75t_R FILLER_273_475 ();
 FILLER_ASAP7_75t_R FILLER_273_481 ();
 DECAPx4_ASAP7_75t_R FILLER_273_491 ();
 FILLER_ASAP7_75t_R FILLER_273_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_513 ();
 FILLER_ASAP7_75t_R FILLER_273_557 ();
 DECAPx4_ASAP7_75t_R FILLER_273_565 ();
 FILLER_ASAP7_75t_R FILLER_273_575 ();
 DECAPx4_ASAP7_75t_R FILLER_273_604 ();
 DECAPx4_ASAP7_75t_R FILLER_273_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_640 ();
 FILLER_ASAP7_75t_R FILLER_273_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_655 ();
 DECAPx2_ASAP7_75t_R FILLER_273_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_681 ();
 DECAPx1_ASAP7_75t_R FILLER_273_685 ();
 DECAPx6_ASAP7_75t_R FILLER_273_695 ();
 FILLER_ASAP7_75t_R FILLER_273_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_728 ();
 DECAPx4_ASAP7_75t_R FILLER_273_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_760 ();
 DECAPx1_ASAP7_75t_R FILLER_273_794 ();
 DECAPx2_ASAP7_75t_R FILLER_273_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_818 ();
 DECAPx2_ASAP7_75t_R FILLER_273_855 ();
 FILLER_ASAP7_75t_R FILLER_273_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_866 ();
 FILLER_ASAP7_75t_R FILLER_273_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_881 ();
 DECAPx4_ASAP7_75t_R FILLER_273_900 ();
 FILLER_ASAP7_75t_R FILLER_273_910 ();
 DECAPx1_ASAP7_75t_R FILLER_273_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_977 ();
 DECAPx2_ASAP7_75t_R FILLER_273_998 ();
 FILLER_ASAP7_75t_R FILLER_273_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_273_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_273_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1365 ();
 DECAPx6_ASAP7_75t_R FILLER_273_1387 ();
 DECAPx1_ASAP7_75t_R FILLER_273_1401 ();
 DECAPx10_ASAP7_75t_R FILLER_274_2 ();
 DECAPx10_ASAP7_75t_R FILLER_274_24 ();
 DECAPx10_ASAP7_75t_R FILLER_274_46 ();
 DECAPx10_ASAP7_75t_R FILLER_274_68 ();
 DECAPx10_ASAP7_75t_R FILLER_274_90 ();
 DECAPx10_ASAP7_75t_R FILLER_274_112 ();
 DECAPx10_ASAP7_75t_R FILLER_274_134 ();
 DECAPx10_ASAP7_75t_R FILLER_274_156 ();
 DECAPx10_ASAP7_75t_R FILLER_274_178 ();
 DECAPx10_ASAP7_75t_R FILLER_274_200 ();
 DECAPx10_ASAP7_75t_R FILLER_274_222 ();
 DECAPx10_ASAP7_75t_R FILLER_274_244 ();
 DECAPx10_ASAP7_75t_R FILLER_274_266 ();
 DECAPx10_ASAP7_75t_R FILLER_274_288 ();
 DECAPx10_ASAP7_75t_R FILLER_274_310 ();
 DECAPx10_ASAP7_75t_R FILLER_274_332 ();
 DECAPx10_ASAP7_75t_R FILLER_274_354 ();
 DECAPx6_ASAP7_75t_R FILLER_274_376 ();
 DECAPx2_ASAP7_75t_R FILLER_274_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_396 ();
 FILLER_ASAP7_75t_R FILLER_274_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_487 ();
 DECAPx10_ASAP7_75t_R FILLER_274_504 ();
 FILLER_ASAP7_75t_R FILLER_274_553 ();
 FILLER_ASAP7_75t_R FILLER_274_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_584 ();
 FILLER_ASAP7_75t_R FILLER_274_591 ();
 FILLER_ASAP7_75t_R FILLER_274_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_600 ();
 DECAPx4_ASAP7_75t_R FILLER_274_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_614 ();
 FILLER_ASAP7_75t_R FILLER_274_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_638 ();
 DECAPx1_ASAP7_75t_R FILLER_274_649 ();
 FILLER_ASAP7_75t_R FILLER_274_674 ();
 DECAPx4_ASAP7_75t_R FILLER_274_682 ();
 FILLER_ASAP7_75t_R FILLER_274_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_694 ();
 FILLER_ASAP7_75t_R FILLER_274_707 ();
 DECAPx4_ASAP7_75t_R FILLER_274_731 ();
 FILLER_ASAP7_75t_R FILLER_274_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_743 ();
 DECAPx2_ASAP7_75t_R FILLER_274_773 ();
 FILLER_ASAP7_75t_R FILLER_274_779 ();
 DECAPx1_ASAP7_75t_R FILLER_274_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_791 ();
 DECAPx4_ASAP7_75t_R FILLER_274_798 ();
 FILLER_ASAP7_75t_R FILLER_274_808 ();
 DECAPx4_ASAP7_75t_R FILLER_274_817 ();
 FILLER_ASAP7_75t_R FILLER_274_827 ();
 DECAPx1_ASAP7_75t_R FILLER_274_844 ();
 FILLER_ASAP7_75t_R FILLER_274_870 ();
 DECAPx6_ASAP7_75t_R FILLER_274_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_976 ();
 DECAPx2_ASAP7_75t_R FILLER_274_983 ();
 FILLER_ASAP7_75t_R FILLER_274_1001 ();
 FILLER_ASAP7_75t_R FILLER_274_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_274_1041 ();
 FILLER_ASAP7_75t_R FILLER_274_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_274_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_274_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_1385 ();
 DECAPx6_ASAP7_75t_R FILLER_274_1388 ();
 FILLER_ASAP7_75t_R FILLER_274_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_275_2 ();
 DECAPx10_ASAP7_75t_R FILLER_275_24 ();
 DECAPx10_ASAP7_75t_R FILLER_275_46 ();
 DECAPx10_ASAP7_75t_R FILLER_275_68 ();
 DECAPx10_ASAP7_75t_R FILLER_275_90 ();
 DECAPx10_ASAP7_75t_R FILLER_275_112 ();
 DECAPx10_ASAP7_75t_R FILLER_275_134 ();
 DECAPx10_ASAP7_75t_R FILLER_275_156 ();
 DECAPx10_ASAP7_75t_R FILLER_275_178 ();
 DECAPx10_ASAP7_75t_R FILLER_275_200 ();
 DECAPx10_ASAP7_75t_R FILLER_275_222 ();
 DECAPx10_ASAP7_75t_R FILLER_275_244 ();
 DECAPx10_ASAP7_75t_R FILLER_275_266 ();
 DECAPx10_ASAP7_75t_R FILLER_275_288 ();
 DECAPx10_ASAP7_75t_R FILLER_275_310 ();
 DECAPx10_ASAP7_75t_R FILLER_275_332 ();
 DECAPx10_ASAP7_75t_R FILLER_275_354 ();
 DECAPx10_ASAP7_75t_R FILLER_275_376 ();
 DECAPx6_ASAP7_75t_R FILLER_275_398 ();
 DECAPx1_ASAP7_75t_R FILLER_275_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_416 ();
 DECAPx2_ASAP7_75t_R FILLER_275_423 ();
 FILLER_ASAP7_75t_R FILLER_275_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_431 ();
 DECAPx1_ASAP7_75t_R FILLER_275_438 ();
 FILLER_ASAP7_75t_R FILLER_275_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_465 ();
 FILLER_ASAP7_75t_R FILLER_275_476 ();
 FILLER_ASAP7_75t_R FILLER_275_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_511 ();
 DECAPx1_ASAP7_75t_R FILLER_275_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_532 ();
 DECAPx6_ASAP7_75t_R FILLER_275_536 ();
 DECAPx1_ASAP7_75t_R FILLER_275_550 ();
 DECAPx4_ASAP7_75t_R FILLER_275_567 ();
 FILLER_ASAP7_75t_R FILLER_275_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_673 ();
 FILLER_ASAP7_75t_R FILLER_275_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_686 ();
 DECAPx6_ASAP7_75t_R FILLER_275_694 ();
 DECAPx2_ASAP7_75t_R FILLER_275_708 ();
 DECAPx10_ASAP7_75t_R FILLER_275_720 ();
 DECAPx6_ASAP7_75t_R FILLER_275_742 ();
 DECAPx1_ASAP7_75t_R FILLER_275_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_760 ();
 DECAPx6_ASAP7_75t_R FILLER_275_770 ();
 DECAPx2_ASAP7_75t_R FILLER_275_791 ();
 DECAPx10_ASAP7_75t_R FILLER_275_822 ();
 DECAPx10_ASAP7_75t_R FILLER_275_844 ();
 DECAPx2_ASAP7_75t_R FILLER_275_866 ();
 FILLER_ASAP7_75t_R FILLER_275_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_874 ();
 DECAPx2_ASAP7_75t_R FILLER_275_881 ();
 FILLER_ASAP7_75t_R FILLER_275_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_889 ();
 DECAPx2_ASAP7_75t_R FILLER_275_902 ();
 DECAPx1_ASAP7_75t_R FILLER_275_920 ();
 DECAPx1_ASAP7_75t_R FILLER_275_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_930 ();
 DECAPx6_ASAP7_75t_R FILLER_275_956 ();
 DECAPx2_ASAP7_75t_R FILLER_275_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_976 ();
 DECAPx4_ASAP7_75t_R FILLER_275_1010 ();
 FILLER_ASAP7_75t_R FILLER_275_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_275_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_275_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_275_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1377 ();
 DECAPx2_ASAP7_75t_R FILLER_275_1399 ();
 DECAPx10_ASAP7_75t_R FILLER_276_2 ();
 DECAPx10_ASAP7_75t_R FILLER_276_24 ();
 DECAPx10_ASAP7_75t_R FILLER_276_46 ();
 DECAPx10_ASAP7_75t_R FILLER_276_68 ();
 DECAPx10_ASAP7_75t_R FILLER_276_90 ();
 DECAPx10_ASAP7_75t_R FILLER_276_112 ();
 DECAPx10_ASAP7_75t_R FILLER_276_134 ();
 DECAPx10_ASAP7_75t_R FILLER_276_156 ();
 DECAPx10_ASAP7_75t_R FILLER_276_178 ();
 DECAPx10_ASAP7_75t_R FILLER_276_200 ();
 DECAPx10_ASAP7_75t_R FILLER_276_222 ();
 DECAPx10_ASAP7_75t_R FILLER_276_244 ();
 DECAPx10_ASAP7_75t_R FILLER_276_266 ();
 DECAPx10_ASAP7_75t_R FILLER_276_288 ();
 DECAPx10_ASAP7_75t_R FILLER_276_310 ();
 DECAPx10_ASAP7_75t_R FILLER_276_332 ();
 DECAPx10_ASAP7_75t_R FILLER_276_354 ();
 DECAPx10_ASAP7_75t_R FILLER_276_376 ();
 DECAPx10_ASAP7_75t_R FILLER_276_398 ();
 DECAPx4_ASAP7_75t_R FILLER_276_420 ();
 DECAPx10_ASAP7_75t_R FILLER_276_440 ();
 DECAPx10_ASAP7_75t_R FILLER_276_464 ();
 DECAPx2_ASAP7_75t_R FILLER_276_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_530 ();
 DECAPx4_ASAP7_75t_R FILLER_276_543 ();
 FILLER_ASAP7_75t_R FILLER_276_553 ();
 DECAPx4_ASAP7_75t_R FILLER_276_567 ();
 FILLER_ASAP7_75t_R FILLER_276_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_601 ();
 DECAPx1_ASAP7_75t_R FILLER_276_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_712 ();
 DECAPx10_ASAP7_75t_R FILLER_276_739 ();
 DECAPx4_ASAP7_75t_R FILLER_276_761 ();
 DECAPx4_ASAP7_75t_R FILLER_276_796 ();
 FILLER_ASAP7_75t_R FILLER_276_806 ();
 DECAPx4_ASAP7_75t_R FILLER_276_820 ();
 FILLER_ASAP7_75t_R FILLER_276_830 ();
 DECAPx10_ASAP7_75t_R FILLER_276_851 ();
 DECAPx10_ASAP7_75t_R FILLER_276_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_895 ();
 DECAPx10_ASAP7_75t_R FILLER_276_902 ();
 DECAPx1_ASAP7_75t_R FILLER_276_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_928 ();
 DECAPx10_ASAP7_75t_R FILLER_276_940 ();
 DECAPx2_ASAP7_75t_R FILLER_276_962 ();
 DECAPx10_ASAP7_75t_R FILLER_276_982 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_276_1048 ();
 FILLER_ASAP7_75t_R FILLER_276_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_276_1071 ();
 FILLER_ASAP7_75t_R FILLER_276_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_276_1382 ();
 DECAPx6_ASAP7_75t_R FILLER_276_1388 ();
 FILLER_ASAP7_75t_R FILLER_276_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_277_2 ();
 DECAPx10_ASAP7_75t_R FILLER_277_24 ();
 DECAPx10_ASAP7_75t_R FILLER_277_46 ();
 DECAPx10_ASAP7_75t_R FILLER_277_68 ();
 DECAPx10_ASAP7_75t_R FILLER_277_90 ();
 DECAPx10_ASAP7_75t_R FILLER_277_112 ();
 DECAPx10_ASAP7_75t_R FILLER_277_134 ();
 DECAPx10_ASAP7_75t_R FILLER_277_156 ();
 DECAPx10_ASAP7_75t_R FILLER_277_178 ();
 DECAPx10_ASAP7_75t_R FILLER_277_200 ();
 DECAPx10_ASAP7_75t_R FILLER_277_222 ();
 DECAPx10_ASAP7_75t_R FILLER_277_244 ();
 DECAPx10_ASAP7_75t_R FILLER_277_266 ();
 DECAPx10_ASAP7_75t_R FILLER_277_288 ();
 DECAPx10_ASAP7_75t_R FILLER_277_310 ();
 DECAPx10_ASAP7_75t_R FILLER_277_332 ();
 DECAPx10_ASAP7_75t_R FILLER_277_354 ();
 DECAPx10_ASAP7_75t_R FILLER_277_376 ();
 DECAPx10_ASAP7_75t_R FILLER_277_398 ();
 DECAPx4_ASAP7_75t_R FILLER_277_420 ();
 FILLER_ASAP7_75t_R FILLER_277_430 ();
 DECAPx2_ASAP7_75t_R FILLER_277_442 ();
 FILLER_ASAP7_75t_R FILLER_277_448 ();
 DECAPx2_ASAP7_75t_R FILLER_277_464 ();
 DECAPx10_ASAP7_75t_R FILLER_277_478 ();
 DECAPx6_ASAP7_75t_R FILLER_277_500 ();
 FILLER_ASAP7_75t_R FILLER_277_514 ();
 DECAPx2_ASAP7_75t_R FILLER_277_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_528 ();
 DECAPx1_ASAP7_75t_R FILLER_277_539 ();
 FILLER_ASAP7_75t_R FILLER_277_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_568 ();
 FILLER_ASAP7_75t_R FILLER_277_581 ();
 DECAPx1_ASAP7_75t_R FILLER_277_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_621 ();
 DECAPx1_ASAP7_75t_R FILLER_277_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_664 ();
 FILLER_ASAP7_75t_R FILLER_277_675 ();
 DECAPx4_ASAP7_75t_R FILLER_277_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_693 ();
 DECAPx4_ASAP7_75t_R FILLER_277_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_716 ();
 DECAPx6_ASAP7_75t_R FILLER_277_727 ();
 FILLER_ASAP7_75t_R FILLER_277_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_743 ();
 FILLER_ASAP7_75t_R FILLER_277_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_793 ();
 DECAPx2_ASAP7_75t_R FILLER_277_809 ();
 FILLER_ASAP7_75t_R FILLER_277_815 ();
 DECAPx2_ASAP7_75t_R FILLER_277_824 ();
 DECAPx2_ASAP7_75t_R FILLER_277_855 ();
 FILLER_ASAP7_75t_R FILLER_277_861 ();
 FILLER_ASAP7_75t_R FILLER_277_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_878 ();
 FILLER_ASAP7_75t_R FILLER_277_891 ();
 FILLER_ASAP7_75t_R FILLER_277_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_901 ();
 DECAPx2_ASAP7_75t_R FILLER_277_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_991 ();
 DECAPx2_ASAP7_75t_R FILLER_277_1005 ();
 FILLER_ASAP7_75t_R FILLER_277_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_1013 ();
 FILLER_ASAP7_75t_R FILLER_277_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_1029 ();
 FILLER_ASAP7_75t_R FILLER_277_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1357 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1379 ();
 DECAPx1_ASAP7_75t_R FILLER_277_1401 ();
 DECAPx10_ASAP7_75t_R FILLER_278_2 ();
 DECAPx10_ASAP7_75t_R FILLER_278_24 ();
 DECAPx10_ASAP7_75t_R FILLER_278_46 ();
 DECAPx10_ASAP7_75t_R FILLER_278_68 ();
 DECAPx10_ASAP7_75t_R FILLER_278_90 ();
 DECAPx10_ASAP7_75t_R FILLER_278_112 ();
 DECAPx10_ASAP7_75t_R FILLER_278_134 ();
 DECAPx10_ASAP7_75t_R FILLER_278_156 ();
 DECAPx10_ASAP7_75t_R FILLER_278_178 ();
 DECAPx10_ASAP7_75t_R FILLER_278_200 ();
 DECAPx10_ASAP7_75t_R FILLER_278_222 ();
 DECAPx10_ASAP7_75t_R FILLER_278_244 ();
 DECAPx10_ASAP7_75t_R FILLER_278_266 ();
 DECAPx10_ASAP7_75t_R FILLER_278_288 ();
 DECAPx10_ASAP7_75t_R FILLER_278_310 ();
 DECAPx10_ASAP7_75t_R FILLER_278_332 ();
 DECAPx10_ASAP7_75t_R FILLER_278_354 ();
 DECAPx10_ASAP7_75t_R FILLER_278_376 ();
 DECAPx6_ASAP7_75t_R FILLER_278_398 ();
 DECAPx2_ASAP7_75t_R FILLER_278_412 ();
 DECAPx1_ASAP7_75t_R FILLER_278_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_430 ();
 DECAPx1_ASAP7_75t_R FILLER_278_441 ();
 DECAPx1_ASAP7_75t_R FILLER_278_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_483 ();
 DECAPx4_ASAP7_75t_R FILLER_278_497 ();
 FILLER_ASAP7_75t_R FILLER_278_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_522 ();
 FILLER_ASAP7_75t_R FILLER_278_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_598 ();
 FILLER_ASAP7_75t_R FILLER_278_612 ();
 FILLER_ASAP7_75t_R FILLER_278_632 ();
 FILLER_ASAP7_75t_R FILLER_278_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_683 ();
 DECAPx2_ASAP7_75t_R FILLER_278_714 ();
 FILLER_ASAP7_75t_R FILLER_278_741 ();
 FILLER_ASAP7_75t_R FILLER_278_801 ();
 FILLER_ASAP7_75t_R FILLER_278_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_835 ();
 DECAPx2_ASAP7_75t_R FILLER_278_846 ();
 FILLER_ASAP7_75t_R FILLER_278_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_876 ();
 FILLER_ASAP7_75t_R FILLER_278_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_892 ();
 FILLER_ASAP7_75t_R FILLER_278_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_969 ();
 FILLER_ASAP7_75t_R FILLER_278_977 ();
 DECAPx1_ASAP7_75t_R FILLER_278_987 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1340 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1362 ();
 FILLER_ASAP7_75t_R FILLER_278_1384 ();
 DECAPx6_ASAP7_75t_R FILLER_278_1388 ();
 FILLER_ASAP7_75t_R FILLER_278_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_1404 ();
 DECAPx10_ASAP7_75t_R FILLER_279_2 ();
 DECAPx10_ASAP7_75t_R FILLER_279_24 ();
 DECAPx10_ASAP7_75t_R FILLER_279_46 ();
 DECAPx10_ASAP7_75t_R FILLER_279_68 ();
 DECAPx10_ASAP7_75t_R FILLER_279_90 ();
 DECAPx10_ASAP7_75t_R FILLER_279_112 ();
 DECAPx10_ASAP7_75t_R FILLER_279_134 ();
 DECAPx10_ASAP7_75t_R FILLER_279_156 ();
 DECAPx10_ASAP7_75t_R FILLER_279_178 ();
 DECAPx10_ASAP7_75t_R FILLER_279_200 ();
 DECAPx10_ASAP7_75t_R FILLER_279_222 ();
 DECAPx10_ASAP7_75t_R FILLER_279_244 ();
 DECAPx10_ASAP7_75t_R FILLER_279_266 ();
 DECAPx10_ASAP7_75t_R FILLER_279_288 ();
 DECAPx10_ASAP7_75t_R FILLER_279_310 ();
 DECAPx10_ASAP7_75t_R FILLER_279_332 ();
 DECAPx10_ASAP7_75t_R FILLER_279_354 ();
 DECAPx10_ASAP7_75t_R FILLER_279_376 ();
 DECAPx10_ASAP7_75t_R FILLER_279_398 ();
 DECAPx6_ASAP7_75t_R FILLER_279_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_434 ();
 FILLER_ASAP7_75t_R FILLER_279_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_686 ();
 DECAPx10_ASAP7_75t_R FILLER_279_729 ();
 FILLER_ASAP7_75t_R FILLER_279_751 ();
 DECAPx1_ASAP7_75t_R FILLER_279_758 ();
 DECAPx1_ASAP7_75t_R FILLER_279_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_850 ();
 FILLER_ASAP7_75t_R FILLER_279_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_895 ();
 DECAPx1_ASAP7_75t_R FILLER_279_903 ();
 DECAPx1_ASAP7_75t_R FILLER_279_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_990 ();
 DECAPx1_ASAP7_75t_R FILLER_279_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_279_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1349 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1371 ();
 DECAPx4_ASAP7_75t_R FILLER_279_1393 ();
 FILLER_ASAP7_75t_R FILLER_279_1403 ();
 DECAPx10_ASAP7_75t_R FILLER_280_2 ();
 DECAPx10_ASAP7_75t_R FILLER_280_24 ();
 DECAPx10_ASAP7_75t_R FILLER_280_46 ();
 DECAPx10_ASAP7_75t_R FILLER_280_68 ();
 DECAPx10_ASAP7_75t_R FILLER_280_90 ();
 DECAPx10_ASAP7_75t_R FILLER_280_112 ();
 DECAPx10_ASAP7_75t_R FILLER_280_134 ();
 DECAPx10_ASAP7_75t_R FILLER_280_156 ();
 DECAPx10_ASAP7_75t_R FILLER_280_178 ();
 DECAPx10_ASAP7_75t_R FILLER_280_200 ();
 DECAPx10_ASAP7_75t_R FILLER_280_222 ();
 DECAPx10_ASAP7_75t_R FILLER_280_244 ();
 DECAPx10_ASAP7_75t_R FILLER_280_266 ();
 DECAPx10_ASAP7_75t_R FILLER_280_288 ();
 DECAPx10_ASAP7_75t_R FILLER_280_310 ();
 DECAPx10_ASAP7_75t_R FILLER_280_332 ();
 DECAPx10_ASAP7_75t_R FILLER_280_354 ();
 DECAPx10_ASAP7_75t_R FILLER_280_376 ();
 DECAPx10_ASAP7_75t_R FILLER_280_398 ();
 DECAPx10_ASAP7_75t_R FILLER_280_420 ();
 DECAPx6_ASAP7_75t_R FILLER_280_442 ();
 DECAPx2_ASAP7_75t_R FILLER_280_456 ();
 DECAPx10_ASAP7_75t_R FILLER_280_464 ();
 FILLER_ASAP7_75t_R FILLER_280_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_538 ();
 FILLER_ASAP7_75t_R FILLER_280_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_587 ();
 FILLER_ASAP7_75t_R FILLER_280_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_679 ();
 FILLER_ASAP7_75t_R FILLER_280_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_694 ();
 FILLER_ASAP7_75t_R FILLER_280_701 ();
 DECAPx2_ASAP7_75t_R FILLER_280_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_886 ();
 FILLER_ASAP7_75t_R FILLER_280_897 ();
 DECAPx1_ASAP7_75t_R FILLER_280_920 ();
 FILLER_ASAP7_75t_R FILLER_280_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_928 ();
 DECAPx1_ASAP7_75t_R FILLER_280_967 ();
 DECAPx10_ASAP7_75t_R FILLER_280_997 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1019 ();
 FILLER_ASAP7_75t_R FILLER_280_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1354 ();
 DECAPx4_ASAP7_75t_R FILLER_280_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_280_1388 ();
 FILLER_ASAP7_75t_R FILLER_280_1402 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_1404 ();
endmodule
