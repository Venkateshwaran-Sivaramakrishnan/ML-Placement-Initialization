module miter (
  input  [  0:0] \__pi_clk ,
  input  [127:0] \__pi_key ,
  input  [  0:0] \__pi_ld ,
  input  [  0:0] \__pi_rst ,
  input  [127:0] \__pi_text_in ,
`ifdef DIRECT_CROSS_POINTS
`else
`endif
  output [  0:0] \__mp_clkbuf_0_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_0_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.Y__gold ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.A__gold ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.Y__gold ,
  output [  0:0] \__mp_clkload0.A__gold ,
  output [  0:0] \__mp_clkload0.Y__gold ,
  output [  0:0] \__mp_clkload1.A__gold ,
  output [  0:0] \__mp_clkload10.A__gold ,
  output [  0:0] \__mp_clkload11.A__gold ,
  output [  0:0] \__mp_clkload12.A__gold ,
  output [  0:0] \__mp_clkload13.A__gold ,
  output [  0:0] \__mp_clkload14.A__gold ,
  output [  0:0] \__mp_clkload15.A__gold ,
  output [  0:0] \__mp_clkload16.A__gold ,
  output [  0:0] \__mp_clkload17.A__gold ,
  output [  0:0] \__mp_clkload18.A__gold ,
  output [  0:0] \__mp_clkload18.Y__gold ,
  output [  0:0] \__mp_clkload19.A__gold ,
  output [  0:0] \__mp_clkload2.A__gold ,
  output [  0:0] \__mp_clkload20.A__gold ,
  output [  0:0] \__mp_clkload21.A__gold ,
  output [  0:0] \__mp_clkload22.A__gold ,
  output [  0:0] \__mp_clkload23.A__gold ,
  output [  0:0] \__mp_clkload24.A__gold ,
  output [  0:0] \__mp_clkload25.A__gold ,
  output [  0:0] \__mp_clkload26.A__gold ,
  output [  0:0] \__mp_clkload27.A__gold ,
  output [  0:0] \__mp_clkload28.A__gold ,
  output [  0:0] \__mp_clkload29.A__gold ,
  output [  0:0] \__mp_clkload3.A__gold ,
  output [  0:0] \__mp_clkload30.A__gold ,
  output [  0:0] \__mp_clkload31.A__gold ,
  output [  0:0] \__mp_clkload31.Y__gold ,
  output [  0:0] \__mp_clkload32.A__gold ,
  output [  0:0] \__mp_clkload4.A__gold ,
  output [  0:0] \__mp_clkload5.A__gold ,
  output [  0:0] \__mp_clkload6.A__gold ,
  output [  0:0] \__mp_clkload7.A__gold ,
  output [  0:0] \__mp_clkload8.A__gold ,
  output [  0:0] \__mp_clkload9.A__gold ,
  output [  0:0] \__mp_clknet_0_clk__gold ,
  output [  0:0] \__mp_clknet_2_0_0_clk__gold ,
  output [  0:0] \__mp_clknet_2_1_0_clk__gold ,
  output [  0:0] \__mp_clknet_2_2_0_clk__gold ,
  output [  0:0] \__mp_clknet_2_3_0_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_0_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_10_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_11_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_12_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_13_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_14_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_15_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_16_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_17_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_18_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_19_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_1_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_20_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_21_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_22_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_23_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_24_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_25_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_26_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_27_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_28_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_29_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_2_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_30_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_31_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_32_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_33_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_3_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_4_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_5_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_6_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_7_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_8_clk__gold ,
  output [  0:0] \__mp_clknet_leaf_9_clk__gold ,
  output [  0:0] \__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gold ,
  output [  0:0] \__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gold ,
  output [  0:0] \__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gold ,
  output [  0:0] \__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gold ,
  output [  0:0] \__mp_done$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_done$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_done$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_input1.A__gold ,
  output [  0:0] \__mp_input1.Y__gold ,
  output [  0:0] \__mp_input10.A__gold ,
  output [  0:0] \__mp_input10.Y__gold ,
  output [  0:0] \__mp_input100.A__gold ,
  output [  0:0] \__mp_input100.Y__gold ,
  output [  0:0] \__mp_input101.A__gold ,
  output [  0:0] \__mp_input101.Y__gold ,
  output [  0:0] \__mp_input102.A__gold ,
  output [  0:0] \__mp_input102.Y__gold ,
  output [  0:0] \__mp_input103.A__gold ,
  output [  0:0] \__mp_input103.Y__gold ,
  output [  0:0] \__mp_input104.A__gold ,
  output [  0:0] \__mp_input104.Y__gold ,
  output [  0:0] \__mp_input105.A__gold ,
  output [  0:0] \__mp_input105.Y__gold ,
  output [  0:0] \__mp_input106.A__gold ,
  output [  0:0] \__mp_input106.Y__gold ,
  output [  0:0] \__mp_input107.A__gold ,
  output [  0:0] \__mp_input107.Y__gold ,
  output [  0:0] \__mp_input108.A__gold ,
  output [  0:0] \__mp_input108.Y__gold ,
  output [  0:0] \__mp_input109.A__gold ,
  output [  0:0] \__mp_input109.Y__gold ,
  output [  0:0] \__mp_input11.A__gold ,
  output [  0:0] \__mp_input11.Y__gold ,
  output [  0:0] \__mp_input110.A__gold ,
  output [  0:0] \__mp_input110.Y__gold ,
  output [  0:0] \__mp_input111.A__gold ,
  output [  0:0] \__mp_input111.Y__gold ,
  output [  0:0] \__mp_input112.A__gold ,
  output [  0:0] \__mp_input112.Y__gold ,
  output [  0:0] \__mp_input113.A__gold ,
  output [  0:0] \__mp_input113.Y__gold ,
  output [  0:0] \__mp_input114.A__gold ,
  output [  0:0] \__mp_input114.Y__gold ,
  output [  0:0] \__mp_input115.A__gold ,
  output [  0:0] \__mp_input115.Y__gold ,
  output [  0:0] \__mp_input116.A__gold ,
  output [  0:0] \__mp_input116.Y__gold ,
  output [  0:0] \__mp_input117.A__gold ,
  output [  0:0] \__mp_input117.Y__gold ,
  output [  0:0] \__mp_input118.A__gold ,
  output [  0:0] \__mp_input118.Y__gold ,
  output [  0:0] \__mp_input119.A__gold ,
  output [  0:0] \__mp_input119.Y__gold ,
  output [  0:0] \__mp_input12.A__gold ,
  output [  0:0] \__mp_input12.Y__gold ,
  output [  0:0] \__mp_input120.A__gold ,
  output [  0:0] \__mp_input120.Y__gold ,
  output [  0:0] \__mp_input121.A__gold ,
  output [  0:0] \__mp_input121.Y__gold ,
  output [  0:0] \__mp_input122.A__gold ,
  output [  0:0] \__mp_input122.Y__gold ,
  output [  0:0] \__mp_input123.A__gold ,
  output [  0:0] \__mp_input123.Y__gold ,
  output [  0:0] \__mp_input124.A__gold ,
  output [  0:0] \__mp_input124.Y__gold ,
  output [  0:0] \__mp_input125.A__gold ,
  output [  0:0] \__mp_input125.Y__gold ,
  output [  0:0] \__mp_input126.A__gold ,
  output [  0:0] \__mp_input126.Y__gold ,
  output [  0:0] \__mp_input127.A__gold ,
  output [  0:0] \__mp_input127.Y__gold ,
  output [  0:0] \__mp_input128.A__gold ,
  output [  0:0] \__mp_input128.Y__gold ,
  output [  0:0] \__mp_input129.A__gold ,
  output [  0:0] \__mp_input129.Y__gold ,
  output [  0:0] \__mp_input13.A__gold ,
  output [  0:0] \__mp_input13.Y__gold ,
  output [  0:0] \__mp_input130.A__gold ,
  output [  0:0] \__mp_input130.Y__gold ,
  output [  0:0] \__mp_input131.A__gold ,
  output [  0:0] \__mp_input131.Y__gold ,
  output [  0:0] \__mp_input132.A__gold ,
  output [  0:0] \__mp_input132.Y__gold ,
  output [  0:0] \__mp_input133.A__gold ,
  output [  0:0] \__mp_input133.Y__gold ,
  output [  0:0] \__mp_input134.A__gold ,
  output [  0:0] \__mp_input134.Y__gold ,
  output [  0:0] \__mp_input135.A__gold ,
  output [  0:0] \__mp_input135.Y__gold ,
  output [  0:0] \__mp_input136.A__gold ,
  output [  0:0] \__mp_input136.Y__gold ,
  output [  0:0] \__mp_input137.A__gold ,
  output [  0:0] \__mp_input137.Y__gold ,
  output [  0:0] \__mp_input138.A__gold ,
  output [  0:0] \__mp_input138.Y__gold ,
  output [  0:0] \__mp_input139.A__gold ,
  output [  0:0] \__mp_input139.Y__gold ,
  output [  0:0] \__mp_input14.A__gold ,
  output [  0:0] \__mp_input14.Y__gold ,
  output [  0:0] \__mp_input140.A__gold ,
  output [  0:0] \__mp_input140.Y__gold ,
  output [  0:0] \__mp_input141.A__gold ,
  output [  0:0] \__mp_input141.Y__gold ,
  output [  0:0] \__mp_input142.A__gold ,
  output [  0:0] \__mp_input142.Y__gold ,
  output [  0:0] \__mp_input143.A__gold ,
  output [  0:0] \__mp_input143.Y__gold ,
  output [  0:0] \__mp_input144.A__gold ,
  output [  0:0] \__mp_input144.Y__gold ,
  output [  0:0] \__mp_input145.A__gold ,
  output [  0:0] \__mp_input145.Y__gold ,
  output [  0:0] \__mp_input146.A__gold ,
  output [  0:0] \__mp_input146.Y__gold ,
  output [  0:0] \__mp_input147.A__gold ,
  output [  0:0] \__mp_input147.Y__gold ,
  output [  0:0] \__mp_input148.A__gold ,
  output [  0:0] \__mp_input148.Y__gold ,
  output [  0:0] \__mp_input149.A__gold ,
  output [  0:0] \__mp_input149.Y__gold ,
  output [  0:0] \__mp_input15.A__gold ,
  output [  0:0] \__mp_input15.Y__gold ,
  output [  0:0] \__mp_input150.A__gold ,
  output [  0:0] \__mp_input150.Y__gold ,
  output [  0:0] \__mp_input151.A__gold ,
  output [  0:0] \__mp_input151.Y__gold ,
  output [  0:0] \__mp_input152.A__gold ,
  output [  0:0] \__mp_input152.Y__gold ,
  output [  0:0] \__mp_input153.A__gold ,
  output [  0:0] \__mp_input153.Y__gold ,
  output [  0:0] \__mp_input154.A__gold ,
  output [  0:0] \__mp_input154.Y__gold ,
  output [  0:0] \__mp_input155.A__gold ,
  output [  0:0] \__mp_input155.Y__gold ,
  output [  0:0] \__mp_input156.A__gold ,
  output [  0:0] \__mp_input156.Y__gold ,
  output [  0:0] \__mp_input157.A__gold ,
  output [  0:0] \__mp_input157.Y__gold ,
  output [  0:0] \__mp_input158.A__gold ,
  output [  0:0] \__mp_input158.Y__gold ,
  output [  0:0] \__mp_input159.A__gold ,
  output [  0:0] \__mp_input159.Y__gold ,
  output [  0:0] \__mp_input16.A__gold ,
  output [  0:0] \__mp_input16.Y__gold ,
  output [  0:0] \__mp_input160.A__gold ,
  output [  0:0] \__mp_input160.Y__gold ,
  output [  0:0] \__mp_input161.A__gold ,
  output [  0:0] \__mp_input161.Y__gold ,
  output [  0:0] \__mp_input162.A__gold ,
  output [  0:0] \__mp_input162.Y__gold ,
  output [  0:0] \__mp_input163.A__gold ,
  output [  0:0] \__mp_input163.Y__gold ,
  output [  0:0] \__mp_input164.A__gold ,
  output [  0:0] \__mp_input164.Y__gold ,
  output [  0:0] \__mp_input165.A__gold ,
  output [  0:0] \__mp_input165.Y__gold ,
  output [  0:0] \__mp_input166.A__gold ,
  output [  0:0] \__mp_input166.Y__gold ,
  output [  0:0] \__mp_input167.A__gold ,
  output [  0:0] \__mp_input167.Y__gold ,
  output [  0:0] \__mp_input168.A__gold ,
  output [  0:0] \__mp_input168.Y__gold ,
  output [  0:0] \__mp_input169.A__gold ,
  output [  0:0] \__mp_input169.Y__gold ,
  output [  0:0] \__mp_input17.A__gold ,
  output [  0:0] \__mp_input17.Y__gold ,
  output [  0:0] \__mp_input170.A__gold ,
  output [  0:0] \__mp_input170.Y__gold ,
  output [  0:0] \__mp_input171.A__gold ,
  output [  0:0] \__mp_input171.Y__gold ,
  output [  0:0] \__mp_input172.A__gold ,
  output [  0:0] \__mp_input172.Y__gold ,
  output [  0:0] \__mp_input173.A__gold ,
  output [  0:0] \__mp_input173.Y__gold ,
  output [  0:0] \__mp_input174.A__gold ,
  output [  0:0] \__mp_input174.Y__gold ,
  output [  0:0] \__mp_input175.A__gold ,
  output [  0:0] \__mp_input175.Y__gold ,
  output [  0:0] \__mp_input176.A__gold ,
  output [  0:0] \__mp_input176.Y__gold ,
  output [  0:0] \__mp_input177.A__gold ,
  output [  0:0] \__mp_input177.Y__gold ,
  output [  0:0] \__mp_input178.A__gold ,
  output [  0:0] \__mp_input178.Y__gold ,
  output [  0:0] \__mp_input179.A__gold ,
  output [  0:0] \__mp_input179.Y__gold ,
  output [  0:0] \__mp_input18.A__gold ,
  output [  0:0] \__mp_input18.Y__gold ,
  output [  0:0] \__mp_input180.A__gold ,
  output [  0:0] \__mp_input180.Y__gold ,
  output [  0:0] \__mp_input181.A__gold ,
  output [  0:0] \__mp_input181.Y__gold ,
  output [  0:0] \__mp_input182.A__gold ,
  output [  0:0] \__mp_input182.Y__gold ,
  output [  0:0] \__mp_input183.A__gold ,
  output [  0:0] \__mp_input183.Y__gold ,
  output [  0:0] \__mp_input184.A__gold ,
  output [  0:0] \__mp_input184.Y__gold ,
  output [  0:0] \__mp_input185.A__gold ,
  output [  0:0] \__mp_input185.Y__gold ,
  output [  0:0] \__mp_input186.A__gold ,
  output [  0:0] \__mp_input186.Y__gold ,
  output [  0:0] \__mp_input187.A__gold ,
  output [  0:0] \__mp_input187.Y__gold ,
  output [  0:0] \__mp_input188.A__gold ,
  output [  0:0] \__mp_input188.Y__gold ,
  output [  0:0] \__mp_input189.A__gold ,
  output [  0:0] \__mp_input189.Y__gold ,
  output [  0:0] \__mp_input19.A__gold ,
  output [  0:0] \__mp_input19.Y__gold ,
  output [  0:0] \__mp_input190.A__gold ,
  output [  0:0] \__mp_input190.Y__gold ,
  output [  0:0] \__mp_input191.A__gold ,
  output [  0:0] \__mp_input191.Y__gold ,
  output [  0:0] \__mp_input192.A__gold ,
  output [  0:0] \__mp_input192.Y__gold ,
  output [  0:0] \__mp_input193.A__gold ,
  output [  0:0] \__mp_input193.Y__gold ,
  output [  0:0] \__mp_input194.A__gold ,
  output [  0:0] \__mp_input194.Y__gold ,
  output [  0:0] \__mp_input195.A__gold ,
  output [  0:0] \__mp_input195.Y__gold ,
  output [  0:0] \__mp_input196.A__gold ,
  output [  0:0] \__mp_input196.Y__gold ,
  output [  0:0] \__mp_input197.A__gold ,
  output [  0:0] \__mp_input197.Y__gold ,
  output [  0:0] \__mp_input198.A__gold ,
  output [  0:0] \__mp_input198.Y__gold ,
  output [  0:0] \__mp_input199.A__gold ,
  output [  0:0] \__mp_input199.Y__gold ,
  output [  0:0] \__mp_input2.A__gold ,
  output [  0:0] \__mp_input2.Y__gold ,
  output [  0:0] \__mp_input20.A__gold ,
  output [  0:0] \__mp_input20.Y__gold ,
  output [  0:0] \__mp_input200.A__gold ,
  output [  0:0] \__mp_input200.Y__gold ,
  output [  0:0] \__mp_input201.A__gold ,
  output [  0:0] \__mp_input201.Y__gold ,
  output [  0:0] \__mp_input202.A__gold ,
  output [  0:0] \__mp_input202.Y__gold ,
  output [  0:0] \__mp_input203.A__gold ,
  output [  0:0] \__mp_input203.Y__gold ,
  output [  0:0] \__mp_input204.A__gold ,
  output [  0:0] \__mp_input204.Y__gold ,
  output [  0:0] \__mp_input205.A__gold ,
  output [  0:0] \__mp_input205.Y__gold ,
  output [  0:0] \__mp_input206.A__gold ,
  output [  0:0] \__mp_input206.Y__gold ,
  output [  0:0] \__mp_input207.A__gold ,
  output [  0:0] \__mp_input207.Y__gold ,
  output [  0:0] \__mp_input208.A__gold ,
  output [  0:0] \__mp_input208.Y__gold ,
  output [  0:0] \__mp_input209.A__gold ,
  output [  0:0] \__mp_input209.Y__gold ,
  output [  0:0] \__mp_input21.A__gold ,
  output [  0:0] \__mp_input21.Y__gold ,
  output [  0:0] \__mp_input210.A__gold ,
  output [  0:0] \__mp_input210.Y__gold ,
  output [  0:0] \__mp_input211.A__gold ,
  output [  0:0] \__mp_input211.Y__gold ,
  output [  0:0] \__mp_input212.A__gold ,
  output [  0:0] \__mp_input212.Y__gold ,
  output [  0:0] \__mp_input213.A__gold ,
  output [  0:0] \__mp_input213.Y__gold ,
  output [  0:0] \__mp_input214.A__gold ,
  output [  0:0] \__mp_input214.Y__gold ,
  output [  0:0] \__mp_input215.A__gold ,
  output [  0:0] \__mp_input215.Y__gold ,
  output [  0:0] \__mp_input216.A__gold ,
  output [  0:0] \__mp_input216.Y__gold ,
  output [  0:0] \__mp_input217.A__gold ,
  output [  0:0] \__mp_input217.Y__gold ,
  output [  0:0] \__mp_input218.A__gold ,
  output [  0:0] \__mp_input218.Y__gold ,
  output [  0:0] \__mp_input219.A__gold ,
  output [  0:0] \__mp_input219.Y__gold ,
  output [  0:0] \__mp_input22.A__gold ,
  output [  0:0] \__mp_input22.Y__gold ,
  output [  0:0] \__mp_input220.A__gold ,
  output [  0:0] \__mp_input220.Y__gold ,
  output [  0:0] \__mp_input221.A__gold ,
  output [  0:0] \__mp_input221.Y__gold ,
  output [  0:0] \__mp_input222.A__gold ,
  output [  0:0] \__mp_input222.Y__gold ,
  output [  0:0] \__mp_input223.A__gold ,
  output [  0:0] \__mp_input223.Y__gold ,
  output [  0:0] \__mp_input224.A__gold ,
  output [  0:0] \__mp_input224.Y__gold ,
  output [  0:0] \__mp_input225.A__gold ,
  output [  0:0] \__mp_input225.Y__gold ,
  output [  0:0] \__mp_input226.A__gold ,
  output [  0:0] \__mp_input226.Y__gold ,
  output [  0:0] \__mp_input227.A__gold ,
  output [  0:0] \__mp_input227.Y__gold ,
  output [  0:0] \__mp_input228.A__gold ,
  output [  0:0] \__mp_input228.Y__gold ,
  output [  0:0] \__mp_input229.A__gold ,
  output [  0:0] \__mp_input229.Y__gold ,
  output [  0:0] \__mp_input23.A__gold ,
  output [  0:0] \__mp_input23.Y__gold ,
  output [  0:0] \__mp_input230.A__gold ,
  output [  0:0] \__mp_input230.Y__gold ,
  output [  0:0] \__mp_input231.A__gold ,
  output [  0:0] \__mp_input231.Y__gold ,
  output [  0:0] \__mp_input232.A__gold ,
  output [  0:0] \__mp_input232.Y__gold ,
  output [  0:0] \__mp_input233.A__gold ,
  output [  0:0] \__mp_input233.Y__gold ,
  output [  0:0] \__mp_input234.A__gold ,
  output [  0:0] \__mp_input234.Y__gold ,
  output [  0:0] \__mp_input235.A__gold ,
  output [  0:0] \__mp_input235.Y__gold ,
  output [  0:0] \__mp_input236.A__gold ,
  output [  0:0] \__mp_input236.Y__gold ,
  output [  0:0] \__mp_input237.A__gold ,
  output [  0:0] \__mp_input237.Y__gold ,
  output [  0:0] \__mp_input238.A__gold ,
  output [  0:0] \__mp_input238.Y__gold ,
  output [  0:0] \__mp_input239.A__gold ,
  output [  0:0] \__mp_input239.Y__gold ,
  output [  0:0] \__mp_input24.A__gold ,
  output [  0:0] \__mp_input24.Y__gold ,
  output [  0:0] \__mp_input240.A__gold ,
  output [  0:0] \__mp_input240.Y__gold ,
  output [  0:0] \__mp_input241.A__gold ,
  output [  0:0] \__mp_input241.Y__gold ,
  output [  0:0] \__mp_input242.A__gold ,
  output [  0:0] \__mp_input242.Y__gold ,
  output [  0:0] \__mp_input243.A__gold ,
  output [  0:0] \__mp_input243.Y__gold ,
  output [  0:0] \__mp_input244.A__gold ,
  output [  0:0] \__mp_input244.Y__gold ,
  output [  0:0] \__mp_input245.A__gold ,
  output [  0:0] \__mp_input245.Y__gold ,
  output [  0:0] \__mp_input246.A__gold ,
  output [  0:0] \__mp_input246.Y__gold ,
  output [  0:0] \__mp_input247.A__gold ,
  output [  0:0] \__mp_input247.Y__gold ,
  output [  0:0] \__mp_input248.A__gold ,
  output [  0:0] \__mp_input248.Y__gold ,
  output [  0:0] \__mp_input249.A__gold ,
  output [  0:0] \__mp_input249.Y__gold ,
  output [  0:0] \__mp_input25.A__gold ,
  output [  0:0] \__mp_input25.Y__gold ,
  output [  0:0] \__mp_input250.A__gold ,
  output [  0:0] \__mp_input250.Y__gold ,
  output [  0:0] \__mp_input251.A__gold ,
  output [  0:0] \__mp_input251.Y__gold ,
  output [  0:0] \__mp_input252.A__gold ,
  output [  0:0] \__mp_input252.Y__gold ,
  output [  0:0] \__mp_input253.A__gold ,
  output [  0:0] \__mp_input253.Y__gold ,
  output [  0:0] \__mp_input254.A__gold ,
  output [  0:0] \__mp_input254.Y__gold ,
  output [  0:0] \__mp_input255.A__gold ,
  output [  0:0] \__mp_input255.Y__gold ,
  output [  0:0] \__mp_input256.A__gold ,
  output [  0:0] \__mp_input256.Y__gold ,
  output [  0:0] \__mp_input257.A__gold ,
  output [  0:0] \__mp_input257.Y__gold ,
  output [  0:0] \__mp_input258.A__gold ,
  output [  0:0] \__mp_input258.Y__gold ,
  output [  0:0] \__mp_input26.A__gold ,
  output [  0:0] \__mp_input26.Y__gold ,
  output [  0:0] \__mp_input27.A__gold ,
  output [  0:0] \__mp_input27.Y__gold ,
  output [  0:0] \__mp_input28.A__gold ,
  output [  0:0] \__mp_input28.Y__gold ,
  output [  0:0] \__mp_input29.A__gold ,
  output [  0:0] \__mp_input29.Y__gold ,
  output [  0:0] \__mp_input3.A__gold ,
  output [  0:0] \__mp_input3.Y__gold ,
  output [  0:0] \__mp_input30.A__gold ,
  output [  0:0] \__mp_input30.Y__gold ,
  output [  0:0] \__mp_input31.A__gold ,
  output [  0:0] \__mp_input31.Y__gold ,
  output [  0:0] \__mp_input32.A__gold ,
  output [  0:0] \__mp_input32.Y__gold ,
  output [  0:0] \__mp_input33.A__gold ,
  output [  0:0] \__mp_input33.Y__gold ,
  output [  0:0] \__mp_input34.A__gold ,
  output [  0:0] \__mp_input34.Y__gold ,
  output [  0:0] \__mp_input35.A__gold ,
  output [  0:0] \__mp_input35.Y__gold ,
  output [  0:0] \__mp_input36.A__gold ,
  output [  0:0] \__mp_input36.Y__gold ,
  output [  0:0] \__mp_input37.A__gold ,
  output [  0:0] \__mp_input37.Y__gold ,
  output [  0:0] \__mp_input38.A__gold ,
  output [  0:0] \__mp_input38.Y__gold ,
  output [  0:0] \__mp_input39.A__gold ,
  output [  0:0] \__mp_input39.Y__gold ,
  output [  0:0] \__mp_input4.A__gold ,
  output [  0:0] \__mp_input4.Y__gold ,
  output [  0:0] \__mp_input40.A__gold ,
  output [  0:0] \__mp_input40.Y__gold ,
  output [  0:0] \__mp_input41.A__gold ,
  output [  0:0] \__mp_input41.Y__gold ,
  output [  0:0] \__mp_input42.A__gold ,
  output [  0:0] \__mp_input42.Y__gold ,
  output [  0:0] \__mp_input43.A__gold ,
  output [  0:0] \__mp_input43.Y__gold ,
  output [  0:0] \__mp_input44.A__gold ,
  output [  0:0] \__mp_input44.Y__gold ,
  output [  0:0] \__mp_input45.A__gold ,
  output [  0:0] \__mp_input45.Y__gold ,
  output [  0:0] \__mp_input46.A__gold ,
  output [  0:0] \__mp_input46.Y__gold ,
  output [  0:0] \__mp_input47.A__gold ,
  output [  0:0] \__mp_input47.Y__gold ,
  output [  0:0] \__mp_input48.A__gold ,
  output [  0:0] \__mp_input48.Y__gold ,
  output [  0:0] \__mp_input49.A__gold ,
  output [  0:0] \__mp_input49.Y__gold ,
  output [  0:0] \__mp_input5.A__gold ,
  output [  0:0] \__mp_input5.Y__gold ,
  output [  0:0] \__mp_input50.A__gold ,
  output [  0:0] \__mp_input50.Y__gold ,
  output [  0:0] \__mp_input51.A__gold ,
  output [  0:0] \__mp_input51.Y__gold ,
  output [  0:0] \__mp_input52.A__gold ,
  output [  0:0] \__mp_input52.Y__gold ,
  output [  0:0] \__mp_input53.A__gold ,
  output [  0:0] \__mp_input53.Y__gold ,
  output [  0:0] \__mp_input54.A__gold ,
  output [  0:0] \__mp_input54.Y__gold ,
  output [  0:0] \__mp_input55.A__gold ,
  output [  0:0] \__mp_input55.Y__gold ,
  output [  0:0] \__mp_input56.A__gold ,
  output [  0:0] \__mp_input56.Y__gold ,
  output [  0:0] \__mp_input57.A__gold ,
  output [  0:0] \__mp_input57.Y__gold ,
  output [  0:0] \__mp_input58.A__gold ,
  output [  0:0] \__mp_input58.Y__gold ,
  output [  0:0] \__mp_input59.A__gold ,
  output [  0:0] \__mp_input59.Y__gold ,
  output [  0:0] \__mp_input6.A__gold ,
  output [  0:0] \__mp_input6.Y__gold ,
  output [  0:0] \__mp_input60.A__gold ,
  output [  0:0] \__mp_input60.Y__gold ,
  output [  0:0] \__mp_input61.A__gold ,
  output [  0:0] \__mp_input61.Y__gold ,
  output [  0:0] \__mp_input62.A__gold ,
  output [  0:0] \__mp_input62.Y__gold ,
  output [  0:0] \__mp_input63.A__gold ,
  output [  0:0] \__mp_input63.Y__gold ,
  output [  0:0] \__mp_input64.A__gold ,
  output [  0:0] \__mp_input64.Y__gold ,
  output [  0:0] \__mp_input65.A__gold ,
  output [  0:0] \__mp_input65.Y__gold ,
  output [  0:0] \__mp_input66.A__gold ,
  output [  0:0] \__mp_input66.Y__gold ,
  output [  0:0] \__mp_input67.A__gold ,
  output [  0:0] \__mp_input67.Y__gold ,
  output [  0:0] \__mp_input68.A__gold ,
  output [  0:0] \__mp_input68.Y__gold ,
  output [  0:0] \__mp_input69.A__gold ,
  output [  0:0] \__mp_input69.Y__gold ,
  output [  0:0] \__mp_input7.A__gold ,
  output [  0:0] \__mp_input7.Y__gold ,
  output [  0:0] \__mp_input70.A__gold ,
  output [  0:0] \__mp_input70.Y__gold ,
  output [  0:0] \__mp_input71.A__gold ,
  output [  0:0] \__mp_input71.Y__gold ,
  output [  0:0] \__mp_input72.A__gold ,
  output [  0:0] \__mp_input72.Y__gold ,
  output [  0:0] \__mp_input73.A__gold ,
  output [  0:0] \__mp_input73.Y__gold ,
  output [  0:0] \__mp_input74.A__gold ,
  output [  0:0] \__mp_input74.Y__gold ,
  output [  0:0] \__mp_input75.A__gold ,
  output [  0:0] \__mp_input75.Y__gold ,
  output [  0:0] \__mp_input76.A__gold ,
  output [  0:0] \__mp_input76.Y__gold ,
  output [  0:0] \__mp_input77.A__gold ,
  output [  0:0] \__mp_input77.Y__gold ,
  output [  0:0] \__mp_input78.A__gold ,
  output [  0:0] \__mp_input78.Y__gold ,
  output [  0:0] \__mp_input79.A__gold ,
  output [  0:0] \__mp_input79.Y__gold ,
  output [  0:0] \__mp_input8.A__gold ,
  output [  0:0] \__mp_input8.Y__gold ,
  output [  0:0] \__mp_input80.A__gold ,
  output [  0:0] \__mp_input80.Y__gold ,
  output [  0:0] \__mp_input81.A__gold ,
  output [  0:0] \__mp_input81.Y__gold ,
  output [  0:0] \__mp_input82.A__gold ,
  output [  0:0] \__mp_input82.Y__gold ,
  output [  0:0] \__mp_input83.A__gold ,
  output [  0:0] \__mp_input83.Y__gold ,
  output [  0:0] \__mp_input84.A__gold ,
  output [  0:0] \__mp_input84.Y__gold ,
  output [  0:0] \__mp_input85.A__gold ,
  output [  0:0] \__mp_input85.Y__gold ,
  output [  0:0] \__mp_input86.A__gold ,
  output [  0:0] \__mp_input86.Y__gold ,
  output [  0:0] \__mp_input87.A__gold ,
  output [  0:0] \__mp_input87.Y__gold ,
  output [  0:0] \__mp_input88.A__gold ,
  output [  0:0] \__mp_input88.Y__gold ,
  output [  0:0] \__mp_input89.A__gold ,
  output [  0:0] \__mp_input89.Y__gold ,
  output [  0:0] \__mp_input9.A__gold ,
  output [  0:0] \__mp_input9.Y__gold ,
  output [  0:0] \__mp_input90.A__gold ,
  output [  0:0] \__mp_input90.Y__gold ,
  output [  0:0] \__mp_input91.A__gold ,
  output [  0:0] \__mp_input91.Y__gold ,
  output [  0:0] \__mp_input92.A__gold ,
  output [  0:0] \__mp_input92.Y__gold ,
  output [  0:0] \__mp_input93.A__gold ,
  output [  0:0] \__mp_input93.Y__gold ,
  output [  0:0] \__mp_input94.A__gold ,
  output [  0:0] \__mp_input94.Y__gold ,
  output [  0:0] \__mp_input95.A__gold ,
  output [  0:0] \__mp_input95.Y__gold ,
  output [  0:0] \__mp_input96.A__gold ,
  output [  0:0] \__mp_input96.Y__gold ,
  output [  0:0] \__mp_input97.A__gold ,
  output [  0:0] \__mp_input97.Y__gold ,
  output [  0:0] \__mp_input98.A__gold ,
  output [  0:0] \__mp_input98.Y__gold ,
  output [  0:0] \__mp_input99.A__gold ,
  output [  0:0] \__mp_input99.Y__gold ,
  output [  0:0] \__mp_ld_r$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_ld_r$_DFF_P_.D__gold ,
  output [  0:0] \__mp_output259.A__gold ,
  output [  0:0] \__mp_output259.Y__gold ,
  output [  0:0] \__mp_output260.A__gold ,
  output [  0:0] \__mp_output260.Y__gold ,
  output [  0:0] \__mp_output261.A__gold ,
  output [  0:0] \__mp_output261.Y__gold ,
  output [  0:0] \__mp_output262.A__gold ,
  output [  0:0] \__mp_output262.Y__gold ,
  output [  0:0] \__mp_output263.A__gold ,
  output [  0:0] \__mp_output263.Y__gold ,
  output [  0:0] \__mp_output264.A__gold ,
  output [  0:0] \__mp_output264.Y__gold ,
  output [  0:0] \__mp_output265.A__gold ,
  output [  0:0] \__mp_output265.Y__gold ,
  output [  0:0] \__mp_output266.A__gold ,
  output [  0:0] \__mp_output266.Y__gold ,
  output [  0:0] \__mp_output267.A__gold ,
  output [  0:0] \__mp_output267.Y__gold ,
  output [  0:0] \__mp_output268.A__gold ,
  output [  0:0] \__mp_output268.Y__gold ,
  output [  0:0] \__mp_output269.A__gold ,
  output [  0:0] \__mp_output269.Y__gold ,
  output [  0:0] \__mp_output270.A__gold ,
  output [  0:0] \__mp_output270.Y__gold ,
  output [  0:0] \__mp_output271.A__gold ,
  output [  0:0] \__mp_output271.Y__gold ,
  output [  0:0] \__mp_output272.A__gold ,
  output [  0:0] \__mp_output272.Y__gold ,
  output [  0:0] \__mp_output273.A__gold ,
  output [  0:0] \__mp_output273.Y__gold ,
  output [  0:0] \__mp_output274.A__gold ,
  output [  0:0] \__mp_output274.Y__gold ,
  output [  0:0] \__mp_output275.A__gold ,
  output [  0:0] \__mp_output275.Y__gold ,
  output [  0:0] \__mp_output276.A__gold ,
  output [  0:0] \__mp_output276.Y__gold ,
  output [  0:0] \__mp_output277.A__gold ,
  output [  0:0] \__mp_output277.Y__gold ,
  output [  0:0] \__mp_output278.A__gold ,
  output [  0:0] \__mp_output278.Y__gold ,
  output [  0:0] \__mp_output279.A__gold ,
  output [  0:0] \__mp_output279.Y__gold ,
  output [  0:0] \__mp_output280.A__gold ,
  output [  0:0] \__mp_output280.Y__gold ,
  output [  0:0] \__mp_output281.A__gold ,
  output [  0:0] \__mp_output281.Y__gold ,
  output [  0:0] \__mp_output282.A__gold ,
  output [  0:0] \__mp_output282.Y__gold ,
  output [  0:0] \__mp_output283.A__gold ,
  output [  0:0] \__mp_output283.Y__gold ,
  output [  0:0] \__mp_output284.A__gold ,
  output [  0:0] \__mp_output284.Y__gold ,
  output [  0:0] \__mp_output285.A__gold ,
  output [  0:0] \__mp_output285.Y__gold ,
  output [  0:0] \__mp_output286.A__gold ,
  output [  0:0] \__mp_output286.Y__gold ,
  output [  0:0] \__mp_output287.A__gold ,
  output [  0:0] \__mp_output287.Y__gold ,
  output [  0:0] \__mp_output288.A__gold ,
  output [  0:0] \__mp_output288.Y__gold ,
  output [  0:0] \__mp_output289.A__gold ,
  output [  0:0] \__mp_output289.Y__gold ,
  output [  0:0] \__mp_output290.A__gold ,
  output [  0:0] \__mp_output290.Y__gold ,
  output [  0:0] \__mp_output291.A__gold ,
  output [  0:0] \__mp_output291.Y__gold ,
  output [  0:0] \__mp_output292.A__gold ,
  output [  0:0] \__mp_output292.Y__gold ,
  output [  0:0] \__mp_output293.A__gold ,
  output [  0:0] \__mp_output293.Y__gold ,
  output [  0:0] \__mp_output294.A__gold ,
  output [  0:0] \__mp_output294.Y__gold ,
  output [  0:0] \__mp_output295.A__gold ,
  output [  0:0] \__mp_output295.Y__gold ,
  output [  0:0] \__mp_output296.A__gold ,
  output [  0:0] \__mp_output296.Y__gold ,
  output [  0:0] \__mp_output297.A__gold ,
  output [  0:0] \__mp_output297.Y__gold ,
  output [  0:0] \__mp_output298.A__gold ,
  output [  0:0] \__mp_output298.Y__gold ,
  output [  0:0] \__mp_output299.A__gold ,
  output [  0:0] \__mp_output299.Y__gold ,
  output [  0:0] \__mp_output300.A__gold ,
  output [  0:0] \__mp_output300.Y__gold ,
  output [  0:0] \__mp_output301.A__gold ,
  output [  0:0] \__mp_output301.Y__gold ,
  output [  0:0] \__mp_output302.A__gold ,
  output [  0:0] \__mp_output302.Y__gold ,
  output [  0:0] \__mp_output303.A__gold ,
  output [  0:0] \__mp_output303.Y__gold ,
  output [  0:0] \__mp_output304.A__gold ,
  output [  0:0] \__mp_output304.Y__gold ,
  output [  0:0] \__mp_output305.A__gold ,
  output [  0:0] \__mp_output305.Y__gold ,
  output [  0:0] \__mp_output306.A__gold ,
  output [  0:0] \__mp_output306.Y__gold ,
  output [  0:0] \__mp_output307.A__gold ,
  output [  0:0] \__mp_output307.Y__gold ,
  output [  0:0] \__mp_output308.A__gold ,
  output [  0:0] \__mp_output308.Y__gold ,
  output [  0:0] \__mp_output309.A__gold ,
  output [  0:0] \__mp_output309.Y__gold ,
  output [  0:0] \__mp_output310.A__gold ,
  output [  0:0] \__mp_output310.Y__gold ,
  output [  0:0] \__mp_output311.A__gold ,
  output [  0:0] \__mp_output311.Y__gold ,
  output [  0:0] \__mp_output312.A__gold ,
  output [  0:0] \__mp_output312.Y__gold ,
  output [  0:0] \__mp_output313.A__gold ,
  output [  0:0] \__mp_output313.Y__gold ,
  output [  0:0] \__mp_output314.A__gold ,
  output [  0:0] \__mp_output314.Y__gold ,
  output [  0:0] \__mp_output315.A__gold ,
  output [  0:0] \__mp_output315.Y__gold ,
  output [  0:0] \__mp_output316.A__gold ,
  output [  0:0] \__mp_output316.Y__gold ,
  output [  0:0] \__mp_output317.A__gold ,
  output [  0:0] \__mp_output317.Y__gold ,
  output [  0:0] \__mp_output318.A__gold ,
  output [  0:0] \__mp_output318.Y__gold ,
  output [  0:0] \__mp_output319.A__gold ,
  output [  0:0] \__mp_output319.Y__gold ,
  output [  0:0] \__mp_output320.A__gold ,
  output [  0:0] \__mp_output320.Y__gold ,
  output [  0:0] \__mp_output321.A__gold ,
  output [  0:0] \__mp_output321.Y__gold ,
  output [  0:0] \__mp_output322.A__gold ,
  output [  0:0] \__mp_output322.Y__gold ,
  output [  0:0] \__mp_output323.A__gold ,
  output [  0:0] \__mp_output323.Y__gold ,
  output [  0:0] \__mp_output324.A__gold ,
  output [  0:0] \__mp_output324.Y__gold ,
  output [  0:0] \__mp_output325.A__gold ,
  output [  0:0] \__mp_output325.Y__gold ,
  output [  0:0] \__mp_output326.A__gold ,
  output [  0:0] \__mp_output326.Y__gold ,
  output [  0:0] \__mp_output327.A__gold ,
  output [  0:0] \__mp_output327.Y__gold ,
  output [  0:0] \__mp_output328.A__gold ,
  output [  0:0] \__mp_output328.Y__gold ,
  output [  0:0] \__mp_output329.A__gold ,
  output [  0:0] \__mp_output329.Y__gold ,
  output [  0:0] \__mp_output330.A__gold ,
  output [  0:0] \__mp_output330.Y__gold ,
  output [  0:0] \__mp_output331.A__gold ,
  output [  0:0] \__mp_output331.Y__gold ,
  output [  0:0] \__mp_output332.A__gold ,
  output [  0:0] \__mp_output332.Y__gold ,
  output [  0:0] \__mp_output333.A__gold ,
  output [  0:0] \__mp_output333.Y__gold ,
  output [  0:0] \__mp_output334.A__gold ,
  output [  0:0] \__mp_output334.Y__gold ,
  output [  0:0] \__mp_output335.A__gold ,
  output [  0:0] \__mp_output335.Y__gold ,
  output [  0:0] \__mp_output336.A__gold ,
  output [  0:0] \__mp_output336.Y__gold ,
  output [  0:0] \__mp_output337.A__gold ,
  output [  0:0] \__mp_output337.Y__gold ,
  output [  0:0] \__mp_output338.A__gold ,
  output [  0:0] \__mp_output338.Y__gold ,
  output [  0:0] \__mp_output339.A__gold ,
  output [  0:0] \__mp_output339.Y__gold ,
  output [  0:0] \__mp_output340.A__gold ,
  output [  0:0] \__mp_output340.Y__gold ,
  output [  0:0] \__mp_output341.A__gold ,
  output [  0:0] \__mp_output341.Y__gold ,
  output [  0:0] \__mp_output342.A__gold ,
  output [  0:0] \__mp_output342.Y__gold ,
  output [  0:0] \__mp_output343.A__gold ,
  output [  0:0] \__mp_output343.Y__gold ,
  output [  0:0] \__mp_output344.A__gold ,
  output [  0:0] \__mp_output344.Y__gold ,
  output [  0:0] \__mp_output345.A__gold ,
  output [  0:0] \__mp_output345.Y__gold ,
  output [  0:0] \__mp_output346.A__gold ,
  output [  0:0] \__mp_output346.Y__gold ,
  output [  0:0] \__mp_output347.A__gold ,
  output [  0:0] \__mp_output347.Y__gold ,
  output [  0:0] \__mp_output348.A__gold ,
  output [  0:0] \__mp_output348.Y__gold ,
  output [  0:0] \__mp_output349.A__gold ,
  output [  0:0] \__mp_output349.Y__gold ,
  output [  0:0] \__mp_output350.A__gold ,
  output [  0:0] \__mp_output350.Y__gold ,
  output [  0:0] \__mp_output351.A__gold ,
  output [  0:0] \__mp_output351.Y__gold ,
  output [  0:0] \__mp_output352.A__gold ,
  output [  0:0] \__mp_output352.Y__gold ,
  output [  0:0] \__mp_output353.A__gold ,
  output [  0:0] \__mp_output353.Y__gold ,
  output [  0:0] \__mp_output354.A__gold ,
  output [  0:0] \__mp_output354.Y__gold ,
  output [  0:0] \__mp_output355.A__gold ,
  output [  0:0] \__mp_output355.Y__gold ,
  output [  0:0] \__mp_output356.A__gold ,
  output [  0:0] \__mp_output356.Y__gold ,
  output [  0:0] \__mp_output357.A__gold ,
  output [  0:0] \__mp_output357.Y__gold ,
  output [  0:0] \__mp_output358.A__gold ,
  output [  0:0] \__mp_output358.Y__gold ,
  output [  0:0] \__mp_output359.A__gold ,
  output [  0:0] \__mp_output359.Y__gold ,
  output [  0:0] \__mp_output360.A__gold ,
  output [  0:0] \__mp_output360.Y__gold ,
  output [  0:0] \__mp_output361.A__gold ,
  output [  0:0] \__mp_output361.Y__gold ,
  output [  0:0] \__mp_output362.A__gold ,
  output [  0:0] \__mp_output362.Y__gold ,
  output [  0:0] \__mp_output363.A__gold ,
  output [  0:0] \__mp_output363.Y__gold ,
  output [  0:0] \__mp_output364.A__gold ,
  output [  0:0] \__mp_output364.Y__gold ,
  output [  0:0] \__mp_output365.A__gold ,
  output [  0:0] \__mp_output365.Y__gold ,
  output [  0:0] \__mp_output366.A__gold ,
  output [  0:0] \__mp_output366.Y__gold ,
  output [  0:0] \__mp_output367.A__gold ,
  output [  0:0] \__mp_output367.Y__gold ,
  output [  0:0] \__mp_output368.A__gold ,
  output [  0:0] \__mp_output368.Y__gold ,
  output [  0:0] \__mp_output369.A__gold ,
  output [  0:0] \__mp_output369.Y__gold ,
  output [  0:0] \__mp_output370.A__gold ,
  output [  0:0] \__mp_output370.Y__gold ,
  output [  0:0] \__mp_output371.A__gold ,
  output [  0:0] \__mp_output371.Y__gold ,
  output [  0:0] \__mp_output372.A__gold ,
  output [  0:0] \__mp_output372.Y__gold ,
  output [  0:0] \__mp_output373.A__gold ,
  output [  0:0] \__mp_output373.Y__gold ,
  output [  0:0] \__mp_output374.A__gold ,
  output [  0:0] \__mp_output374.Y__gold ,
  output [  0:0] \__mp_output375.A__gold ,
  output [  0:0] \__mp_output375.Y__gold ,
  output [  0:0] \__mp_output376.A__gold ,
  output [  0:0] \__mp_output376.Y__gold ,
  output [  0:0] \__mp_output377.A__gold ,
  output [  0:0] \__mp_output377.Y__gold ,
  output [  0:0] \__mp_output378.A__gold ,
  output [  0:0] \__mp_output378.Y__gold ,
  output [  0:0] \__mp_output379.A__gold ,
  output [  0:0] \__mp_output379.Y__gold ,
  output [  0:0] \__mp_output380.A__gold ,
  output [  0:0] \__mp_output380.Y__gold ,
  output [  0:0] \__mp_output381.A__gold ,
  output [  0:0] \__mp_output381.Y__gold ,
  output [  0:0] \__mp_output382.A__gold ,
  output [  0:0] \__mp_output382.Y__gold ,
  output [  0:0] \__mp_output383.A__gold ,
  output [  0:0] \__mp_output383.Y__gold ,
  output [  0:0] \__mp_output384.A__gold ,
  output [  0:0] \__mp_output384.Y__gold ,
  output [  0:0] \__mp_output385.A__gold ,
  output [  0:0] \__mp_output385.Y__gold ,
  output [  0:0] \__mp_output386.A__gold ,
  output [  0:0] \__mp_output386.Y__gold ,
  output [  0:0] \__mp_output387.A__gold ,
  output [  0:0] \__mp_output387.Y__gold ,
  output [  0:0] \__mp_sa00_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa00_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa00_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa00_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa00_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa00_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa00_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa00_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa01_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa02_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa03_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa10_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa11_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa12_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa13_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa20_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa21_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa22_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa23_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa30_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa31_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa32_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_sa33_sr[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[0]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[100]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[101]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[102]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[103]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[104]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[105]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[106]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[107]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[108]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[109]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[10]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[110]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[111]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[112]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[113]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[114]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[115]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[116]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[117]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[118]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[119]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[11]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[120]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[121]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[122]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[123]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[124]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[125]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[126]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[127]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[12]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[13]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[14]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[15]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[16]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[17]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[18]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[19]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[1]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[20]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[21]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[22]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[23]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[24]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[25]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[26]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[27]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[28]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[29]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[2]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[30]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[31]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[32]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[33]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[34]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[35]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[36]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[37]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[38]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[39]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[3]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[40]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[41]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[42]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[43]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[44]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[45]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[46]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[47]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[48]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[49]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[4]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[50]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[51]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[52]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[53]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[54]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[55]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[56]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[57]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[58]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[59]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[5]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[60]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[61]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[62]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[63]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[64]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[65]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[66]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[67]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[68]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[69]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[6]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[70]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[71]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[72]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[73]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[74]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[75]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[76]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[77]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[78]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[79]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[7]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[80]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[81]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[82]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[83]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[84]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[85]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[86]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[87]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[88]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[89]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[8]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[90]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[91]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[92]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[93]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[94]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[95]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[96]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[97]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[98]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[99]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_in_r[9]$_DFFE_PP_.CLK__gold ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.QN__gold ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gold ,
  output [  0:0] \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u0.d[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u1.d[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u2.d[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.u3.d[7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][10]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][11]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][12]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][13]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][14]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][15]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][16]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][17]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][18]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][19]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][20]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][21]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][22]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][23]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][24]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][25]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][26]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][27]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][28]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][29]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][30]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][31]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][8]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[0][9]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][10]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][11]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][12]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][13]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][14]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][15]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][16]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][17]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][18]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][19]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][20]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][21]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][22]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][23]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][24]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][25]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][26]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][27]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][28]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][29]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][30]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][31]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][8]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[1][9]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][10]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][11]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][12]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][13]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][14]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][15]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][16]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][17]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][18]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][19]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][20]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][21]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][22]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][23]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][24]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][25]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][26]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][27]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][28]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][29]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][30]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][31]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][8]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[2][9]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][0]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][10]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][11]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][12]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][13]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][14]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][15]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][16]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][17]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][18]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][19]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][1]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][20]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][21]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][22]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][23]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][24]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][25]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][26]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][27]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][28]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][29]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][2]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][30]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][31]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][3]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][4]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][5]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][6]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][7]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][8]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_u0.w[3][9]$_DFF_P_.CLK__gold ,
  output [  0:0] \__mp_clkbuf_0_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_0_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.Y__gate ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.A__gate ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.Y__gate ,
  output [  0:0] \__mp_clkload0.A__gate ,
  output [  0:0] \__mp_clkload0.Y__gate ,
  output [  0:0] \__mp_clkload1.A__gate ,
  output [  0:0] \__mp_clkload10.A__gate ,
  output [  0:0] \__mp_clkload11.A__gate ,
  output [  0:0] \__mp_clkload12.A__gate ,
  output [  0:0] \__mp_clkload13.A__gate ,
  output [  0:0] \__mp_clkload14.A__gate ,
  output [  0:0] \__mp_clkload15.A__gate ,
  output [  0:0] \__mp_clkload16.A__gate ,
  output [  0:0] \__mp_clkload17.A__gate ,
  output [  0:0] \__mp_clkload18.A__gate ,
  output [  0:0] \__mp_clkload18.Y__gate ,
  output [  0:0] \__mp_clkload19.A__gate ,
  output [  0:0] \__mp_clkload2.A__gate ,
  output [  0:0] \__mp_clkload20.A__gate ,
  output [  0:0] \__mp_clkload21.A__gate ,
  output [  0:0] \__mp_clkload22.A__gate ,
  output [  0:0] \__mp_clkload23.A__gate ,
  output [  0:0] \__mp_clkload24.A__gate ,
  output [  0:0] \__mp_clkload25.A__gate ,
  output [  0:0] \__mp_clkload26.A__gate ,
  output [  0:0] \__mp_clkload27.A__gate ,
  output [  0:0] \__mp_clkload28.A__gate ,
  output [  0:0] \__mp_clkload29.A__gate ,
  output [  0:0] \__mp_clkload3.A__gate ,
  output [  0:0] \__mp_clkload30.A__gate ,
  output [  0:0] \__mp_clkload31.A__gate ,
  output [  0:0] \__mp_clkload31.Y__gate ,
  output [  0:0] \__mp_clkload32.A__gate ,
  output [  0:0] \__mp_clkload4.A__gate ,
  output [  0:0] \__mp_clkload5.A__gate ,
  output [  0:0] \__mp_clkload6.A__gate ,
  output [  0:0] \__mp_clkload7.A__gate ,
  output [  0:0] \__mp_clkload8.A__gate ,
  output [  0:0] \__mp_clkload9.A__gate ,
  output [  0:0] \__mp_clknet_0_clk__gate ,
  output [  0:0] \__mp_clknet_2_0_0_clk__gate ,
  output [  0:0] \__mp_clknet_2_1_0_clk__gate ,
  output [  0:0] \__mp_clknet_2_2_0_clk__gate ,
  output [  0:0] \__mp_clknet_2_3_0_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_0_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_10_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_11_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_12_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_13_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_14_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_15_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_16_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_17_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_18_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_19_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_1_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_20_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_21_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_22_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_23_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_24_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_25_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_26_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_27_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_28_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_29_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_2_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_30_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_31_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_32_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_33_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_3_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_4_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_5_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_6_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_7_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_8_clk__gate ,
  output [  0:0] \__mp_clknet_leaf_9_clk__gate ,
  output [  0:0] \__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gate ,
  output [  0:0] \__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gate ,
  output [  0:0] \__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gate ,
  output [  0:0] \__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gate ,
  output [  0:0] \__mp_done$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_done$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_done$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_input1.A__gate ,
  output [  0:0] \__mp_input1.Y__gate ,
  output [  0:0] \__mp_input10.A__gate ,
  output [  0:0] \__mp_input10.Y__gate ,
  output [  0:0] \__mp_input100.A__gate ,
  output [  0:0] \__mp_input100.Y__gate ,
  output [  0:0] \__mp_input101.A__gate ,
  output [  0:0] \__mp_input101.Y__gate ,
  output [  0:0] \__mp_input102.A__gate ,
  output [  0:0] \__mp_input102.Y__gate ,
  output [  0:0] \__mp_input103.A__gate ,
  output [  0:0] \__mp_input103.Y__gate ,
  output [  0:0] \__mp_input104.A__gate ,
  output [  0:0] \__mp_input104.Y__gate ,
  output [  0:0] \__mp_input105.A__gate ,
  output [  0:0] \__mp_input105.Y__gate ,
  output [  0:0] \__mp_input106.A__gate ,
  output [  0:0] \__mp_input106.Y__gate ,
  output [  0:0] \__mp_input107.A__gate ,
  output [  0:0] \__mp_input107.Y__gate ,
  output [  0:0] \__mp_input108.A__gate ,
  output [  0:0] \__mp_input108.Y__gate ,
  output [  0:0] \__mp_input109.A__gate ,
  output [  0:0] \__mp_input109.Y__gate ,
  output [  0:0] \__mp_input11.A__gate ,
  output [  0:0] \__mp_input11.Y__gate ,
  output [  0:0] \__mp_input110.A__gate ,
  output [  0:0] \__mp_input110.Y__gate ,
  output [  0:0] \__mp_input111.A__gate ,
  output [  0:0] \__mp_input111.Y__gate ,
  output [  0:0] \__mp_input112.A__gate ,
  output [  0:0] \__mp_input112.Y__gate ,
  output [  0:0] \__mp_input113.A__gate ,
  output [  0:0] \__mp_input113.Y__gate ,
  output [  0:0] \__mp_input114.A__gate ,
  output [  0:0] \__mp_input114.Y__gate ,
  output [  0:0] \__mp_input115.A__gate ,
  output [  0:0] \__mp_input115.Y__gate ,
  output [  0:0] \__mp_input116.A__gate ,
  output [  0:0] \__mp_input116.Y__gate ,
  output [  0:0] \__mp_input117.A__gate ,
  output [  0:0] \__mp_input117.Y__gate ,
  output [  0:0] \__mp_input118.A__gate ,
  output [  0:0] \__mp_input118.Y__gate ,
  output [  0:0] \__mp_input119.A__gate ,
  output [  0:0] \__mp_input119.Y__gate ,
  output [  0:0] \__mp_input12.A__gate ,
  output [  0:0] \__mp_input12.Y__gate ,
  output [  0:0] \__mp_input120.A__gate ,
  output [  0:0] \__mp_input120.Y__gate ,
  output [  0:0] \__mp_input121.A__gate ,
  output [  0:0] \__mp_input121.Y__gate ,
  output [  0:0] \__mp_input122.A__gate ,
  output [  0:0] \__mp_input122.Y__gate ,
  output [  0:0] \__mp_input123.A__gate ,
  output [  0:0] \__mp_input123.Y__gate ,
  output [  0:0] \__mp_input124.A__gate ,
  output [  0:0] \__mp_input124.Y__gate ,
  output [  0:0] \__mp_input125.A__gate ,
  output [  0:0] \__mp_input125.Y__gate ,
  output [  0:0] \__mp_input126.A__gate ,
  output [  0:0] \__mp_input126.Y__gate ,
  output [  0:0] \__mp_input127.A__gate ,
  output [  0:0] \__mp_input127.Y__gate ,
  output [  0:0] \__mp_input128.A__gate ,
  output [  0:0] \__mp_input128.Y__gate ,
  output [  0:0] \__mp_input129.A__gate ,
  output [  0:0] \__mp_input129.Y__gate ,
  output [  0:0] \__mp_input13.A__gate ,
  output [  0:0] \__mp_input13.Y__gate ,
  output [  0:0] \__mp_input130.A__gate ,
  output [  0:0] \__mp_input130.Y__gate ,
  output [  0:0] \__mp_input131.A__gate ,
  output [  0:0] \__mp_input131.Y__gate ,
  output [  0:0] \__mp_input132.A__gate ,
  output [  0:0] \__mp_input132.Y__gate ,
  output [  0:0] \__mp_input133.A__gate ,
  output [  0:0] \__mp_input133.Y__gate ,
  output [  0:0] \__mp_input134.A__gate ,
  output [  0:0] \__mp_input134.Y__gate ,
  output [  0:0] \__mp_input135.A__gate ,
  output [  0:0] \__mp_input135.Y__gate ,
  output [  0:0] \__mp_input136.A__gate ,
  output [  0:0] \__mp_input136.Y__gate ,
  output [  0:0] \__mp_input137.A__gate ,
  output [  0:0] \__mp_input137.Y__gate ,
  output [  0:0] \__mp_input138.A__gate ,
  output [  0:0] \__mp_input138.Y__gate ,
  output [  0:0] \__mp_input139.A__gate ,
  output [  0:0] \__mp_input139.Y__gate ,
  output [  0:0] \__mp_input14.A__gate ,
  output [  0:0] \__mp_input14.Y__gate ,
  output [  0:0] \__mp_input140.A__gate ,
  output [  0:0] \__mp_input140.Y__gate ,
  output [  0:0] \__mp_input141.A__gate ,
  output [  0:0] \__mp_input141.Y__gate ,
  output [  0:0] \__mp_input142.A__gate ,
  output [  0:0] \__mp_input142.Y__gate ,
  output [  0:0] \__mp_input143.A__gate ,
  output [  0:0] \__mp_input143.Y__gate ,
  output [  0:0] \__mp_input144.A__gate ,
  output [  0:0] \__mp_input144.Y__gate ,
  output [  0:0] \__mp_input145.A__gate ,
  output [  0:0] \__mp_input145.Y__gate ,
  output [  0:0] \__mp_input146.A__gate ,
  output [  0:0] \__mp_input146.Y__gate ,
  output [  0:0] \__mp_input147.A__gate ,
  output [  0:0] \__mp_input147.Y__gate ,
  output [  0:0] \__mp_input148.A__gate ,
  output [  0:0] \__mp_input148.Y__gate ,
  output [  0:0] \__mp_input149.A__gate ,
  output [  0:0] \__mp_input149.Y__gate ,
  output [  0:0] \__mp_input15.A__gate ,
  output [  0:0] \__mp_input15.Y__gate ,
  output [  0:0] \__mp_input150.A__gate ,
  output [  0:0] \__mp_input150.Y__gate ,
  output [  0:0] \__mp_input151.A__gate ,
  output [  0:0] \__mp_input151.Y__gate ,
  output [  0:0] \__mp_input152.A__gate ,
  output [  0:0] \__mp_input152.Y__gate ,
  output [  0:0] \__mp_input153.A__gate ,
  output [  0:0] \__mp_input153.Y__gate ,
  output [  0:0] \__mp_input154.A__gate ,
  output [  0:0] \__mp_input154.Y__gate ,
  output [  0:0] \__mp_input155.A__gate ,
  output [  0:0] \__mp_input155.Y__gate ,
  output [  0:0] \__mp_input156.A__gate ,
  output [  0:0] \__mp_input156.Y__gate ,
  output [  0:0] \__mp_input157.A__gate ,
  output [  0:0] \__mp_input157.Y__gate ,
  output [  0:0] \__mp_input158.A__gate ,
  output [  0:0] \__mp_input158.Y__gate ,
  output [  0:0] \__mp_input159.A__gate ,
  output [  0:0] \__mp_input159.Y__gate ,
  output [  0:0] \__mp_input16.A__gate ,
  output [  0:0] \__mp_input16.Y__gate ,
  output [  0:0] \__mp_input160.A__gate ,
  output [  0:0] \__mp_input160.Y__gate ,
  output [  0:0] \__mp_input161.A__gate ,
  output [  0:0] \__mp_input161.Y__gate ,
  output [  0:0] \__mp_input162.A__gate ,
  output [  0:0] \__mp_input162.Y__gate ,
  output [  0:0] \__mp_input163.A__gate ,
  output [  0:0] \__mp_input163.Y__gate ,
  output [  0:0] \__mp_input164.A__gate ,
  output [  0:0] \__mp_input164.Y__gate ,
  output [  0:0] \__mp_input165.A__gate ,
  output [  0:0] \__mp_input165.Y__gate ,
  output [  0:0] \__mp_input166.A__gate ,
  output [  0:0] \__mp_input166.Y__gate ,
  output [  0:0] \__mp_input167.A__gate ,
  output [  0:0] \__mp_input167.Y__gate ,
  output [  0:0] \__mp_input168.A__gate ,
  output [  0:0] \__mp_input168.Y__gate ,
  output [  0:0] \__mp_input169.A__gate ,
  output [  0:0] \__mp_input169.Y__gate ,
  output [  0:0] \__mp_input17.A__gate ,
  output [  0:0] \__mp_input17.Y__gate ,
  output [  0:0] \__mp_input170.A__gate ,
  output [  0:0] \__mp_input170.Y__gate ,
  output [  0:0] \__mp_input171.A__gate ,
  output [  0:0] \__mp_input171.Y__gate ,
  output [  0:0] \__mp_input172.A__gate ,
  output [  0:0] \__mp_input172.Y__gate ,
  output [  0:0] \__mp_input173.A__gate ,
  output [  0:0] \__mp_input173.Y__gate ,
  output [  0:0] \__mp_input174.A__gate ,
  output [  0:0] \__mp_input174.Y__gate ,
  output [  0:0] \__mp_input175.A__gate ,
  output [  0:0] \__mp_input175.Y__gate ,
  output [  0:0] \__mp_input176.A__gate ,
  output [  0:0] \__mp_input176.Y__gate ,
  output [  0:0] \__mp_input177.A__gate ,
  output [  0:0] \__mp_input177.Y__gate ,
  output [  0:0] \__mp_input178.A__gate ,
  output [  0:0] \__mp_input178.Y__gate ,
  output [  0:0] \__mp_input179.A__gate ,
  output [  0:0] \__mp_input179.Y__gate ,
  output [  0:0] \__mp_input18.A__gate ,
  output [  0:0] \__mp_input18.Y__gate ,
  output [  0:0] \__mp_input180.A__gate ,
  output [  0:0] \__mp_input180.Y__gate ,
  output [  0:0] \__mp_input181.A__gate ,
  output [  0:0] \__mp_input181.Y__gate ,
  output [  0:0] \__mp_input182.A__gate ,
  output [  0:0] \__mp_input182.Y__gate ,
  output [  0:0] \__mp_input183.A__gate ,
  output [  0:0] \__mp_input183.Y__gate ,
  output [  0:0] \__mp_input184.A__gate ,
  output [  0:0] \__mp_input184.Y__gate ,
  output [  0:0] \__mp_input185.A__gate ,
  output [  0:0] \__mp_input185.Y__gate ,
  output [  0:0] \__mp_input186.A__gate ,
  output [  0:0] \__mp_input186.Y__gate ,
  output [  0:0] \__mp_input187.A__gate ,
  output [  0:0] \__mp_input187.Y__gate ,
  output [  0:0] \__mp_input188.A__gate ,
  output [  0:0] \__mp_input188.Y__gate ,
  output [  0:0] \__mp_input189.A__gate ,
  output [  0:0] \__mp_input189.Y__gate ,
  output [  0:0] \__mp_input19.A__gate ,
  output [  0:0] \__mp_input19.Y__gate ,
  output [  0:0] \__mp_input190.A__gate ,
  output [  0:0] \__mp_input190.Y__gate ,
  output [  0:0] \__mp_input191.A__gate ,
  output [  0:0] \__mp_input191.Y__gate ,
  output [  0:0] \__mp_input192.A__gate ,
  output [  0:0] \__mp_input192.Y__gate ,
  output [  0:0] \__mp_input193.A__gate ,
  output [  0:0] \__mp_input193.Y__gate ,
  output [  0:0] \__mp_input194.A__gate ,
  output [  0:0] \__mp_input194.Y__gate ,
  output [  0:0] \__mp_input195.A__gate ,
  output [  0:0] \__mp_input195.Y__gate ,
  output [  0:0] \__mp_input196.A__gate ,
  output [  0:0] \__mp_input196.Y__gate ,
  output [  0:0] \__mp_input197.A__gate ,
  output [  0:0] \__mp_input197.Y__gate ,
  output [  0:0] \__mp_input198.A__gate ,
  output [  0:0] \__mp_input198.Y__gate ,
  output [  0:0] \__mp_input199.A__gate ,
  output [  0:0] \__mp_input199.Y__gate ,
  output [  0:0] \__mp_input2.A__gate ,
  output [  0:0] \__mp_input2.Y__gate ,
  output [  0:0] \__mp_input20.A__gate ,
  output [  0:0] \__mp_input20.Y__gate ,
  output [  0:0] \__mp_input200.A__gate ,
  output [  0:0] \__mp_input200.Y__gate ,
  output [  0:0] \__mp_input201.A__gate ,
  output [  0:0] \__mp_input201.Y__gate ,
  output [  0:0] \__mp_input202.A__gate ,
  output [  0:0] \__mp_input202.Y__gate ,
  output [  0:0] \__mp_input203.A__gate ,
  output [  0:0] \__mp_input203.Y__gate ,
  output [  0:0] \__mp_input204.A__gate ,
  output [  0:0] \__mp_input204.Y__gate ,
  output [  0:0] \__mp_input205.A__gate ,
  output [  0:0] \__mp_input205.Y__gate ,
  output [  0:0] \__mp_input206.A__gate ,
  output [  0:0] \__mp_input206.Y__gate ,
  output [  0:0] \__mp_input207.A__gate ,
  output [  0:0] \__mp_input207.Y__gate ,
  output [  0:0] \__mp_input208.A__gate ,
  output [  0:0] \__mp_input208.Y__gate ,
  output [  0:0] \__mp_input209.A__gate ,
  output [  0:0] \__mp_input209.Y__gate ,
  output [  0:0] \__mp_input21.A__gate ,
  output [  0:0] \__mp_input21.Y__gate ,
  output [  0:0] \__mp_input210.A__gate ,
  output [  0:0] \__mp_input210.Y__gate ,
  output [  0:0] \__mp_input211.A__gate ,
  output [  0:0] \__mp_input211.Y__gate ,
  output [  0:0] \__mp_input212.A__gate ,
  output [  0:0] \__mp_input212.Y__gate ,
  output [  0:0] \__mp_input213.A__gate ,
  output [  0:0] \__mp_input213.Y__gate ,
  output [  0:0] \__mp_input214.A__gate ,
  output [  0:0] \__mp_input214.Y__gate ,
  output [  0:0] \__mp_input215.A__gate ,
  output [  0:0] \__mp_input215.Y__gate ,
  output [  0:0] \__mp_input216.A__gate ,
  output [  0:0] \__mp_input216.Y__gate ,
  output [  0:0] \__mp_input217.A__gate ,
  output [  0:0] \__mp_input217.Y__gate ,
  output [  0:0] \__mp_input218.A__gate ,
  output [  0:0] \__mp_input218.Y__gate ,
  output [  0:0] \__mp_input219.A__gate ,
  output [  0:0] \__mp_input219.Y__gate ,
  output [  0:0] \__mp_input22.A__gate ,
  output [  0:0] \__mp_input22.Y__gate ,
  output [  0:0] \__mp_input220.A__gate ,
  output [  0:0] \__mp_input220.Y__gate ,
  output [  0:0] \__mp_input221.A__gate ,
  output [  0:0] \__mp_input221.Y__gate ,
  output [  0:0] \__mp_input222.A__gate ,
  output [  0:0] \__mp_input222.Y__gate ,
  output [  0:0] \__mp_input223.A__gate ,
  output [  0:0] \__mp_input223.Y__gate ,
  output [  0:0] \__mp_input224.A__gate ,
  output [  0:0] \__mp_input224.Y__gate ,
  output [  0:0] \__mp_input225.A__gate ,
  output [  0:0] \__mp_input225.Y__gate ,
  output [  0:0] \__mp_input226.A__gate ,
  output [  0:0] \__mp_input226.Y__gate ,
  output [  0:0] \__mp_input227.A__gate ,
  output [  0:0] \__mp_input227.Y__gate ,
  output [  0:0] \__mp_input228.A__gate ,
  output [  0:0] \__mp_input228.Y__gate ,
  output [  0:0] \__mp_input229.A__gate ,
  output [  0:0] \__mp_input229.Y__gate ,
  output [  0:0] \__mp_input23.A__gate ,
  output [  0:0] \__mp_input23.Y__gate ,
  output [  0:0] \__mp_input230.A__gate ,
  output [  0:0] \__mp_input230.Y__gate ,
  output [  0:0] \__mp_input231.A__gate ,
  output [  0:0] \__mp_input231.Y__gate ,
  output [  0:0] \__mp_input232.A__gate ,
  output [  0:0] \__mp_input232.Y__gate ,
  output [  0:0] \__mp_input233.A__gate ,
  output [  0:0] \__mp_input233.Y__gate ,
  output [  0:0] \__mp_input234.A__gate ,
  output [  0:0] \__mp_input234.Y__gate ,
  output [  0:0] \__mp_input235.A__gate ,
  output [  0:0] \__mp_input235.Y__gate ,
  output [  0:0] \__mp_input236.A__gate ,
  output [  0:0] \__mp_input236.Y__gate ,
  output [  0:0] \__mp_input237.A__gate ,
  output [  0:0] \__mp_input237.Y__gate ,
  output [  0:0] \__mp_input238.A__gate ,
  output [  0:0] \__mp_input238.Y__gate ,
  output [  0:0] \__mp_input239.A__gate ,
  output [  0:0] \__mp_input239.Y__gate ,
  output [  0:0] \__mp_input24.A__gate ,
  output [  0:0] \__mp_input24.Y__gate ,
  output [  0:0] \__mp_input240.A__gate ,
  output [  0:0] \__mp_input240.Y__gate ,
  output [  0:0] \__mp_input241.A__gate ,
  output [  0:0] \__mp_input241.Y__gate ,
  output [  0:0] \__mp_input242.A__gate ,
  output [  0:0] \__mp_input242.Y__gate ,
  output [  0:0] \__mp_input243.A__gate ,
  output [  0:0] \__mp_input243.Y__gate ,
  output [  0:0] \__mp_input244.A__gate ,
  output [  0:0] \__mp_input244.Y__gate ,
  output [  0:0] \__mp_input245.A__gate ,
  output [  0:0] \__mp_input245.Y__gate ,
  output [  0:0] \__mp_input246.A__gate ,
  output [  0:0] \__mp_input246.Y__gate ,
  output [  0:0] \__mp_input247.A__gate ,
  output [  0:0] \__mp_input247.Y__gate ,
  output [  0:0] \__mp_input248.A__gate ,
  output [  0:0] \__mp_input248.Y__gate ,
  output [  0:0] \__mp_input249.A__gate ,
  output [  0:0] \__mp_input249.Y__gate ,
  output [  0:0] \__mp_input25.A__gate ,
  output [  0:0] \__mp_input25.Y__gate ,
  output [  0:0] \__mp_input250.A__gate ,
  output [  0:0] \__mp_input250.Y__gate ,
  output [  0:0] \__mp_input251.A__gate ,
  output [  0:0] \__mp_input251.Y__gate ,
  output [  0:0] \__mp_input252.A__gate ,
  output [  0:0] \__mp_input252.Y__gate ,
  output [  0:0] \__mp_input253.A__gate ,
  output [  0:0] \__mp_input253.Y__gate ,
  output [  0:0] \__mp_input254.A__gate ,
  output [  0:0] \__mp_input254.Y__gate ,
  output [  0:0] \__mp_input255.A__gate ,
  output [  0:0] \__mp_input255.Y__gate ,
  output [  0:0] \__mp_input256.A__gate ,
  output [  0:0] \__mp_input256.Y__gate ,
  output [  0:0] \__mp_input257.A__gate ,
  output [  0:0] \__mp_input257.Y__gate ,
  output [  0:0] \__mp_input258.A__gate ,
  output [  0:0] \__mp_input258.Y__gate ,
  output [  0:0] \__mp_input26.A__gate ,
  output [  0:0] \__mp_input26.Y__gate ,
  output [  0:0] \__mp_input27.A__gate ,
  output [  0:0] \__mp_input27.Y__gate ,
  output [  0:0] \__mp_input28.A__gate ,
  output [  0:0] \__mp_input28.Y__gate ,
  output [  0:0] \__mp_input29.A__gate ,
  output [  0:0] \__mp_input29.Y__gate ,
  output [  0:0] \__mp_input3.A__gate ,
  output [  0:0] \__mp_input3.Y__gate ,
  output [  0:0] \__mp_input30.A__gate ,
  output [  0:0] \__mp_input30.Y__gate ,
  output [  0:0] \__mp_input31.A__gate ,
  output [  0:0] \__mp_input31.Y__gate ,
  output [  0:0] \__mp_input32.A__gate ,
  output [  0:0] \__mp_input32.Y__gate ,
  output [  0:0] \__mp_input33.A__gate ,
  output [  0:0] \__mp_input33.Y__gate ,
  output [  0:0] \__mp_input34.A__gate ,
  output [  0:0] \__mp_input34.Y__gate ,
  output [  0:0] \__mp_input35.A__gate ,
  output [  0:0] \__mp_input35.Y__gate ,
  output [  0:0] \__mp_input36.A__gate ,
  output [  0:0] \__mp_input36.Y__gate ,
  output [  0:0] \__mp_input37.A__gate ,
  output [  0:0] \__mp_input37.Y__gate ,
  output [  0:0] \__mp_input38.A__gate ,
  output [  0:0] \__mp_input38.Y__gate ,
  output [  0:0] \__mp_input39.A__gate ,
  output [  0:0] \__mp_input39.Y__gate ,
  output [  0:0] \__mp_input4.A__gate ,
  output [  0:0] \__mp_input4.Y__gate ,
  output [  0:0] \__mp_input40.A__gate ,
  output [  0:0] \__mp_input40.Y__gate ,
  output [  0:0] \__mp_input41.A__gate ,
  output [  0:0] \__mp_input41.Y__gate ,
  output [  0:0] \__mp_input42.A__gate ,
  output [  0:0] \__mp_input42.Y__gate ,
  output [  0:0] \__mp_input43.A__gate ,
  output [  0:0] \__mp_input43.Y__gate ,
  output [  0:0] \__mp_input44.A__gate ,
  output [  0:0] \__mp_input44.Y__gate ,
  output [  0:0] \__mp_input45.A__gate ,
  output [  0:0] \__mp_input45.Y__gate ,
  output [  0:0] \__mp_input46.A__gate ,
  output [  0:0] \__mp_input46.Y__gate ,
  output [  0:0] \__mp_input47.A__gate ,
  output [  0:0] \__mp_input47.Y__gate ,
  output [  0:0] \__mp_input48.A__gate ,
  output [  0:0] \__mp_input48.Y__gate ,
  output [  0:0] \__mp_input49.A__gate ,
  output [  0:0] \__mp_input49.Y__gate ,
  output [  0:0] \__mp_input5.A__gate ,
  output [  0:0] \__mp_input5.Y__gate ,
  output [  0:0] \__mp_input50.A__gate ,
  output [  0:0] \__mp_input50.Y__gate ,
  output [  0:0] \__mp_input51.A__gate ,
  output [  0:0] \__mp_input51.Y__gate ,
  output [  0:0] \__mp_input52.A__gate ,
  output [  0:0] \__mp_input52.Y__gate ,
  output [  0:0] \__mp_input53.A__gate ,
  output [  0:0] \__mp_input53.Y__gate ,
  output [  0:0] \__mp_input54.A__gate ,
  output [  0:0] \__mp_input54.Y__gate ,
  output [  0:0] \__mp_input55.A__gate ,
  output [  0:0] \__mp_input55.Y__gate ,
  output [  0:0] \__mp_input56.A__gate ,
  output [  0:0] \__mp_input56.Y__gate ,
  output [  0:0] \__mp_input57.A__gate ,
  output [  0:0] \__mp_input57.Y__gate ,
  output [  0:0] \__mp_input58.A__gate ,
  output [  0:0] \__mp_input58.Y__gate ,
  output [  0:0] \__mp_input59.A__gate ,
  output [  0:0] \__mp_input59.Y__gate ,
  output [  0:0] \__mp_input6.A__gate ,
  output [  0:0] \__mp_input6.Y__gate ,
  output [  0:0] \__mp_input60.A__gate ,
  output [  0:0] \__mp_input60.Y__gate ,
  output [  0:0] \__mp_input61.A__gate ,
  output [  0:0] \__mp_input61.Y__gate ,
  output [  0:0] \__mp_input62.A__gate ,
  output [  0:0] \__mp_input62.Y__gate ,
  output [  0:0] \__mp_input63.A__gate ,
  output [  0:0] \__mp_input63.Y__gate ,
  output [  0:0] \__mp_input64.A__gate ,
  output [  0:0] \__mp_input64.Y__gate ,
  output [  0:0] \__mp_input65.A__gate ,
  output [  0:0] \__mp_input65.Y__gate ,
  output [  0:0] \__mp_input66.A__gate ,
  output [  0:0] \__mp_input66.Y__gate ,
  output [  0:0] \__mp_input67.A__gate ,
  output [  0:0] \__mp_input67.Y__gate ,
  output [  0:0] \__mp_input68.A__gate ,
  output [  0:0] \__mp_input68.Y__gate ,
  output [  0:0] \__mp_input69.A__gate ,
  output [  0:0] \__mp_input69.Y__gate ,
  output [  0:0] \__mp_input7.A__gate ,
  output [  0:0] \__mp_input7.Y__gate ,
  output [  0:0] \__mp_input70.A__gate ,
  output [  0:0] \__mp_input70.Y__gate ,
  output [  0:0] \__mp_input71.A__gate ,
  output [  0:0] \__mp_input71.Y__gate ,
  output [  0:0] \__mp_input72.A__gate ,
  output [  0:0] \__mp_input72.Y__gate ,
  output [  0:0] \__mp_input73.A__gate ,
  output [  0:0] \__mp_input73.Y__gate ,
  output [  0:0] \__mp_input74.A__gate ,
  output [  0:0] \__mp_input74.Y__gate ,
  output [  0:0] \__mp_input75.A__gate ,
  output [  0:0] \__mp_input75.Y__gate ,
  output [  0:0] \__mp_input76.A__gate ,
  output [  0:0] \__mp_input76.Y__gate ,
  output [  0:0] \__mp_input77.A__gate ,
  output [  0:0] \__mp_input77.Y__gate ,
  output [  0:0] \__mp_input78.A__gate ,
  output [  0:0] \__mp_input78.Y__gate ,
  output [  0:0] \__mp_input79.A__gate ,
  output [  0:0] \__mp_input79.Y__gate ,
  output [  0:0] \__mp_input8.A__gate ,
  output [  0:0] \__mp_input8.Y__gate ,
  output [  0:0] \__mp_input80.A__gate ,
  output [  0:0] \__mp_input80.Y__gate ,
  output [  0:0] \__mp_input81.A__gate ,
  output [  0:0] \__mp_input81.Y__gate ,
  output [  0:0] \__mp_input82.A__gate ,
  output [  0:0] \__mp_input82.Y__gate ,
  output [  0:0] \__mp_input83.A__gate ,
  output [  0:0] \__mp_input83.Y__gate ,
  output [  0:0] \__mp_input84.A__gate ,
  output [  0:0] \__mp_input84.Y__gate ,
  output [  0:0] \__mp_input85.A__gate ,
  output [  0:0] \__mp_input85.Y__gate ,
  output [  0:0] \__mp_input86.A__gate ,
  output [  0:0] \__mp_input86.Y__gate ,
  output [  0:0] \__mp_input87.A__gate ,
  output [  0:0] \__mp_input87.Y__gate ,
  output [  0:0] \__mp_input88.A__gate ,
  output [  0:0] \__mp_input88.Y__gate ,
  output [  0:0] \__mp_input89.A__gate ,
  output [  0:0] \__mp_input89.Y__gate ,
  output [  0:0] \__mp_input9.A__gate ,
  output [  0:0] \__mp_input9.Y__gate ,
  output [  0:0] \__mp_input90.A__gate ,
  output [  0:0] \__mp_input90.Y__gate ,
  output [  0:0] \__mp_input91.A__gate ,
  output [  0:0] \__mp_input91.Y__gate ,
  output [  0:0] \__mp_input92.A__gate ,
  output [  0:0] \__mp_input92.Y__gate ,
  output [  0:0] \__mp_input93.A__gate ,
  output [  0:0] \__mp_input93.Y__gate ,
  output [  0:0] \__mp_input94.A__gate ,
  output [  0:0] \__mp_input94.Y__gate ,
  output [  0:0] \__mp_input95.A__gate ,
  output [  0:0] \__mp_input95.Y__gate ,
  output [  0:0] \__mp_input96.A__gate ,
  output [  0:0] \__mp_input96.Y__gate ,
  output [  0:0] \__mp_input97.A__gate ,
  output [  0:0] \__mp_input97.Y__gate ,
  output [  0:0] \__mp_input98.A__gate ,
  output [  0:0] \__mp_input98.Y__gate ,
  output [  0:0] \__mp_input99.A__gate ,
  output [  0:0] \__mp_input99.Y__gate ,
  output [  0:0] \__mp_ld_r$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_ld_r$_DFF_P_.D__gate ,
  output [  0:0] \__mp_output259.A__gate ,
  output [  0:0] \__mp_output259.Y__gate ,
  output [  0:0] \__mp_output260.A__gate ,
  output [  0:0] \__mp_output260.Y__gate ,
  output [  0:0] \__mp_output261.A__gate ,
  output [  0:0] \__mp_output261.Y__gate ,
  output [  0:0] \__mp_output262.A__gate ,
  output [  0:0] \__mp_output262.Y__gate ,
  output [  0:0] \__mp_output263.A__gate ,
  output [  0:0] \__mp_output263.Y__gate ,
  output [  0:0] \__mp_output264.A__gate ,
  output [  0:0] \__mp_output264.Y__gate ,
  output [  0:0] \__mp_output265.A__gate ,
  output [  0:0] \__mp_output265.Y__gate ,
  output [  0:0] \__mp_output266.A__gate ,
  output [  0:0] \__mp_output266.Y__gate ,
  output [  0:0] \__mp_output267.A__gate ,
  output [  0:0] \__mp_output267.Y__gate ,
  output [  0:0] \__mp_output268.A__gate ,
  output [  0:0] \__mp_output268.Y__gate ,
  output [  0:0] \__mp_output269.A__gate ,
  output [  0:0] \__mp_output269.Y__gate ,
  output [  0:0] \__mp_output270.A__gate ,
  output [  0:0] \__mp_output270.Y__gate ,
  output [  0:0] \__mp_output271.A__gate ,
  output [  0:0] \__mp_output271.Y__gate ,
  output [  0:0] \__mp_output272.A__gate ,
  output [  0:0] \__mp_output272.Y__gate ,
  output [  0:0] \__mp_output273.A__gate ,
  output [  0:0] \__mp_output273.Y__gate ,
  output [  0:0] \__mp_output274.A__gate ,
  output [  0:0] \__mp_output274.Y__gate ,
  output [  0:0] \__mp_output275.A__gate ,
  output [  0:0] \__mp_output275.Y__gate ,
  output [  0:0] \__mp_output276.A__gate ,
  output [  0:0] \__mp_output276.Y__gate ,
  output [  0:0] \__mp_output277.A__gate ,
  output [  0:0] \__mp_output277.Y__gate ,
  output [  0:0] \__mp_output278.A__gate ,
  output [  0:0] \__mp_output278.Y__gate ,
  output [  0:0] \__mp_output279.A__gate ,
  output [  0:0] \__mp_output279.Y__gate ,
  output [  0:0] \__mp_output280.A__gate ,
  output [  0:0] \__mp_output280.Y__gate ,
  output [  0:0] \__mp_output281.A__gate ,
  output [  0:0] \__mp_output281.Y__gate ,
  output [  0:0] \__mp_output282.A__gate ,
  output [  0:0] \__mp_output282.Y__gate ,
  output [  0:0] \__mp_output283.A__gate ,
  output [  0:0] \__mp_output283.Y__gate ,
  output [  0:0] \__mp_output284.A__gate ,
  output [  0:0] \__mp_output284.Y__gate ,
  output [  0:0] \__mp_output285.A__gate ,
  output [  0:0] \__mp_output285.Y__gate ,
  output [  0:0] \__mp_output286.A__gate ,
  output [  0:0] \__mp_output286.Y__gate ,
  output [  0:0] \__mp_output287.A__gate ,
  output [  0:0] \__mp_output287.Y__gate ,
  output [  0:0] \__mp_output288.A__gate ,
  output [  0:0] \__mp_output288.Y__gate ,
  output [  0:0] \__mp_output289.A__gate ,
  output [  0:0] \__mp_output289.Y__gate ,
  output [  0:0] \__mp_output290.A__gate ,
  output [  0:0] \__mp_output290.Y__gate ,
  output [  0:0] \__mp_output291.A__gate ,
  output [  0:0] \__mp_output291.Y__gate ,
  output [  0:0] \__mp_output292.A__gate ,
  output [  0:0] \__mp_output292.Y__gate ,
  output [  0:0] \__mp_output293.A__gate ,
  output [  0:0] \__mp_output293.Y__gate ,
  output [  0:0] \__mp_output294.A__gate ,
  output [  0:0] \__mp_output294.Y__gate ,
  output [  0:0] \__mp_output295.A__gate ,
  output [  0:0] \__mp_output295.Y__gate ,
  output [  0:0] \__mp_output296.A__gate ,
  output [  0:0] \__mp_output296.Y__gate ,
  output [  0:0] \__mp_output297.A__gate ,
  output [  0:0] \__mp_output297.Y__gate ,
  output [  0:0] \__mp_output298.A__gate ,
  output [  0:0] \__mp_output298.Y__gate ,
  output [  0:0] \__mp_output299.A__gate ,
  output [  0:0] \__mp_output299.Y__gate ,
  output [  0:0] \__mp_output300.A__gate ,
  output [  0:0] \__mp_output300.Y__gate ,
  output [  0:0] \__mp_output301.A__gate ,
  output [  0:0] \__mp_output301.Y__gate ,
  output [  0:0] \__mp_output302.A__gate ,
  output [  0:0] \__mp_output302.Y__gate ,
  output [  0:0] \__mp_output303.A__gate ,
  output [  0:0] \__mp_output303.Y__gate ,
  output [  0:0] \__mp_output304.A__gate ,
  output [  0:0] \__mp_output304.Y__gate ,
  output [  0:0] \__mp_output305.A__gate ,
  output [  0:0] \__mp_output305.Y__gate ,
  output [  0:0] \__mp_output306.A__gate ,
  output [  0:0] \__mp_output306.Y__gate ,
  output [  0:0] \__mp_output307.A__gate ,
  output [  0:0] \__mp_output307.Y__gate ,
  output [  0:0] \__mp_output308.A__gate ,
  output [  0:0] \__mp_output308.Y__gate ,
  output [  0:0] \__mp_output309.A__gate ,
  output [  0:0] \__mp_output309.Y__gate ,
  output [  0:0] \__mp_output310.A__gate ,
  output [  0:0] \__mp_output310.Y__gate ,
  output [  0:0] \__mp_output311.A__gate ,
  output [  0:0] \__mp_output311.Y__gate ,
  output [  0:0] \__mp_output312.A__gate ,
  output [  0:0] \__mp_output312.Y__gate ,
  output [  0:0] \__mp_output313.A__gate ,
  output [  0:0] \__mp_output313.Y__gate ,
  output [  0:0] \__mp_output314.A__gate ,
  output [  0:0] \__mp_output314.Y__gate ,
  output [  0:0] \__mp_output315.A__gate ,
  output [  0:0] \__mp_output315.Y__gate ,
  output [  0:0] \__mp_output316.A__gate ,
  output [  0:0] \__mp_output316.Y__gate ,
  output [  0:0] \__mp_output317.A__gate ,
  output [  0:0] \__mp_output317.Y__gate ,
  output [  0:0] \__mp_output318.A__gate ,
  output [  0:0] \__mp_output318.Y__gate ,
  output [  0:0] \__mp_output319.A__gate ,
  output [  0:0] \__mp_output319.Y__gate ,
  output [  0:0] \__mp_output320.A__gate ,
  output [  0:0] \__mp_output320.Y__gate ,
  output [  0:0] \__mp_output321.A__gate ,
  output [  0:0] \__mp_output321.Y__gate ,
  output [  0:0] \__mp_output322.A__gate ,
  output [  0:0] \__mp_output322.Y__gate ,
  output [  0:0] \__mp_output323.A__gate ,
  output [  0:0] \__mp_output323.Y__gate ,
  output [  0:0] \__mp_output324.A__gate ,
  output [  0:0] \__mp_output324.Y__gate ,
  output [  0:0] \__mp_output325.A__gate ,
  output [  0:0] \__mp_output325.Y__gate ,
  output [  0:0] \__mp_output326.A__gate ,
  output [  0:0] \__mp_output326.Y__gate ,
  output [  0:0] \__mp_output327.A__gate ,
  output [  0:0] \__mp_output327.Y__gate ,
  output [  0:0] \__mp_output328.A__gate ,
  output [  0:0] \__mp_output328.Y__gate ,
  output [  0:0] \__mp_output329.A__gate ,
  output [  0:0] \__mp_output329.Y__gate ,
  output [  0:0] \__mp_output330.A__gate ,
  output [  0:0] \__mp_output330.Y__gate ,
  output [  0:0] \__mp_output331.A__gate ,
  output [  0:0] \__mp_output331.Y__gate ,
  output [  0:0] \__mp_output332.A__gate ,
  output [  0:0] \__mp_output332.Y__gate ,
  output [  0:0] \__mp_output333.A__gate ,
  output [  0:0] \__mp_output333.Y__gate ,
  output [  0:0] \__mp_output334.A__gate ,
  output [  0:0] \__mp_output334.Y__gate ,
  output [  0:0] \__mp_output335.A__gate ,
  output [  0:0] \__mp_output335.Y__gate ,
  output [  0:0] \__mp_output336.A__gate ,
  output [  0:0] \__mp_output336.Y__gate ,
  output [  0:0] \__mp_output337.A__gate ,
  output [  0:0] \__mp_output337.Y__gate ,
  output [  0:0] \__mp_output338.A__gate ,
  output [  0:0] \__mp_output338.Y__gate ,
  output [  0:0] \__mp_output339.A__gate ,
  output [  0:0] \__mp_output339.Y__gate ,
  output [  0:0] \__mp_output340.A__gate ,
  output [  0:0] \__mp_output340.Y__gate ,
  output [  0:0] \__mp_output341.A__gate ,
  output [  0:0] \__mp_output341.Y__gate ,
  output [  0:0] \__mp_output342.A__gate ,
  output [  0:0] \__mp_output342.Y__gate ,
  output [  0:0] \__mp_output343.A__gate ,
  output [  0:0] \__mp_output343.Y__gate ,
  output [  0:0] \__mp_output344.A__gate ,
  output [  0:0] \__mp_output344.Y__gate ,
  output [  0:0] \__mp_output345.A__gate ,
  output [  0:0] \__mp_output345.Y__gate ,
  output [  0:0] \__mp_output346.A__gate ,
  output [  0:0] \__mp_output346.Y__gate ,
  output [  0:0] \__mp_output347.A__gate ,
  output [  0:0] \__mp_output347.Y__gate ,
  output [  0:0] \__mp_output348.A__gate ,
  output [  0:0] \__mp_output348.Y__gate ,
  output [  0:0] \__mp_output349.A__gate ,
  output [  0:0] \__mp_output349.Y__gate ,
  output [  0:0] \__mp_output350.A__gate ,
  output [  0:0] \__mp_output350.Y__gate ,
  output [  0:0] \__mp_output351.A__gate ,
  output [  0:0] \__mp_output351.Y__gate ,
  output [  0:0] \__mp_output352.A__gate ,
  output [  0:0] \__mp_output352.Y__gate ,
  output [  0:0] \__mp_output353.A__gate ,
  output [  0:0] \__mp_output353.Y__gate ,
  output [  0:0] \__mp_output354.A__gate ,
  output [  0:0] \__mp_output354.Y__gate ,
  output [  0:0] \__mp_output355.A__gate ,
  output [  0:0] \__mp_output355.Y__gate ,
  output [  0:0] \__mp_output356.A__gate ,
  output [  0:0] \__mp_output356.Y__gate ,
  output [  0:0] \__mp_output357.A__gate ,
  output [  0:0] \__mp_output357.Y__gate ,
  output [  0:0] \__mp_output358.A__gate ,
  output [  0:0] \__mp_output358.Y__gate ,
  output [  0:0] \__mp_output359.A__gate ,
  output [  0:0] \__mp_output359.Y__gate ,
  output [  0:0] \__mp_output360.A__gate ,
  output [  0:0] \__mp_output360.Y__gate ,
  output [  0:0] \__mp_output361.A__gate ,
  output [  0:0] \__mp_output361.Y__gate ,
  output [  0:0] \__mp_output362.A__gate ,
  output [  0:0] \__mp_output362.Y__gate ,
  output [  0:0] \__mp_output363.A__gate ,
  output [  0:0] \__mp_output363.Y__gate ,
  output [  0:0] \__mp_output364.A__gate ,
  output [  0:0] \__mp_output364.Y__gate ,
  output [  0:0] \__mp_output365.A__gate ,
  output [  0:0] \__mp_output365.Y__gate ,
  output [  0:0] \__mp_output366.A__gate ,
  output [  0:0] \__mp_output366.Y__gate ,
  output [  0:0] \__mp_output367.A__gate ,
  output [  0:0] \__mp_output367.Y__gate ,
  output [  0:0] \__mp_output368.A__gate ,
  output [  0:0] \__mp_output368.Y__gate ,
  output [  0:0] \__mp_output369.A__gate ,
  output [  0:0] \__mp_output369.Y__gate ,
  output [  0:0] \__mp_output370.A__gate ,
  output [  0:0] \__mp_output370.Y__gate ,
  output [  0:0] \__mp_output371.A__gate ,
  output [  0:0] \__mp_output371.Y__gate ,
  output [  0:0] \__mp_output372.A__gate ,
  output [  0:0] \__mp_output372.Y__gate ,
  output [  0:0] \__mp_output373.A__gate ,
  output [  0:0] \__mp_output373.Y__gate ,
  output [  0:0] \__mp_output374.A__gate ,
  output [  0:0] \__mp_output374.Y__gate ,
  output [  0:0] \__mp_output375.A__gate ,
  output [  0:0] \__mp_output375.Y__gate ,
  output [  0:0] \__mp_output376.A__gate ,
  output [  0:0] \__mp_output376.Y__gate ,
  output [  0:0] \__mp_output377.A__gate ,
  output [  0:0] \__mp_output377.Y__gate ,
  output [  0:0] \__mp_output378.A__gate ,
  output [  0:0] \__mp_output378.Y__gate ,
  output [  0:0] \__mp_output379.A__gate ,
  output [  0:0] \__mp_output379.Y__gate ,
  output [  0:0] \__mp_output380.A__gate ,
  output [  0:0] \__mp_output380.Y__gate ,
  output [  0:0] \__mp_output381.A__gate ,
  output [  0:0] \__mp_output381.Y__gate ,
  output [  0:0] \__mp_output382.A__gate ,
  output [  0:0] \__mp_output382.Y__gate ,
  output [  0:0] \__mp_output383.A__gate ,
  output [  0:0] \__mp_output383.Y__gate ,
  output [  0:0] \__mp_output384.A__gate ,
  output [  0:0] \__mp_output384.Y__gate ,
  output [  0:0] \__mp_output385.A__gate ,
  output [  0:0] \__mp_output385.Y__gate ,
  output [  0:0] \__mp_output386.A__gate ,
  output [  0:0] \__mp_output386.Y__gate ,
  output [  0:0] \__mp_output387.A__gate ,
  output [  0:0] \__mp_output387.Y__gate ,
  output [  0:0] \__mp_sa00_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa00_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa00_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa00_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa00_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa00_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa00_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa00_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa01_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa02_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa03_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa10_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa11_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa12_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa13_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa20_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa21_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa22_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa23_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa30_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa31_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa32_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_sa33_sr[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[0]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[100]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[101]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[102]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[103]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[104]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[105]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[106]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[107]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[108]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[109]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[10]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[110]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[111]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[112]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[113]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[114]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[115]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[116]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[117]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[118]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[119]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[11]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[120]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[121]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[122]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[123]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[124]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[125]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[126]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[127]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[12]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[13]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[14]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[15]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[16]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[17]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[18]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[19]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[1]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[20]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[21]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[22]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[23]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[24]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[25]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[26]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[27]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[28]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[29]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[2]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[30]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[31]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[32]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[33]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[34]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[35]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[36]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[37]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[38]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[39]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[3]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[40]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[41]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[42]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[43]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[44]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[45]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[46]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[47]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[48]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[49]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[4]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[50]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[51]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[52]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[53]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[54]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[55]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[56]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[57]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[58]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[59]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[5]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[60]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[61]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[62]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[63]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[64]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[65]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[66]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[67]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[68]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[69]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[6]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[70]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[71]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[72]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[73]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[74]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[75]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[76]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[77]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[78]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[79]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[7]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[80]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[81]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[82]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[83]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[84]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[85]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[86]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[87]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[88]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[89]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[8]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[90]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[91]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[92]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[93]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[94]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[95]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[96]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[97]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[98]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[99]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_in_r[9]$_DFFE_PP_.CLK__gate ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.QN__gate ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gate ,
  output [  0:0] \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u0.d[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u1.d[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u2.d[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.u3.d[7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][10]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][11]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][12]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][13]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][14]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][15]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][16]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][17]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][18]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][19]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][20]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][21]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][22]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][23]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][24]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][25]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][26]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][27]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][28]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][29]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][30]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][31]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][8]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[0][9]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][10]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][11]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][12]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][13]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][14]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][15]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][16]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][17]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][18]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][19]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][20]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][21]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][22]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][23]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][24]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][25]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][26]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][27]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][28]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][29]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][30]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][31]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][8]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[1][9]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][10]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][11]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][12]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][13]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][14]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][15]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][16]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][17]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][18]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][19]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][20]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][21]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][22]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][23]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][24]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][25]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][26]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][27]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][28]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][29]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][30]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][31]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][8]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[2][9]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][0]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][10]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][11]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][12]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][13]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][14]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][15]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][16]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][17]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][18]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][19]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][1]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][20]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][21]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][22]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][23]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][24]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][25]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][26]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][27]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][28]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][29]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][2]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][30]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][31]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][3]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][4]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][5]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][6]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][7]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][8]$_DFF_P_.CLK__gate ,
  output [  0:0] \__mp_u0.w[3][9]$_DFF_P_.CLK__gate ,
  output [  0:0] \__po_done__gold ,
  output [127:0] \__po_text_out__gold ,
  output [  0:0] \__po_done__gate ,
  output [127:0] \__po_text_out__gate
);
  \gold.aes_cipher_top gold (
    .\__pi_clk (\__pi_clk ),
    .\__pi_key (\__pi_key ),
    .\__pi_ld (\__pi_ld ),
    .\__pi_rst (\__pi_rst ),
    .\__pi_text_in (\__pi_text_in ),
`ifdef DIRECT_CROSS_POINTS
`else
`endif
    .\__mp_clkbuf_0_clk.A (\__mp_clkbuf_0_clk.A__gold ),
    .\__mp_clkbuf_0_clk.Y (\__mp_clkbuf_0_clk.Y__gold ),
    .\__mp_clkbuf_2_0_0_clk.A (\__mp_clkbuf_2_0_0_clk.A__gold ),
    .\__mp_clkbuf_2_0_0_clk.Y (\__mp_clkbuf_2_0_0_clk.Y__gold ),
    .\__mp_clkbuf_2_1_0_clk.A (\__mp_clkbuf_2_1_0_clk.A__gold ),
    .\__mp_clkbuf_2_1_0_clk.Y (\__mp_clkbuf_2_1_0_clk.Y__gold ),
    .\__mp_clkbuf_2_2_0_clk.A (\__mp_clkbuf_2_2_0_clk.A__gold ),
    .\__mp_clkbuf_2_2_0_clk.Y (\__mp_clkbuf_2_2_0_clk.Y__gold ),
    .\__mp_clkbuf_2_3_0_clk.A (\__mp_clkbuf_2_3_0_clk.A__gold ),
    .\__mp_clkbuf_2_3_0_clk.Y (\__mp_clkbuf_2_3_0_clk.Y__gold ),
    .\__mp_clkbuf_leaf_0_clk.A (\__mp_clkbuf_leaf_0_clk.A__gold ),
    .\__mp_clkbuf_leaf_0_clk.Y (\__mp_clkbuf_leaf_0_clk.Y__gold ),
    .\__mp_clkbuf_leaf_10_clk.A (\__mp_clkbuf_leaf_10_clk.A__gold ),
    .\__mp_clkbuf_leaf_10_clk.Y (\__mp_clkbuf_leaf_10_clk.Y__gold ),
    .\__mp_clkbuf_leaf_11_clk.A (\__mp_clkbuf_leaf_11_clk.A__gold ),
    .\__mp_clkbuf_leaf_11_clk.Y (\__mp_clkbuf_leaf_11_clk.Y__gold ),
    .\__mp_clkbuf_leaf_12_clk.A (\__mp_clkbuf_leaf_12_clk.A__gold ),
    .\__mp_clkbuf_leaf_12_clk.Y (\__mp_clkbuf_leaf_12_clk.Y__gold ),
    .\__mp_clkbuf_leaf_13_clk.A (\__mp_clkbuf_leaf_13_clk.A__gold ),
    .\__mp_clkbuf_leaf_13_clk.Y (\__mp_clkbuf_leaf_13_clk.Y__gold ),
    .\__mp_clkbuf_leaf_14_clk.A (\__mp_clkbuf_leaf_14_clk.A__gold ),
    .\__mp_clkbuf_leaf_14_clk.Y (\__mp_clkbuf_leaf_14_clk.Y__gold ),
    .\__mp_clkbuf_leaf_15_clk.A (\__mp_clkbuf_leaf_15_clk.A__gold ),
    .\__mp_clkbuf_leaf_15_clk.Y (\__mp_clkbuf_leaf_15_clk.Y__gold ),
    .\__mp_clkbuf_leaf_16_clk.A (\__mp_clkbuf_leaf_16_clk.A__gold ),
    .\__mp_clkbuf_leaf_16_clk.Y (\__mp_clkbuf_leaf_16_clk.Y__gold ),
    .\__mp_clkbuf_leaf_17_clk.A (\__mp_clkbuf_leaf_17_clk.A__gold ),
    .\__mp_clkbuf_leaf_17_clk.Y (\__mp_clkbuf_leaf_17_clk.Y__gold ),
    .\__mp_clkbuf_leaf_18_clk.A (\__mp_clkbuf_leaf_18_clk.A__gold ),
    .\__mp_clkbuf_leaf_18_clk.Y (\__mp_clkbuf_leaf_18_clk.Y__gold ),
    .\__mp_clkbuf_leaf_19_clk.A (\__mp_clkbuf_leaf_19_clk.A__gold ),
    .\__mp_clkbuf_leaf_19_clk.Y (\__mp_clkbuf_leaf_19_clk.Y__gold ),
    .\__mp_clkbuf_leaf_1_clk.A (\__mp_clkbuf_leaf_1_clk.A__gold ),
    .\__mp_clkbuf_leaf_1_clk.Y (\__mp_clkbuf_leaf_1_clk.Y__gold ),
    .\__mp_clkbuf_leaf_20_clk.A (\__mp_clkbuf_leaf_20_clk.A__gold ),
    .\__mp_clkbuf_leaf_20_clk.Y (\__mp_clkbuf_leaf_20_clk.Y__gold ),
    .\__mp_clkbuf_leaf_21_clk.A (\__mp_clkbuf_leaf_21_clk.A__gold ),
    .\__mp_clkbuf_leaf_21_clk.Y (\__mp_clkbuf_leaf_21_clk.Y__gold ),
    .\__mp_clkbuf_leaf_22_clk.A (\__mp_clkbuf_leaf_22_clk.A__gold ),
    .\__mp_clkbuf_leaf_22_clk.Y (\__mp_clkbuf_leaf_22_clk.Y__gold ),
    .\__mp_clkbuf_leaf_23_clk.A (\__mp_clkbuf_leaf_23_clk.A__gold ),
    .\__mp_clkbuf_leaf_23_clk.Y (\__mp_clkbuf_leaf_23_clk.Y__gold ),
    .\__mp_clkbuf_leaf_24_clk.A (\__mp_clkbuf_leaf_24_clk.A__gold ),
    .\__mp_clkbuf_leaf_24_clk.Y (\__mp_clkbuf_leaf_24_clk.Y__gold ),
    .\__mp_clkbuf_leaf_25_clk.A (\__mp_clkbuf_leaf_25_clk.A__gold ),
    .\__mp_clkbuf_leaf_25_clk.Y (\__mp_clkbuf_leaf_25_clk.Y__gold ),
    .\__mp_clkbuf_leaf_26_clk.A (\__mp_clkbuf_leaf_26_clk.A__gold ),
    .\__mp_clkbuf_leaf_26_clk.Y (\__mp_clkbuf_leaf_26_clk.Y__gold ),
    .\__mp_clkbuf_leaf_27_clk.A (\__mp_clkbuf_leaf_27_clk.A__gold ),
    .\__mp_clkbuf_leaf_27_clk.Y (\__mp_clkbuf_leaf_27_clk.Y__gold ),
    .\__mp_clkbuf_leaf_28_clk.A (\__mp_clkbuf_leaf_28_clk.A__gold ),
    .\__mp_clkbuf_leaf_28_clk.Y (\__mp_clkbuf_leaf_28_clk.Y__gold ),
    .\__mp_clkbuf_leaf_29_clk.A (\__mp_clkbuf_leaf_29_clk.A__gold ),
    .\__mp_clkbuf_leaf_29_clk.Y (\__mp_clkbuf_leaf_29_clk.Y__gold ),
    .\__mp_clkbuf_leaf_2_clk.A (\__mp_clkbuf_leaf_2_clk.A__gold ),
    .\__mp_clkbuf_leaf_2_clk.Y (\__mp_clkbuf_leaf_2_clk.Y__gold ),
    .\__mp_clkbuf_leaf_30_clk.A (\__mp_clkbuf_leaf_30_clk.A__gold ),
    .\__mp_clkbuf_leaf_30_clk.Y (\__mp_clkbuf_leaf_30_clk.Y__gold ),
    .\__mp_clkbuf_leaf_31_clk.A (\__mp_clkbuf_leaf_31_clk.A__gold ),
    .\__mp_clkbuf_leaf_31_clk.Y (\__mp_clkbuf_leaf_31_clk.Y__gold ),
    .\__mp_clkbuf_leaf_32_clk.A (\__mp_clkbuf_leaf_32_clk.A__gold ),
    .\__mp_clkbuf_leaf_32_clk.Y (\__mp_clkbuf_leaf_32_clk.Y__gold ),
    .\__mp_clkbuf_leaf_33_clk.A (\__mp_clkbuf_leaf_33_clk.A__gold ),
    .\__mp_clkbuf_leaf_33_clk.Y (\__mp_clkbuf_leaf_33_clk.Y__gold ),
    .\__mp_clkbuf_leaf_3_clk.A (\__mp_clkbuf_leaf_3_clk.A__gold ),
    .\__mp_clkbuf_leaf_3_clk.Y (\__mp_clkbuf_leaf_3_clk.Y__gold ),
    .\__mp_clkbuf_leaf_4_clk.A (\__mp_clkbuf_leaf_4_clk.A__gold ),
    .\__mp_clkbuf_leaf_4_clk.Y (\__mp_clkbuf_leaf_4_clk.Y__gold ),
    .\__mp_clkbuf_leaf_5_clk.A (\__mp_clkbuf_leaf_5_clk.A__gold ),
    .\__mp_clkbuf_leaf_5_clk.Y (\__mp_clkbuf_leaf_5_clk.Y__gold ),
    .\__mp_clkbuf_leaf_6_clk.A (\__mp_clkbuf_leaf_6_clk.A__gold ),
    .\__mp_clkbuf_leaf_6_clk.Y (\__mp_clkbuf_leaf_6_clk.Y__gold ),
    .\__mp_clkbuf_leaf_7_clk.A (\__mp_clkbuf_leaf_7_clk.A__gold ),
    .\__mp_clkbuf_leaf_7_clk.Y (\__mp_clkbuf_leaf_7_clk.Y__gold ),
    .\__mp_clkbuf_leaf_8_clk.A (\__mp_clkbuf_leaf_8_clk.A__gold ),
    .\__mp_clkbuf_leaf_8_clk.Y (\__mp_clkbuf_leaf_8_clk.Y__gold ),
    .\__mp_clkbuf_leaf_9_clk.A (\__mp_clkbuf_leaf_9_clk.A__gold ),
    .\__mp_clkbuf_leaf_9_clk.Y (\__mp_clkbuf_leaf_9_clk.Y__gold ),
    .\__mp_clkload0.A (\__mp_clkload0.A__gold ),
    .\__mp_clkload0.Y (\__mp_clkload0.Y__gold ),
    .\__mp_clkload1.A (\__mp_clkload1.A__gold ),
    .\__mp_clkload10.A (\__mp_clkload10.A__gold ),
    .\__mp_clkload11.A (\__mp_clkload11.A__gold ),
    .\__mp_clkload12.A (\__mp_clkload12.A__gold ),
    .\__mp_clkload13.A (\__mp_clkload13.A__gold ),
    .\__mp_clkload14.A (\__mp_clkload14.A__gold ),
    .\__mp_clkload15.A (\__mp_clkload15.A__gold ),
    .\__mp_clkload16.A (\__mp_clkload16.A__gold ),
    .\__mp_clkload17.A (\__mp_clkload17.A__gold ),
    .\__mp_clkload18.A (\__mp_clkload18.A__gold ),
    .\__mp_clkload18.Y (\__mp_clkload18.Y__gold ),
    .\__mp_clkload19.A (\__mp_clkload19.A__gold ),
    .\__mp_clkload2.A (\__mp_clkload2.A__gold ),
    .\__mp_clkload20.A (\__mp_clkload20.A__gold ),
    .\__mp_clkload21.A (\__mp_clkload21.A__gold ),
    .\__mp_clkload22.A (\__mp_clkload22.A__gold ),
    .\__mp_clkload23.A (\__mp_clkload23.A__gold ),
    .\__mp_clkload24.A (\__mp_clkload24.A__gold ),
    .\__mp_clkload25.A (\__mp_clkload25.A__gold ),
    .\__mp_clkload26.A (\__mp_clkload26.A__gold ),
    .\__mp_clkload27.A (\__mp_clkload27.A__gold ),
    .\__mp_clkload28.A (\__mp_clkload28.A__gold ),
    .\__mp_clkload29.A (\__mp_clkload29.A__gold ),
    .\__mp_clkload3.A (\__mp_clkload3.A__gold ),
    .\__mp_clkload30.A (\__mp_clkload30.A__gold ),
    .\__mp_clkload31.A (\__mp_clkload31.A__gold ),
    .\__mp_clkload31.Y (\__mp_clkload31.Y__gold ),
    .\__mp_clkload32.A (\__mp_clkload32.A__gold ),
    .\__mp_clkload4.A (\__mp_clkload4.A__gold ),
    .\__mp_clkload5.A (\__mp_clkload5.A__gold ),
    .\__mp_clkload6.A (\__mp_clkload6.A__gold ),
    .\__mp_clkload7.A (\__mp_clkload7.A__gold ),
    .\__mp_clkload8.A (\__mp_clkload8.A__gold ),
    .\__mp_clkload9.A (\__mp_clkload9.A__gold ),
    .\__mp_clknet_0_clk (\__mp_clknet_0_clk__gold ),
    .\__mp_clknet_2_0_0_clk (\__mp_clknet_2_0_0_clk__gold ),
    .\__mp_clknet_2_1_0_clk (\__mp_clknet_2_1_0_clk__gold ),
    .\__mp_clknet_2_2_0_clk (\__mp_clknet_2_2_0_clk__gold ),
    .\__mp_clknet_2_3_0_clk (\__mp_clknet_2_3_0_clk__gold ),
    .\__mp_clknet_leaf_0_clk (\__mp_clknet_leaf_0_clk__gold ),
    .\__mp_clknet_leaf_10_clk (\__mp_clknet_leaf_10_clk__gold ),
    .\__mp_clknet_leaf_11_clk (\__mp_clknet_leaf_11_clk__gold ),
    .\__mp_clknet_leaf_12_clk (\__mp_clknet_leaf_12_clk__gold ),
    .\__mp_clknet_leaf_13_clk (\__mp_clknet_leaf_13_clk__gold ),
    .\__mp_clknet_leaf_14_clk (\__mp_clknet_leaf_14_clk__gold ),
    .\__mp_clknet_leaf_15_clk (\__mp_clknet_leaf_15_clk__gold ),
    .\__mp_clknet_leaf_16_clk (\__mp_clknet_leaf_16_clk__gold ),
    .\__mp_clknet_leaf_17_clk (\__mp_clknet_leaf_17_clk__gold ),
    .\__mp_clknet_leaf_18_clk (\__mp_clknet_leaf_18_clk__gold ),
    .\__mp_clknet_leaf_19_clk (\__mp_clknet_leaf_19_clk__gold ),
    .\__mp_clknet_leaf_1_clk (\__mp_clknet_leaf_1_clk__gold ),
    .\__mp_clknet_leaf_20_clk (\__mp_clknet_leaf_20_clk__gold ),
    .\__mp_clknet_leaf_21_clk (\__mp_clknet_leaf_21_clk__gold ),
    .\__mp_clknet_leaf_22_clk (\__mp_clknet_leaf_22_clk__gold ),
    .\__mp_clknet_leaf_23_clk (\__mp_clknet_leaf_23_clk__gold ),
    .\__mp_clknet_leaf_24_clk (\__mp_clknet_leaf_24_clk__gold ),
    .\__mp_clknet_leaf_25_clk (\__mp_clknet_leaf_25_clk__gold ),
    .\__mp_clknet_leaf_26_clk (\__mp_clknet_leaf_26_clk__gold ),
    .\__mp_clknet_leaf_27_clk (\__mp_clknet_leaf_27_clk__gold ),
    .\__mp_clknet_leaf_28_clk (\__mp_clknet_leaf_28_clk__gold ),
    .\__mp_clknet_leaf_29_clk (\__mp_clknet_leaf_29_clk__gold ),
    .\__mp_clknet_leaf_2_clk (\__mp_clknet_leaf_2_clk__gold ),
    .\__mp_clknet_leaf_30_clk (\__mp_clknet_leaf_30_clk__gold ),
    .\__mp_clknet_leaf_31_clk (\__mp_clknet_leaf_31_clk__gold ),
    .\__mp_clknet_leaf_32_clk (\__mp_clknet_leaf_32_clk__gold ),
    .\__mp_clknet_leaf_33_clk (\__mp_clknet_leaf_33_clk__gold ),
    .\__mp_clknet_leaf_3_clk (\__mp_clknet_leaf_3_clk__gold ),
    .\__mp_clknet_leaf_4_clk (\__mp_clknet_leaf_4_clk__gold ),
    .\__mp_clknet_leaf_5_clk (\__mp_clknet_leaf_5_clk__gold ),
    .\__mp_clknet_leaf_6_clk (\__mp_clknet_leaf_6_clk__gold ),
    .\__mp_clknet_leaf_7_clk (\__mp_clknet_leaf_7_clk__gold ),
    .\__mp_clknet_leaf_8_clk (\__mp_clknet_leaf_8_clk__gold ),
    .\__mp_clknet_leaf_9_clk (\__mp_clknet_leaf_9_clk__gold ),
    .\__mp_dcnt[0]$_SDFFE_PN0P_.CLK (\__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gold ),
    .\__mp_dcnt[1]$_SDFFE_PN0P_.CLK (\__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gold ),
    .\__mp_dcnt[2]$_SDFFE_PP0P_.CLK (\__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gold ),
    .\__mp_dcnt[3]$_SDFFE_PN0P_.CLK (\__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gold ),
    .\__mp_done$_DFF_P_.CLK (\__mp_done$_DFF_P_.CLK__gold ),
    .\__mp_done$_DFF_P_.QN (\__mp_done$_DFF_P_.QN__gold ),
    .\__mp_done$_DFF_P_.int_fwire_IQN (\__mp_done$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_input1.A (\__mp_input1.A__gold ),
    .\__mp_input1.Y (\__mp_input1.Y__gold ),
    .\__mp_input10.A (\__mp_input10.A__gold ),
    .\__mp_input10.Y (\__mp_input10.Y__gold ),
    .\__mp_input100.A (\__mp_input100.A__gold ),
    .\__mp_input100.Y (\__mp_input100.Y__gold ),
    .\__mp_input101.A (\__mp_input101.A__gold ),
    .\__mp_input101.Y (\__mp_input101.Y__gold ),
    .\__mp_input102.A (\__mp_input102.A__gold ),
    .\__mp_input102.Y (\__mp_input102.Y__gold ),
    .\__mp_input103.A (\__mp_input103.A__gold ),
    .\__mp_input103.Y (\__mp_input103.Y__gold ),
    .\__mp_input104.A (\__mp_input104.A__gold ),
    .\__mp_input104.Y (\__mp_input104.Y__gold ),
    .\__mp_input105.A (\__mp_input105.A__gold ),
    .\__mp_input105.Y (\__mp_input105.Y__gold ),
    .\__mp_input106.A (\__mp_input106.A__gold ),
    .\__mp_input106.Y (\__mp_input106.Y__gold ),
    .\__mp_input107.A (\__mp_input107.A__gold ),
    .\__mp_input107.Y (\__mp_input107.Y__gold ),
    .\__mp_input108.A (\__mp_input108.A__gold ),
    .\__mp_input108.Y (\__mp_input108.Y__gold ),
    .\__mp_input109.A (\__mp_input109.A__gold ),
    .\__mp_input109.Y (\__mp_input109.Y__gold ),
    .\__mp_input11.A (\__mp_input11.A__gold ),
    .\__mp_input11.Y (\__mp_input11.Y__gold ),
    .\__mp_input110.A (\__mp_input110.A__gold ),
    .\__mp_input110.Y (\__mp_input110.Y__gold ),
    .\__mp_input111.A (\__mp_input111.A__gold ),
    .\__mp_input111.Y (\__mp_input111.Y__gold ),
    .\__mp_input112.A (\__mp_input112.A__gold ),
    .\__mp_input112.Y (\__mp_input112.Y__gold ),
    .\__mp_input113.A (\__mp_input113.A__gold ),
    .\__mp_input113.Y (\__mp_input113.Y__gold ),
    .\__mp_input114.A (\__mp_input114.A__gold ),
    .\__mp_input114.Y (\__mp_input114.Y__gold ),
    .\__mp_input115.A (\__mp_input115.A__gold ),
    .\__mp_input115.Y (\__mp_input115.Y__gold ),
    .\__mp_input116.A (\__mp_input116.A__gold ),
    .\__mp_input116.Y (\__mp_input116.Y__gold ),
    .\__mp_input117.A (\__mp_input117.A__gold ),
    .\__mp_input117.Y (\__mp_input117.Y__gold ),
    .\__mp_input118.A (\__mp_input118.A__gold ),
    .\__mp_input118.Y (\__mp_input118.Y__gold ),
    .\__mp_input119.A (\__mp_input119.A__gold ),
    .\__mp_input119.Y (\__mp_input119.Y__gold ),
    .\__mp_input12.A (\__mp_input12.A__gold ),
    .\__mp_input12.Y (\__mp_input12.Y__gold ),
    .\__mp_input120.A (\__mp_input120.A__gold ),
    .\__mp_input120.Y (\__mp_input120.Y__gold ),
    .\__mp_input121.A (\__mp_input121.A__gold ),
    .\__mp_input121.Y (\__mp_input121.Y__gold ),
    .\__mp_input122.A (\__mp_input122.A__gold ),
    .\__mp_input122.Y (\__mp_input122.Y__gold ),
    .\__mp_input123.A (\__mp_input123.A__gold ),
    .\__mp_input123.Y (\__mp_input123.Y__gold ),
    .\__mp_input124.A (\__mp_input124.A__gold ),
    .\__mp_input124.Y (\__mp_input124.Y__gold ),
    .\__mp_input125.A (\__mp_input125.A__gold ),
    .\__mp_input125.Y (\__mp_input125.Y__gold ),
    .\__mp_input126.A (\__mp_input126.A__gold ),
    .\__mp_input126.Y (\__mp_input126.Y__gold ),
    .\__mp_input127.A (\__mp_input127.A__gold ),
    .\__mp_input127.Y (\__mp_input127.Y__gold ),
    .\__mp_input128.A (\__mp_input128.A__gold ),
    .\__mp_input128.Y (\__mp_input128.Y__gold ),
    .\__mp_input129.A (\__mp_input129.A__gold ),
    .\__mp_input129.Y (\__mp_input129.Y__gold ),
    .\__mp_input13.A (\__mp_input13.A__gold ),
    .\__mp_input13.Y (\__mp_input13.Y__gold ),
    .\__mp_input130.A (\__mp_input130.A__gold ),
    .\__mp_input130.Y (\__mp_input130.Y__gold ),
    .\__mp_input131.A (\__mp_input131.A__gold ),
    .\__mp_input131.Y (\__mp_input131.Y__gold ),
    .\__mp_input132.A (\__mp_input132.A__gold ),
    .\__mp_input132.Y (\__mp_input132.Y__gold ),
    .\__mp_input133.A (\__mp_input133.A__gold ),
    .\__mp_input133.Y (\__mp_input133.Y__gold ),
    .\__mp_input134.A (\__mp_input134.A__gold ),
    .\__mp_input134.Y (\__mp_input134.Y__gold ),
    .\__mp_input135.A (\__mp_input135.A__gold ),
    .\__mp_input135.Y (\__mp_input135.Y__gold ),
    .\__mp_input136.A (\__mp_input136.A__gold ),
    .\__mp_input136.Y (\__mp_input136.Y__gold ),
    .\__mp_input137.A (\__mp_input137.A__gold ),
    .\__mp_input137.Y (\__mp_input137.Y__gold ),
    .\__mp_input138.A (\__mp_input138.A__gold ),
    .\__mp_input138.Y (\__mp_input138.Y__gold ),
    .\__mp_input139.A (\__mp_input139.A__gold ),
    .\__mp_input139.Y (\__mp_input139.Y__gold ),
    .\__mp_input14.A (\__mp_input14.A__gold ),
    .\__mp_input14.Y (\__mp_input14.Y__gold ),
    .\__mp_input140.A (\__mp_input140.A__gold ),
    .\__mp_input140.Y (\__mp_input140.Y__gold ),
    .\__mp_input141.A (\__mp_input141.A__gold ),
    .\__mp_input141.Y (\__mp_input141.Y__gold ),
    .\__mp_input142.A (\__mp_input142.A__gold ),
    .\__mp_input142.Y (\__mp_input142.Y__gold ),
    .\__mp_input143.A (\__mp_input143.A__gold ),
    .\__mp_input143.Y (\__mp_input143.Y__gold ),
    .\__mp_input144.A (\__mp_input144.A__gold ),
    .\__mp_input144.Y (\__mp_input144.Y__gold ),
    .\__mp_input145.A (\__mp_input145.A__gold ),
    .\__mp_input145.Y (\__mp_input145.Y__gold ),
    .\__mp_input146.A (\__mp_input146.A__gold ),
    .\__mp_input146.Y (\__mp_input146.Y__gold ),
    .\__mp_input147.A (\__mp_input147.A__gold ),
    .\__mp_input147.Y (\__mp_input147.Y__gold ),
    .\__mp_input148.A (\__mp_input148.A__gold ),
    .\__mp_input148.Y (\__mp_input148.Y__gold ),
    .\__mp_input149.A (\__mp_input149.A__gold ),
    .\__mp_input149.Y (\__mp_input149.Y__gold ),
    .\__mp_input15.A (\__mp_input15.A__gold ),
    .\__mp_input15.Y (\__mp_input15.Y__gold ),
    .\__mp_input150.A (\__mp_input150.A__gold ),
    .\__mp_input150.Y (\__mp_input150.Y__gold ),
    .\__mp_input151.A (\__mp_input151.A__gold ),
    .\__mp_input151.Y (\__mp_input151.Y__gold ),
    .\__mp_input152.A (\__mp_input152.A__gold ),
    .\__mp_input152.Y (\__mp_input152.Y__gold ),
    .\__mp_input153.A (\__mp_input153.A__gold ),
    .\__mp_input153.Y (\__mp_input153.Y__gold ),
    .\__mp_input154.A (\__mp_input154.A__gold ),
    .\__mp_input154.Y (\__mp_input154.Y__gold ),
    .\__mp_input155.A (\__mp_input155.A__gold ),
    .\__mp_input155.Y (\__mp_input155.Y__gold ),
    .\__mp_input156.A (\__mp_input156.A__gold ),
    .\__mp_input156.Y (\__mp_input156.Y__gold ),
    .\__mp_input157.A (\__mp_input157.A__gold ),
    .\__mp_input157.Y (\__mp_input157.Y__gold ),
    .\__mp_input158.A (\__mp_input158.A__gold ),
    .\__mp_input158.Y (\__mp_input158.Y__gold ),
    .\__mp_input159.A (\__mp_input159.A__gold ),
    .\__mp_input159.Y (\__mp_input159.Y__gold ),
    .\__mp_input16.A (\__mp_input16.A__gold ),
    .\__mp_input16.Y (\__mp_input16.Y__gold ),
    .\__mp_input160.A (\__mp_input160.A__gold ),
    .\__mp_input160.Y (\__mp_input160.Y__gold ),
    .\__mp_input161.A (\__mp_input161.A__gold ),
    .\__mp_input161.Y (\__mp_input161.Y__gold ),
    .\__mp_input162.A (\__mp_input162.A__gold ),
    .\__mp_input162.Y (\__mp_input162.Y__gold ),
    .\__mp_input163.A (\__mp_input163.A__gold ),
    .\__mp_input163.Y (\__mp_input163.Y__gold ),
    .\__mp_input164.A (\__mp_input164.A__gold ),
    .\__mp_input164.Y (\__mp_input164.Y__gold ),
    .\__mp_input165.A (\__mp_input165.A__gold ),
    .\__mp_input165.Y (\__mp_input165.Y__gold ),
    .\__mp_input166.A (\__mp_input166.A__gold ),
    .\__mp_input166.Y (\__mp_input166.Y__gold ),
    .\__mp_input167.A (\__mp_input167.A__gold ),
    .\__mp_input167.Y (\__mp_input167.Y__gold ),
    .\__mp_input168.A (\__mp_input168.A__gold ),
    .\__mp_input168.Y (\__mp_input168.Y__gold ),
    .\__mp_input169.A (\__mp_input169.A__gold ),
    .\__mp_input169.Y (\__mp_input169.Y__gold ),
    .\__mp_input17.A (\__mp_input17.A__gold ),
    .\__mp_input17.Y (\__mp_input17.Y__gold ),
    .\__mp_input170.A (\__mp_input170.A__gold ),
    .\__mp_input170.Y (\__mp_input170.Y__gold ),
    .\__mp_input171.A (\__mp_input171.A__gold ),
    .\__mp_input171.Y (\__mp_input171.Y__gold ),
    .\__mp_input172.A (\__mp_input172.A__gold ),
    .\__mp_input172.Y (\__mp_input172.Y__gold ),
    .\__mp_input173.A (\__mp_input173.A__gold ),
    .\__mp_input173.Y (\__mp_input173.Y__gold ),
    .\__mp_input174.A (\__mp_input174.A__gold ),
    .\__mp_input174.Y (\__mp_input174.Y__gold ),
    .\__mp_input175.A (\__mp_input175.A__gold ),
    .\__mp_input175.Y (\__mp_input175.Y__gold ),
    .\__mp_input176.A (\__mp_input176.A__gold ),
    .\__mp_input176.Y (\__mp_input176.Y__gold ),
    .\__mp_input177.A (\__mp_input177.A__gold ),
    .\__mp_input177.Y (\__mp_input177.Y__gold ),
    .\__mp_input178.A (\__mp_input178.A__gold ),
    .\__mp_input178.Y (\__mp_input178.Y__gold ),
    .\__mp_input179.A (\__mp_input179.A__gold ),
    .\__mp_input179.Y (\__mp_input179.Y__gold ),
    .\__mp_input18.A (\__mp_input18.A__gold ),
    .\__mp_input18.Y (\__mp_input18.Y__gold ),
    .\__mp_input180.A (\__mp_input180.A__gold ),
    .\__mp_input180.Y (\__mp_input180.Y__gold ),
    .\__mp_input181.A (\__mp_input181.A__gold ),
    .\__mp_input181.Y (\__mp_input181.Y__gold ),
    .\__mp_input182.A (\__mp_input182.A__gold ),
    .\__mp_input182.Y (\__mp_input182.Y__gold ),
    .\__mp_input183.A (\__mp_input183.A__gold ),
    .\__mp_input183.Y (\__mp_input183.Y__gold ),
    .\__mp_input184.A (\__mp_input184.A__gold ),
    .\__mp_input184.Y (\__mp_input184.Y__gold ),
    .\__mp_input185.A (\__mp_input185.A__gold ),
    .\__mp_input185.Y (\__mp_input185.Y__gold ),
    .\__mp_input186.A (\__mp_input186.A__gold ),
    .\__mp_input186.Y (\__mp_input186.Y__gold ),
    .\__mp_input187.A (\__mp_input187.A__gold ),
    .\__mp_input187.Y (\__mp_input187.Y__gold ),
    .\__mp_input188.A (\__mp_input188.A__gold ),
    .\__mp_input188.Y (\__mp_input188.Y__gold ),
    .\__mp_input189.A (\__mp_input189.A__gold ),
    .\__mp_input189.Y (\__mp_input189.Y__gold ),
    .\__mp_input19.A (\__mp_input19.A__gold ),
    .\__mp_input19.Y (\__mp_input19.Y__gold ),
    .\__mp_input190.A (\__mp_input190.A__gold ),
    .\__mp_input190.Y (\__mp_input190.Y__gold ),
    .\__mp_input191.A (\__mp_input191.A__gold ),
    .\__mp_input191.Y (\__mp_input191.Y__gold ),
    .\__mp_input192.A (\__mp_input192.A__gold ),
    .\__mp_input192.Y (\__mp_input192.Y__gold ),
    .\__mp_input193.A (\__mp_input193.A__gold ),
    .\__mp_input193.Y (\__mp_input193.Y__gold ),
    .\__mp_input194.A (\__mp_input194.A__gold ),
    .\__mp_input194.Y (\__mp_input194.Y__gold ),
    .\__mp_input195.A (\__mp_input195.A__gold ),
    .\__mp_input195.Y (\__mp_input195.Y__gold ),
    .\__mp_input196.A (\__mp_input196.A__gold ),
    .\__mp_input196.Y (\__mp_input196.Y__gold ),
    .\__mp_input197.A (\__mp_input197.A__gold ),
    .\__mp_input197.Y (\__mp_input197.Y__gold ),
    .\__mp_input198.A (\__mp_input198.A__gold ),
    .\__mp_input198.Y (\__mp_input198.Y__gold ),
    .\__mp_input199.A (\__mp_input199.A__gold ),
    .\__mp_input199.Y (\__mp_input199.Y__gold ),
    .\__mp_input2.A (\__mp_input2.A__gold ),
    .\__mp_input2.Y (\__mp_input2.Y__gold ),
    .\__mp_input20.A (\__mp_input20.A__gold ),
    .\__mp_input20.Y (\__mp_input20.Y__gold ),
    .\__mp_input200.A (\__mp_input200.A__gold ),
    .\__mp_input200.Y (\__mp_input200.Y__gold ),
    .\__mp_input201.A (\__mp_input201.A__gold ),
    .\__mp_input201.Y (\__mp_input201.Y__gold ),
    .\__mp_input202.A (\__mp_input202.A__gold ),
    .\__mp_input202.Y (\__mp_input202.Y__gold ),
    .\__mp_input203.A (\__mp_input203.A__gold ),
    .\__mp_input203.Y (\__mp_input203.Y__gold ),
    .\__mp_input204.A (\__mp_input204.A__gold ),
    .\__mp_input204.Y (\__mp_input204.Y__gold ),
    .\__mp_input205.A (\__mp_input205.A__gold ),
    .\__mp_input205.Y (\__mp_input205.Y__gold ),
    .\__mp_input206.A (\__mp_input206.A__gold ),
    .\__mp_input206.Y (\__mp_input206.Y__gold ),
    .\__mp_input207.A (\__mp_input207.A__gold ),
    .\__mp_input207.Y (\__mp_input207.Y__gold ),
    .\__mp_input208.A (\__mp_input208.A__gold ),
    .\__mp_input208.Y (\__mp_input208.Y__gold ),
    .\__mp_input209.A (\__mp_input209.A__gold ),
    .\__mp_input209.Y (\__mp_input209.Y__gold ),
    .\__mp_input21.A (\__mp_input21.A__gold ),
    .\__mp_input21.Y (\__mp_input21.Y__gold ),
    .\__mp_input210.A (\__mp_input210.A__gold ),
    .\__mp_input210.Y (\__mp_input210.Y__gold ),
    .\__mp_input211.A (\__mp_input211.A__gold ),
    .\__mp_input211.Y (\__mp_input211.Y__gold ),
    .\__mp_input212.A (\__mp_input212.A__gold ),
    .\__mp_input212.Y (\__mp_input212.Y__gold ),
    .\__mp_input213.A (\__mp_input213.A__gold ),
    .\__mp_input213.Y (\__mp_input213.Y__gold ),
    .\__mp_input214.A (\__mp_input214.A__gold ),
    .\__mp_input214.Y (\__mp_input214.Y__gold ),
    .\__mp_input215.A (\__mp_input215.A__gold ),
    .\__mp_input215.Y (\__mp_input215.Y__gold ),
    .\__mp_input216.A (\__mp_input216.A__gold ),
    .\__mp_input216.Y (\__mp_input216.Y__gold ),
    .\__mp_input217.A (\__mp_input217.A__gold ),
    .\__mp_input217.Y (\__mp_input217.Y__gold ),
    .\__mp_input218.A (\__mp_input218.A__gold ),
    .\__mp_input218.Y (\__mp_input218.Y__gold ),
    .\__mp_input219.A (\__mp_input219.A__gold ),
    .\__mp_input219.Y (\__mp_input219.Y__gold ),
    .\__mp_input22.A (\__mp_input22.A__gold ),
    .\__mp_input22.Y (\__mp_input22.Y__gold ),
    .\__mp_input220.A (\__mp_input220.A__gold ),
    .\__mp_input220.Y (\__mp_input220.Y__gold ),
    .\__mp_input221.A (\__mp_input221.A__gold ),
    .\__mp_input221.Y (\__mp_input221.Y__gold ),
    .\__mp_input222.A (\__mp_input222.A__gold ),
    .\__mp_input222.Y (\__mp_input222.Y__gold ),
    .\__mp_input223.A (\__mp_input223.A__gold ),
    .\__mp_input223.Y (\__mp_input223.Y__gold ),
    .\__mp_input224.A (\__mp_input224.A__gold ),
    .\__mp_input224.Y (\__mp_input224.Y__gold ),
    .\__mp_input225.A (\__mp_input225.A__gold ),
    .\__mp_input225.Y (\__mp_input225.Y__gold ),
    .\__mp_input226.A (\__mp_input226.A__gold ),
    .\__mp_input226.Y (\__mp_input226.Y__gold ),
    .\__mp_input227.A (\__mp_input227.A__gold ),
    .\__mp_input227.Y (\__mp_input227.Y__gold ),
    .\__mp_input228.A (\__mp_input228.A__gold ),
    .\__mp_input228.Y (\__mp_input228.Y__gold ),
    .\__mp_input229.A (\__mp_input229.A__gold ),
    .\__mp_input229.Y (\__mp_input229.Y__gold ),
    .\__mp_input23.A (\__mp_input23.A__gold ),
    .\__mp_input23.Y (\__mp_input23.Y__gold ),
    .\__mp_input230.A (\__mp_input230.A__gold ),
    .\__mp_input230.Y (\__mp_input230.Y__gold ),
    .\__mp_input231.A (\__mp_input231.A__gold ),
    .\__mp_input231.Y (\__mp_input231.Y__gold ),
    .\__mp_input232.A (\__mp_input232.A__gold ),
    .\__mp_input232.Y (\__mp_input232.Y__gold ),
    .\__mp_input233.A (\__mp_input233.A__gold ),
    .\__mp_input233.Y (\__mp_input233.Y__gold ),
    .\__mp_input234.A (\__mp_input234.A__gold ),
    .\__mp_input234.Y (\__mp_input234.Y__gold ),
    .\__mp_input235.A (\__mp_input235.A__gold ),
    .\__mp_input235.Y (\__mp_input235.Y__gold ),
    .\__mp_input236.A (\__mp_input236.A__gold ),
    .\__mp_input236.Y (\__mp_input236.Y__gold ),
    .\__mp_input237.A (\__mp_input237.A__gold ),
    .\__mp_input237.Y (\__mp_input237.Y__gold ),
    .\__mp_input238.A (\__mp_input238.A__gold ),
    .\__mp_input238.Y (\__mp_input238.Y__gold ),
    .\__mp_input239.A (\__mp_input239.A__gold ),
    .\__mp_input239.Y (\__mp_input239.Y__gold ),
    .\__mp_input24.A (\__mp_input24.A__gold ),
    .\__mp_input24.Y (\__mp_input24.Y__gold ),
    .\__mp_input240.A (\__mp_input240.A__gold ),
    .\__mp_input240.Y (\__mp_input240.Y__gold ),
    .\__mp_input241.A (\__mp_input241.A__gold ),
    .\__mp_input241.Y (\__mp_input241.Y__gold ),
    .\__mp_input242.A (\__mp_input242.A__gold ),
    .\__mp_input242.Y (\__mp_input242.Y__gold ),
    .\__mp_input243.A (\__mp_input243.A__gold ),
    .\__mp_input243.Y (\__mp_input243.Y__gold ),
    .\__mp_input244.A (\__mp_input244.A__gold ),
    .\__mp_input244.Y (\__mp_input244.Y__gold ),
    .\__mp_input245.A (\__mp_input245.A__gold ),
    .\__mp_input245.Y (\__mp_input245.Y__gold ),
    .\__mp_input246.A (\__mp_input246.A__gold ),
    .\__mp_input246.Y (\__mp_input246.Y__gold ),
    .\__mp_input247.A (\__mp_input247.A__gold ),
    .\__mp_input247.Y (\__mp_input247.Y__gold ),
    .\__mp_input248.A (\__mp_input248.A__gold ),
    .\__mp_input248.Y (\__mp_input248.Y__gold ),
    .\__mp_input249.A (\__mp_input249.A__gold ),
    .\__mp_input249.Y (\__mp_input249.Y__gold ),
    .\__mp_input25.A (\__mp_input25.A__gold ),
    .\__mp_input25.Y (\__mp_input25.Y__gold ),
    .\__mp_input250.A (\__mp_input250.A__gold ),
    .\__mp_input250.Y (\__mp_input250.Y__gold ),
    .\__mp_input251.A (\__mp_input251.A__gold ),
    .\__mp_input251.Y (\__mp_input251.Y__gold ),
    .\__mp_input252.A (\__mp_input252.A__gold ),
    .\__mp_input252.Y (\__mp_input252.Y__gold ),
    .\__mp_input253.A (\__mp_input253.A__gold ),
    .\__mp_input253.Y (\__mp_input253.Y__gold ),
    .\__mp_input254.A (\__mp_input254.A__gold ),
    .\__mp_input254.Y (\__mp_input254.Y__gold ),
    .\__mp_input255.A (\__mp_input255.A__gold ),
    .\__mp_input255.Y (\__mp_input255.Y__gold ),
    .\__mp_input256.A (\__mp_input256.A__gold ),
    .\__mp_input256.Y (\__mp_input256.Y__gold ),
    .\__mp_input257.A (\__mp_input257.A__gold ),
    .\__mp_input257.Y (\__mp_input257.Y__gold ),
    .\__mp_input258.A (\__mp_input258.A__gold ),
    .\__mp_input258.Y (\__mp_input258.Y__gold ),
    .\__mp_input26.A (\__mp_input26.A__gold ),
    .\__mp_input26.Y (\__mp_input26.Y__gold ),
    .\__mp_input27.A (\__mp_input27.A__gold ),
    .\__mp_input27.Y (\__mp_input27.Y__gold ),
    .\__mp_input28.A (\__mp_input28.A__gold ),
    .\__mp_input28.Y (\__mp_input28.Y__gold ),
    .\__mp_input29.A (\__mp_input29.A__gold ),
    .\__mp_input29.Y (\__mp_input29.Y__gold ),
    .\__mp_input3.A (\__mp_input3.A__gold ),
    .\__mp_input3.Y (\__mp_input3.Y__gold ),
    .\__mp_input30.A (\__mp_input30.A__gold ),
    .\__mp_input30.Y (\__mp_input30.Y__gold ),
    .\__mp_input31.A (\__mp_input31.A__gold ),
    .\__mp_input31.Y (\__mp_input31.Y__gold ),
    .\__mp_input32.A (\__mp_input32.A__gold ),
    .\__mp_input32.Y (\__mp_input32.Y__gold ),
    .\__mp_input33.A (\__mp_input33.A__gold ),
    .\__mp_input33.Y (\__mp_input33.Y__gold ),
    .\__mp_input34.A (\__mp_input34.A__gold ),
    .\__mp_input34.Y (\__mp_input34.Y__gold ),
    .\__mp_input35.A (\__mp_input35.A__gold ),
    .\__mp_input35.Y (\__mp_input35.Y__gold ),
    .\__mp_input36.A (\__mp_input36.A__gold ),
    .\__mp_input36.Y (\__mp_input36.Y__gold ),
    .\__mp_input37.A (\__mp_input37.A__gold ),
    .\__mp_input37.Y (\__mp_input37.Y__gold ),
    .\__mp_input38.A (\__mp_input38.A__gold ),
    .\__mp_input38.Y (\__mp_input38.Y__gold ),
    .\__mp_input39.A (\__mp_input39.A__gold ),
    .\__mp_input39.Y (\__mp_input39.Y__gold ),
    .\__mp_input4.A (\__mp_input4.A__gold ),
    .\__mp_input4.Y (\__mp_input4.Y__gold ),
    .\__mp_input40.A (\__mp_input40.A__gold ),
    .\__mp_input40.Y (\__mp_input40.Y__gold ),
    .\__mp_input41.A (\__mp_input41.A__gold ),
    .\__mp_input41.Y (\__mp_input41.Y__gold ),
    .\__mp_input42.A (\__mp_input42.A__gold ),
    .\__mp_input42.Y (\__mp_input42.Y__gold ),
    .\__mp_input43.A (\__mp_input43.A__gold ),
    .\__mp_input43.Y (\__mp_input43.Y__gold ),
    .\__mp_input44.A (\__mp_input44.A__gold ),
    .\__mp_input44.Y (\__mp_input44.Y__gold ),
    .\__mp_input45.A (\__mp_input45.A__gold ),
    .\__mp_input45.Y (\__mp_input45.Y__gold ),
    .\__mp_input46.A (\__mp_input46.A__gold ),
    .\__mp_input46.Y (\__mp_input46.Y__gold ),
    .\__mp_input47.A (\__mp_input47.A__gold ),
    .\__mp_input47.Y (\__mp_input47.Y__gold ),
    .\__mp_input48.A (\__mp_input48.A__gold ),
    .\__mp_input48.Y (\__mp_input48.Y__gold ),
    .\__mp_input49.A (\__mp_input49.A__gold ),
    .\__mp_input49.Y (\__mp_input49.Y__gold ),
    .\__mp_input5.A (\__mp_input5.A__gold ),
    .\__mp_input5.Y (\__mp_input5.Y__gold ),
    .\__mp_input50.A (\__mp_input50.A__gold ),
    .\__mp_input50.Y (\__mp_input50.Y__gold ),
    .\__mp_input51.A (\__mp_input51.A__gold ),
    .\__mp_input51.Y (\__mp_input51.Y__gold ),
    .\__mp_input52.A (\__mp_input52.A__gold ),
    .\__mp_input52.Y (\__mp_input52.Y__gold ),
    .\__mp_input53.A (\__mp_input53.A__gold ),
    .\__mp_input53.Y (\__mp_input53.Y__gold ),
    .\__mp_input54.A (\__mp_input54.A__gold ),
    .\__mp_input54.Y (\__mp_input54.Y__gold ),
    .\__mp_input55.A (\__mp_input55.A__gold ),
    .\__mp_input55.Y (\__mp_input55.Y__gold ),
    .\__mp_input56.A (\__mp_input56.A__gold ),
    .\__mp_input56.Y (\__mp_input56.Y__gold ),
    .\__mp_input57.A (\__mp_input57.A__gold ),
    .\__mp_input57.Y (\__mp_input57.Y__gold ),
    .\__mp_input58.A (\__mp_input58.A__gold ),
    .\__mp_input58.Y (\__mp_input58.Y__gold ),
    .\__mp_input59.A (\__mp_input59.A__gold ),
    .\__mp_input59.Y (\__mp_input59.Y__gold ),
    .\__mp_input6.A (\__mp_input6.A__gold ),
    .\__mp_input6.Y (\__mp_input6.Y__gold ),
    .\__mp_input60.A (\__mp_input60.A__gold ),
    .\__mp_input60.Y (\__mp_input60.Y__gold ),
    .\__mp_input61.A (\__mp_input61.A__gold ),
    .\__mp_input61.Y (\__mp_input61.Y__gold ),
    .\__mp_input62.A (\__mp_input62.A__gold ),
    .\__mp_input62.Y (\__mp_input62.Y__gold ),
    .\__mp_input63.A (\__mp_input63.A__gold ),
    .\__mp_input63.Y (\__mp_input63.Y__gold ),
    .\__mp_input64.A (\__mp_input64.A__gold ),
    .\__mp_input64.Y (\__mp_input64.Y__gold ),
    .\__mp_input65.A (\__mp_input65.A__gold ),
    .\__mp_input65.Y (\__mp_input65.Y__gold ),
    .\__mp_input66.A (\__mp_input66.A__gold ),
    .\__mp_input66.Y (\__mp_input66.Y__gold ),
    .\__mp_input67.A (\__mp_input67.A__gold ),
    .\__mp_input67.Y (\__mp_input67.Y__gold ),
    .\__mp_input68.A (\__mp_input68.A__gold ),
    .\__mp_input68.Y (\__mp_input68.Y__gold ),
    .\__mp_input69.A (\__mp_input69.A__gold ),
    .\__mp_input69.Y (\__mp_input69.Y__gold ),
    .\__mp_input7.A (\__mp_input7.A__gold ),
    .\__mp_input7.Y (\__mp_input7.Y__gold ),
    .\__mp_input70.A (\__mp_input70.A__gold ),
    .\__mp_input70.Y (\__mp_input70.Y__gold ),
    .\__mp_input71.A (\__mp_input71.A__gold ),
    .\__mp_input71.Y (\__mp_input71.Y__gold ),
    .\__mp_input72.A (\__mp_input72.A__gold ),
    .\__mp_input72.Y (\__mp_input72.Y__gold ),
    .\__mp_input73.A (\__mp_input73.A__gold ),
    .\__mp_input73.Y (\__mp_input73.Y__gold ),
    .\__mp_input74.A (\__mp_input74.A__gold ),
    .\__mp_input74.Y (\__mp_input74.Y__gold ),
    .\__mp_input75.A (\__mp_input75.A__gold ),
    .\__mp_input75.Y (\__mp_input75.Y__gold ),
    .\__mp_input76.A (\__mp_input76.A__gold ),
    .\__mp_input76.Y (\__mp_input76.Y__gold ),
    .\__mp_input77.A (\__mp_input77.A__gold ),
    .\__mp_input77.Y (\__mp_input77.Y__gold ),
    .\__mp_input78.A (\__mp_input78.A__gold ),
    .\__mp_input78.Y (\__mp_input78.Y__gold ),
    .\__mp_input79.A (\__mp_input79.A__gold ),
    .\__mp_input79.Y (\__mp_input79.Y__gold ),
    .\__mp_input8.A (\__mp_input8.A__gold ),
    .\__mp_input8.Y (\__mp_input8.Y__gold ),
    .\__mp_input80.A (\__mp_input80.A__gold ),
    .\__mp_input80.Y (\__mp_input80.Y__gold ),
    .\__mp_input81.A (\__mp_input81.A__gold ),
    .\__mp_input81.Y (\__mp_input81.Y__gold ),
    .\__mp_input82.A (\__mp_input82.A__gold ),
    .\__mp_input82.Y (\__mp_input82.Y__gold ),
    .\__mp_input83.A (\__mp_input83.A__gold ),
    .\__mp_input83.Y (\__mp_input83.Y__gold ),
    .\__mp_input84.A (\__mp_input84.A__gold ),
    .\__mp_input84.Y (\__mp_input84.Y__gold ),
    .\__mp_input85.A (\__mp_input85.A__gold ),
    .\__mp_input85.Y (\__mp_input85.Y__gold ),
    .\__mp_input86.A (\__mp_input86.A__gold ),
    .\__mp_input86.Y (\__mp_input86.Y__gold ),
    .\__mp_input87.A (\__mp_input87.A__gold ),
    .\__mp_input87.Y (\__mp_input87.Y__gold ),
    .\__mp_input88.A (\__mp_input88.A__gold ),
    .\__mp_input88.Y (\__mp_input88.Y__gold ),
    .\__mp_input89.A (\__mp_input89.A__gold ),
    .\__mp_input89.Y (\__mp_input89.Y__gold ),
    .\__mp_input9.A (\__mp_input9.A__gold ),
    .\__mp_input9.Y (\__mp_input9.Y__gold ),
    .\__mp_input90.A (\__mp_input90.A__gold ),
    .\__mp_input90.Y (\__mp_input90.Y__gold ),
    .\__mp_input91.A (\__mp_input91.A__gold ),
    .\__mp_input91.Y (\__mp_input91.Y__gold ),
    .\__mp_input92.A (\__mp_input92.A__gold ),
    .\__mp_input92.Y (\__mp_input92.Y__gold ),
    .\__mp_input93.A (\__mp_input93.A__gold ),
    .\__mp_input93.Y (\__mp_input93.Y__gold ),
    .\__mp_input94.A (\__mp_input94.A__gold ),
    .\__mp_input94.Y (\__mp_input94.Y__gold ),
    .\__mp_input95.A (\__mp_input95.A__gold ),
    .\__mp_input95.Y (\__mp_input95.Y__gold ),
    .\__mp_input96.A (\__mp_input96.A__gold ),
    .\__mp_input96.Y (\__mp_input96.Y__gold ),
    .\__mp_input97.A (\__mp_input97.A__gold ),
    .\__mp_input97.Y (\__mp_input97.Y__gold ),
    .\__mp_input98.A (\__mp_input98.A__gold ),
    .\__mp_input98.Y (\__mp_input98.Y__gold ),
    .\__mp_input99.A (\__mp_input99.A__gold ),
    .\__mp_input99.Y (\__mp_input99.Y__gold ),
    .\__mp_ld_r$_DFF_P_.CLK (\__mp_ld_r$_DFF_P_.CLK__gold ),
    .\__mp_ld_r$_DFF_P_.D (\__mp_ld_r$_DFF_P_.D__gold ),
    .\__mp_output259.A (\__mp_output259.A__gold ),
    .\__mp_output259.Y (\__mp_output259.Y__gold ),
    .\__mp_output260.A (\__mp_output260.A__gold ),
    .\__mp_output260.Y (\__mp_output260.Y__gold ),
    .\__mp_output261.A (\__mp_output261.A__gold ),
    .\__mp_output261.Y (\__mp_output261.Y__gold ),
    .\__mp_output262.A (\__mp_output262.A__gold ),
    .\__mp_output262.Y (\__mp_output262.Y__gold ),
    .\__mp_output263.A (\__mp_output263.A__gold ),
    .\__mp_output263.Y (\__mp_output263.Y__gold ),
    .\__mp_output264.A (\__mp_output264.A__gold ),
    .\__mp_output264.Y (\__mp_output264.Y__gold ),
    .\__mp_output265.A (\__mp_output265.A__gold ),
    .\__mp_output265.Y (\__mp_output265.Y__gold ),
    .\__mp_output266.A (\__mp_output266.A__gold ),
    .\__mp_output266.Y (\__mp_output266.Y__gold ),
    .\__mp_output267.A (\__mp_output267.A__gold ),
    .\__mp_output267.Y (\__mp_output267.Y__gold ),
    .\__mp_output268.A (\__mp_output268.A__gold ),
    .\__mp_output268.Y (\__mp_output268.Y__gold ),
    .\__mp_output269.A (\__mp_output269.A__gold ),
    .\__mp_output269.Y (\__mp_output269.Y__gold ),
    .\__mp_output270.A (\__mp_output270.A__gold ),
    .\__mp_output270.Y (\__mp_output270.Y__gold ),
    .\__mp_output271.A (\__mp_output271.A__gold ),
    .\__mp_output271.Y (\__mp_output271.Y__gold ),
    .\__mp_output272.A (\__mp_output272.A__gold ),
    .\__mp_output272.Y (\__mp_output272.Y__gold ),
    .\__mp_output273.A (\__mp_output273.A__gold ),
    .\__mp_output273.Y (\__mp_output273.Y__gold ),
    .\__mp_output274.A (\__mp_output274.A__gold ),
    .\__mp_output274.Y (\__mp_output274.Y__gold ),
    .\__mp_output275.A (\__mp_output275.A__gold ),
    .\__mp_output275.Y (\__mp_output275.Y__gold ),
    .\__mp_output276.A (\__mp_output276.A__gold ),
    .\__mp_output276.Y (\__mp_output276.Y__gold ),
    .\__mp_output277.A (\__mp_output277.A__gold ),
    .\__mp_output277.Y (\__mp_output277.Y__gold ),
    .\__mp_output278.A (\__mp_output278.A__gold ),
    .\__mp_output278.Y (\__mp_output278.Y__gold ),
    .\__mp_output279.A (\__mp_output279.A__gold ),
    .\__mp_output279.Y (\__mp_output279.Y__gold ),
    .\__mp_output280.A (\__mp_output280.A__gold ),
    .\__mp_output280.Y (\__mp_output280.Y__gold ),
    .\__mp_output281.A (\__mp_output281.A__gold ),
    .\__mp_output281.Y (\__mp_output281.Y__gold ),
    .\__mp_output282.A (\__mp_output282.A__gold ),
    .\__mp_output282.Y (\__mp_output282.Y__gold ),
    .\__mp_output283.A (\__mp_output283.A__gold ),
    .\__mp_output283.Y (\__mp_output283.Y__gold ),
    .\__mp_output284.A (\__mp_output284.A__gold ),
    .\__mp_output284.Y (\__mp_output284.Y__gold ),
    .\__mp_output285.A (\__mp_output285.A__gold ),
    .\__mp_output285.Y (\__mp_output285.Y__gold ),
    .\__mp_output286.A (\__mp_output286.A__gold ),
    .\__mp_output286.Y (\__mp_output286.Y__gold ),
    .\__mp_output287.A (\__mp_output287.A__gold ),
    .\__mp_output287.Y (\__mp_output287.Y__gold ),
    .\__mp_output288.A (\__mp_output288.A__gold ),
    .\__mp_output288.Y (\__mp_output288.Y__gold ),
    .\__mp_output289.A (\__mp_output289.A__gold ),
    .\__mp_output289.Y (\__mp_output289.Y__gold ),
    .\__mp_output290.A (\__mp_output290.A__gold ),
    .\__mp_output290.Y (\__mp_output290.Y__gold ),
    .\__mp_output291.A (\__mp_output291.A__gold ),
    .\__mp_output291.Y (\__mp_output291.Y__gold ),
    .\__mp_output292.A (\__mp_output292.A__gold ),
    .\__mp_output292.Y (\__mp_output292.Y__gold ),
    .\__mp_output293.A (\__mp_output293.A__gold ),
    .\__mp_output293.Y (\__mp_output293.Y__gold ),
    .\__mp_output294.A (\__mp_output294.A__gold ),
    .\__mp_output294.Y (\__mp_output294.Y__gold ),
    .\__mp_output295.A (\__mp_output295.A__gold ),
    .\__mp_output295.Y (\__mp_output295.Y__gold ),
    .\__mp_output296.A (\__mp_output296.A__gold ),
    .\__mp_output296.Y (\__mp_output296.Y__gold ),
    .\__mp_output297.A (\__mp_output297.A__gold ),
    .\__mp_output297.Y (\__mp_output297.Y__gold ),
    .\__mp_output298.A (\__mp_output298.A__gold ),
    .\__mp_output298.Y (\__mp_output298.Y__gold ),
    .\__mp_output299.A (\__mp_output299.A__gold ),
    .\__mp_output299.Y (\__mp_output299.Y__gold ),
    .\__mp_output300.A (\__mp_output300.A__gold ),
    .\__mp_output300.Y (\__mp_output300.Y__gold ),
    .\__mp_output301.A (\__mp_output301.A__gold ),
    .\__mp_output301.Y (\__mp_output301.Y__gold ),
    .\__mp_output302.A (\__mp_output302.A__gold ),
    .\__mp_output302.Y (\__mp_output302.Y__gold ),
    .\__mp_output303.A (\__mp_output303.A__gold ),
    .\__mp_output303.Y (\__mp_output303.Y__gold ),
    .\__mp_output304.A (\__mp_output304.A__gold ),
    .\__mp_output304.Y (\__mp_output304.Y__gold ),
    .\__mp_output305.A (\__mp_output305.A__gold ),
    .\__mp_output305.Y (\__mp_output305.Y__gold ),
    .\__mp_output306.A (\__mp_output306.A__gold ),
    .\__mp_output306.Y (\__mp_output306.Y__gold ),
    .\__mp_output307.A (\__mp_output307.A__gold ),
    .\__mp_output307.Y (\__mp_output307.Y__gold ),
    .\__mp_output308.A (\__mp_output308.A__gold ),
    .\__mp_output308.Y (\__mp_output308.Y__gold ),
    .\__mp_output309.A (\__mp_output309.A__gold ),
    .\__mp_output309.Y (\__mp_output309.Y__gold ),
    .\__mp_output310.A (\__mp_output310.A__gold ),
    .\__mp_output310.Y (\__mp_output310.Y__gold ),
    .\__mp_output311.A (\__mp_output311.A__gold ),
    .\__mp_output311.Y (\__mp_output311.Y__gold ),
    .\__mp_output312.A (\__mp_output312.A__gold ),
    .\__mp_output312.Y (\__mp_output312.Y__gold ),
    .\__mp_output313.A (\__mp_output313.A__gold ),
    .\__mp_output313.Y (\__mp_output313.Y__gold ),
    .\__mp_output314.A (\__mp_output314.A__gold ),
    .\__mp_output314.Y (\__mp_output314.Y__gold ),
    .\__mp_output315.A (\__mp_output315.A__gold ),
    .\__mp_output315.Y (\__mp_output315.Y__gold ),
    .\__mp_output316.A (\__mp_output316.A__gold ),
    .\__mp_output316.Y (\__mp_output316.Y__gold ),
    .\__mp_output317.A (\__mp_output317.A__gold ),
    .\__mp_output317.Y (\__mp_output317.Y__gold ),
    .\__mp_output318.A (\__mp_output318.A__gold ),
    .\__mp_output318.Y (\__mp_output318.Y__gold ),
    .\__mp_output319.A (\__mp_output319.A__gold ),
    .\__mp_output319.Y (\__mp_output319.Y__gold ),
    .\__mp_output320.A (\__mp_output320.A__gold ),
    .\__mp_output320.Y (\__mp_output320.Y__gold ),
    .\__mp_output321.A (\__mp_output321.A__gold ),
    .\__mp_output321.Y (\__mp_output321.Y__gold ),
    .\__mp_output322.A (\__mp_output322.A__gold ),
    .\__mp_output322.Y (\__mp_output322.Y__gold ),
    .\__mp_output323.A (\__mp_output323.A__gold ),
    .\__mp_output323.Y (\__mp_output323.Y__gold ),
    .\__mp_output324.A (\__mp_output324.A__gold ),
    .\__mp_output324.Y (\__mp_output324.Y__gold ),
    .\__mp_output325.A (\__mp_output325.A__gold ),
    .\__mp_output325.Y (\__mp_output325.Y__gold ),
    .\__mp_output326.A (\__mp_output326.A__gold ),
    .\__mp_output326.Y (\__mp_output326.Y__gold ),
    .\__mp_output327.A (\__mp_output327.A__gold ),
    .\__mp_output327.Y (\__mp_output327.Y__gold ),
    .\__mp_output328.A (\__mp_output328.A__gold ),
    .\__mp_output328.Y (\__mp_output328.Y__gold ),
    .\__mp_output329.A (\__mp_output329.A__gold ),
    .\__mp_output329.Y (\__mp_output329.Y__gold ),
    .\__mp_output330.A (\__mp_output330.A__gold ),
    .\__mp_output330.Y (\__mp_output330.Y__gold ),
    .\__mp_output331.A (\__mp_output331.A__gold ),
    .\__mp_output331.Y (\__mp_output331.Y__gold ),
    .\__mp_output332.A (\__mp_output332.A__gold ),
    .\__mp_output332.Y (\__mp_output332.Y__gold ),
    .\__mp_output333.A (\__mp_output333.A__gold ),
    .\__mp_output333.Y (\__mp_output333.Y__gold ),
    .\__mp_output334.A (\__mp_output334.A__gold ),
    .\__mp_output334.Y (\__mp_output334.Y__gold ),
    .\__mp_output335.A (\__mp_output335.A__gold ),
    .\__mp_output335.Y (\__mp_output335.Y__gold ),
    .\__mp_output336.A (\__mp_output336.A__gold ),
    .\__mp_output336.Y (\__mp_output336.Y__gold ),
    .\__mp_output337.A (\__mp_output337.A__gold ),
    .\__mp_output337.Y (\__mp_output337.Y__gold ),
    .\__mp_output338.A (\__mp_output338.A__gold ),
    .\__mp_output338.Y (\__mp_output338.Y__gold ),
    .\__mp_output339.A (\__mp_output339.A__gold ),
    .\__mp_output339.Y (\__mp_output339.Y__gold ),
    .\__mp_output340.A (\__mp_output340.A__gold ),
    .\__mp_output340.Y (\__mp_output340.Y__gold ),
    .\__mp_output341.A (\__mp_output341.A__gold ),
    .\__mp_output341.Y (\__mp_output341.Y__gold ),
    .\__mp_output342.A (\__mp_output342.A__gold ),
    .\__mp_output342.Y (\__mp_output342.Y__gold ),
    .\__mp_output343.A (\__mp_output343.A__gold ),
    .\__mp_output343.Y (\__mp_output343.Y__gold ),
    .\__mp_output344.A (\__mp_output344.A__gold ),
    .\__mp_output344.Y (\__mp_output344.Y__gold ),
    .\__mp_output345.A (\__mp_output345.A__gold ),
    .\__mp_output345.Y (\__mp_output345.Y__gold ),
    .\__mp_output346.A (\__mp_output346.A__gold ),
    .\__mp_output346.Y (\__mp_output346.Y__gold ),
    .\__mp_output347.A (\__mp_output347.A__gold ),
    .\__mp_output347.Y (\__mp_output347.Y__gold ),
    .\__mp_output348.A (\__mp_output348.A__gold ),
    .\__mp_output348.Y (\__mp_output348.Y__gold ),
    .\__mp_output349.A (\__mp_output349.A__gold ),
    .\__mp_output349.Y (\__mp_output349.Y__gold ),
    .\__mp_output350.A (\__mp_output350.A__gold ),
    .\__mp_output350.Y (\__mp_output350.Y__gold ),
    .\__mp_output351.A (\__mp_output351.A__gold ),
    .\__mp_output351.Y (\__mp_output351.Y__gold ),
    .\__mp_output352.A (\__mp_output352.A__gold ),
    .\__mp_output352.Y (\__mp_output352.Y__gold ),
    .\__mp_output353.A (\__mp_output353.A__gold ),
    .\__mp_output353.Y (\__mp_output353.Y__gold ),
    .\__mp_output354.A (\__mp_output354.A__gold ),
    .\__mp_output354.Y (\__mp_output354.Y__gold ),
    .\__mp_output355.A (\__mp_output355.A__gold ),
    .\__mp_output355.Y (\__mp_output355.Y__gold ),
    .\__mp_output356.A (\__mp_output356.A__gold ),
    .\__mp_output356.Y (\__mp_output356.Y__gold ),
    .\__mp_output357.A (\__mp_output357.A__gold ),
    .\__mp_output357.Y (\__mp_output357.Y__gold ),
    .\__mp_output358.A (\__mp_output358.A__gold ),
    .\__mp_output358.Y (\__mp_output358.Y__gold ),
    .\__mp_output359.A (\__mp_output359.A__gold ),
    .\__mp_output359.Y (\__mp_output359.Y__gold ),
    .\__mp_output360.A (\__mp_output360.A__gold ),
    .\__mp_output360.Y (\__mp_output360.Y__gold ),
    .\__mp_output361.A (\__mp_output361.A__gold ),
    .\__mp_output361.Y (\__mp_output361.Y__gold ),
    .\__mp_output362.A (\__mp_output362.A__gold ),
    .\__mp_output362.Y (\__mp_output362.Y__gold ),
    .\__mp_output363.A (\__mp_output363.A__gold ),
    .\__mp_output363.Y (\__mp_output363.Y__gold ),
    .\__mp_output364.A (\__mp_output364.A__gold ),
    .\__mp_output364.Y (\__mp_output364.Y__gold ),
    .\__mp_output365.A (\__mp_output365.A__gold ),
    .\__mp_output365.Y (\__mp_output365.Y__gold ),
    .\__mp_output366.A (\__mp_output366.A__gold ),
    .\__mp_output366.Y (\__mp_output366.Y__gold ),
    .\__mp_output367.A (\__mp_output367.A__gold ),
    .\__mp_output367.Y (\__mp_output367.Y__gold ),
    .\__mp_output368.A (\__mp_output368.A__gold ),
    .\__mp_output368.Y (\__mp_output368.Y__gold ),
    .\__mp_output369.A (\__mp_output369.A__gold ),
    .\__mp_output369.Y (\__mp_output369.Y__gold ),
    .\__mp_output370.A (\__mp_output370.A__gold ),
    .\__mp_output370.Y (\__mp_output370.Y__gold ),
    .\__mp_output371.A (\__mp_output371.A__gold ),
    .\__mp_output371.Y (\__mp_output371.Y__gold ),
    .\__mp_output372.A (\__mp_output372.A__gold ),
    .\__mp_output372.Y (\__mp_output372.Y__gold ),
    .\__mp_output373.A (\__mp_output373.A__gold ),
    .\__mp_output373.Y (\__mp_output373.Y__gold ),
    .\__mp_output374.A (\__mp_output374.A__gold ),
    .\__mp_output374.Y (\__mp_output374.Y__gold ),
    .\__mp_output375.A (\__mp_output375.A__gold ),
    .\__mp_output375.Y (\__mp_output375.Y__gold ),
    .\__mp_output376.A (\__mp_output376.A__gold ),
    .\__mp_output376.Y (\__mp_output376.Y__gold ),
    .\__mp_output377.A (\__mp_output377.A__gold ),
    .\__mp_output377.Y (\__mp_output377.Y__gold ),
    .\__mp_output378.A (\__mp_output378.A__gold ),
    .\__mp_output378.Y (\__mp_output378.Y__gold ),
    .\__mp_output379.A (\__mp_output379.A__gold ),
    .\__mp_output379.Y (\__mp_output379.Y__gold ),
    .\__mp_output380.A (\__mp_output380.A__gold ),
    .\__mp_output380.Y (\__mp_output380.Y__gold ),
    .\__mp_output381.A (\__mp_output381.A__gold ),
    .\__mp_output381.Y (\__mp_output381.Y__gold ),
    .\__mp_output382.A (\__mp_output382.A__gold ),
    .\__mp_output382.Y (\__mp_output382.Y__gold ),
    .\__mp_output383.A (\__mp_output383.A__gold ),
    .\__mp_output383.Y (\__mp_output383.Y__gold ),
    .\__mp_output384.A (\__mp_output384.A__gold ),
    .\__mp_output384.Y (\__mp_output384.Y__gold ),
    .\__mp_output385.A (\__mp_output385.A__gold ),
    .\__mp_output385.Y (\__mp_output385.Y__gold ),
    .\__mp_output386.A (\__mp_output386.A__gold ),
    .\__mp_output386.Y (\__mp_output386.Y__gold ),
    .\__mp_output387.A (\__mp_output387.A__gold ),
    .\__mp_output387.Y (\__mp_output387.Y__gold ),
    .\__mp_sa00_sr[0]$_DFF_P_.CLK (\__mp_sa00_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa00_sr[1]$_DFF_P_.CLK (\__mp_sa00_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa00_sr[2]$_DFF_P_.CLK (\__mp_sa00_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa00_sr[3]$_DFF_P_.CLK (\__mp_sa00_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa00_sr[4]$_DFF_P_.CLK (\__mp_sa00_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa00_sr[5]$_DFF_P_.CLK (\__mp_sa00_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa00_sr[6]$_DFF_P_.CLK (\__mp_sa00_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa00_sr[7]$_DFF_P_.CLK (\__mp_sa00_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[0]$_DFF_P_.CLK (\__mp_sa01_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[1]$_DFF_P_.CLK (\__mp_sa01_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[2]$_DFF_P_.CLK (\__mp_sa01_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[3]$_DFF_P_.CLK (\__mp_sa01_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[4]$_DFF_P_.CLK (\__mp_sa01_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[5]$_DFF_P_.CLK (\__mp_sa01_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[6]$_DFF_P_.CLK (\__mp_sa01_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa01_sr[7]$_DFF_P_.CLK (\__mp_sa01_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[0]$_DFF_P_.CLK (\__mp_sa02_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[1]$_DFF_P_.CLK (\__mp_sa02_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[2]$_DFF_P_.CLK (\__mp_sa02_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[3]$_DFF_P_.CLK (\__mp_sa02_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[4]$_DFF_P_.CLK (\__mp_sa02_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[5]$_DFF_P_.CLK (\__mp_sa02_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[6]$_DFF_P_.CLK (\__mp_sa02_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa02_sr[7]$_DFF_P_.CLK (\__mp_sa02_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[0]$_DFF_P_.CLK (\__mp_sa03_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[1]$_DFF_P_.CLK (\__mp_sa03_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[2]$_DFF_P_.CLK (\__mp_sa03_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[3]$_DFF_P_.CLK (\__mp_sa03_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[4]$_DFF_P_.CLK (\__mp_sa03_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[5]$_DFF_P_.CLK (\__mp_sa03_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[6]$_DFF_P_.CLK (\__mp_sa03_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa03_sr[7]$_DFF_P_.CLK (\__mp_sa03_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[0]$_DFF_P_.CLK (\__mp_sa10_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[1]$_DFF_P_.CLK (\__mp_sa10_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[2]$_DFF_P_.CLK (\__mp_sa10_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[3]$_DFF_P_.CLK (\__mp_sa10_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[4]$_DFF_P_.CLK (\__mp_sa10_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[5]$_DFF_P_.CLK (\__mp_sa10_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[6]$_DFF_P_.CLK (\__mp_sa10_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa10_sr[7]$_DFF_P_.CLK (\__mp_sa10_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[0]$_DFF_P_.CLK (\__mp_sa11_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[1]$_DFF_P_.CLK (\__mp_sa11_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[2]$_DFF_P_.CLK (\__mp_sa11_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[3]$_DFF_P_.CLK (\__mp_sa11_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[4]$_DFF_P_.CLK (\__mp_sa11_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[5]$_DFF_P_.CLK (\__mp_sa11_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[6]$_DFF_P_.CLK (\__mp_sa11_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa11_sr[7]$_DFF_P_.CLK (\__mp_sa11_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[0]$_DFF_P_.CLK (\__mp_sa12_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[1]$_DFF_P_.CLK (\__mp_sa12_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[2]$_DFF_P_.CLK (\__mp_sa12_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[3]$_DFF_P_.CLK (\__mp_sa12_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[4]$_DFF_P_.CLK (\__mp_sa12_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[5]$_DFF_P_.CLK (\__mp_sa12_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[6]$_DFF_P_.CLK (\__mp_sa12_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa12_sr[7]$_DFF_P_.CLK (\__mp_sa12_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[0]$_DFF_P_.CLK (\__mp_sa13_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[1]$_DFF_P_.CLK (\__mp_sa13_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[2]$_DFF_P_.CLK (\__mp_sa13_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[3]$_DFF_P_.CLK (\__mp_sa13_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[4]$_DFF_P_.CLK (\__mp_sa13_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[5]$_DFF_P_.CLK (\__mp_sa13_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[6]$_DFF_P_.CLK (\__mp_sa13_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa13_sr[7]$_DFF_P_.CLK (\__mp_sa13_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[0]$_DFF_P_.CLK (\__mp_sa20_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[1]$_DFF_P_.CLK (\__mp_sa20_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[2]$_DFF_P_.CLK (\__mp_sa20_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[3]$_DFF_P_.CLK (\__mp_sa20_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[4]$_DFF_P_.CLK (\__mp_sa20_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[5]$_DFF_P_.CLK (\__mp_sa20_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[6]$_DFF_P_.CLK (\__mp_sa20_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa20_sr[7]$_DFF_P_.CLK (\__mp_sa20_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[0]$_DFF_P_.CLK (\__mp_sa21_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[1]$_DFF_P_.CLK (\__mp_sa21_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[2]$_DFF_P_.CLK (\__mp_sa21_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[3]$_DFF_P_.CLK (\__mp_sa21_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[4]$_DFF_P_.CLK (\__mp_sa21_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[5]$_DFF_P_.CLK (\__mp_sa21_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[6]$_DFF_P_.CLK (\__mp_sa21_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa21_sr[7]$_DFF_P_.CLK (\__mp_sa21_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[0]$_DFF_P_.CLK (\__mp_sa22_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[1]$_DFF_P_.CLK (\__mp_sa22_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[2]$_DFF_P_.CLK (\__mp_sa22_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[3]$_DFF_P_.CLK (\__mp_sa22_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[4]$_DFF_P_.CLK (\__mp_sa22_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[5]$_DFF_P_.CLK (\__mp_sa22_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[6]$_DFF_P_.CLK (\__mp_sa22_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa22_sr[7]$_DFF_P_.CLK (\__mp_sa22_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[0]$_DFF_P_.CLK (\__mp_sa23_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[1]$_DFF_P_.CLK (\__mp_sa23_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[2]$_DFF_P_.CLK (\__mp_sa23_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[3]$_DFF_P_.CLK (\__mp_sa23_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[4]$_DFF_P_.CLK (\__mp_sa23_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[5]$_DFF_P_.CLK (\__mp_sa23_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[6]$_DFF_P_.CLK (\__mp_sa23_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa23_sr[7]$_DFF_P_.CLK (\__mp_sa23_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[0]$_DFF_P_.CLK (\__mp_sa30_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[1]$_DFF_P_.CLK (\__mp_sa30_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[2]$_DFF_P_.CLK (\__mp_sa30_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[3]$_DFF_P_.CLK (\__mp_sa30_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[4]$_DFF_P_.CLK (\__mp_sa30_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[5]$_DFF_P_.CLK (\__mp_sa30_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[6]$_DFF_P_.CLK (\__mp_sa30_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa30_sr[7]$_DFF_P_.CLK (\__mp_sa30_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[0]$_DFF_P_.CLK (\__mp_sa31_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[1]$_DFF_P_.CLK (\__mp_sa31_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[2]$_DFF_P_.CLK (\__mp_sa31_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[3]$_DFF_P_.CLK (\__mp_sa31_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[4]$_DFF_P_.CLK (\__mp_sa31_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[5]$_DFF_P_.CLK (\__mp_sa31_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[6]$_DFF_P_.CLK (\__mp_sa31_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa31_sr[7]$_DFF_P_.CLK (\__mp_sa31_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[0]$_DFF_P_.CLK (\__mp_sa32_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[1]$_DFF_P_.CLK (\__mp_sa32_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[2]$_DFF_P_.CLK (\__mp_sa32_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[3]$_DFF_P_.CLK (\__mp_sa32_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[4]$_DFF_P_.CLK (\__mp_sa32_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[5]$_DFF_P_.CLK (\__mp_sa32_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[6]$_DFF_P_.CLK (\__mp_sa32_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa32_sr[7]$_DFF_P_.CLK (\__mp_sa32_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[0]$_DFF_P_.CLK (\__mp_sa33_sr[0]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[1]$_DFF_P_.CLK (\__mp_sa33_sr[1]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[2]$_DFF_P_.CLK (\__mp_sa33_sr[2]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[3]$_DFF_P_.CLK (\__mp_sa33_sr[3]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[4]$_DFF_P_.CLK (\__mp_sa33_sr[4]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[5]$_DFF_P_.CLK (\__mp_sa33_sr[5]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[6]$_DFF_P_.CLK (\__mp_sa33_sr[6]$_DFF_P_.CLK__gold ),
    .\__mp_sa33_sr[7]$_DFF_P_.CLK (\__mp_sa33_sr[7]$_DFF_P_.CLK__gold ),
    .\__mp_text_in_r[0]$_DFFE_PP_.CLK (\__mp_text_in_r[0]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[100]$_DFFE_PP_.CLK (\__mp_text_in_r[100]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[101]$_DFFE_PP_.CLK (\__mp_text_in_r[101]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[102]$_DFFE_PP_.CLK (\__mp_text_in_r[102]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[103]$_DFFE_PP_.CLK (\__mp_text_in_r[103]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[104]$_DFFE_PP_.CLK (\__mp_text_in_r[104]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[105]$_DFFE_PP_.CLK (\__mp_text_in_r[105]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[106]$_DFFE_PP_.CLK (\__mp_text_in_r[106]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[107]$_DFFE_PP_.CLK (\__mp_text_in_r[107]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[108]$_DFFE_PP_.CLK (\__mp_text_in_r[108]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[109]$_DFFE_PP_.CLK (\__mp_text_in_r[109]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[10]$_DFFE_PP_.CLK (\__mp_text_in_r[10]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[110]$_DFFE_PP_.CLK (\__mp_text_in_r[110]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[111]$_DFFE_PP_.CLK (\__mp_text_in_r[111]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[112]$_DFFE_PP_.CLK (\__mp_text_in_r[112]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[113]$_DFFE_PP_.CLK (\__mp_text_in_r[113]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[114]$_DFFE_PP_.CLK (\__mp_text_in_r[114]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[115]$_DFFE_PP_.CLK (\__mp_text_in_r[115]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[116]$_DFFE_PP_.CLK (\__mp_text_in_r[116]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[117]$_DFFE_PP_.CLK (\__mp_text_in_r[117]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[118]$_DFFE_PP_.CLK (\__mp_text_in_r[118]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[119]$_DFFE_PP_.CLK (\__mp_text_in_r[119]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[11]$_DFFE_PP_.CLK (\__mp_text_in_r[11]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[120]$_DFFE_PP_.CLK (\__mp_text_in_r[120]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[121]$_DFFE_PP_.CLK (\__mp_text_in_r[121]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[122]$_DFFE_PP_.CLK (\__mp_text_in_r[122]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[123]$_DFFE_PP_.CLK (\__mp_text_in_r[123]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[124]$_DFFE_PP_.CLK (\__mp_text_in_r[124]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[125]$_DFFE_PP_.CLK (\__mp_text_in_r[125]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[126]$_DFFE_PP_.CLK (\__mp_text_in_r[126]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[127]$_DFFE_PP_.CLK (\__mp_text_in_r[127]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[12]$_DFFE_PP_.CLK (\__mp_text_in_r[12]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[13]$_DFFE_PP_.CLK (\__mp_text_in_r[13]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[14]$_DFFE_PP_.CLK (\__mp_text_in_r[14]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[15]$_DFFE_PP_.CLK (\__mp_text_in_r[15]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[16]$_DFFE_PP_.CLK (\__mp_text_in_r[16]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[17]$_DFFE_PP_.CLK (\__mp_text_in_r[17]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[18]$_DFFE_PP_.CLK (\__mp_text_in_r[18]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[19]$_DFFE_PP_.CLK (\__mp_text_in_r[19]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[1]$_DFFE_PP_.CLK (\__mp_text_in_r[1]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[20]$_DFFE_PP_.CLK (\__mp_text_in_r[20]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[21]$_DFFE_PP_.CLK (\__mp_text_in_r[21]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[22]$_DFFE_PP_.CLK (\__mp_text_in_r[22]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[23]$_DFFE_PP_.CLK (\__mp_text_in_r[23]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[24]$_DFFE_PP_.CLK (\__mp_text_in_r[24]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[25]$_DFFE_PP_.CLK (\__mp_text_in_r[25]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[26]$_DFFE_PP_.CLK (\__mp_text_in_r[26]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[27]$_DFFE_PP_.CLK (\__mp_text_in_r[27]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[28]$_DFFE_PP_.CLK (\__mp_text_in_r[28]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[29]$_DFFE_PP_.CLK (\__mp_text_in_r[29]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[2]$_DFFE_PP_.CLK (\__mp_text_in_r[2]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[30]$_DFFE_PP_.CLK (\__mp_text_in_r[30]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[31]$_DFFE_PP_.CLK (\__mp_text_in_r[31]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[32]$_DFFE_PP_.CLK (\__mp_text_in_r[32]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[33]$_DFFE_PP_.CLK (\__mp_text_in_r[33]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[34]$_DFFE_PP_.CLK (\__mp_text_in_r[34]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[35]$_DFFE_PP_.CLK (\__mp_text_in_r[35]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[36]$_DFFE_PP_.CLK (\__mp_text_in_r[36]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[37]$_DFFE_PP_.CLK (\__mp_text_in_r[37]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[38]$_DFFE_PP_.CLK (\__mp_text_in_r[38]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[39]$_DFFE_PP_.CLK (\__mp_text_in_r[39]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[3]$_DFFE_PP_.CLK (\__mp_text_in_r[3]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[40]$_DFFE_PP_.CLK (\__mp_text_in_r[40]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[41]$_DFFE_PP_.CLK (\__mp_text_in_r[41]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[42]$_DFFE_PP_.CLK (\__mp_text_in_r[42]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[43]$_DFFE_PP_.CLK (\__mp_text_in_r[43]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[44]$_DFFE_PP_.CLK (\__mp_text_in_r[44]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[45]$_DFFE_PP_.CLK (\__mp_text_in_r[45]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[46]$_DFFE_PP_.CLK (\__mp_text_in_r[46]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[47]$_DFFE_PP_.CLK (\__mp_text_in_r[47]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[48]$_DFFE_PP_.CLK (\__mp_text_in_r[48]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[49]$_DFFE_PP_.CLK (\__mp_text_in_r[49]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[4]$_DFFE_PP_.CLK (\__mp_text_in_r[4]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[50]$_DFFE_PP_.CLK (\__mp_text_in_r[50]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[51]$_DFFE_PP_.CLK (\__mp_text_in_r[51]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[52]$_DFFE_PP_.CLK (\__mp_text_in_r[52]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[53]$_DFFE_PP_.CLK (\__mp_text_in_r[53]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[54]$_DFFE_PP_.CLK (\__mp_text_in_r[54]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[55]$_DFFE_PP_.CLK (\__mp_text_in_r[55]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[56]$_DFFE_PP_.CLK (\__mp_text_in_r[56]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[57]$_DFFE_PP_.CLK (\__mp_text_in_r[57]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[58]$_DFFE_PP_.CLK (\__mp_text_in_r[58]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[59]$_DFFE_PP_.CLK (\__mp_text_in_r[59]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[5]$_DFFE_PP_.CLK (\__mp_text_in_r[5]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[60]$_DFFE_PP_.CLK (\__mp_text_in_r[60]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[61]$_DFFE_PP_.CLK (\__mp_text_in_r[61]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[62]$_DFFE_PP_.CLK (\__mp_text_in_r[62]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[63]$_DFFE_PP_.CLK (\__mp_text_in_r[63]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[64]$_DFFE_PP_.CLK (\__mp_text_in_r[64]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[65]$_DFFE_PP_.CLK (\__mp_text_in_r[65]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[66]$_DFFE_PP_.CLK (\__mp_text_in_r[66]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[67]$_DFFE_PP_.CLK (\__mp_text_in_r[67]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[68]$_DFFE_PP_.CLK (\__mp_text_in_r[68]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[69]$_DFFE_PP_.CLK (\__mp_text_in_r[69]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[6]$_DFFE_PP_.CLK (\__mp_text_in_r[6]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[70]$_DFFE_PP_.CLK (\__mp_text_in_r[70]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[71]$_DFFE_PP_.CLK (\__mp_text_in_r[71]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[72]$_DFFE_PP_.CLK (\__mp_text_in_r[72]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[73]$_DFFE_PP_.CLK (\__mp_text_in_r[73]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[74]$_DFFE_PP_.CLK (\__mp_text_in_r[74]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[75]$_DFFE_PP_.CLK (\__mp_text_in_r[75]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[76]$_DFFE_PP_.CLK (\__mp_text_in_r[76]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[77]$_DFFE_PP_.CLK (\__mp_text_in_r[77]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[78]$_DFFE_PP_.CLK (\__mp_text_in_r[78]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[79]$_DFFE_PP_.CLK (\__mp_text_in_r[79]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[7]$_DFFE_PP_.CLK (\__mp_text_in_r[7]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[80]$_DFFE_PP_.CLK (\__mp_text_in_r[80]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[81]$_DFFE_PP_.CLK (\__mp_text_in_r[81]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[82]$_DFFE_PP_.CLK (\__mp_text_in_r[82]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[83]$_DFFE_PP_.CLK (\__mp_text_in_r[83]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[84]$_DFFE_PP_.CLK (\__mp_text_in_r[84]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[85]$_DFFE_PP_.CLK (\__mp_text_in_r[85]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[86]$_DFFE_PP_.CLK (\__mp_text_in_r[86]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[87]$_DFFE_PP_.CLK (\__mp_text_in_r[87]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[88]$_DFFE_PP_.CLK (\__mp_text_in_r[88]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[89]$_DFFE_PP_.CLK (\__mp_text_in_r[89]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[8]$_DFFE_PP_.CLK (\__mp_text_in_r[8]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[90]$_DFFE_PP_.CLK (\__mp_text_in_r[90]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[91]$_DFFE_PP_.CLK (\__mp_text_in_r[91]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[92]$_DFFE_PP_.CLK (\__mp_text_in_r[92]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[93]$_DFFE_PP_.CLK (\__mp_text_in_r[93]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[94]$_DFFE_PP_.CLK (\__mp_text_in_r[94]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[95]$_DFFE_PP_.CLK (\__mp_text_in_r[95]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[96]$_DFFE_PP_.CLK (\__mp_text_in_r[96]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[97]$_DFFE_PP_.CLK (\__mp_text_in_r[97]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[98]$_DFFE_PP_.CLK (\__mp_text_in_r[98]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[99]$_DFFE_PP_.CLK (\__mp_text_in_r[99]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_in_r[9]$_DFFE_PP_.CLK (\__mp_text_in_r[9]$_DFFE_PP_.CLK__gold ),
    .\__mp_text_out[0]$_DFF_P_.CLK (\__mp_text_out[0]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[0]$_DFF_P_.QN (\__mp_text_out[0]$_DFF_P_.QN__gold ),
    .\__mp_text_out[0]$_DFF_P_.int_fwire_IQN (\__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[100]$_DFF_P_.CLK (\__mp_text_out[100]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[100]$_DFF_P_.QN (\__mp_text_out[100]$_DFF_P_.QN__gold ),
    .\__mp_text_out[100]$_DFF_P_.int_fwire_IQN (\__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[101]$_DFF_P_.CLK (\__mp_text_out[101]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[101]$_DFF_P_.QN (\__mp_text_out[101]$_DFF_P_.QN__gold ),
    .\__mp_text_out[101]$_DFF_P_.int_fwire_IQN (\__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[102]$_DFF_P_.CLK (\__mp_text_out[102]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[102]$_DFF_P_.QN (\__mp_text_out[102]$_DFF_P_.QN__gold ),
    .\__mp_text_out[102]$_DFF_P_.int_fwire_IQN (\__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[103]$_DFF_P_.CLK (\__mp_text_out[103]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[103]$_DFF_P_.QN (\__mp_text_out[103]$_DFF_P_.QN__gold ),
    .\__mp_text_out[103]$_DFF_P_.int_fwire_IQN (\__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[104]$_DFF_P_.CLK (\__mp_text_out[104]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[104]$_DFF_P_.QN (\__mp_text_out[104]$_DFF_P_.QN__gold ),
    .\__mp_text_out[104]$_DFF_P_.int_fwire_IQN (\__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[105]$_DFF_P_.CLK (\__mp_text_out[105]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[105]$_DFF_P_.QN (\__mp_text_out[105]$_DFF_P_.QN__gold ),
    .\__mp_text_out[105]$_DFF_P_.int_fwire_IQN (\__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[106]$_DFF_P_.CLK (\__mp_text_out[106]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[106]$_DFF_P_.QN (\__mp_text_out[106]$_DFF_P_.QN__gold ),
    .\__mp_text_out[106]$_DFF_P_.int_fwire_IQN (\__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[107]$_DFF_P_.CLK (\__mp_text_out[107]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[107]$_DFF_P_.QN (\__mp_text_out[107]$_DFF_P_.QN__gold ),
    .\__mp_text_out[107]$_DFF_P_.int_fwire_IQN (\__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[108]$_DFF_P_.CLK (\__mp_text_out[108]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[108]$_DFF_P_.QN (\__mp_text_out[108]$_DFF_P_.QN__gold ),
    .\__mp_text_out[108]$_DFF_P_.int_fwire_IQN (\__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[109]$_DFF_P_.CLK (\__mp_text_out[109]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[109]$_DFF_P_.QN (\__mp_text_out[109]$_DFF_P_.QN__gold ),
    .\__mp_text_out[109]$_DFF_P_.int_fwire_IQN (\__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[10]$_DFF_P_.CLK (\__mp_text_out[10]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[10]$_DFF_P_.QN (\__mp_text_out[10]$_DFF_P_.QN__gold ),
    .\__mp_text_out[10]$_DFF_P_.int_fwire_IQN (\__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[110]$_DFF_P_.CLK (\__mp_text_out[110]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[110]$_DFF_P_.QN (\__mp_text_out[110]$_DFF_P_.QN__gold ),
    .\__mp_text_out[110]$_DFF_P_.int_fwire_IQN (\__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[111]$_DFF_P_.CLK (\__mp_text_out[111]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[111]$_DFF_P_.QN (\__mp_text_out[111]$_DFF_P_.QN__gold ),
    .\__mp_text_out[111]$_DFF_P_.int_fwire_IQN (\__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[112]$_DFF_P_.CLK (\__mp_text_out[112]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[112]$_DFF_P_.QN (\__mp_text_out[112]$_DFF_P_.QN__gold ),
    .\__mp_text_out[112]$_DFF_P_.int_fwire_IQN (\__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[113]$_DFF_P_.CLK (\__mp_text_out[113]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[113]$_DFF_P_.QN (\__mp_text_out[113]$_DFF_P_.QN__gold ),
    .\__mp_text_out[113]$_DFF_P_.int_fwire_IQN (\__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[114]$_DFF_P_.CLK (\__mp_text_out[114]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[114]$_DFF_P_.QN (\__mp_text_out[114]$_DFF_P_.QN__gold ),
    .\__mp_text_out[114]$_DFF_P_.int_fwire_IQN (\__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[115]$_DFF_P_.CLK (\__mp_text_out[115]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[115]$_DFF_P_.QN (\__mp_text_out[115]$_DFF_P_.QN__gold ),
    .\__mp_text_out[115]$_DFF_P_.int_fwire_IQN (\__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[116]$_DFF_P_.CLK (\__mp_text_out[116]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[116]$_DFF_P_.QN (\__mp_text_out[116]$_DFF_P_.QN__gold ),
    .\__mp_text_out[116]$_DFF_P_.int_fwire_IQN (\__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[117]$_DFF_P_.CLK (\__mp_text_out[117]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[117]$_DFF_P_.QN (\__mp_text_out[117]$_DFF_P_.QN__gold ),
    .\__mp_text_out[117]$_DFF_P_.int_fwire_IQN (\__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[118]$_DFF_P_.CLK (\__mp_text_out[118]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[118]$_DFF_P_.QN (\__mp_text_out[118]$_DFF_P_.QN__gold ),
    .\__mp_text_out[118]$_DFF_P_.int_fwire_IQN (\__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[119]$_DFF_P_.CLK (\__mp_text_out[119]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[119]$_DFF_P_.QN (\__mp_text_out[119]$_DFF_P_.QN__gold ),
    .\__mp_text_out[119]$_DFF_P_.int_fwire_IQN (\__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[11]$_DFF_P_.CLK (\__mp_text_out[11]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[11]$_DFF_P_.QN (\__mp_text_out[11]$_DFF_P_.QN__gold ),
    .\__mp_text_out[11]$_DFF_P_.int_fwire_IQN (\__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[120]$_DFF_P_.CLK (\__mp_text_out[120]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[120]$_DFF_P_.QN (\__mp_text_out[120]$_DFF_P_.QN__gold ),
    .\__mp_text_out[120]$_DFF_P_.int_fwire_IQN (\__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[121]$_DFF_P_.CLK (\__mp_text_out[121]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[121]$_DFF_P_.QN (\__mp_text_out[121]$_DFF_P_.QN__gold ),
    .\__mp_text_out[121]$_DFF_P_.int_fwire_IQN (\__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[122]$_DFF_P_.CLK (\__mp_text_out[122]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[122]$_DFF_P_.QN (\__mp_text_out[122]$_DFF_P_.QN__gold ),
    .\__mp_text_out[122]$_DFF_P_.int_fwire_IQN (\__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[123]$_DFF_P_.CLK (\__mp_text_out[123]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[123]$_DFF_P_.QN (\__mp_text_out[123]$_DFF_P_.QN__gold ),
    .\__mp_text_out[123]$_DFF_P_.int_fwire_IQN (\__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[124]$_DFF_P_.CLK (\__mp_text_out[124]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[124]$_DFF_P_.QN (\__mp_text_out[124]$_DFF_P_.QN__gold ),
    .\__mp_text_out[124]$_DFF_P_.int_fwire_IQN (\__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[125]$_DFF_P_.CLK (\__mp_text_out[125]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[125]$_DFF_P_.QN (\__mp_text_out[125]$_DFF_P_.QN__gold ),
    .\__mp_text_out[125]$_DFF_P_.int_fwire_IQN (\__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[126]$_DFF_P_.CLK (\__mp_text_out[126]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[126]$_DFF_P_.QN (\__mp_text_out[126]$_DFF_P_.QN__gold ),
    .\__mp_text_out[126]$_DFF_P_.int_fwire_IQN (\__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[127]$_DFF_P_.CLK (\__mp_text_out[127]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[127]$_DFF_P_.QN (\__mp_text_out[127]$_DFF_P_.QN__gold ),
    .\__mp_text_out[127]$_DFF_P_.int_fwire_IQN (\__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[12]$_DFF_P_.CLK (\__mp_text_out[12]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[12]$_DFF_P_.QN (\__mp_text_out[12]$_DFF_P_.QN__gold ),
    .\__mp_text_out[12]$_DFF_P_.int_fwire_IQN (\__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[13]$_DFF_P_.CLK (\__mp_text_out[13]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[13]$_DFF_P_.QN (\__mp_text_out[13]$_DFF_P_.QN__gold ),
    .\__mp_text_out[13]$_DFF_P_.int_fwire_IQN (\__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[14]$_DFF_P_.CLK (\__mp_text_out[14]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[14]$_DFF_P_.QN (\__mp_text_out[14]$_DFF_P_.QN__gold ),
    .\__mp_text_out[14]$_DFF_P_.int_fwire_IQN (\__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[15]$_DFF_P_.CLK (\__mp_text_out[15]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[15]$_DFF_P_.QN (\__mp_text_out[15]$_DFF_P_.QN__gold ),
    .\__mp_text_out[15]$_DFF_P_.int_fwire_IQN (\__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[16]$_DFF_P_.CLK (\__mp_text_out[16]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[16]$_DFF_P_.QN (\__mp_text_out[16]$_DFF_P_.QN__gold ),
    .\__mp_text_out[16]$_DFF_P_.int_fwire_IQN (\__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[17]$_DFF_P_.CLK (\__mp_text_out[17]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[17]$_DFF_P_.QN (\__mp_text_out[17]$_DFF_P_.QN__gold ),
    .\__mp_text_out[17]$_DFF_P_.int_fwire_IQN (\__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[18]$_DFF_P_.CLK (\__mp_text_out[18]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[18]$_DFF_P_.QN (\__mp_text_out[18]$_DFF_P_.QN__gold ),
    .\__mp_text_out[18]$_DFF_P_.int_fwire_IQN (\__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[19]$_DFF_P_.CLK (\__mp_text_out[19]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[19]$_DFF_P_.QN (\__mp_text_out[19]$_DFF_P_.QN__gold ),
    .\__mp_text_out[19]$_DFF_P_.int_fwire_IQN (\__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[1]$_DFF_P_.CLK (\__mp_text_out[1]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[1]$_DFF_P_.QN (\__mp_text_out[1]$_DFF_P_.QN__gold ),
    .\__mp_text_out[1]$_DFF_P_.int_fwire_IQN (\__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[20]$_DFF_P_.CLK (\__mp_text_out[20]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[20]$_DFF_P_.QN (\__mp_text_out[20]$_DFF_P_.QN__gold ),
    .\__mp_text_out[20]$_DFF_P_.int_fwire_IQN (\__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[21]$_DFF_P_.CLK (\__mp_text_out[21]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[21]$_DFF_P_.QN (\__mp_text_out[21]$_DFF_P_.QN__gold ),
    .\__mp_text_out[21]$_DFF_P_.int_fwire_IQN (\__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[22]$_DFF_P_.CLK (\__mp_text_out[22]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[22]$_DFF_P_.QN (\__mp_text_out[22]$_DFF_P_.QN__gold ),
    .\__mp_text_out[22]$_DFF_P_.int_fwire_IQN (\__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[23]$_DFF_P_.CLK (\__mp_text_out[23]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[23]$_DFF_P_.QN (\__mp_text_out[23]$_DFF_P_.QN__gold ),
    .\__mp_text_out[23]$_DFF_P_.int_fwire_IQN (\__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[24]$_DFF_P_.CLK (\__mp_text_out[24]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[24]$_DFF_P_.QN (\__mp_text_out[24]$_DFF_P_.QN__gold ),
    .\__mp_text_out[24]$_DFF_P_.int_fwire_IQN (\__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[25]$_DFF_P_.CLK (\__mp_text_out[25]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[25]$_DFF_P_.QN (\__mp_text_out[25]$_DFF_P_.QN__gold ),
    .\__mp_text_out[25]$_DFF_P_.int_fwire_IQN (\__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[26]$_DFF_P_.CLK (\__mp_text_out[26]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[26]$_DFF_P_.QN (\__mp_text_out[26]$_DFF_P_.QN__gold ),
    .\__mp_text_out[26]$_DFF_P_.int_fwire_IQN (\__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[27]$_DFF_P_.CLK (\__mp_text_out[27]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[27]$_DFF_P_.QN (\__mp_text_out[27]$_DFF_P_.QN__gold ),
    .\__mp_text_out[27]$_DFF_P_.int_fwire_IQN (\__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[28]$_DFF_P_.CLK (\__mp_text_out[28]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[28]$_DFF_P_.QN (\__mp_text_out[28]$_DFF_P_.QN__gold ),
    .\__mp_text_out[28]$_DFF_P_.int_fwire_IQN (\__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[29]$_DFF_P_.CLK (\__mp_text_out[29]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[29]$_DFF_P_.QN (\__mp_text_out[29]$_DFF_P_.QN__gold ),
    .\__mp_text_out[29]$_DFF_P_.int_fwire_IQN (\__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[2]$_DFF_P_.CLK (\__mp_text_out[2]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[2]$_DFF_P_.QN (\__mp_text_out[2]$_DFF_P_.QN__gold ),
    .\__mp_text_out[2]$_DFF_P_.int_fwire_IQN (\__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[30]$_DFF_P_.CLK (\__mp_text_out[30]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[30]$_DFF_P_.QN (\__mp_text_out[30]$_DFF_P_.QN__gold ),
    .\__mp_text_out[30]$_DFF_P_.int_fwire_IQN (\__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[31]$_DFF_P_.CLK (\__mp_text_out[31]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[31]$_DFF_P_.QN (\__mp_text_out[31]$_DFF_P_.QN__gold ),
    .\__mp_text_out[31]$_DFF_P_.int_fwire_IQN (\__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[32]$_DFF_P_.CLK (\__mp_text_out[32]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[32]$_DFF_P_.QN (\__mp_text_out[32]$_DFF_P_.QN__gold ),
    .\__mp_text_out[32]$_DFF_P_.int_fwire_IQN (\__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[33]$_DFF_P_.CLK (\__mp_text_out[33]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[33]$_DFF_P_.QN (\__mp_text_out[33]$_DFF_P_.QN__gold ),
    .\__mp_text_out[33]$_DFF_P_.int_fwire_IQN (\__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[34]$_DFF_P_.CLK (\__mp_text_out[34]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[34]$_DFF_P_.QN (\__mp_text_out[34]$_DFF_P_.QN__gold ),
    .\__mp_text_out[34]$_DFF_P_.int_fwire_IQN (\__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[35]$_DFF_P_.CLK (\__mp_text_out[35]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[35]$_DFF_P_.QN (\__mp_text_out[35]$_DFF_P_.QN__gold ),
    .\__mp_text_out[35]$_DFF_P_.int_fwire_IQN (\__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[36]$_DFF_P_.CLK (\__mp_text_out[36]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[36]$_DFF_P_.QN (\__mp_text_out[36]$_DFF_P_.QN__gold ),
    .\__mp_text_out[36]$_DFF_P_.int_fwire_IQN (\__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[37]$_DFF_P_.CLK (\__mp_text_out[37]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[37]$_DFF_P_.QN (\__mp_text_out[37]$_DFF_P_.QN__gold ),
    .\__mp_text_out[37]$_DFF_P_.int_fwire_IQN (\__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[38]$_DFF_P_.CLK (\__mp_text_out[38]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[38]$_DFF_P_.QN (\__mp_text_out[38]$_DFF_P_.QN__gold ),
    .\__mp_text_out[38]$_DFF_P_.int_fwire_IQN (\__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[39]$_DFF_P_.CLK (\__mp_text_out[39]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[39]$_DFF_P_.QN (\__mp_text_out[39]$_DFF_P_.QN__gold ),
    .\__mp_text_out[39]$_DFF_P_.int_fwire_IQN (\__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[3]$_DFF_P_.CLK (\__mp_text_out[3]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[3]$_DFF_P_.QN (\__mp_text_out[3]$_DFF_P_.QN__gold ),
    .\__mp_text_out[3]$_DFF_P_.int_fwire_IQN (\__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[40]$_DFF_P_.CLK (\__mp_text_out[40]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[40]$_DFF_P_.QN (\__mp_text_out[40]$_DFF_P_.QN__gold ),
    .\__mp_text_out[40]$_DFF_P_.int_fwire_IQN (\__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[41]$_DFF_P_.CLK (\__mp_text_out[41]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[41]$_DFF_P_.QN (\__mp_text_out[41]$_DFF_P_.QN__gold ),
    .\__mp_text_out[41]$_DFF_P_.int_fwire_IQN (\__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[42]$_DFF_P_.CLK (\__mp_text_out[42]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[42]$_DFF_P_.QN (\__mp_text_out[42]$_DFF_P_.QN__gold ),
    .\__mp_text_out[42]$_DFF_P_.int_fwire_IQN (\__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[43]$_DFF_P_.CLK (\__mp_text_out[43]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[43]$_DFF_P_.QN (\__mp_text_out[43]$_DFF_P_.QN__gold ),
    .\__mp_text_out[43]$_DFF_P_.int_fwire_IQN (\__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[44]$_DFF_P_.CLK (\__mp_text_out[44]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[44]$_DFF_P_.QN (\__mp_text_out[44]$_DFF_P_.QN__gold ),
    .\__mp_text_out[44]$_DFF_P_.int_fwire_IQN (\__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[45]$_DFF_P_.CLK (\__mp_text_out[45]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[45]$_DFF_P_.QN (\__mp_text_out[45]$_DFF_P_.QN__gold ),
    .\__mp_text_out[45]$_DFF_P_.int_fwire_IQN (\__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[46]$_DFF_P_.CLK (\__mp_text_out[46]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[46]$_DFF_P_.QN (\__mp_text_out[46]$_DFF_P_.QN__gold ),
    .\__mp_text_out[46]$_DFF_P_.int_fwire_IQN (\__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[47]$_DFF_P_.CLK (\__mp_text_out[47]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[47]$_DFF_P_.QN (\__mp_text_out[47]$_DFF_P_.QN__gold ),
    .\__mp_text_out[47]$_DFF_P_.int_fwire_IQN (\__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[48]$_DFF_P_.CLK (\__mp_text_out[48]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[48]$_DFF_P_.QN (\__mp_text_out[48]$_DFF_P_.QN__gold ),
    .\__mp_text_out[48]$_DFF_P_.int_fwire_IQN (\__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[49]$_DFF_P_.CLK (\__mp_text_out[49]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[49]$_DFF_P_.QN (\__mp_text_out[49]$_DFF_P_.QN__gold ),
    .\__mp_text_out[49]$_DFF_P_.int_fwire_IQN (\__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[4]$_DFF_P_.CLK (\__mp_text_out[4]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[4]$_DFF_P_.QN (\__mp_text_out[4]$_DFF_P_.QN__gold ),
    .\__mp_text_out[4]$_DFF_P_.int_fwire_IQN (\__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[50]$_DFF_P_.CLK (\__mp_text_out[50]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[50]$_DFF_P_.QN (\__mp_text_out[50]$_DFF_P_.QN__gold ),
    .\__mp_text_out[50]$_DFF_P_.int_fwire_IQN (\__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[51]$_DFF_P_.CLK (\__mp_text_out[51]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[51]$_DFF_P_.QN (\__mp_text_out[51]$_DFF_P_.QN__gold ),
    .\__mp_text_out[51]$_DFF_P_.int_fwire_IQN (\__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[52]$_DFF_P_.CLK (\__mp_text_out[52]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[52]$_DFF_P_.QN (\__mp_text_out[52]$_DFF_P_.QN__gold ),
    .\__mp_text_out[52]$_DFF_P_.int_fwire_IQN (\__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[53]$_DFF_P_.CLK (\__mp_text_out[53]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[53]$_DFF_P_.QN (\__mp_text_out[53]$_DFF_P_.QN__gold ),
    .\__mp_text_out[53]$_DFF_P_.int_fwire_IQN (\__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[54]$_DFF_P_.CLK (\__mp_text_out[54]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[54]$_DFF_P_.QN (\__mp_text_out[54]$_DFF_P_.QN__gold ),
    .\__mp_text_out[54]$_DFF_P_.int_fwire_IQN (\__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[55]$_DFF_P_.CLK (\__mp_text_out[55]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[55]$_DFF_P_.QN (\__mp_text_out[55]$_DFF_P_.QN__gold ),
    .\__mp_text_out[55]$_DFF_P_.int_fwire_IQN (\__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[56]$_DFF_P_.CLK (\__mp_text_out[56]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[56]$_DFF_P_.QN (\__mp_text_out[56]$_DFF_P_.QN__gold ),
    .\__mp_text_out[56]$_DFF_P_.int_fwire_IQN (\__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[57]$_DFF_P_.CLK (\__mp_text_out[57]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[57]$_DFF_P_.QN (\__mp_text_out[57]$_DFF_P_.QN__gold ),
    .\__mp_text_out[57]$_DFF_P_.int_fwire_IQN (\__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[58]$_DFF_P_.CLK (\__mp_text_out[58]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[58]$_DFF_P_.QN (\__mp_text_out[58]$_DFF_P_.QN__gold ),
    .\__mp_text_out[58]$_DFF_P_.int_fwire_IQN (\__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[59]$_DFF_P_.CLK (\__mp_text_out[59]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[59]$_DFF_P_.QN (\__mp_text_out[59]$_DFF_P_.QN__gold ),
    .\__mp_text_out[59]$_DFF_P_.int_fwire_IQN (\__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[5]$_DFF_P_.CLK (\__mp_text_out[5]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[5]$_DFF_P_.QN (\__mp_text_out[5]$_DFF_P_.QN__gold ),
    .\__mp_text_out[5]$_DFF_P_.int_fwire_IQN (\__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[60]$_DFF_P_.CLK (\__mp_text_out[60]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[60]$_DFF_P_.QN (\__mp_text_out[60]$_DFF_P_.QN__gold ),
    .\__mp_text_out[60]$_DFF_P_.int_fwire_IQN (\__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[61]$_DFF_P_.CLK (\__mp_text_out[61]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[61]$_DFF_P_.QN (\__mp_text_out[61]$_DFF_P_.QN__gold ),
    .\__mp_text_out[61]$_DFF_P_.int_fwire_IQN (\__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[62]$_DFF_P_.CLK (\__mp_text_out[62]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[62]$_DFF_P_.QN (\__mp_text_out[62]$_DFF_P_.QN__gold ),
    .\__mp_text_out[62]$_DFF_P_.int_fwire_IQN (\__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[63]$_DFF_P_.CLK (\__mp_text_out[63]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[63]$_DFF_P_.QN (\__mp_text_out[63]$_DFF_P_.QN__gold ),
    .\__mp_text_out[63]$_DFF_P_.int_fwire_IQN (\__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[64]$_DFF_P_.CLK (\__mp_text_out[64]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[64]$_DFF_P_.QN (\__mp_text_out[64]$_DFF_P_.QN__gold ),
    .\__mp_text_out[64]$_DFF_P_.int_fwire_IQN (\__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[65]$_DFF_P_.CLK (\__mp_text_out[65]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[65]$_DFF_P_.QN (\__mp_text_out[65]$_DFF_P_.QN__gold ),
    .\__mp_text_out[65]$_DFF_P_.int_fwire_IQN (\__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[66]$_DFF_P_.CLK (\__mp_text_out[66]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[66]$_DFF_P_.QN (\__mp_text_out[66]$_DFF_P_.QN__gold ),
    .\__mp_text_out[66]$_DFF_P_.int_fwire_IQN (\__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[67]$_DFF_P_.CLK (\__mp_text_out[67]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[67]$_DFF_P_.QN (\__mp_text_out[67]$_DFF_P_.QN__gold ),
    .\__mp_text_out[67]$_DFF_P_.int_fwire_IQN (\__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[68]$_DFF_P_.CLK (\__mp_text_out[68]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[68]$_DFF_P_.QN (\__mp_text_out[68]$_DFF_P_.QN__gold ),
    .\__mp_text_out[68]$_DFF_P_.int_fwire_IQN (\__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[69]$_DFF_P_.CLK (\__mp_text_out[69]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[69]$_DFF_P_.QN (\__mp_text_out[69]$_DFF_P_.QN__gold ),
    .\__mp_text_out[69]$_DFF_P_.int_fwire_IQN (\__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[6]$_DFF_P_.CLK (\__mp_text_out[6]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[6]$_DFF_P_.QN (\__mp_text_out[6]$_DFF_P_.QN__gold ),
    .\__mp_text_out[6]$_DFF_P_.int_fwire_IQN (\__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[70]$_DFF_P_.CLK (\__mp_text_out[70]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[70]$_DFF_P_.QN (\__mp_text_out[70]$_DFF_P_.QN__gold ),
    .\__mp_text_out[70]$_DFF_P_.int_fwire_IQN (\__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[71]$_DFF_P_.CLK (\__mp_text_out[71]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[71]$_DFF_P_.QN (\__mp_text_out[71]$_DFF_P_.QN__gold ),
    .\__mp_text_out[71]$_DFF_P_.int_fwire_IQN (\__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[72]$_DFF_P_.CLK (\__mp_text_out[72]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[72]$_DFF_P_.QN (\__mp_text_out[72]$_DFF_P_.QN__gold ),
    .\__mp_text_out[72]$_DFF_P_.int_fwire_IQN (\__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[73]$_DFF_P_.CLK (\__mp_text_out[73]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[73]$_DFF_P_.QN (\__mp_text_out[73]$_DFF_P_.QN__gold ),
    .\__mp_text_out[73]$_DFF_P_.int_fwire_IQN (\__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[74]$_DFF_P_.CLK (\__mp_text_out[74]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[74]$_DFF_P_.QN (\__mp_text_out[74]$_DFF_P_.QN__gold ),
    .\__mp_text_out[74]$_DFF_P_.int_fwire_IQN (\__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[75]$_DFF_P_.CLK (\__mp_text_out[75]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[75]$_DFF_P_.QN (\__mp_text_out[75]$_DFF_P_.QN__gold ),
    .\__mp_text_out[75]$_DFF_P_.int_fwire_IQN (\__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[76]$_DFF_P_.CLK (\__mp_text_out[76]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[76]$_DFF_P_.QN (\__mp_text_out[76]$_DFF_P_.QN__gold ),
    .\__mp_text_out[76]$_DFF_P_.int_fwire_IQN (\__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[77]$_DFF_P_.CLK (\__mp_text_out[77]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[77]$_DFF_P_.QN (\__mp_text_out[77]$_DFF_P_.QN__gold ),
    .\__mp_text_out[77]$_DFF_P_.int_fwire_IQN (\__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[78]$_DFF_P_.CLK (\__mp_text_out[78]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[78]$_DFF_P_.QN (\__mp_text_out[78]$_DFF_P_.QN__gold ),
    .\__mp_text_out[78]$_DFF_P_.int_fwire_IQN (\__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[79]$_DFF_P_.CLK (\__mp_text_out[79]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[79]$_DFF_P_.QN (\__mp_text_out[79]$_DFF_P_.QN__gold ),
    .\__mp_text_out[79]$_DFF_P_.int_fwire_IQN (\__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[7]$_DFF_P_.CLK (\__mp_text_out[7]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[7]$_DFF_P_.QN (\__mp_text_out[7]$_DFF_P_.QN__gold ),
    .\__mp_text_out[7]$_DFF_P_.int_fwire_IQN (\__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[80]$_DFF_P_.CLK (\__mp_text_out[80]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[80]$_DFF_P_.QN (\__mp_text_out[80]$_DFF_P_.QN__gold ),
    .\__mp_text_out[80]$_DFF_P_.int_fwire_IQN (\__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[81]$_DFF_P_.CLK (\__mp_text_out[81]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[81]$_DFF_P_.QN (\__mp_text_out[81]$_DFF_P_.QN__gold ),
    .\__mp_text_out[81]$_DFF_P_.int_fwire_IQN (\__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[82]$_DFF_P_.CLK (\__mp_text_out[82]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[82]$_DFF_P_.QN (\__mp_text_out[82]$_DFF_P_.QN__gold ),
    .\__mp_text_out[82]$_DFF_P_.int_fwire_IQN (\__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[83]$_DFF_P_.CLK (\__mp_text_out[83]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[83]$_DFF_P_.QN (\__mp_text_out[83]$_DFF_P_.QN__gold ),
    .\__mp_text_out[83]$_DFF_P_.int_fwire_IQN (\__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[84]$_DFF_P_.CLK (\__mp_text_out[84]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[84]$_DFF_P_.QN (\__mp_text_out[84]$_DFF_P_.QN__gold ),
    .\__mp_text_out[84]$_DFF_P_.int_fwire_IQN (\__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[85]$_DFF_P_.CLK (\__mp_text_out[85]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[85]$_DFF_P_.QN (\__mp_text_out[85]$_DFF_P_.QN__gold ),
    .\__mp_text_out[85]$_DFF_P_.int_fwire_IQN (\__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[86]$_DFF_P_.CLK (\__mp_text_out[86]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[86]$_DFF_P_.QN (\__mp_text_out[86]$_DFF_P_.QN__gold ),
    .\__mp_text_out[86]$_DFF_P_.int_fwire_IQN (\__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[87]$_DFF_P_.CLK (\__mp_text_out[87]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[87]$_DFF_P_.QN (\__mp_text_out[87]$_DFF_P_.QN__gold ),
    .\__mp_text_out[87]$_DFF_P_.int_fwire_IQN (\__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[88]$_DFF_P_.CLK (\__mp_text_out[88]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[88]$_DFF_P_.QN (\__mp_text_out[88]$_DFF_P_.QN__gold ),
    .\__mp_text_out[88]$_DFF_P_.int_fwire_IQN (\__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[89]$_DFF_P_.CLK (\__mp_text_out[89]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[89]$_DFF_P_.QN (\__mp_text_out[89]$_DFF_P_.QN__gold ),
    .\__mp_text_out[89]$_DFF_P_.int_fwire_IQN (\__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[8]$_DFF_P_.CLK (\__mp_text_out[8]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[8]$_DFF_P_.QN (\__mp_text_out[8]$_DFF_P_.QN__gold ),
    .\__mp_text_out[8]$_DFF_P_.int_fwire_IQN (\__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[90]$_DFF_P_.CLK (\__mp_text_out[90]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[90]$_DFF_P_.QN (\__mp_text_out[90]$_DFF_P_.QN__gold ),
    .\__mp_text_out[90]$_DFF_P_.int_fwire_IQN (\__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[91]$_DFF_P_.CLK (\__mp_text_out[91]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[91]$_DFF_P_.QN (\__mp_text_out[91]$_DFF_P_.QN__gold ),
    .\__mp_text_out[91]$_DFF_P_.int_fwire_IQN (\__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[92]$_DFF_P_.CLK (\__mp_text_out[92]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[92]$_DFF_P_.QN (\__mp_text_out[92]$_DFF_P_.QN__gold ),
    .\__mp_text_out[92]$_DFF_P_.int_fwire_IQN (\__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[93]$_DFF_P_.CLK (\__mp_text_out[93]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[93]$_DFF_P_.QN (\__mp_text_out[93]$_DFF_P_.QN__gold ),
    .\__mp_text_out[93]$_DFF_P_.int_fwire_IQN (\__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[94]$_DFF_P_.CLK (\__mp_text_out[94]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[94]$_DFF_P_.QN (\__mp_text_out[94]$_DFF_P_.QN__gold ),
    .\__mp_text_out[94]$_DFF_P_.int_fwire_IQN (\__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[95]$_DFF_P_.CLK (\__mp_text_out[95]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[95]$_DFF_P_.QN (\__mp_text_out[95]$_DFF_P_.QN__gold ),
    .\__mp_text_out[95]$_DFF_P_.int_fwire_IQN (\__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[96]$_DFF_P_.CLK (\__mp_text_out[96]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[96]$_DFF_P_.QN (\__mp_text_out[96]$_DFF_P_.QN__gold ),
    .\__mp_text_out[96]$_DFF_P_.int_fwire_IQN (\__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[97]$_DFF_P_.CLK (\__mp_text_out[97]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[97]$_DFF_P_.QN (\__mp_text_out[97]$_DFF_P_.QN__gold ),
    .\__mp_text_out[97]$_DFF_P_.int_fwire_IQN (\__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[98]$_DFF_P_.CLK (\__mp_text_out[98]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[98]$_DFF_P_.QN (\__mp_text_out[98]$_DFF_P_.QN__gold ),
    .\__mp_text_out[98]$_DFF_P_.int_fwire_IQN (\__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[99]$_DFF_P_.CLK (\__mp_text_out[99]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[99]$_DFF_P_.QN (\__mp_text_out[99]$_DFF_P_.QN__gold ),
    .\__mp_text_out[99]$_DFF_P_.int_fwire_IQN (\__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_text_out[9]$_DFF_P_.CLK (\__mp_text_out[9]$_DFF_P_.CLK__gold ),
    .\__mp_text_out[9]$_DFF_P_.QN (\__mp_text_out[9]$_DFF_P_.QN__gold ),
    .\__mp_text_out[9]$_DFF_P_.int_fwire_IQN (\__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gold ),
    .\__mp_u0.r0.out[24]$_SDFF_PP1_.CLK (\__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gold ),
    .\__mp_u0.r0.out[25]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.out[26]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.out[27]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.out[28]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.out[29]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.out[30]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.out[31]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gold ),
    .\__mp_u0.u0.d[0]$_DFF_P_.CLK (\__mp_u0.u0.d[0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u0.d[1]$_DFF_P_.CLK (\__mp_u0.u0.d[1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u0.d[2]$_DFF_P_.CLK (\__mp_u0.u0.d[2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u0.d[3]$_DFF_P_.CLK (\__mp_u0.u0.d[3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u0.d[4]$_DFF_P_.CLK (\__mp_u0.u0.d[4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u0.d[5]$_DFF_P_.CLK (\__mp_u0.u0.d[5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u0.d[6]$_DFF_P_.CLK (\__mp_u0.u0.d[6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u0.d[7]$_DFF_P_.CLK (\__mp_u0.u0.d[7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[0]$_DFF_P_.CLK (\__mp_u0.u1.d[0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[1]$_DFF_P_.CLK (\__mp_u0.u1.d[1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[2]$_DFF_P_.CLK (\__mp_u0.u1.d[2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[3]$_DFF_P_.CLK (\__mp_u0.u1.d[3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[4]$_DFF_P_.CLK (\__mp_u0.u1.d[4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[5]$_DFF_P_.CLK (\__mp_u0.u1.d[5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[6]$_DFF_P_.CLK (\__mp_u0.u1.d[6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u1.d[7]$_DFF_P_.CLK (\__mp_u0.u1.d[7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[0]$_DFF_P_.CLK (\__mp_u0.u2.d[0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[1]$_DFF_P_.CLK (\__mp_u0.u2.d[1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[2]$_DFF_P_.CLK (\__mp_u0.u2.d[2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[3]$_DFF_P_.CLK (\__mp_u0.u2.d[3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[4]$_DFF_P_.CLK (\__mp_u0.u2.d[4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[5]$_DFF_P_.CLK (\__mp_u0.u2.d[5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[6]$_DFF_P_.CLK (\__mp_u0.u2.d[6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u2.d[7]$_DFF_P_.CLK (\__mp_u0.u2.d[7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[0]$_DFF_P_.CLK (\__mp_u0.u3.d[0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[1]$_DFF_P_.CLK (\__mp_u0.u3.d[1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[2]$_DFF_P_.CLK (\__mp_u0.u3.d[2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[3]$_DFF_P_.CLK (\__mp_u0.u3.d[3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[4]$_DFF_P_.CLK (\__mp_u0.u3.d[4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[5]$_DFF_P_.CLK (\__mp_u0.u3.d[5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[6]$_DFF_P_.CLK (\__mp_u0.u3.d[6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.u3.d[7]$_DFF_P_.CLK (\__mp_u0.u3.d[7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][0]$_DFF_P_.CLK (\__mp_u0.w[0][0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][10]$_DFF_P_.CLK (\__mp_u0.w[0][10]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][11]$_DFF_P_.CLK (\__mp_u0.w[0][11]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][12]$_DFF_P_.CLK (\__mp_u0.w[0][12]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][13]$_DFF_P_.CLK (\__mp_u0.w[0][13]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][14]$_DFF_P_.CLK (\__mp_u0.w[0][14]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][15]$_DFF_P_.CLK (\__mp_u0.w[0][15]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][16]$_DFF_P_.CLK (\__mp_u0.w[0][16]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][17]$_DFF_P_.CLK (\__mp_u0.w[0][17]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][18]$_DFF_P_.CLK (\__mp_u0.w[0][18]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][19]$_DFF_P_.CLK (\__mp_u0.w[0][19]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][1]$_DFF_P_.CLK (\__mp_u0.w[0][1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][20]$_DFF_P_.CLK (\__mp_u0.w[0][20]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][21]$_DFF_P_.CLK (\__mp_u0.w[0][21]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][22]$_DFF_P_.CLK (\__mp_u0.w[0][22]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][23]$_DFF_P_.CLK (\__mp_u0.w[0][23]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][24]$_DFF_P_.CLK (\__mp_u0.w[0][24]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][25]$_DFF_P_.CLK (\__mp_u0.w[0][25]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][26]$_DFF_P_.CLK (\__mp_u0.w[0][26]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][27]$_DFF_P_.CLK (\__mp_u0.w[0][27]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][28]$_DFF_P_.CLK (\__mp_u0.w[0][28]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][29]$_DFF_P_.CLK (\__mp_u0.w[0][29]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][2]$_DFF_P_.CLK (\__mp_u0.w[0][2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][30]$_DFF_P_.CLK (\__mp_u0.w[0][30]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][31]$_DFF_P_.CLK (\__mp_u0.w[0][31]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][3]$_DFF_P_.CLK (\__mp_u0.w[0][3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][4]$_DFF_P_.CLK (\__mp_u0.w[0][4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][5]$_DFF_P_.CLK (\__mp_u0.w[0][5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][6]$_DFF_P_.CLK (\__mp_u0.w[0][6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][7]$_DFF_P_.CLK (\__mp_u0.w[0][7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][8]$_DFF_P_.CLK (\__mp_u0.w[0][8]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[0][9]$_DFF_P_.CLK (\__mp_u0.w[0][9]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][0]$_DFF_P_.CLK (\__mp_u0.w[1][0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][10]$_DFF_P_.CLK (\__mp_u0.w[1][10]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][11]$_DFF_P_.CLK (\__mp_u0.w[1][11]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][12]$_DFF_P_.CLK (\__mp_u0.w[1][12]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][13]$_DFF_P_.CLK (\__mp_u0.w[1][13]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][14]$_DFF_P_.CLK (\__mp_u0.w[1][14]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][15]$_DFF_P_.CLK (\__mp_u0.w[1][15]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][16]$_DFF_P_.CLK (\__mp_u0.w[1][16]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][17]$_DFF_P_.CLK (\__mp_u0.w[1][17]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][18]$_DFF_P_.CLK (\__mp_u0.w[1][18]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][19]$_DFF_P_.CLK (\__mp_u0.w[1][19]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][1]$_DFF_P_.CLK (\__mp_u0.w[1][1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][20]$_DFF_P_.CLK (\__mp_u0.w[1][20]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][21]$_DFF_P_.CLK (\__mp_u0.w[1][21]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][22]$_DFF_P_.CLK (\__mp_u0.w[1][22]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][23]$_DFF_P_.CLK (\__mp_u0.w[1][23]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][24]$_DFF_P_.CLK (\__mp_u0.w[1][24]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][25]$_DFF_P_.CLK (\__mp_u0.w[1][25]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][26]$_DFF_P_.CLK (\__mp_u0.w[1][26]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][27]$_DFF_P_.CLK (\__mp_u0.w[1][27]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][28]$_DFF_P_.CLK (\__mp_u0.w[1][28]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][29]$_DFF_P_.CLK (\__mp_u0.w[1][29]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][2]$_DFF_P_.CLK (\__mp_u0.w[1][2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][30]$_DFF_P_.CLK (\__mp_u0.w[1][30]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][31]$_DFF_P_.CLK (\__mp_u0.w[1][31]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][3]$_DFF_P_.CLK (\__mp_u0.w[1][3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][4]$_DFF_P_.CLK (\__mp_u0.w[1][4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][5]$_DFF_P_.CLK (\__mp_u0.w[1][5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][6]$_DFF_P_.CLK (\__mp_u0.w[1][6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][7]$_DFF_P_.CLK (\__mp_u0.w[1][7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][8]$_DFF_P_.CLK (\__mp_u0.w[1][8]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[1][9]$_DFF_P_.CLK (\__mp_u0.w[1][9]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][0]$_DFF_P_.CLK (\__mp_u0.w[2][0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][10]$_DFF_P_.CLK (\__mp_u0.w[2][10]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][11]$_DFF_P_.CLK (\__mp_u0.w[2][11]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][12]$_DFF_P_.CLK (\__mp_u0.w[2][12]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][13]$_DFF_P_.CLK (\__mp_u0.w[2][13]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][14]$_DFF_P_.CLK (\__mp_u0.w[2][14]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][15]$_DFF_P_.CLK (\__mp_u0.w[2][15]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][16]$_DFF_P_.CLK (\__mp_u0.w[2][16]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][17]$_DFF_P_.CLK (\__mp_u0.w[2][17]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][18]$_DFF_P_.CLK (\__mp_u0.w[2][18]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][19]$_DFF_P_.CLK (\__mp_u0.w[2][19]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][1]$_DFF_P_.CLK (\__mp_u0.w[2][1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][20]$_DFF_P_.CLK (\__mp_u0.w[2][20]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][21]$_DFF_P_.CLK (\__mp_u0.w[2][21]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][22]$_DFF_P_.CLK (\__mp_u0.w[2][22]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][23]$_DFF_P_.CLK (\__mp_u0.w[2][23]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][24]$_DFF_P_.CLK (\__mp_u0.w[2][24]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][25]$_DFF_P_.CLK (\__mp_u0.w[2][25]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][26]$_DFF_P_.CLK (\__mp_u0.w[2][26]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][27]$_DFF_P_.CLK (\__mp_u0.w[2][27]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][28]$_DFF_P_.CLK (\__mp_u0.w[2][28]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][29]$_DFF_P_.CLK (\__mp_u0.w[2][29]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][2]$_DFF_P_.CLK (\__mp_u0.w[2][2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][30]$_DFF_P_.CLK (\__mp_u0.w[2][30]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][31]$_DFF_P_.CLK (\__mp_u0.w[2][31]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][3]$_DFF_P_.CLK (\__mp_u0.w[2][3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][4]$_DFF_P_.CLK (\__mp_u0.w[2][4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][5]$_DFF_P_.CLK (\__mp_u0.w[2][5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][6]$_DFF_P_.CLK (\__mp_u0.w[2][6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][7]$_DFF_P_.CLK (\__mp_u0.w[2][7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][8]$_DFF_P_.CLK (\__mp_u0.w[2][8]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[2][9]$_DFF_P_.CLK (\__mp_u0.w[2][9]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][0]$_DFF_P_.CLK (\__mp_u0.w[3][0]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][10]$_DFF_P_.CLK (\__mp_u0.w[3][10]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][11]$_DFF_P_.CLK (\__mp_u0.w[3][11]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][12]$_DFF_P_.CLK (\__mp_u0.w[3][12]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][13]$_DFF_P_.CLK (\__mp_u0.w[3][13]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][14]$_DFF_P_.CLK (\__mp_u0.w[3][14]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][15]$_DFF_P_.CLK (\__mp_u0.w[3][15]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][16]$_DFF_P_.CLK (\__mp_u0.w[3][16]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][17]$_DFF_P_.CLK (\__mp_u0.w[3][17]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][18]$_DFF_P_.CLK (\__mp_u0.w[3][18]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][19]$_DFF_P_.CLK (\__mp_u0.w[3][19]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][1]$_DFF_P_.CLK (\__mp_u0.w[3][1]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][20]$_DFF_P_.CLK (\__mp_u0.w[3][20]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][21]$_DFF_P_.CLK (\__mp_u0.w[3][21]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][22]$_DFF_P_.CLK (\__mp_u0.w[3][22]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][23]$_DFF_P_.CLK (\__mp_u0.w[3][23]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][24]$_DFF_P_.CLK (\__mp_u0.w[3][24]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][25]$_DFF_P_.CLK (\__mp_u0.w[3][25]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][26]$_DFF_P_.CLK (\__mp_u0.w[3][26]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][27]$_DFF_P_.CLK (\__mp_u0.w[3][27]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][28]$_DFF_P_.CLK (\__mp_u0.w[3][28]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][29]$_DFF_P_.CLK (\__mp_u0.w[3][29]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][2]$_DFF_P_.CLK (\__mp_u0.w[3][2]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][30]$_DFF_P_.CLK (\__mp_u0.w[3][30]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][31]$_DFF_P_.CLK (\__mp_u0.w[3][31]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][3]$_DFF_P_.CLK (\__mp_u0.w[3][3]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][4]$_DFF_P_.CLK (\__mp_u0.w[3][4]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][5]$_DFF_P_.CLK (\__mp_u0.w[3][5]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][6]$_DFF_P_.CLK (\__mp_u0.w[3][6]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][7]$_DFF_P_.CLK (\__mp_u0.w[3][7]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][8]$_DFF_P_.CLK (\__mp_u0.w[3][8]$_DFF_P_.CLK__gold ),
    .\__mp_u0.w[3][9]$_DFF_P_.CLK (\__mp_u0.w[3][9]$_DFF_P_.CLK__gold ),
    .\__po_done (\__po_done__gold ),
    .\__po_text_out (\__po_text_out__gold )
  );
  \gate.aes_cipher_top gate (
    .\__pi_clk (\__pi_clk ),
    .\__pi_key (\__pi_key ),
    .\__pi_ld (\__pi_ld ),
    .\__pi_rst (\__pi_rst ),
    .\__pi_text_in (\__pi_text_in ),
`ifdef DIRECT_CROSS_POINTS
`else
`endif
    .\__mp_clkbuf_0_clk.A (\__mp_clkbuf_0_clk.A__gate ),
    .\__mp_clkbuf_0_clk.Y (\__mp_clkbuf_0_clk.Y__gate ),
    .\__mp_clkbuf_2_0_0_clk.A (\__mp_clkbuf_2_0_0_clk.A__gate ),
    .\__mp_clkbuf_2_0_0_clk.Y (\__mp_clkbuf_2_0_0_clk.Y__gate ),
    .\__mp_clkbuf_2_1_0_clk.A (\__mp_clkbuf_2_1_0_clk.A__gate ),
    .\__mp_clkbuf_2_1_0_clk.Y (\__mp_clkbuf_2_1_0_clk.Y__gate ),
    .\__mp_clkbuf_2_2_0_clk.A (\__mp_clkbuf_2_2_0_clk.A__gate ),
    .\__mp_clkbuf_2_2_0_clk.Y (\__mp_clkbuf_2_2_0_clk.Y__gate ),
    .\__mp_clkbuf_2_3_0_clk.A (\__mp_clkbuf_2_3_0_clk.A__gate ),
    .\__mp_clkbuf_2_3_0_clk.Y (\__mp_clkbuf_2_3_0_clk.Y__gate ),
    .\__mp_clkbuf_leaf_0_clk.A (\__mp_clkbuf_leaf_0_clk.A__gate ),
    .\__mp_clkbuf_leaf_0_clk.Y (\__mp_clkbuf_leaf_0_clk.Y__gate ),
    .\__mp_clkbuf_leaf_10_clk.A (\__mp_clkbuf_leaf_10_clk.A__gate ),
    .\__mp_clkbuf_leaf_10_clk.Y (\__mp_clkbuf_leaf_10_clk.Y__gate ),
    .\__mp_clkbuf_leaf_11_clk.A (\__mp_clkbuf_leaf_11_clk.A__gate ),
    .\__mp_clkbuf_leaf_11_clk.Y (\__mp_clkbuf_leaf_11_clk.Y__gate ),
    .\__mp_clkbuf_leaf_12_clk.A (\__mp_clkbuf_leaf_12_clk.A__gate ),
    .\__mp_clkbuf_leaf_12_clk.Y (\__mp_clkbuf_leaf_12_clk.Y__gate ),
    .\__mp_clkbuf_leaf_13_clk.A (\__mp_clkbuf_leaf_13_clk.A__gate ),
    .\__mp_clkbuf_leaf_13_clk.Y (\__mp_clkbuf_leaf_13_clk.Y__gate ),
    .\__mp_clkbuf_leaf_14_clk.A (\__mp_clkbuf_leaf_14_clk.A__gate ),
    .\__mp_clkbuf_leaf_14_clk.Y (\__mp_clkbuf_leaf_14_clk.Y__gate ),
    .\__mp_clkbuf_leaf_15_clk.A (\__mp_clkbuf_leaf_15_clk.A__gate ),
    .\__mp_clkbuf_leaf_15_clk.Y (\__mp_clkbuf_leaf_15_clk.Y__gate ),
    .\__mp_clkbuf_leaf_16_clk.A (\__mp_clkbuf_leaf_16_clk.A__gate ),
    .\__mp_clkbuf_leaf_16_clk.Y (\__mp_clkbuf_leaf_16_clk.Y__gate ),
    .\__mp_clkbuf_leaf_17_clk.A (\__mp_clkbuf_leaf_17_clk.A__gate ),
    .\__mp_clkbuf_leaf_17_clk.Y (\__mp_clkbuf_leaf_17_clk.Y__gate ),
    .\__mp_clkbuf_leaf_18_clk.A (\__mp_clkbuf_leaf_18_clk.A__gate ),
    .\__mp_clkbuf_leaf_18_clk.Y (\__mp_clkbuf_leaf_18_clk.Y__gate ),
    .\__mp_clkbuf_leaf_19_clk.A (\__mp_clkbuf_leaf_19_clk.A__gate ),
    .\__mp_clkbuf_leaf_19_clk.Y (\__mp_clkbuf_leaf_19_clk.Y__gate ),
    .\__mp_clkbuf_leaf_1_clk.A (\__mp_clkbuf_leaf_1_clk.A__gate ),
    .\__mp_clkbuf_leaf_1_clk.Y (\__mp_clkbuf_leaf_1_clk.Y__gate ),
    .\__mp_clkbuf_leaf_20_clk.A (\__mp_clkbuf_leaf_20_clk.A__gate ),
    .\__mp_clkbuf_leaf_20_clk.Y (\__mp_clkbuf_leaf_20_clk.Y__gate ),
    .\__mp_clkbuf_leaf_21_clk.A (\__mp_clkbuf_leaf_21_clk.A__gate ),
    .\__mp_clkbuf_leaf_21_clk.Y (\__mp_clkbuf_leaf_21_clk.Y__gate ),
    .\__mp_clkbuf_leaf_22_clk.A (\__mp_clkbuf_leaf_22_clk.A__gate ),
    .\__mp_clkbuf_leaf_22_clk.Y (\__mp_clkbuf_leaf_22_clk.Y__gate ),
    .\__mp_clkbuf_leaf_23_clk.A (\__mp_clkbuf_leaf_23_clk.A__gate ),
    .\__mp_clkbuf_leaf_23_clk.Y (\__mp_clkbuf_leaf_23_clk.Y__gate ),
    .\__mp_clkbuf_leaf_24_clk.A (\__mp_clkbuf_leaf_24_clk.A__gate ),
    .\__mp_clkbuf_leaf_24_clk.Y (\__mp_clkbuf_leaf_24_clk.Y__gate ),
    .\__mp_clkbuf_leaf_25_clk.A (\__mp_clkbuf_leaf_25_clk.A__gate ),
    .\__mp_clkbuf_leaf_25_clk.Y (\__mp_clkbuf_leaf_25_clk.Y__gate ),
    .\__mp_clkbuf_leaf_26_clk.A (\__mp_clkbuf_leaf_26_clk.A__gate ),
    .\__mp_clkbuf_leaf_26_clk.Y (\__mp_clkbuf_leaf_26_clk.Y__gate ),
    .\__mp_clkbuf_leaf_27_clk.A (\__mp_clkbuf_leaf_27_clk.A__gate ),
    .\__mp_clkbuf_leaf_27_clk.Y (\__mp_clkbuf_leaf_27_clk.Y__gate ),
    .\__mp_clkbuf_leaf_28_clk.A (\__mp_clkbuf_leaf_28_clk.A__gate ),
    .\__mp_clkbuf_leaf_28_clk.Y (\__mp_clkbuf_leaf_28_clk.Y__gate ),
    .\__mp_clkbuf_leaf_29_clk.A (\__mp_clkbuf_leaf_29_clk.A__gate ),
    .\__mp_clkbuf_leaf_29_clk.Y (\__mp_clkbuf_leaf_29_clk.Y__gate ),
    .\__mp_clkbuf_leaf_2_clk.A (\__mp_clkbuf_leaf_2_clk.A__gate ),
    .\__mp_clkbuf_leaf_2_clk.Y (\__mp_clkbuf_leaf_2_clk.Y__gate ),
    .\__mp_clkbuf_leaf_30_clk.A (\__mp_clkbuf_leaf_30_clk.A__gate ),
    .\__mp_clkbuf_leaf_30_clk.Y (\__mp_clkbuf_leaf_30_clk.Y__gate ),
    .\__mp_clkbuf_leaf_31_clk.A (\__mp_clkbuf_leaf_31_clk.A__gate ),
    .\__mp_clkbuf_leaf_31_clk.Y (\__mp_clkbuf_leaf_31_clk.Y__gate ),
    .\__mp_clkbuf_leaf_32_clk.A (\__mp_clkbuf_leaf_32_clk.A__gate ),
    .\__mp_clkbuf_leaf_32_clk.Y (\__mp_clkbuf_leaf_32_clk.Y__gate ),
    .\__mp_clkbuf_leaf_33_clk.A (\__mp_clkbuf_leaf_33_clk.A__gate ),
    .\__mp_clkbuf_leaf_33_clk.Y (\__mp_clkbuf_leaf_33_clk.Y__gate ),
    .\__mp_clkbuf_leaf_3_clk.A (\__mp_clkbuf_leaf_3_clk.A__gate ),
    .\__mp_clkbuf_leaf_3_clk.Y (\__mp_clkbuf_leaf_3_clk.Y__gate ),
    .\__mp_clkbuf_leaf_4_clk.A (\__mp_clkbuf_leaf_4_clk.A__gate ),
    .\__mp_clkbuf_leaf_4_clk.Y (\__mp_clkbuf_leaf_4_clk.Y__gate ),
    .\__mp_clkbuf_leaf_5_clk.A (\__mp_clkbuf_leaf_5_clk.A__gate ),
    .\__mp_clkbuf_leaf_5_clk.Y (\__mp_clkbuf_leaf_5_clk.Y__gate ),
    .\__mp_clkbuf_leaf_6_clk.A (\__mp_clkbuf_leaf_6_clk.A__gate ),
    .\__mp_clkbuf_leaf_6_clk.Y (\__mp_clkbuf_leaf_6_clk.Y__gate ),
    .\__mp_clkbuf_leaf_7_clk.A (\__mp_clkbuf_leaf_7_clk.A__gate ),
    .\__mp_clkbuf_leaf_7_clk.Y (\__mp_clkbuf_leaf_7_clk.Y__gate ),
    .\__mp_clkbuf_leaf_8_clk.A (\__mp_clkbuf_leaf_8_clk.A__gate ),
    .\__mp_clkbuf_leaf_8_clk.Y (\__mp_clkbuf_leaf_8_clk.Y__gate ),
    .\__mp_clkbuf_leaf_9_clk.A (\__mp_clkbuf_leaf_9_clk.A__gate ),
    .\__mp_clkbuf_leaf_9_clk.Y (\__mp_clkbuf_leaf_9_clk.Y__gate ),
    .\__mp_clkload0.A (\__mp_clkload0.A__gate ),
    .\__mp_clkload0.Y (\__mp_clkload0.Y__gate ),
    .\__mp_clkload1.A (\__mp_clkload1.A__gate ),
    .\__mp_clkload10.A (\__mp_clkload10.A__gate ),
    .\__mp_clkload11.A (\__mp_clkload11.A__gate ),
    .\__mp_clkload12.A (\__mp_clkload12.A__gate ),
    .\__mp_clkload13.A (\__mp_clkload13.A__gate ),
    .\__mp_clkload14.A (\__mp_clkload14.A__gate ),
    .\__mp_clkload15.A (\__mp_clkload15.A__gate ),
    .\__mp_clkload16.A (\__mp_clkload16.A__gate ),
    .\__mp_clkload17.A (\__mp_clkload17.A__gate ),
    .\__mp_clkload18.A (\__mp_clkload18.A__gate ),
    .\__mp_clkload18.Y (\__mp_clkload18.Y__gate ),
    .\__mp_clkload19.A (\__mp_clkload19.A__gate ),
    .\__mp_clkload2.A (\__mp_clkload2.A__gate ),
    .\__mp_clkload20.A (\__mp_clkload20.A__gate ),
    .\__mp_clkload21.A (\__mp_clkload21.A__gate ),
    .\__mp_clkload22.A (\__mp_clkload22.A__gate ),
    .\__mp_clkload23.A (\__mp_clkload23.A__gate ),
    .\__mp_clkload24.A (\__mp_clkload24.A__gate ),
    .\__mp_clkload25.A (\__mp_clkload25.A__gate ),
    .\__mp_clkload26.A (\__mp_clkload26.A__gate ),
    .\__mp_clkload27.A (\__mp_clkload27.A__gate ),
    .\__mp_clkload28.A (\__mp_clkload28.A__gate ),
    .\__mp_clkload29.A (\__mp_clkload29.A__gate ),
    .\__mp_clkload3.A (\__mp_clkload3.A__gate ),
    .\__mp_clkload30.A (\__mp_clkload30.A__gate ),
    .\__mp_clkload31.A (\__mp_clkload31.A__gate ),
    .\__mp_clkload31.Y (\__mp_clkload31.Y__gate ),
    .\__mp_clkload32.A (\__mp_clkload32.A__gate ),
    .\__mp_clkload4.A (\__mp_clkload4.A__gate ),
    .\__mp_clkload5.A (\__mp_clkload5.A__gate ),
    .\__mp_clkload6.A (\__mp_clkload6.A__gate ),
    .\__mp_clkload7.A (\__mp_clkload7.A__gate ),
    .\__mp_clkload8.A (\__mp_clkload8.A__gate ),
    .\__mp_clkload9.A (\__mp_clkload9.A__gate ),
    .\__mp_clknet_0_clk (\__mp_clknet_0_clk__gate ),
    .\__mp_clknet_2_0_0_clk (\__mp_clknet_2_0_0_clk__gate ),
    .\__mp_clknet_2_1_0_clk (\__mp_clknet_2_1_0_clk__gate ),
    .\__mp_clknet_2_2_0_clk (\__mp_clknet_2_2_0_clk__gate ),
    .\__mp_clknet_2_3_0_clk (\__mp_clknet_2_3_0_clk__gate ),
    .\__mp_clknet_leaf_0_clk (\__mp_clknet_leaf_0_clk__gate ),
    .\__mp_clknet_leaf_10_clk (\__mp_clknet_leaf_10_clk__gate ),
    .\__mp_clknet_leaf_11_clk (\__mp_clknet_leaf_11_clk__gate ),
    .\__mp_clknet_leaf_12_clk (\__mp_clknet_leaf_12_clk__gate ),
    .\__mp_clknet_leaf_13_clk (\__mp_clknet_leaf_13_clk__gate ),
    .\__mp_clknet_leaf_14_clk (\__mp_clknet_leaf_14_clk__gate ),
    .\__mp_clknet_leaf_15_clk (\__mp_clknet_leaf_15_clk__gate ),
    .\__mp_clknet_leaf_16_clk (\__mp_clknet_leaf_16_clk__gate ),
    .\__mp_clknet_leaf_17_clk (\__mp_clknet_leaf_17_clk__gate ),
    .\__mp_clknet_leaf_18_clk (\__mp_clknet_leaf_18_clk__gate ),
    .\__mp_clknet_leaf_19_clk (\__mp_clknet_leaf_19_clk__gate ),
    .\__mp_clknet_leaf_1_clk (\__mp_clknet_leaf_1_clk__gate ),
    .\__mp_clknet_leaf_20_clk (\__mp_clknet_leaf_20_clk__gate ),
    .\__mp_clknet_leaf_21_clk (\__mp_clknet_leaf_21_clk__gate ),
    .\__mp_clknet_leaf_22_clk (\__mp_clknet_leaf_22_clk__gate ),
    .\__mp_clknet_leaf_23_clk (\__mp_clknet_leaf_23_clk__gate ),
    .\__mp_clknet_leaf_24_clk (\__mp_clknet_leaf_24_clk__gate ),
    .\__mp_clknet_leaf_25_clk (\__mp_clknet_leaf_25_clk__gate ),
    .\__mp_clknet_leaf_26_clk (\__mp_clknet_leaf_26_clk__gate ),
    .\__mp_clknet_leaf_27_clk (\__mp_clknet_leaf_27_clk__gate ),
    .\__mp_clknet_leaf_28_clk (\__mp_clknet_leaf_28_clk__gate ),
    .\__mp_clknet_leaf_29_clk (\__mp_clknet_leaf_29_clk__gate ),
    .\__mp_clknet_leaf_2_clk (\__mp_clknet_leaf_2_clk__gate ),
    .\__mp_clknet_leaf_30_clk (\__mp_clknet_leaf_30_clk__gate ),
    .\__mp_clknet_leaf_31_clk (\__mp_clknet_leaf_31_clk__gate ),
    .\__mp_clknet_leaf_32_clk (\__mp_clknet_leaf_32_clk__gate ),
    .\__mp_clknet_leaf_33_clk (\__mp_clknet_leaf_33_clk__gate ),
    .\__mp_clknet_leaf_3_clk (\__mp_clknet_leaf_3_clk__gate ),
    .\__mp_clknet_leaf_4_clk (\__mp_clknet_leaf_4_clk__gate ),
    .\__mp_clknet_leaf_5_clk (\__mp_clknet_leaf_5_clk__gate ),
    .\__mp_clknet_leaf_6_clk (\__mp_clknet_leaf_6_clk__gate ),
    .\__mp_clknet_leaf_7_clk (\__mp_clknet_leaf_7_clk__gate ),
    .\__mp_clknet_leaf_8_clk (\__mp_clknet_leaf_8_clk__gate ),
    .\__mp_clknet_leaf_9_clk (\__mp_clknet_leaf_9_clk__gate ),
    .\__mp_dcnt[0]$_SDFFE_PN0P_.CLK (\__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gate ),
    .\__mp_dcnt[1]$_SDFFE_PN0P_.CLK (\__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gate ),
    .\__mp_dcnt[2]$_SDFFE_PP0P_.CLK (\__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gate ),
    .\__mp_dcnt[3]$_SDFFE_PN0P_.CLK (\__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gate ),
    .\__mp_done$_DFF_P_.CLK (\__mp_done$_DFF_P_.CLK__gate ),
    .\__mp_done$_DFF_P_.QN (\__mp_done$_DFF_P_.QN__gate ),
    .\__mp_done$_DFF_P_.int_fwire_IQN (\__mp_done$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_input1.A (\__mp_input1.A__gate ),
    .\__mp_input1.Y (\__mp_input1.Y__gate ),
    .\__mp_input10.A (\__mp_input10.A__gate ),
    .\__mp_input10.Y (\__mp_input10.Y__gate ),
    .\__mp_input100.A (\__mp_input100.A__gate ),
    .\__mp_input100.Y (\__mp_input100.Y__gate ),
    .\__mp_input101.A (\__mp_input101.A__gate ),
    .\__mp_input101.Y (\__mp_input101.Y__gate ),
    .\__mp_input102.A (\__mp_input102.A__gate ),
    .\__mp_input102.Y (\__mp_input102.Y__gate ),
    .\__mp_input103.A (\__mp_input103.A__gate ),
    .\__mp_input103.Y (\__mp_input103.Y__gate ),
    .\__mp_input104.A (\__mp_input104.A__gate ),
    .\__mp_input104.Y (\__mp_input104.Y__gate ),
    .\__mp_input105.A (\__mp_input105.A__gate ),
    .\__mp_input105.Y (\__mp_input105.Y__gate ),
    .\__mp_input106.A (\__mp_input106.A__gate ),
    .\__mp_input106.Y (\__mp_input106.Y__gate ),
    .\__mp_input107.A (\__mp_input107.A__gate ),
    .\__mp_input107.Y (\__mp_input107.Y__gate ),
    .\__mp_input108.A (\__mp_input108.A__gate ),
    .\__mp_input108.Y (\__mp_input108.Y__gate ),
    .\__mp_input109.A (\__mp_input109.A__gate ),
    .\__mp_input109.Y (\__mp_input109.Y__gate ),
    .\__mp_input11.A (\__mp_input11.A__gate ),
    .\__mp_input11.Y (\__mp_input11.Y__gate ),
    .\__mp_input110.A (\__mp_input110.A__gate ),
    .\__mp_input110.Y (\__mp_input110.Y__gate ),
    .\__mp_input111.A (\__mp_input111.A__gate ),
    .\__mp_input111.Y (\__mp_input111.Y__gate ),
    .\__mp_input112.A (\__mp_input112.A__gate ),
    .\__mp_input112.Y (\__mp_input112.Y__gate ),
    .\__mp_input113.A (\__mp_input113.A__gate ),
    .\__mp_input113.Y (\__mp_input113.Y__gate ),
    .\__mp_input114.A (\__mp_input114.A__gate ),
    .\__mp_input114.Y (\__mp_input114.Y__gate ),
    .\__mp_input115.A (\__mp_input115.A__gate ),
    .\__mp_input115.Y (\__mp_input115.Y__gate ),
    .\__mp_input116.A (\__mp_input116.A__gate ),
    .\__mp_input116.Y (\__mp_input116.Y__gate ),
    .\__mp_input117.A (\__mp_input117.A__gate ),
    .\__mp_input117.Y (\__mp_input117.Y__gate ),
    .\__mp_input118.A (\__mp_input118.A__gate ),
    .\__mp_input118.Y (\__mp_input118.Y__gate ),
    .\__mp_input119.A (\__mp_input119.A__gate ),
    .\__mp_input119.Y (\__mp_input119.Y__gate ),
    .\__mp_input12.A (\__mp_input12.A__gate ),
    .\__mp_input12.Y (\__mp_input12.Y__gate ),
    .\__mp_input120.A (\__mp_input120.A__gate ),
    .\__mp_input120.Y (\__mp_input120.Y__gate ),
    .\__mp_input121.A (\__mp_input121.A__gate ),
    .\__mp_input121.Y (\__mp_input121.Y__gate ),
    .\__mp_input122.A (\__mp_input122.A__gate ),
    .\__mp_input122.Y (\__mp_input122.Y__gate ),
    .\__mp_input123.A (\__mp_input123.A__gate ),
    .\__mp_input123.Y (\__mp_input123.Y__gate ),
    .\__mp_input124.A (\__mp_input124.A__gate ),
    .\__mp_input124.Y (\__mp_input124.Y__gate ),
    .\__mp_input125.A (\__mp_input125.A__gate ),
    .\__mp_input125.Y (\__mp_input125.Y__gate ),
    .\__mp_input126.A (\__mp_input126.A__gate ),
    .\__mp_input126.Y (\__mp_input126.Y__gate ),
    .\__mp_input127.A (\__mp_input127.A__gate ),
    .\__mp_input127.Y (\__mp_input127.Y__gate ),
    .\__mp_input128.A (\__mp_input128.A__gate ),
    .\__mp_input128.Y (\__mp_input128.Y__gate ),
    .\__mp_input129.A (\__mp_input129.A__gate ),
    .\__mp_input129.Y (\__mp_input129.Y__gate ),
    .\__mp_input13.A (\__mp_input13.A__gate ),
    .\__mp_input13.Y (\__mp_input13.Y__gate ),
    .\__mp_input130.A (\__mp_input130.A__gate ),
    .\__mp_input130.Y (\__mp_input130.Y__gate ),
    .\__mp_input131.A (\__mp_input131.A__gate ),
    .\__mp_input131.Y (\__mp_input131.Y__gate ),
    .\__mp_input132.A (\__mp_input132.A__gate ),
    .\__mp_input132.Y (\__mp_input132.Y__gate ),
    .\__mp_input133.A (\__mp_input133.A__gate ),
    .\__mp_input133.Y (\__mp_input133.Y__gate ),
    .\__mp_input134.A (\__mp_input134.A__gate ),
    .\__mp_input134.Y (\__mp_input134.Y__gate ),
    .\__mp_input135.A (\__mp_input135.A__gate ),
    .\__mp_input135.Y (\__mp_input135.Y__gate ),
    .\__mp_input136.A (\__mp_input136.A__gate ),
    .\__mp_input136.Y (\__mp_input136.Y__gate ),
    .\__mp_input137.A (\__mp_input137.A__gate ),
    .\__mp_input137.Y (\__mp_input137.Y__gate ),
    .\__mp_input138.A (\__mp_input138.A__gate ),
    .\__mp_input138.Y (\__mp_input138.Y__gate ),
    .\__mp_input139.A (\__mp_input139.A__gate ),
    .\__mp_input139.Y (\__mp_input139.Y__gate ),
    .\__mp_input14.A (\__mp_input14.A__gate ),
    .\__mp_input14.Y (\__mp_input14.Y__gate ),
    .\__mp_input140.A (\__mp_input140.A__gate ),
    .\__mp_input140.Y (\__mp_input140.Y__gate ),
    .\__mp_input141.A (\__mp_input141.A__gate ),
    .\__mp_input141.Y (\__mp_input141.Y__gate ),
    .\__mp_input142.A (\__mp_input142.A__gate ),
    .\__mp_input142.Y (\__mp_input142.Y__gate ),
    .\__mp_input143.A (\__mp_input143.A__gate ),
    .\__mp_input143.Y (\__mp_input143.Y__gate ),
    .\__mp_input144.A (\__mp_input144.A__gate ),
    .\__mp_input144.Y (\__mp_input144.Y__gate ),
    .\__mp_input145.A (\__mp_input145.A__gate ),
    .\__mp_input145.Y (\__mp_input145.Y__gate ),
    .\__mp_input146.A (\__mp_input146.A__gate ),
    .\__mp_input146.Y (\__mp_input146.Y__gate ),
    .\__mp_input147.A (\__mp_input147.A__gate ),
    .\__mp_input147.Y (\__mp_input147.Y__gate ),
    .\__mp_input148.A (\__mp_input148.A__gate ),
    .\__mp_input148.Y (\__mp_input148.Y__gate ),
    .\__mp_input149.A (\__mp_input149.A__gate ),
    .\__mp_input149.Y (\__mp_input149.Y__gate ),
    .\__mp_input15.A (\__mp_input15.A__gate ),
    .\__mp_input15.Y (\__mp_input15.Y__gate ),
    .\__mp_input150.A (\__mp_input150.A__gate ),
    .\__mp_input150.Y (\__mp_input150.Y__gate ),
    .\__mp_input151.A (\__mp_input151.A__gate ),
    .\__mp_input151.Y (\__mp_input151.Y__gate ),
    .\__mp_input152.A (\__mp_input152.A__gate ),
    .\__mp_input152.Y (\__mp_input152.Y__gate ),
    .\__mp_input153.A (\__mp_input153.A__gate ),
    .\__mp_input153.Y (\__mp_input153.Y__gate ),
    .\__mp_input154.A (\__mp_input154.A__gate ),
    .\__mp_input154.Y (\__mp_input154.Y__gate ),
    .\__mp_input155.A (\__mp_input155.A__gate ),
    .\__mp_input155.Y (\__mp_input155.Y__gate ),
    .\__mp_input156.A (\__mp_input156.A__gate ),
    .\__mp_input156.Y (\__mp_input156.Y__gate ),
    .\__mp_input157.A (\__mp_input157.A__gate ),
    .\__mp_input157.Y (\__mp_input157.Y__gate ),
    .\__mp_input158.A (\__mp_input158.A__gate ),
    .\__mp_input158.Y (\__mp_input158.Y__gate ),
    .\__mp_input159.A (\__mp_input159.A__gate ),
    .\__mp_input159.Y (\__mp_input159.Y__gate ),
    .\__mp_input16.A (\__mp_input16.A__gate ),
    .\__mp_input16.Y (\__mp_input16.Y__gate ),
    .\__mp_input160.A (\__mp_input160.A__gate ),
    .\__mp_input160.Y (\__mp_input160.Y__gate ),
    .\__mp_input161.A (\__mp_input161.A__gate ),
    .\__mp_input161.Y (\__mp_input161.Y__gate ),
    .\__mp_input162.A (\__mp_input162.A__gate ),
    .\__mp_input162.Y (\__mp_input162.Y__gate ),
    .\__mp_input163.A (\__mp_input163.A__gate ),
    .\__mp_input163.Y (\__mp_input163.Y__gate ),
    .\__mp_input164.A (\__mp_input164.A__gate ),
    .\__mp_input164.Y (\__mp_input164.Y__gate ),
    .\__mp_input165.A (\__mp_input165.A__gate ),
    .\__mp_input165.Y (\__mp_input165.Y__gate ),
    .\__mp_input166.A (\__mp_input166.A__gate ),
    .\__mp_input166.Y (\__mp_input166.Y__gate ),
    .\__mp_input167.A (\__mp_input167.A__gate ),
    .\__mp_input167.Y (\__mp_input167.Y__gate ),
    .\__mp_input168.A (\__mp_input168.A__gate ),
    .\__mp_input168.Y (\__mp_input168.Y__gate ),
    .\__mp_input169.A (\__mp_input169.A__gate ),
    .\__mp_input169.Y (\__mp_input169.Y__gate ),
    .\__mp_input17.A (\__mp_input17.A__gate ),
    .\__mp_input17.Y (\__mp_input17.Y__gate ),
    .\__mp_input170.A (\__mp_input170.A__gate ),
    .\__mp_input170.Y (\__mp_input170.Y__gate ),
    .\__mp_input171.A (\__mp_input171.A__gate ),
    .\__mp_input171.Y (\__mp_input171.Y__gate ),
    .\__mp_input172.A (\__mp_input172.A__gate ),
    .\__mp_input172.Y (\__mp_input172.Y__gate ),
    .\__mp_input173.A (\__mp_input173.A__gate ),
    .\__mp_input173.Y (\__mp_input173.Y__gate ),
    .\__mp_input174.A (\__mp_input174.A__gate ),
    .\__mp_input174.Y (\__mp_input174.Y__gate ),
    .\__mp_input175.A (\__mp_input175.A__gate ),
    .\__mp_input175.Y (\__mp_input175.Y__gate ),
    .\__mp_input176.A (\__mp_input176.A__gate ),
    .\__mp_input176.Y (\__mp_input176.Y__gate ),
    .\__mp_input177.A (\__mp_input177.A__gate ),
    .\__mp_input177.Y (\__mp_input177.Y__gate ),
    .\__mp_input178.A (\__mp_input178.A__gate ),
    .\__mp_input178.Y (\__mp_input178.Y__gate ),
    .\__mp_input179.A (\__mp_input179.A__gate ),
    .\__mp_input179.Y (\__mp_input179.Y__gate ),
    .\__mp_input18.A (\__mp_input18.A__gate ),
    .\__mp_input18.Y (\__mp_input18.Y__gate ),
    .\__mp_input180.A (\__mp_input180.A__gate ),
    .\__mp_input180.Y (\__mp_input180.Y__gate ),
    .\__mp_input181.A (\__mp_input181.A__gate ),
    .\__mp_input181.Y (\__mp_input181.Y__gate ),
    .\__mp_input182.A (\__mp_input182.A__gate ),
    .\__mp_input182.Y (\__mp_input182.Y__gate ),
    .\__mp_input183.A (\__mp_input183.A__gate ),
    .\__mp_input183.Y (\__mp_input183.Y__gate ),
    .\__mp_input184.A (\__mp_input184.A__gate ),
    .\__mp_input184.Y (\__mp_input184.Y__gate ),
    .\__mp_input185.A (\__mp_input185.A__gate ),
    .\__mp_input185.Y (\__mp_input185.Y__gate ),
    .\__mp_input186.A (\__mp_input186.A__gate ),
    .\__mp_input186.Y (\__mp_input186.Y__gate ),
    .\__mp_input187.A (\__mp_input187.A__gate ),
    .\__mp_input187.Y (\__mp_input187.Y__gate ),
    .\__mp_input188.A (\__mp_input188.A__gate ),
    .\__mp_input188.Y (\__mp_input188.Y__gate ),
    .\__mp_input189.A (\__mp_input189.A__gate ),
    .\__mp_input189.Y (\__mp_input189.Y__gate ),
    .\__mp_input19.A (\__mp_input19.A__gate ),
    .\__mp_input19.Y (\__mp_input19.Y__gate ),
    .\__mp_input190.A (\__mp_input190.A__gate ),
    .\__mp_input190.Y (\__mp_input190.Y__gate ),
    .\__mp_input191.A (\__mp_input191.A__gate ),
    .\__mp_input191.Y (\__mp_input191.Y__gate ),
    .\__mp_input192.A (\__mp_input192.A__gate ),
    .\__mp_input192.Y (\__mp_input192.Y__gate ),
    .\__mp_input193.A (\__mp_input193.A__gate ),
    .\__mp_input193.Y (\__mp_input193.Y__gate ),
    .\__mp_input194.A (\__mp_input194.A__gate ),
    .\__mp_input194.Y (\__mp_input194.Y__gate ),
    .\__mp_input195.A (\__mp_input195.A__gate ),
    .\__mp_input195.Y (\__mp_input195.Y__gate ),
    .\__mp_input196.A (\__mp_input196.A__gate ),
    .\__mp_input196.Y (\__mp_input196.Y__gate ),
    .\__mp_input197.A (\__mp_input197.A__gate ),
    .\__mp_input197.Y (\__mp_input197.Y__gate ),
    .\__mp_input198.A (\__mp_input198.A__gate ),
    .\__mp_input198.Y (\__mp_input198.Y__gate ),
    .\__mp_input199.A (\__mp_input199.A__gate ),
    .\__mp_input199.Y (\__mp_input199.Y__gate ),
    .\__mp_input2.A (\__mp_input2.A__gate ),
    .\__mp_input2.Y (\__mp_input2.Y__gate ),
    .\__mp_input20.A (\__mp_input20.A__gate ),
    .\__mp_input20.Y (\__mp_input20.Y__gate ),
    .\__mp_input200.A (\__mp_input200.A__gate ),
    .\__mp_input200.Y (\__mp_input200.Y__gate ),
    .\__mp_input201.A (\__mp_input201.A__gate ),
    .\__mp_input201.Y (\__mp_input201.Y__gate ),
    .\__mp_input202.A (\__mp_input202.A__gate ),
    .\__mp_input202.Y (\__mp_input202.Y__gate ),
    .\__mp_input203.A (\__mp_input203.A__gate ),
    .\__mp_input203.Y (\__mp_input203.Y__gate ),
    .\__mp_input204.A (\__mp_input204.A__gate ),
    .\__mp_input204.Y (\__mp_input204.Y__gate ),
    .\__mp_input205.A (\__mp_input205.A__gate ),
    .\__mp_input205.Y (\__mp_input205.Y__gate ),
    .\__mp_input206.A (\__mp_input206.A__gate ),
    .\__mp_input206.Y (\__mp_input206.Y__gate ),
    .\__mp_input207.A (\__mp_input207.A__gate ),
    .\__mp_input207.Y (\__mp_input207.Y__gate ),
    .\__mp_input208.A (\__mp_input208.A__gate ),
    .\__mp_input208.Y (\__mp_input208.Y__gate ),
    .\__mp_input209.A (\__mp_input209.A__gate ),
    .\__mp_input209.Y (\__mp_input209.Y__gate ),
    .\__mp_input21.A (\__mp_input21.A__gate ),
    .\__mp_input21.Y (\__mp_input21.Y__gate ),
    .\__mp_input210.A (\__mp_input210.A__gate ),
    .\__mp_input210.Y (\__mp_input210.Y__gate ),
    .\__mp_input211.A (\__mp_input211.A__gate ),
    .\__mp_input211.Y (\__mp_input211.Y__gate ),
    .\__mp_input212.A (\__mp_input212.A__gate ),
    .\__mp_input212.Y (\__mp_input212.Y__gate ),
    .\__mp_input213.A (\__mp_input213.A__gate ),
    .\__mp_input213.Y (\__mp_input213.Y__gate ),
    .\__mp_input214.A (\__mp_input214.A__gate ),
    .\__mp_input214.Y (\__mp_input214.Y__gate ),
    .\__mp_input215.A (\__mp_input215.A__gate ),
    .\__mp_input215.Y (\__mp_input215.Y__gate ),
    .\__mp_input216.A (\__mp_input216.A__gate ),
    .\__mp_input216.Y (\__mp_input216.Y__gate ),
    .\__mp_input217.A (\__mp_input217.A__gate ),
    .\__mp_input217.Y (\__mp_input217.Y__gate ),
    .\__mp_input218.A (\__mp_input218.A__gate ),
    .\__mp_input218.Y (\__mp_input218.Y__gate ),
    .\__mp_input219.A (\__mp_input219.A__gate ),
    .\__mp_input219.Y (\__mp_input219.Y__gate ),
    .\__mp_input22.A (\__mp_input22.A__gate ),
    .\__mp_input22.Y (\__mp_input22.Y__gate ),
    .\__mp_input220.A (\__mp_input220.A__gate ),
    .\__mp_input220.Y (\__mp_input220.Y__gate ),
    .\__mp_input221.A (\__mp_input221.A__gate ),
    .\__mp_input221.Y (\__mp_input221.Y__gate ),
    .\__mp_input222.A (\__mp_input222.A__gate ),
    .\__mp_input222.Y (\__mp_input222.Y__gate ),
    .\__mp_input223.A (\__mp_input223.A__gate ),
    .\__mp_input223.Y (\__mp_input223.Y__gate ),
    .\__mp_input224.A (\__mp_input224.A__gate ),
    .\__mp_input224.Y (\__mp_input224.Y__gate ),
    .\__mp_input225.A (\__mp_input225.A__gate ),
    .\__mp_input225.Y (\__mp_input225.Y__gate ),
    .\__mp_input226.A (\__mp_input226.A__gate ),
    .\__mp_input226.Y (\__mp_input226.Y__gate ),
    .\__mp_input227.A (\__mp_input227.A__gate ),
    .\__mp_input227.Y (\__mp_input227.Y__gate ),
    .\__mp_input228.A (\__mp_input228.A__gate ),
    .\__mp_input228.Y (\__mp_input228.Y__gate ),
    .\__mp_input229.A (\__mp_input229.A__gate ),
    .\__mp_input229.Y (\__mp_input229.Y__gate ),
    .\__mp_input23.A (\__mp_input23.A__gate ),
    .\__mp_input23.Y (\__mp_input23.Y__gate ),
    .\__mp_input230.A (\__mp_input230.A__gate ),
    .\__mp_input230.Y (\__mp_input230.Y__gate ),
    .\__mp_input231.A (\__mp_input231.A__gate ),
    .\__mp_input231.Y (\__mp_input231.Y__gate ),
    .\__mp_input232.A (\__mp_input232.A__gate ),
    .\__mp_input232.Y (\__mp_input232.Y__gate ),
    .\__mp_input233.A (\__mp_input233.A__gate ),
    .\__mp_input233.Y (\__mp_input233.Y__gate ),
    .\__mp_input234.A (\__mp_input234.A__gate ),
    .\__mp_input234.Y (\__mp_input234.Y__gate ),
    .\__mp_input235.A (\__mp_input235.A__gate ),
    .\__mp_input235.Y (\__mp_input235.Y__gate ),
    .\__mp_input236.A (\__mp_input236.A__gate ),
    .\__mp_input236.Y (\__mp_input236.Y__gate ),
    .\__mp_input237.A (\__mp_input237.A__gate ),
    .\__mp_input237.Y (\__mp_input237.Y__gate ),
    .\__mp_input238.A (\__mp_input238.A__gate ),
    .\__mp_input238.Y (\__mp_input238.Y__gate ),
    .\__mp_input239.A (\__mp_input239.A__gate ),
    .\__mp_input239.Y (\__mp_input239.Y__gate ),
    .\__mp_input24.A (\__mp_input24.A__gate ),
    .\__mp_input24.Y (\__mp_input24.Y__gate ),
    .\__mp_input240.A (\__mp_input240.A__gate ),
    .\__mp_input240.Y (\__mp_input240.Y__gate ),
    .\__mp_input241.A (\__mp_input241.A__gate ),
    .\__mp_input241.Y (\__mp_input241.Y__gate ),
    .\__mp_input242.A (\__mp_input242.A__gate ),
    .\__mp_input242.Y (\__mp_input242.Y__gate ),
    .\__mp_input243.A (\__mp_input243.A__gate ),
    .\__mp_input243.Y (\__mp_input243.Y__gate ),
    .\__mp_input244.A (\__mp_input244.A__gate ),
    .\__mp_input244.Y (\__mp_input244.Y__gate ),
    .\__mp_input245.A (\__mp_input245.A__gate ),
    .\__mp_input245.Y (\__mp_input245.Y__gate ),
    .\__mp_input246.A (\__mp_input246.A__gate ),
    .\__mp_input246.Y (\__mp_input246.Y__gate ),
    .\__mp_input247.A (\__mp_input247.A__gate ),
    .\__mp_input247.Y (\__mp_input247.Y__gate ),
    .\__mp_input248.A (\__mp_input248.A__gate ),
    .\__mp_input248.Y (\__mp_input248.Y__gate ),
    .\__mp_input249.A (\__mp_input249.A__gate ),
    .\__mp_input249.Y (\__mp_input249.Y__gate ),
    .\__mp_input25.A (\__mp_input25.A__gate ),
    .\__mp_input25.Y (\__mp_input25.Y__gate ),
    .\__mp_input250.A (\__mp_input250.A__gate ),
    .\__mp_input250.Y (\__mp_input250.Y__gate ),
    .\__mp_input251.A (\__mp_input251.A__gate ),
    .\__mp_input251.Y (\__mp_input251.Y__gate ),
    .\__mp_input252.A (\__mp_input252.A__gate ),
    .\__mp_input252.Y (\__mp_input252.Y__gate ),
    .\__mp_input253.A (\__mp_input253.A__gate ),
    .\__mp_input253.Y (\__mp_input253.Y__gate ),
    .\__mp_input254.A (\__mp_input254.A__gate ),
    .\__mp_input254.Y (\__mp_input254.Y__gate ),
    .\__mp_input255.A (\__mp_input255.A__gate ),
    .\__mp_input255.Y (\__mp_input255.Y__gate ),
    .\__mp_input256.A (\__mp_input256.A__gate ),
    .\__mp_input256.Y (\__mp_input256.Y__gate ),
    .\__mp_input257.A (\__mp_input257.A__gate ),
    .\__mp_input257.Y (\__mp_input257.Y__gate ),
    .\__mp_input258.A (\__mp_input258.A__gate ),
    .\__mp_input258.Y (\__mp_input258.Y__gate ),
    .\__mp_input26.A (\__mp_input26.A__gate ),
    .\__mp_input26.Y (\__mp_input26.Y__gate ),
    .\__mp_input27.A (\__mp_input27.A__gate ),
    .\__mp_input27.Y (\__mp_input27.Y__gate ),
    .\__mp_input28.A (\__mp_input28.A__gate ),
    .\__mp_input28.Y (\__mp_input28.Y__gate ),
    .\__mp_input29.A (\__mp_input29.A__gate ),
    .\__mp_input29.Y (\__mp_input29.Y__gate ),
    .\__mp_input3.A (\__mp_input3.A__gate ),
    .\__mp_input3.Y (\__mp_input3.Y__gate ),
    .\__mp_input30.A (\__mp_input30.A__gate ),
    .\__mp_input30.Y (\__mp_input30.Y__gate ),
    .\__mp_input31.A (\__mp_input31.A__gate ),
    .\__mp_input31.Y (\__mp_input31.Y__gate ),
    .\__mp_input32.A (\__mp_input32.A__gate ),
    .\__mp_input32.Y (\__mp_input32.Y__gate ),
    .\__mp_input33.A (\__mp_input33.A__gate ),
    .\__mp_input33.Y (\__mp_input33.Y__gate ),
    .\__mp_input34.A (\__mp_input34.A__gate ),
    .\__mp_input34.Y (\__mp_input34.Y__gate ),
    .\__mp_input35.A (\__mp_input35.A__gate ),
    .\__mp_input35.Y (\__mp_input35.Y__gate ),
    .\__mp_input36.A (\__mp_input36.A__gate ),
    .\__mp_input36.Y (\__mp_input36.Y__gate ),
    .\__mp_input37.A (\__mp_input37.A__gate ),
    .\__mp_input37.Y (\__mp_input37.Y__gate ),
    .\__mp_input38.A (\__mp_input38.A__gate ),
    .\__mp_input38.Y (\__mp_input38.Y__gate ),
    .\__mp_input39.A (\__mp_input39.A__gate ),
    .\__mp_input39.Y (\__mp_input39.Y__gate ),
    .\__mp_input4.A (\__mp_input4.A__gate ),
    .\__mp_input4.Y (\__mp_input4.Y__gate ),
    .\__mp_input40.A (\__mp_input40.A__gate ),
    .\__mp_input40.Y (\__mp_input40.Y__gate ),
    .\__mp_input41.A (\__mp_input41.A__gate ),
    .\__mp_input41.Y (\__mp_input41.Y__gate ),
    .\__mp_input42.A (\__mp_input42.A__gate ),
    .\__mp_input42.Y (\__mp_input42.Y__gate ),
    .\__mp_input43.A (\__mp_input43.A__gate ),
    .\__mp_input43.Y (\__mp_input43.Y__gate ),
    .\__mp_input44.A (\__mp_input44.A__gate ),
    .\__mp_input44.Y (\__mp_input44.Y__gate ),
    .\__mp_input45.A (\__mp_input45.A__gate ),
    .\__mp_input45.Y (\__mp_input45.Y__gate ),
    .\__mp_input46.A (\__mp_input46.A__gate ),
    .\__mp_input46.Y (\__mp_input46.Y__gate ),
    .\__mp_input47.A (\__mp_input47.A__gate ),
    .\__mp_input47.Y (\__mp_input47.Y__gate ),
    .\__mp_input48.A (\__mp_input48.A__gate ),
    .\__mp_input48.Y (\__mp_input48.Y__gate ),
    .\__mp_input49.A (\__mp_input49.A__gate ),
    .\__mp_input49.Y (\__mp_input49.Y__gate ),
    .\__mp_input5.A (\__mp_input5.A__gate ),
    .\__mp_input5.Y (\__mp_input5.Y__gate ),
    .\__mp_input50.A (\__mp_input50.A__gate ),
    .\__mp_input50.Y (\__mp_input50.Y__gate ),
    .\__mp_input51.A (\__mp_input51.A__gate ),
    .\__mp_input51.Y (\__mp_input51.Y__gate ),
    .\__mp_input52.A (\__mp_input52.A__gate ),
    .\__mp_input52.Y (\__mp_input52.Y__gate ),
    .\__mp_input53.A (\__mp_input53.A__gate ),
    .\__mp_input53.Y (\__mp_input53.Y__gate ),
    .\__mp_input54.A (\__mp_input54.A__gate ),
    .\__mp_input54.Y (\__mp_input54.Y__gate ),
    .\__mp_input55.A (\__mp_input55.A__gate ),
    .\__mp_input55.Y (\__mp_input55.Y__gate ),
    .\__mp_input56.A (\__mp_input56.A__gate ),
    .\__mp_input56.Y (\__mp_input56.Y__gate ),
    .\__mp_input57.A (\__mp_input57.A__gate ),
    .\__mp_input57.Y (\__mp_input57.Y__gate ),
    .\__mp_input58.A (\__mp_input58.A__gate ),
    .\__mp_input58.Y (\__mp_input58.Y__gate ),
    .\__mp_input59.A (\__mp_input59.A__gate ),
    .\__mp_input59.Y (\__mp_input59.Y__gate ),
    .\__mp_input6.A (\__mp_input6.A__gate ),
    .\__mp_input6.Y (\__mp_input6.Y__gate ),
    .\__mp_input60.A (\__mp_input60.A__gate ),
    .\__mp_input60.Y (\__mp_input60.Y__gate ),
    .\__mp_input61.A (\__mp_input61.A__gate ),
    .\__mp_input61.Y (\__mp_input61.Y__gate ),
    .\__mp_input62.A (\__mp_input62.A__gate ),
    .\__mp_input62.Y (\__mp_input62.Y__gate ),
    .\__mp_input63.A (\__mp_input63.A__gate ),
    .\__mp_input63.Y (\__mp_input63.Y__gate ),
    .\__mp_input64.A (\__mp_input64.A__gate ),
    .\__mp_input64.Y (\__mp_input64.Y__gate ),
    .\__mp_input65.A (\__mp_input65.A__gate ),
    .\__mp_input65.Y (\__mp_input65.Y__gate ),
    .\__mp_input66.A (\__mp_input66.A__gate ),
    .\__mp_input66.Y (\__mp_input66.Y__gate ),
    .\__mp_input67.A (\__mp_input67.A__gate ),
    .\__mp_input67.Y (\__mp_input67.Y__gate ),
    .\__mp_input68.A (\__mp_input68.A__gate ),
    .\__mp_input68.Y (\__mp_input68.Y__gate ),
    .\__mp_input69.A (\__mp_input69.A__gate ),
    .\__mp_input69.Y (\__mp_input69.Y__gate ),
    .\__mp_input7.A (\__mp_input7.A__gate ),
    .\__mp_input7.Y (\__mp_input7.Y__gate ),
    .\__mp_input70.A (\__mp_input70.A__gate ),
    .\__mp_input70.Y (\__mp_input70.Y__gate ),
    .\__mp_input71.A (\__mp_input71.A__gate ),
    .\__mp_input71.Y (\__mp_input71.Y__gate ),
    .\__mp_input72.A (\__mp_input72.A__gate ),
    .\__mp_input72.Y (\__mp_input72.Y__gate ),
    .\__mp_input73.A (\__mp_input73.A__gate ),
    .\__mp_input73.Y (\__mp_input73.Y__gate ),
    .\__mp_input74.A (\__mp_input74.A__gate ),
    .\__mp_input74.Y (\__mp_input74.Y__gate ),
    .\__mp_input75.A (\__mp_input75.A__gate ),
    .\__mp_input75.Y (\__mp_input75.Y__gate ),
    .\__mp_input76.A (\__mp_input76.A__gate ),
    .\__mp_input76.Y (\__mp_input76.Y__gate ),
    .\__mp_input77.A (\__mp_input77.A__gate ),
    .\__mp_input77.Y (\__mp_input77.Y__gate ),
    .\__mp_input78.A (\__mp_input78.A__gate ),
    .\__mp_input78.Y (\__mp_input78.Y__gate ),
    .\__mp_input79.A (\__mp_input79.A__gate ),
    .\__mp_input79.Y (\__mp_input79.Y__gate ),
    .\__mp_input8.A (\__mp_input8.A__gate ),
    .\__mp_input8.Y (\__mp_input8.Y__gate ),
    .\__mp_input80.A (\__mp_input80.A__gate ),
    .\__mp_input80.Y (\__mp_input80.Y__gate ),
    .\__mp_input81.A (\__mp_input81.A__gate ),
    .\__mp_input81.Y (\__mp_input81.Y__gate ),
    .\__mp_input82.A (\__mp_input82.A__gate ),
    .\__mp_input82.Y (\__mp_input82.Y__gate ),
    .\__mp_input83.A (\__mp_input83.A__gate ),
    .\__mp_input83.Y (\__mp_input83.Y__gate ),
    .\__mp_input84.A (\__mp_input84.A__gate ),
    .\__mp_input84.Y (\__mp_input84.Y__gate ),
    .\__mp_input85.A (\__mp_input85.A__gate ),
    .\__mp_input85.Y (\__mp_input85.Y__gate ),
    .\__mp_input86.A (\__mp_input86.A__gate ),
    .\__mp_input86.Y (\__mp_input86.Y__gate ),
    .\__mp_input87.A (\__mp_input87.A__gate ),
    .\__mp_input87.Y (\__mp_input87.Y__gate ),
    .\__mp_input88.A (\__mp_input88.A__gate ),
    .\__mp_input88.Y (\__mp_input88.Y__gate ),
    .\__mp_input89.A (\__mp_input89.A__gate ),
    .\__mp_input89.Y (\__mp_input89.Y__gate ),
    .\__mp_input9.A (\__mp_input9.A__gate ),
    .\__mp_input9.Y (\__mp_input9.Y__gate ),
    .\__mp_input90.A (\__mp_input90.A__gate ),
    .\__mp_input90.Y (\__mp_input90.Y__gate ),
    .\__mp_input91.A (\__mp_input91.A__gate ),
    .\__mp_input91.Y (\__mp_input91.Y__gate ),
    .\__mp_input92.A (\__mp_input92.A__gate ),
    .\__mp_input92.Y (\__mp_input92.Y__gate ),
    .\__mp_input93.A (\__mp_input93.A__gate ),
    .\__mp_input93.Y (\__mp_input93.Y__gate ),
    .\__mp_input94.A (\__mp_input94.A__gate ),
    .\__mp_input94.Y (\__mp_input94.Y__gate ),
    .\__mp_input95.A (\__mp_input95.A__gate ),
    .\__mp_input95.Y (\__mp_input95.Y__gate ),
    .\__mp_input96.A (\__mp_input96.A__gate ),
    .\__mp_input96.Y (\__mp_input96.Y__gate ),
    .\__mp_input97.A (\__mp_input97.A__gate ),
    .\__mp_input97.Y (\__mp_input97.Y__gate ),
    .\__mp_input98.A (\__mp_input98.A__gate ),
    .\__mp_input98.Y (\__mp_input98.Y__gate ),
    .\__mp_input99.A (\__mp_input99.A__gate ),
    .\__mp_input99.Y (\__mp_input99.Y__gate ),
    .\__mp_ld_r$_DFF_P_.CLK (\__mp_ld_r$_DFF_P_.CLK__gate ),
    .\__mp_ld_r$_DFF_P_.D (\__mp_ld_r$_DFF_P_.D__gate ),
    .\__mp_output259.A (\__mp_output259.A__gate ),
    .\__mp_output259.Y (\__mp_output259.Y__gate ),
    .\__mp_output260.A (\__mp_output260.A__gate ),
    .\__mp_output260.Y (\__mp_output260.Y__gate ),
    .\__mp_output261.A (\__mp_output261.A__gate ),
    .\__mp_output261.Y (\__mp_output261.Y__gate ),
    .\__mp_output262.A (\__mp_output262.A__gate ),
    .\__mp_output262.Y (\__mp_output262.Y__gate ),
    .\__mp_output263.A (\__mp_output263.A__gate ),
    .\__mp_output263.Y (\__mp_output263.Y__gate ),
    .\__mp_output264.A (\__mp_output264.A__gate ),
    .\__mp_output264.Y (\__mp_output264.Y__gate ),
    .\__mp_output265.A (\__mp_output265.A__gate ),
    .\__mp_output265.Y (\__mp_output265.Y__gate ),
    .\__mp_output266.A (\__mp_output266.A__gate ),
    .\__mp_output266.Y (\__mp_output266.Y__gate ),
    .\__mp_output267.A (\__mp_output267.A__gate ),
    .\__mp_output267.Y (\__mp_output267.Y__gate ),
    .\__mp_output268.A (\__mp_output268.A__gate ),
    .\__mp_output268.Y (\__mp_output268.Y__gate ),
    .\__mp_output269.A (\__mp_output269.A__gate ),
    .\__mp_output269.Y (\__mp_output269.Y__gate ),
    .\__mp_output270.A (\__mp_output270.A__gate ),
    .\__mp_output270.Y (\__mp_output270.Y__gate ),
    .\__mp_output271.A (\__mp_output271.A__gate ),
    .\__mp_output271.Y (\__mp_output271.Y__gate ),
    .\__mp_output272.A (\__mp_output272.A__gate ),
    .\__mp_output272.Y (\__mp_output272.Y__gate ),
    .\__mp_output273.A (\__mp_output273.A__gate ),
    .\__mp_output273.Y (\__mp_output273.Y__gate ),
    .\__mp_output274.A (\__mp_output274.A__gate ),
    .\__mp_output274.Y (\__mp_output274.Y__gate ),
    .\__mp_output275.A (\__mp_output275.A__gate ),
    .\__mp_output275.Y (\__mp_output275.Y__gate ),
    .\__mp_output276.A (\__mp_output276.A__gate ),
    .\__mp_output276.Y (\__mp_output276.Y__gate ),
    .\__mp_output277.A (\__mp_output277.A__gate ),
    .\__mp_output277.Y (\__mp_output277.Y__gate ),
    .\__mp_output278.A (\__mp_output278.A__gate ),
    .\__mp_output278.Y (\__mp_output278.Y__gate ),
    .\__mp_output279.A (\__mp_output279.A__gate ),
    .\__mp_output279.Y (\__mp_output279.Y__gate ),
    .\__mp_output280.A (\__mp_output280.A__gate ),
    .\__mp_output280.Y (\__mp_output280.Y__gate ),
    .\__mp_output281.A (\__mp_output281.A__gate ),
    .\__mp_output281.Y (\__mp_output281.Y__gate ),
    .\__mp_output282.A (\__mp_output282.A__gate ),
    .\__mp_output282.Y (\__mp_output282.Y__gate ),
    .\__mp_output283.A (\__mp_output283.A__gate ),
    .\__mp_output283.Y (\__mp_output283.Y__gate ),
    .\__mp_output284.A (\__mp_output284.A__gate ),
    .\__mp_output284.Y (\__mp_output284.Y__gate ),
    .\__mp_output285.A (\__mp_output285.A__gate ),
    .\__mp_output285.Y (\__mp_output285.Y__gate ),
    .\__mp_output286.A (\__mp_output286.A__gate ),
    .\__mp_output286.Y (\__mp_output286.Y__gate ),
    .\__mp_output287.A (\__mp_output287.A__gate ),
    .\__mp_output287.Y (\__mp_output287.Y__gate ),
    .\__mp_output288.A (\__mp_output288.A__gate ),
    .\__mp_output288.Y (\__mp_output288.Y__gate ),
    .\__mp_output289.A (\__mp_output289.A__gate ),
    .\__mp_output289.Y (\__mp_output289.Y__gate ),
    .\__mp_output290.A (\__mp_output290.A__gate ),
    .\__mp_output290.Y (\__mp_output290.Y__gate ),
    .\__mp_output291.A (\__mp_output291.A__gate ),
    .\__mp_output291.Y (\__mp_output291.Y__gate ),
    .\__mp_output292.A (\__mp_output292.A__gate ),
    .\__mp_output292.Y (\__mp_output292.Y__gate ),
    .\__mp_output293.A (\__mp_output293.A__gate ),
    .\__mp_output293.Y (\__mp_output293.Y__gate ),
    .\__mp_output294.A (\__mp_output294.A__gate ),
    .\__mp_output294.Y (\__mp_output294.Y__gate ),
    .\__mp_output295.A (\__mp_output295.A__gate ),
    .\__mp_output295.Y (\__mp_output295.Y__gate ),
    .\__mp_output296.A (\__mp_output296.A__gate ),
    .\__mp_output296.Y (\__mp_output296.Y__gate ),
    .\__mp_output297.A (\__mp_output297.A__gate ),
    .\__mp_output297.Y (\__mp_output297.Y__gate ),
    .\__mp_output298.A (\__mp_output298.A__gate ),
    .\__mp_output298.Y (\__mp_output298.Y__gate ),
    .\__mp_output299.A (\__mp_output299.A__gate ),
    .\__mp_output299.Y (\__mp_output299.Y__gate ),
    .\__mp_output300.A (\__mp_output300.A__gate ),
    .\__mp_output300.Y (\__mp_output300.Y__gate ),
    .\__mp_output301.A (\__mp_output301.A__gate ),
    .\__mp_output301.Y (\__mp_output301.Y__gate ),
    .\__mp_output302.A (\__mp_output302.A__gate ),
    .\__mp_output302.Y (\__mp_output302.Y__gate ),
    .\__mp_output303.A (\__mp_output303.A__gate ),
    .\__mp_output303.Y (\__mp_output303.Y__gate ),
    .\__mp_output304.A (\__mp_output304.A__gate ),
    .\__mp_output304.Y (\__mp_output304.Y__gate ),
    .\__mp_output305.A (\__mp_output305.A__gate ),
    .\__mp_output305.Y (\__mp_output305.Y__gate ),
    .\__mp_output306.A (\__mp_output306.A__gate ),
    .\__mp_output306.Y (\__mp_output306.Y__gate ),
    .\__mp_output307.A (\__mp_output307.A__gate ),
    .\__mp_output307.Y (\__mp_output307.Y__gate ),
    .\__mp_output308.A (\__mp_output308.A__gate ),
    .\__mp_output308.Y (\__mp_output308.Y__gate ),
    .\__mp_output309.A (\__mp_output309.A__gate ),
    .\__mp_output309.Y (\__mp_output309.Y__gate ),
    .\__mp_output310.A (\__mp_output310.A__gate ),
    .\__mp_output310.Y (\__mp_output310.Y__gate ),
    .\__mp_output311.A (\__mp_output311.A__gate ),
    .\__mp_output311.Y (\__mp_output311.Y__gate ),
    .\__mp_output312.A (\__mp_output312.A__gate ),
    .\__mp_output312.Y (\__mp_output312.Y__gate ),
    .\__mp_output313.A (\__mp_output313.A__gate ),
    .\__mp_output313.Y (\__mp_output313.Y__gate ),
    .\__mp_output314.A (\__mp_output314.A__gate ),
    .\__mp_output314.Y (\__mp_output314.Y__gate ),
    .\__mp_output315.A (\__mp_output315.A__gate ),
    .\__mp_output315.Y (\__mp_output315.Y__gate ),
    .\__mp_output316.A (\__mp_output316.A__gate ),
    .\__mp_output316.Y (\__mp_output316.Y__gate ),
    .\__mp_output317.A (\__mp_output317.A__gate ),
    .\__mp_output317.Y (\__mp_output317.Y__gate ),
    .\__mp_output318.A (\__mp_output318.A__gate ),
    .\__mp_output318.Y (\__mp_output318.Y__gate ),
    .\__mp_output319.A (\__mp_output319.A__gate ),
    .\__mp_output319.Y (\__mp_output319.Y__gate ),
    .\__mp_output320.A (\__mp_output320.A__gate ),
    .\__mp_output320.Y (\__mp_output320.Y__gate ),
    .\__mp_output321.A (\__mp_output321.A__gate ),
    .\__mp_output321.Y (\__mp_output321.Y__gate ),
    .\__mp_output322.A (\__mp_output322.A__gate ),
    .\__mp_output322.Y (\__mp_output322.Y__gate ),
    .\__mp_output323.A (\__mp_output323.A__gate ),
    .\__mp_output323.Y (\__mp_output323.Y__gate ),
    .\__mp_output324.A (\__mp_output324.A__gate ),
    .\__mp_output324.Y (\__mp_output324.Y__gate ),
    .\__mp_output325.A (\__mp_output325.A__gate ),
    .\__mp_output325.Y (\__mp_output325.Y__gate ),
    .\__mp_output326.A (\__mp_output326.A__gate ),
    .\__mp_output326.Y (\__mp_output326.Y__gate ),
    .\__mp_output327.A (\__mp_output327.A__gate ),
    .\__mp_output327.Y (\__mp_output327.Y__gate ),
    .\__mp_output328.A (\__mp_output328.A__gate ),
    .\__mp_output328.Y (\__mp_output328.Y__gate ),
    .\__mp_output329.A (\__mp_output329.A__gate ),
    .\__mp_output329.Y (\__mp_output329.Y__gate ),
    .\__mp_output330.A (\__mp_output330.A__gate ),
    .\__mp_output330.Y (\__mp_output330.Y__gate ),
    .\__mp_output331.A (\__mp_output331.A__gate ),
    .\__mp_output331.Y (\__mp_output331.Y__gate ),
    .\__mp_output332.A (\__mp_output332.A__gate ),
    .\__mp_output332.Y (\__mp_output332.Y__gate ),
    .\__mp_output333.A (\__mp_output333.A__gate ),
    .\__mp_output333.Y (\__mp_output333.Y__gate ),
    .\__mp_output334.A (\__mp_output334.A__gate ),
    .\__mp_output334.Y (\__mp_output334.Y__gate ),
    .\__mp_output335.A (\__mp_output335.A__gate ),
    .\__mp_output335.Y (\__mp_output335.Y__gate ),
    .\__mp_output336.A (\__mp_output336.A__gate ),
    .\__mp_output336.Y (\__mp_output336.Y__gate ),
    .\__mp_output337.A (\__mp_output337.A__gate ),
    .\__mp_output337.Y (\__mp_output337.Y__gate ),
    .\__mp_output338.A (\__mp_output338.A__gate ),
    .\__mp_output338.Y (\__mp_output338.Y__gate ),
    .\__mp_output339.A (\__mp_output339.A__gate ),
    .\__mp_output339.Y (\__mp_output339.Y__gate ),
    .\__mp_output340.A (\__mp_output340.A__gate ),
    .\__mp_output340.Y (\__mp_output340.Y__gate ),
    .\__mp_output341.A (\__mp_output341.A__gate ),
    .\__mp_output341.Y (\__mp_output341.Y__gate ),
    .\__mp_output342.A (\__mp_output342.A__gate ),
    .\__mp_output342.Y (\__mp_output342.Y__gate ),
    .\__mp_output343.A (\__mp_output343.A__gate ),
    .\__mp_output343.Y (\__mp_output343.Y__gate ),
    .\__mp_output344.A (\__mp_output344.A__gate ),
    .\__mp_output344.Y (\__mp_output344.Y__gate ),
    .\__mp_output345.A (\__mp_output345.A__gate ),
    .\__mp_output345.Y (\__mp_output345.Y__gate ),
    .\__mp_output346.A (\__mp_output346.A__gate ),
    .\__mp_output346.Y (\__mp_output346.Y__gate ),
    .\__mp_output347.A (\__mp_output347.A__gate ),
    .\__mp_output347.Y (\__mp_output347.Y__gate ),
    .\__mp_output348.A (\__mp_output348.A__gate ),
    .\__mp_output348.Y (\__mp_output348.Y__gate ),
    .\__mp_output349.A (\__mp_output349.A__gate ),
    .\__mp_output349.Y (\__mp_output349.Y__gate ),
    .\__mp_output350.A (\__mp_output350.A__gate ),
    .\__mp_output350.Y (\__mp_output350.Y__gate ),
    .\__mp_output351.A (\__mp_output351.A__gate ),
    .\__mp_output351.Y (\__mp_output351.Y__gate ),
    .\__mp_output352.A (\__mp_output352.A__gate ),
    .\__mp_output352.Y (\__mp_output352.Y__gate ),
    .\__mp_output353.A (\__mp_output353.A__gate ),
    .\__mp_output353.Y (\__mp_output353.Y__gate ),
    .\__mp_output354.A (\__mp_output354.A__gate ),
    .\__mp_output354.Y (\__mp_output354.Y__gate ),
    .\__mp_output355.A (\__mp_output355.A__gate ),
    .\__mp_output355.Y (\__mp_output355.Y__gate ),
    .\__mp_output356.A (\__mp_output356.A__gate ),
    .\__mp_output356.Y (\__mp_output356.Y__gate ),
    .\__mp_output357.A (\__mp_output357.A__gate ),
    .\__mp_output357.Y (\__mp_output357.Y__gate ),
    .\__mp_output358.A (\__mp_output358.A__gate ),
    .\__mp_output358.Y (\__mp_output358.Y__gate ),
    .\__mp_output359.A (\__mp_output359.A__gate ),
    .\__mp_output359.Y (\__mp_output359.Y__gate ),
    .\__mp_output360.A (\__mp_output360.A__gate ),
    .\__mp_output360.Y (\__mp_output360.Y__gate ),
    .\__mp_output361.A (\__mp_output361.A__gate ),
    .\__mp_output361.Y (\__mp_output361.Y__gate ),
    .\__mp_output362.A (\__mp_output362.A__gate ),
    .\__mp_output362.Y (\__mp_output362.Y__gate ),
    .\__mp_output363.A (\__mp_output363.A__gate ),
    .\__mp_output363.Y (\__mp_output363.Y__gate ),
    .\__mp_output364.A (\__mp_output364.A__gate ),
    .\__mp_output364.Y (\__mp_output364.Y__gate ),
    .\__mp_output365.A (\__mp_output365.A__gate ),
    .\__mp_output365.Y (\__mp_output365.Y__gate ),
    .\__mp_output366.A (\__mp_output366.A__gate ),
    .\__mp_output366.Y (\__mp_output366.Y__gate ),
    .\__mp_output367.A (\__mp_output367.A__gate ),
    .\__mp_output367.Y (\__mp_output367.Y__gate ),
    .\__mp_output368.A (\__mp_output368.A__gate ),
    .\__mp_output368.Y (\__mp_output368.Y__gate ),
    .\__mp_output369.A (\__mp_output369.A__gate ),
    .\__mp_output369.Y (\__mp_output369.Y__gate ),
    .\__mp_output370.A (\__mp_output370.A__gate ),
    .\__mp_output370.Y (\__mp_output370.Y__gate ),
    .\__mp_output371.A (\__mp_output371.A__gate ),
    .\__mp_output371.Y (\__mp_output371.Y__gate ),
    .\__mp_output372.A (\__mp_output372.A__gate ),
    .\__mp_output372.Y (\__mp_output372.Y__gate ),
    .\__mp_output373.A (\__mp_output373.A__gate ),
    .\__mp_output373.Y (\__mp_output373.Y__gate ),
    .\__mp_output374.A (\__mp_output374.A__gate ),
    .\__mp_output374.Y (\__mp_output374.Y__gate ),
    .\__mp_output375.A (\__mp_output375.A__gate ),
    .\__mp_output375.Y (\__mp_output375.Y__gate ),
    .\__mp_output376.A (\__mp_output376.A__gate ),
    .\__mp_output376.Y (\__mp_output376.Y__gate ),
    .\__mp_output377.A (\__mp_output377.A__gate ),
    .\__mp_output377.Y (\__mp_output377.Y__gate ),
    .\__mp_output378.A (\__mp_output378.A__gate ),
    .\__mp_output378.Y (\__mp_output378.Y__gate ),
    .\__mp_output379.A (\__mp_output379.A__gate ),
    .\__mp_output379.Y (\__mp_output379.Y__gate ),
    .\__mp_output380.A (\__mp_output380.A__gate ),
    .\__mp_output380.Y (\__mp_output380.Y__gate ),
    .\__mp_output381.A (\__mp_output381.A__gate ),
    .\__mp_output381.Y (\__mp_output381.Y__gate ),
    .\__mp_output382.A (\__mp_output382.A__gate ),
    .\__mp_output382.Y (\__mp_output382.Y__gate ),
    .\__mp_output383.A (\__mp_output383.A__gate ),
    .\__mp_output383.Y (\__mp_output383.Y__gate ),
    .\__mp_output384.A (\__mp_output384.A__gate ),
    .\__mp_output384.Y (\__mp_output384.Y__gate ),
    .\__mp_output385.A (\__mp_output385.A__gate ),
    .\__mp_output385.Y (\__mp_output385.Y__gate ),
    .\__mp_output386.A (\__mp_output386.A__gate ),
    .\__mp_output386.Y (\__mp_output386.Y__gate ),
    .\__mp_output387.A (\__mp_output387.A__gate ),
    .\__mp_output387.Y (\__mp_output387.Y__gate ),
    .\__mp_sa00_sr[0]$_DFF_P_.CLK (\__mp_sa00_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa00_sr[1]$_DFF_P_.CLK (\__mp_sa00_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa00_sr[2]$_DFF_P_.CLK (\__mp_sa00_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa00_sr[3]$_DFF_P_.CLK (\__mp_sa00_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa00_sr[4]$_DFF_P_.CLK (\__mp_sa00_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa00_sr[5]$_DFF_P_.CLK (\__mp_sa00_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa00_sr[6]$_DFF_P_.CLK (\__mp_sa00_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa00_sr[7]$_DFF_P_.CLK (\__mp_sa00_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[0]$_DFF_P_.CLK (\__mp_sa01_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[1]$_DFF_P_.CLK (\__mp_sa01_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[2]$_DFF_P_.CLK (\__mp_sa01_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[3]$_DFF_P_.CLK (\__mp_sa01_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[4]$_DFF_P_.CLK (\__mp_sa01_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[5]$_DFF_P_.CLK (\__mp_sa01_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[6]$_DFF_P_.CLK (\__mp_sa01_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa01_sr[7]$_DFF_P_.CLK (\__mp_sa01_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[0]$_DFF_P_.CLK (\__mp_sa02_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[1]$_DFF_P_.CLK (\__mp_sa02_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[2]$_DFF_P_.CLK (\__mp_sa02_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[3]$_DFF_P_.CLK (\__mp_sa02_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[4]$_DFF_P_.CLK (\__mp_sa02_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[5]$_DFF_P_.CLK (\__mp_sa02_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[6]$_DFF_P_.CLK (\__mp_sa02_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa02_sr[7]$_DFF_P_.CLK (\__mp_sa02_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[0]$_DFF_P_.CLK (\__mp_sa03_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[1]$_DFF_P_.CLK (\__mp_sa03_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[2]$_DFF_P_.CLK (\__mp_sa03_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[3]$_DFF_P_.CLK (\__mp_sa03_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[4]$_DFF_P_.CLK (\__mp_sa03_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[5]$_DFF_P_.CLK (\__mp_sa03_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[6]$_DFF_P_.CLK (\__mp_sa03_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa03_sr[7]$_DFF_P_.CLK (\__mp_sa03_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[0]$_DFF_P_.CLK (\__mp_sa10_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[1]$_DFF_P_.CLK (\__mp_sa10_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[2]$_DFF_P_.CLK (\__mp_sa10_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[3]$_DFF_P_.CLK (\__mp_sa10_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[4]$_DFF_P_.CLK (\__mp_sa10_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[5]$_DFF_P_.CLK (\__mp_sa10_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[6]$_DFF_P_.CLK (\__mp_sa10_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa10_sr[7]$_DFF_P_.CLK (\__mp_sa10_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[0]$_DFF_P_.CLK (\__mp_sa11_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[1]$_DFF_P_.CLK (\__mp_sa11_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[2]$_DFF_P_.CLK (\__mp_sa11_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[3]$_DFF_P_.CLK (\__mp_sa11_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[4]$_DFF_P_.CLK (\__mp_sa11_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[5]$_DFF_P_.CLK (\__mp_sa11_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[6]$_DFF_P_.CLK (\__mp_sa11_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa11_sr[7]$_DFF_P_.CLK (\__mp_sa11_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[0]$_DFF_P_.CLK (\__mp_sa12_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[1]$_DFF_P_.CLK (\__mp_sa12_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[2]$_DFF_P_.CLK (\__mp_sa12_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[3]$_DFF_P_.CLK (\__mp_sa12_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[4]$_DFF_P_.CLK (\__mp_sa12_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[5]$_DFF_P_.CLK (\__mp_sa12_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[6]$_DFF_P_.CLK (\__mp_sa12_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa12_sr[7]$_DFF_P_.CLK (\__mp_sa12_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[0]$_DFF_P_.CLK (\__mp_sa13_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[1]$_DFF_P_.CLK (\__mp_sa13_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[2]$_DFF_P_.CLK (\__mp_sa13_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[3]$_DFF_P_.CLK (\__mp_sa13_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[4]$_DFF_P_.CLK (\__mp_sa13_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[5]$_DFF_P_.CLK (\__mp_sa13_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[6]$_DFF_P_.CLK (\__mp_sa13_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa13_sr[7]$_DFF_P_.CLK (\__mp_sa13_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[0]$_DFF_P_.CLK (\__mp_sa20_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[1]$_DFF_P_.CLK (\__mp_sa20_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[2]$_DFF_P_.CLK (\__mp_sa20_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[3]$_DFF_P_.CLK (\__mp_sa20_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[4]$_DFF_P_.CLK (\__mp_sa20_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[5]$_DFF_P_.CLK (\__mp_sa20_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[6]$_DFF_P_.CLK (\__mp_sa20_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa20_sr[7]$_DFF_P_.CLK (\__mp_sa20_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[0]$_DFF_P_.CLK (\__mp_sa21_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[1]$_DFF_P_.CLK (\__mp_sa21_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[2]$_DFF_P_.CLK (\__mp_sa21_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[3]$_DFF_P_.CLK (\__mp_sa21_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[4]$_DFF_P_.CLK (\__mp_sa21_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[5]$_DFF_P_.CLK (\__mp_sa21_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[6]$_DFF_P_.CLK (\__mp_sa21_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa21_sr[7]$_DFF_P_.CLK (\__mp_sa21_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[0]$_DFF_P_.CLK (\__mp_sa22_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[1]$_DFF_P_.CLK (\__mp_sa22_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[2]$_DFF_P_.CLK (\__mp_sa22_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[3]$_DFF_P_.CLK (\__mp_sa22_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[4]$_DFF_P_.CLK (\__mp_sa22_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[5]$_DFF_P_.CLK (\__mp_sa22_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[6]$_DFF_P_.CLK (\__mp_sa22_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa22_sr[7]$_DFF_P_.CLK (\__mp_sa22_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[0]$_DFF_P_.CLK (\__mp_sa23_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[1]$_DFF_P_.CLK (\__mp_sa23_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[2]$_DFF_P_.CLK (\__mp_sa23_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[3]$_DFF_P_.CLK (\__mp_sa23_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[4]$_DFF_P_.CLK (\__mp_sa23_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[5]$_DFF_P_.CLK (\__mp_sa23_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[6]$_DFF_P_.CLK (\__mp_sa23_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa23_sr[7]$_DFF_P_.CLK (\__mp_sa23_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[0]$_DFF_P_.CLK (\__mp_sa30_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[1]$_DFF_P_.CLK (\__mp_sa30_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[2]$_DFF_P_.CLK (\__mp_sa30_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[3]$_DFF_P_.CLK (\__mp_sa30_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[4]$_DFF_P_.CLK (\__mp_sa30_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[5]$_DFF_P_.CLK (\__mp_sa30_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[6]$_DFF_P_.CLK (\__mp_sa30_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa30_sr[7]$_DFF_P_.CLK (\__mp_sa30_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[0]$_DFF_P_.CLK (\__mp_sa31_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[1]$_DFF_P_.CLK (\__mp_sa31_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[2]$_DFF_P_.CLK (\__mp_sa31_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[3]$_DFF_P_.CLK (\__mp_sa31_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[4]$_DFF_P_.CLK (\__mp_sa31_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[5]$_DFF_P_.CLK (\__mp_sa31_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[6]$_DFF_P_.CLK (\__mp_sa31_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa31_sr[7]$_DFF_P_.CLK (\__mp_sa31_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[0]$_DFF_P_.CLK (\__mp_sa32_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[1]$_DFF_P_.CLK (\__mp_sa32_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[2]$_DFF_P_.CLK (\__mp_sa32_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[3]$_DFF_P_.CLK (\__mp_sa32_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[4]$_DFF_P_.CLK (\__mp_sa32_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[5]$_DFF_P_.CLK (\__mp_sa32_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[6]$_DFF_P_.CLK (\__mp_sa32_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa32_sr[7]$_DFF_P_.CLK (\__mp_sa32_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[0]$_DFF_P_.CLK (\__mp_sa33_sr[0]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[1]$_DFF_P_.CLK (\__mp_sa33_sr[1]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[2]$_DFF_P_.CLK (\__mp_sa33_sr[2]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[3]$_DFF_P_.CLK (\__mp_sa33_sr[3]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[4]$_DFF_P_.CLK (\__mp_sa33_sr[4]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[5]$_DFF_P_.CLK (\__mp_sa33_sr[5]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[6]$_DFF_P_.CLK (\__mp_sa33_sr[6]$_DFF_P_.CLK__gate ),
    .\__mp_sa33_sr[7]$_DFF_P_.CLK (\__mp_sa33_sr[7]$_DFF_P_.CLK__gate ),
    .\__mp_text_in_r[0]$_DFFE_PP_.CLK (\__mp_text_in_r[0]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[100]$_DFFE_PP_.CLK (\__mp_text_in_r[100]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[101]$_DFFE_PP_.CLK (\__mp_text_in_r[101]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[102]$_DFFE_PP_.CLK (\__mp_text_in_r[102]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[103]$_DFFE_PP_.CLK (\__mp_text_in_r[103]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[104]$_DFFE_PP_.CLK (\__mp_text_in_r[104]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[105]$_DFFE_PP_.CLK (\__mp_text_in_r[105]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[106]$_DFFE_PP_.CLK (\__mp_text_in_r[106]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[107]$_DFFE_PP_.CLK (\__mp_text_in_r[107]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[108]$_DFFE_PP_.CLK (\__mp_text_in_r[108]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[109]$_DFFE_PP_.CLK (\__mp_text_in_r[109]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[10]$_DFFE_PP_.CLK (\__mp_text_in_r[10]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[110]$_DFFE_PP_.CLK (\__mp_text_in_r[110]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[111]$_DFFE_PP_.CLK (\__mp_text_in_r[111]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[112]$_DFFE_PP_.CLK (\__mp_text_in_r[112]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[113]$_DFFE_PP_.CLK (\__mp_text_in_r[113]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[114]$_DFFE_PP_.CLK (\__mp_text_in_r[114]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[115]$_DFFE_PP_.CLK (\__mp_text_in_r[115]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[116]$_DFFE_PP_.CLK (\__mp_text_in_r[116]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[117]$_DFFE_PP_.CLK (\__mp_text_in_r[117]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[118]$_DFFE_PP_.CLK (\__mp_text_in_r[118]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[119]$_DFFE_PP_.CLK (\__mp_text_in_r[119]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[11]$_DFFE_PP_.CLK (\__mp_text_in_r[11]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[120]$_DFFE_PP_.CLK (\__mp_text_in_r[120]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[121]$_DFFE_PP_.CLK (\__mp_text_in_r[121]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[122]$_DFFE_PP_.CLK (\__mp_text_in_r[122]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[123]$_DFFE_PP_.CLK (\__mp_text_in_r[123]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[124]$_DFFE_PP_.CLK (\__mp_text_in_r[124]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[125]$_DFFE_PP_.CLK (\__mp_text_in_r[125]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[126]$_DFFE_PP_.CLK (\__mp_text_in_r[126]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[127]$_DFFE_PP_.CLK (\__mp_text_in_r[127]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[12]$_DFFE_PP_.CLK (\__mp_text_in_r[12]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[13]$_DFFE_PP_.CLK (\__mp_text_in_r[13]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[14]$_DFFE_PP_.CLK (\__mp_text_in_r[14]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[15]$_DFFE_PP_.CLK (\__mp_text_in_r[15]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[16]$_DFFE_PP_.CLK (\__mp_text_in_r[16]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[17]$_DFFE_PP_.CLK (\__mp_text_in_r[17]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[18]$_DFFE_PP_.CLK (\__mp_text_in_r[18]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[19]$_DFFE_PP_.CLK (\__mp_text_in_r[19]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[1]$_DFFE_PP_.CLK (\__mp_text_in_r[1]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[20]$_DFFE_PP_.CLK (\__mp_text_in_r[20]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[21]$_DFFE_PP_.CLK (\__mp_text_in_r[21]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[22]$_DFFE_PP_.CLK (\__mp_text_in_r[22]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[23]$_DFFE_PP_.CLK (\__mp_text_in_r[23]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[24]$_DFFE_PP_.CLK (\__mp_text_in_r[24]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[25]$_DFFE_PP_.CLK (\__mp_text_in_r[25]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[26]$_DFFE_PP_.CLK (\__mp_text_in_r[26]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[27]$_DFFE_PP_.CLK (\__mp_text_in_r[27]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[28]$_DFFE_PP_.CLK (\__mp_text_in_r[28]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[29]$_DFFE_PP_.CLK (\__mp_text_in_r[29]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[2]$_DFFE_PP_.CLK (\__mp_text_in_r[2]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[30]$_DFFE_PP_.CLK (\__mp_text_in_r[30]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[31]$_DFFE_PP_.CLK (\__mp_text_in_r[31]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[32]$_DFFE_PP_.CLK (\__mp_text_in_r[32]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[33]$_DFFE_PP_.CLK (\__mp_text_in_r[33]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[34]$_DFFE_PP_.CLK (\__mp_text_in_r[34]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[35]$_DFFE_PP_.CLK (\__mp_text_in_r[35]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[36]$_DFFE_PP_.CLK (\__mp_text_in_r[36]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[37]$_DFFE_PP_.CLK (\__mp_text_in_r[37]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[38]$_DFFE_PP_.CLK (\__mp_text_in_r[38]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[39]$_DFFE_PP_.CLK (\__mp_text_in_r[39]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[3]$_DFFE_PP_.CLK (\__mp_text_in_r[3]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[40]$_DFFE_PP_.CLK (\__mp_text_in_r[40]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[41]$_DFFE_PP_.CLK (\__mp_text_in_r[41]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[42]$_DFFE_PP_.CLK (\__mp_text_in_r[42]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[43]$_DFFE_PP_.CLK (\__mp_text_in_r[43]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[44]$_DFFE_PP_.CLK (\__mp_text_in_r[44]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[45]$_DFFE_PP_.CLK (\__mp_text_in_r[45]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[46]$_DFFE_PP_.CLK (\__mp_text_in_r[46]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[47]$_DFFE_PP_.CLK (\__mp_text_in_r[47]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[48]$_DFFE_PP_.CLK (\__mp_text_in_r[48]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[49]$_DFFE_PP_.CLK (\__mp_text_in_r[49]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[4]$_DFFE_PP_.CLK (\__mp_text_in_r[4]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[50]$_DFFE_PP_.CLK (\__mp_text_in_r[50]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[51]$_DFFE_PP_.CLK (\__mp_text_in_r[51]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[52]$_DFFE_PP_.CLK (\__mp_text_in_r[52]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[53]$_DFFE_PP_.CLK (\__mp_text_in_r[53]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[54]$_DFFE_PP_.CLK (\__mp_text_in_r[54]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[55]$_DFFE_PP_.CLK (\__mp_text_in_r[55]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[56]$_DFFE_PP_.CLK (\__mp_text_in_r[56]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[57]$_DFFE_PP_.CLK (\__mp_text_in_r[57]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[58]$_DFFE_PP_.CLK (\__mp_text_in_r[58]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[59]$_DFFE_PP_.CLK (\__mp_text_in_r[59]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[5]$_DFFE_PP_.CLK (\__mp_text_in_r[5]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[60]$_DFFE_PP_.CLK (\__mp_text_in_r[60]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[61]$_DFFE_PP_.CLK (\__mp_text_in_r[61]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[62]$_DFFE_PP_.CLK (\__mp_text_in_r[62]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[63]$_DFFE_PP_.CLK (\__mp_text_in_r[63]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[64]$_DFFE_PP_.CLK (\__mp_text_in_r[64]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[65]$_DFFE_PP_.CLK (\__mp_text_in_r[65]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[66]$_DFFE_PP_.CLK (\__mp_text_in_r[66]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[67]$_DFFE_PP_.CLK (\__mp_text_in_r[67]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[68]$_DFFE_PP_.CLK (\__mp_text_in_r[68]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[69]$_DFFE_PP_.CLK (\__mp_text_in_r[69]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[6]$_DFFE_PP_.CLK (\__mp_text_in_r[6]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[70]$_DFFE_PP_.CLK (\__mp_text_in_r[70]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[71]$_DFFE_PP_.CLK (\__mp_text_in_r[71]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[72]$_DFFE_PP_.CLK (\__mp_text_in_r[72]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[73]$_DFFE_PP_.CLK (\__mp_text_in_r[73]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[74]$_DFFE_PP_.CLK (\__mp_text_in_r[74]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[75]$_DFFE_PP_.CLK (\__mp_text_in_r[75]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[76]$_DFFE_PP_.CLK (\__mp_text_in_r[76]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[77]$_DFFE_PP_.CLK (\__mp_text_in_r[77]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[78]$_DFFE_PP_.CLK (\__mp_text_in_r[78]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[79]$_DFFE_PP_.CLK (\__mp_text_in_r[79]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[7]$_DFFE_PP_.CLK (\__mp_text_in_r[7]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[80]$_DFFE_PP_.CLK (\__mp_text_in_r[80]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[81]$_DFFE_PP_.CLK (\__mp_text_in_r[81]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[82]$_DFFE_PP_.CLK (\__mp_text_in_r[82]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[83]$_DFFE_PP_.CLK (\__mp_text_in_r[83]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[84]$_DFFE_PP_.CLK (\__mp_text_in_r[84]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[85]$_DFFE_PP_.CLK (\__mp_text_in_r[85]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[86]$_DFFE_PP_.CLK (\__mp_text_in_r[86]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[87]$_DFFE_PP_.CLK (\__mp_text_in_r[87]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[88]$_DFFE_PP_.CLK (\__mp_text_in_r[88]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[89]$_DFFE_PP_.CLK (\__mp_text_in_r[89]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[8]$_DFFE_PP_.CLK (\__mp_text_in_r[8]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[90]$_DFFE_PP_.CLK (\__mp_text_in_r[90]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[91]$_DFFE_PP_.CLK (\__mp_text_in_r[91]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[92]$_DFFE_PP_.CLK (\__mp_text_in_r[92]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[93]$_DFFE_PP_.CLK (\__mp_text_in_r[93]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[94]$_DFFE_PP_.CLK (\__mp_text_in_r[94]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[95]$_DFFE_PP_.CLK (\__mp_text_in_r[95]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[96]$_DFFE_PP_.CLK (\__mp_text_in_r[96]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[97]$_DFFE_PP_.CLK (\__mp_text_in_r[97]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[98]$_DFFE_PP_.CLK (\__mp_text_in_r[98]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[99]$_DFFE_PP_.CLK (\__mp_text_in_r[99]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_in_r[9]$_DFFE_PP_.CLK (\__mp_text_in_r[9]$_DFFE_PP_.CLK__gate ),
    .\__mp_text_out[0]$_DFF_P_.CLK (\__mp_text_out[0]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[0]$_DFF_P_.QN (\__mp_text_out[0]$_DFF_P_.QN__gate ),
    .\__mp_text_out[0]$_DFF_P_.int_fwire_IQN (\__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[100]$_DFF_P_.CLK (\__mp_text_out[100]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[100]$_DFF_P_.QN (\__mp_text_out[100]$_DFF_P_.QN__gate ),
    .\__mp_text_out[100]$_DFF_P_.int_fwire_IQN (\__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[101]$_DFF_P_.CLK (\__mp_text_out[101]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[101]$_DFF_P_.QN (\__mp_text_out[101]$_DFF_P_.QN__gate ),
    .\__mp_text_out[101]$_DFF_P_.int_fwire_IQN (\__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[102]$_DFF_P_.CLK (\__mp_text_out[102]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[102]$_DFF_P_.QN (\__mp_text_out[102]$_DFF_P_.QN__gate ),
    .\__mp_text_out[102]$_DFF_P_.int_fwire_IQN (\__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[103]$_DFF_P_.CLK (\__mp_text_out[103]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[103]$_DFF_P_.QN (\__mp_text_out[103]$_DFF_P_.QN__gate ),
    .\__mp_text_out[103]$_DFF_P_.int_fwire_IQN (\__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[104]$_DFF_P_.CLK (\__mp_text_out[104]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[104]$_DFF_P_.QN (\__mp_text_out[104]$_DFF_P_.QN__gate ),
    .\__mp_text_out[104]$_DFF_P_.int_fwire_IQN (\__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[105]$_DFF_P_.CLK (\__mp_text_out[105]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[105]$_DFF_P_.QN (\__mp_text_out[105]$_DFF_P_.QN__gate ),
    .\__mp_text_out[105]$_DFF_P_.int_fwire_IQN (\__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[106]$_DFF_P_.CLK (\__mp_text_out[106]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[106]$_DFF_P_.QN (\__mp_text_out[106]$_DFF_P_.QN__gate ),
    .\__mp_text_out[106]$_DFF_P_.int_fwire_IQN (\__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[107]$_DFF_P_.CLK (\__mp_text_out[107]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[107]$_DFF_P_.QN (\__mp_text_out[107]$_DFF_P_.QN__gate ),
    .\__mp_text_out[107]$_DFF_P_.int_fwire_IQN (\__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[108]$_DFF_P_.CLK (\__mp_text_out[108]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[108]$_DFF_P_.QN (\__mp_text_out[108]$_DFF_P_.QN__gate ),
    .\__mp_text_out[108]$_DFF_P_.int_fwire_IQN (\__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[109]$_DFF_P_.CLK (\__mp_text_out[109]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[109]$_DFF_P_.QN (\__mp_text_out[109]$_DFF_P_.QN__gate ),
    .\__mp_text_out[109]$_DFF_P_.int_fwire_IQN (\__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[10]$_DFF_P_.CLK (\__mp_text_out[10]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[10]$_DFF_P_.QN (\__mp_text_out[10]$_DFF_P_.QN__gate ),
    .\__mp_text_out[10]$_DFF_P_.int_fwire_IQN (\__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[110]$_DFF_P_.CLK (\__mp_text_out[110]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[110]$_DFF_P_.QN (\__mp_text_out[110]$_DFF_P_.QN__gate ),
    .\__mp_text_out[110]$_DFF_P_.int_fwire_IQN (\__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[111]$_DFF_P_.CLK (\__mp_text_out[111]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[111]$_DFF_P_.QN (\__mp_text_out[111]$_DFF_P_.QN__gate ),
    .\__mp_text_out[111]$_DFF_P_.int_fwire_IQN (\__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[112]$_DFF_P_.CLK (\__mp_text_out[112]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[112]$_DFF_P_.QN (\__mp_text_out[112]$_DFF_P_.QN__gate ),
    .\__mp_text_out[112]$_DFF_P_.int_fwire_IQN (\__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[113]$_DFF_P_.CLK (\__mp_text_out[113]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[113]$_DFF_P_.QN (\__mp_text_out[113]$_DFF_P_.QN__gate ),
    .\__mp_text_out[113]$_DFF_P_.int_fwire_IQN (\__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[114]$_DFF_P_.CLK (\__mp_text_out[114]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[114]$_DFF_P_.QN (\__mp_text_out[114]$_DFF_P_.QN__gate ),
    .\__mp_text_out[114]$_DFF_P_.int_fwire_IQN (\__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[115]$_DFF_P_.CLK (\__mp_text_out[115]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[115]$_DFF_P_.QN (\__mp_text_out[115]$_DFF_P_.QN__gate ),
    .\__mp_text_out[115]$_DFF_P_.int_fwire_IQN (\__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[116]$_DFF_P_.CLK (\__mp_text_out[116]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[116]$_DFF_P_.QN (\__mp_text_out[116]$_DFF_P_.QN__gate ),
    .\__mp_text_out[116]$_DFF_P_.int_fwire_IQN (\__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[117]$_DFF_P_.CLK (\__mp_text_out[117]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[117]$_DFF_P_.QN (\__mp_text_out[117]$_DFF_P_.QN__gate ),
    .\__mp_text_out[117]$_DFF_P_.int_fwire_IQN (\__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[118]$_DFF_P_.CLK (\__mp_text_out[118]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[118]$_DFF_P_.QN (\__mp_text_out[118]$_DFF_P_.QN__gate ),
    .\__mp_text_out[118]$_DFF_P_.int_fwire_IQN (\__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[119]$_DFF_P_.CLK (\__mp_text_out[119]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[119]$_DFF_P_.QN (\__mp_text_out[119]$_DFF_P_.QN__gate ),
    .\__mp_text_out[119]$_DFF_P_.int_fwire_IQN (\__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[11]$_DFF_P_.CLK (\__mp_text_out[11]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[11]$_DFF_P_.QN (\__mp_text_out[11]$_DFF_P_.QN__gate ),
    .\__mp_text_out[11]$_DFF_P_.int_fwire_IQN (\__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[120]$_DFF_P_.CLK (\__mp_text_out[120]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[120]$_DFF_P_.QN (\__mp_text_out[120]$_DFF_P_.QN__gate ),
    .\__mp_text_out[120]$_DFF_P_.int_fwire_IQN (\__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[121]$_DFF_P_.CLK (\__mp_text_out[121]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[121]$_DFF_P_.QN (\__mp_text_out[121]$_DFF_P_.QN__gate ),
    .\__mp_text_out[121]$_DFF_P_.int_fwire_IQN (\__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[122]$_DFF_P_.CLK (\__mp_text_out[122]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[122]$_DFF_P_.QN (\__mp_text_out[122]$_DFF_P_.QN__gate ),
    .\__mp_text_out[122]$_DFF_P_.int_fwire_IQN (\__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[123]$_DFF_P_.CLK (\__mp_text_out[123]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[123]$_DFF_P_.QN (\__mp_text_out[123]$_DFF_P_.QN__gate ),
    .\__mp_text_out[123]$_DFF_P_.int_fwire_IQN (\__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[124]$_DFF_P_.CLK (\__mp_text_out[124]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[124]$_DFF_P_.QN (\__mp_text_out[124]$_DFF_P_.QN__gate ),
    .\__mp_text_out[124]$_DFF_P_.int_fwire_IQN (\__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[125]$_DFF_P_.CLK (\__mp_text_out[125]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[125]$_DFF_P_.QN (\__mp_text_out[125]$_DFF_P_.QN__gate ),
    .\__mp_text_out[125]$_DFF_P_.int_fwire_IQN (\__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[126]$_DFF_P_.CLK (\__mp_text_out[126]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[126]$_DFF_P_.QN (\__mp_text_out[126]$_DFF_P_.QN__gate ),
    .\__mp_text_out[126]$_DFF_P_.int_fwire_IQN (\__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[127]$_DFF_P_.CLK (\__mp_text_out[127]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[127]$_DFF_P_.QN (\__mp_text_out[127]$_DFF_P_.QN__gate ),
    .\__mp_text_out[127]$_DFF_P_.int_fwire_IQN (\__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[12]$_DFF_P_.CLK (\__mp_text_out[12]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[12]$_DFF_P_.QN (\__mp_text_out[12]$_DFF_P_.QN__gate ),
    .\__mp_text_out[12]$_DFF_P_.int_fwire_IQN (\__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[13]$_DFF_P_.CLK (\__mp_text_out[13]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[13]$_DFF_P_.QN (\__mp_text_out[13]$_DFF_P_.QN__gate ),
    .\__mp_text_out[13]$_DFF_P_.int_fwire_IQN (\__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[14]$_DFF_P_.CLK (\__mp_text_out[14]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[14]$_DFF_P_.QN (\__mp_text_out[14]$_DFF_P_.QN__gate ),
    .\__mp_text_out[14]$_DFF_P_.int_fwire_IQN (\__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[15]$_DFF_P_.CLK (\__mp_text_out[15]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[15]$_DFF_P_.QN (\__mp_text_out[15]$_DFF_P_.QN__gate ),
    .\__mp_text_out[15]$_DFF_P_.int_fwire_IQN (\__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[16]$_DFF_P_.CLK (\__mp_text_out[16]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[16]$_DFF_P_.QN (\__mp_text_out[16]$_DFF_P_.QN__gate ),
    .\__mp_text_out[16]$_DFF_P_.int_fwire_IQN (\__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[17]$_DFF_P_.CLK (\__mp_text_out[17]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[17]$_DFF_P_.QN (\__mp_text_out[17]$_DFF_P_.QN__gate ),
    .\__mp_text_out[17]$_DFF_P_.int_fwire_IQN (\__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[18]$_DFF_P_.CLK (\__mp_text_out[18]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[18]$_DFF_P_.QN (\__mp_text_out[18]$_DFF_P_.QN__gate ),
    .\__mp_text_out[18]$_DFF_P_.int_fwire_IQN (\__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[19]$_DFF_P_.CLK (\__mp_text_out[19]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[19]$_DFF_P_.QN (\__mp_text_out[19]$_DFF_P_.QN__gate ),
    .\__mp_text_out[19]$_DFF_P_.int_fwire_IQN (\__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[1]$_DFF_P_.CLK (\__mp_text_out[1]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[1]$_DFF_P_.QN (\__mp_text_out[1]$_DFF_P_.QN__gate ),
    .\__mp_text_out[1]$_DFF_P_.int_fwire_IQN (\__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[20]$_DFF_P_.CLK (\__mp_text_out[20]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[20]$_DFF_P_.QN (\__mp_text_out[20]$_DFF_P_.QN__gate ),
    .\__mp_text_out[20]$_DFF_P_.int_fwire_IQN (\__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[21]$_DFF_P_.CLK (\__mp_text_out[21]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[21]$_DFF_P_.QN (\__mp_text_out[21]$_DFF_P_.QN__gate ),
    .\__mp_text_out[21]$_DFF_P_.int_fwire_IQN (\__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[22]$_DFF_P_.CLK (\__mp_text_out[22]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[22]$_DFF_P_.QN (\__mp_text_out[22]$_DFF_P_.QN__gate ),
    .\__mp_text_out[22]$_DFF_P_.int_fwire_IQN (\__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[23]$_DFF_P_.CLK (\__mp_text_out[23]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[23]$_DFF_P_.QN (\__mp_text_out[23]$_DFF_P_.QN__gate ),
    .\__mp_text_out[23]$_DFF_P_.int_fwire_IQN (\__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[24]$_DFF_P_.CLK (\__mp_text_out[24]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[24]$_DFF_P_.QN (\__mp_text_out[24]$_DFF_P_.QN__gate ),
    .\__mp_text_out[24]$_DFF_P_.int_fwire_IQN (\__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[25]$_DFF_P_.CLK (\__mp_text_out[25]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[25]$_DFF_P_.QN (\__mp_text_out[25]$_DFF_P_.QN__gate ),
    .\__mp_text_out[25]$_DFF_P_.int_fwire_IQN (\__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[26]$_DFF_P_.CLK (\__mp_text_out[26]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[26]$_DFF_P_.QN (\__mp_text_out[26]$_DFF_P_.QN__gate ),
    .\__mp_text_out[26]$_DFF_P_.int_fwire_IQN (\__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[27]$_DFF_P_.CLK (\__mp_text_out[27]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[27]$_DFF_P_.QN (\__mp_text_out[27]$_DFF_P_.QN__gate ),
    .\__mp_text_out[27]$_DFF_P_.int_fwire_IQN (\__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[28]$_DFF_P_.CLK (\__mp_text_out[28]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[28]$_DFF_P_.QN (\__mp_text_out[28]$_DFF_P_.QN__gate ),
    .\__mp_text_out[28]$_DFF_P_.int_fwire_IQN (\__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[29]$_DFF_P_.CLK (\__mp_text_out[29]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[29]$_DFF_P_.QN (\__mp_text_out[29]$_DFF_P_.QN__gate ),
    .\__mp_text_out[29]$_DFF_P_.int_fwire_IQN (\__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[2]$_DFF_P_.CLK (\__mp_text_out[2]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[2]$_DFF_P_.QN (\__mp_text_out[2]$_DFF_P_.QN__gate ),
    .\__mp_text_out[2]$_DFF_P_.int_fwire_IQN (\__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[30]$_DFF_P_.CLK (\__mp_text_out[30]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[30]$_DFF_P_.QN (\__mp_text_out[30]$_DFF_P_.QN__gate ),
    .\__mp_text_out[30]$_DFF_P_.int_fwire_IQN (\__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[31]$_DFF_P_.CLK (\__mp_text_out[31]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[31]$_DFF_P_.QN (\__mp_text_out[31]$_DFF_P_.QN__gate ),
    .\__mp_text_out[31]$_DFF_P_.int_fwire_IQN (\__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[32]$_DFF_P_.CLK (\__mp_text_out[32]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[32]$_DFF_P_.QN (\__mp_text_out[32]$_DFF_P_.QN__gate ),
    .\__mp_text_out[32]$_DFF_P_.int_fwire_IQN (\__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[33]$_DFF_P_.CLK (\__mp_text_out[33]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[33]$_DFF_P_.QN (\__mp_text_out[33]$_DFF_P_.QN__gate ),
    .\__mp_text_out[33]$_DFF_P_.int_fwire_IQN (\__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[34]$_DFF_P_.CLK (\__mp_text_out[34]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[34]$_DFF_P_.QN (\__mp_text_out[34]$_DFF_P_.QN__gate ),
    .\__mp_text_out[34]$_DFF_P_.int_fwire_IQN (\__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[35]$_DFF_P_.CLK (\__mp_text_out[35]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[35]$_DFF_P_.QN (\__mp_text_out[35]$_DFF_P_.QN__gate ),
    .\__mp_text_out[35]$_DFF_P_.int_fwire_IQN (\__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[36]$_DFF_P_.CLK (\__mp_text_out[36]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[36]$_DFF_P_.QN (\__mp_text_out[36]$_DFF_P_.QN__gate ),
    .\__mp_text_out[36]$_DFF_P_.int_fwire_IQN (\__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[37]$_DFF_P_.CLK (\__mp_text_out[37]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[37]$_DFF_P_.QN (\__mp_text_out[37]$_DFF_P_.QN__gate ),
    .\__mp_text_out[37]$_DFF_P_.int_fwire_IQN (\__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[38]$_DFF_P_.CLK (\__mp_text_out[38]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[38]$_DFF_P_.QN (\__mp_text_out[38]$_DFF_P_.QN__gate ),
    .\__mp_text_out[38]$_DFF_P_.int_fwire_IQN (\__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[39]$_DFF_P_.CLK (\__mp_text_out[39]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[39]$_DFF_P_.QN (\__mp_text_out[39]$_DFF_P_.QN__gate ),
    .\__mp_text_out[39]$_DFF_P_.int_fwire_IQN (\__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[3]$_DFF_P_.CLK (\__mp_text_out[3]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[3]$_DFF_P_.QN (\__mp_text_out[3]$_DFF_P_.QN__gate ),
    .\__mp_text_out[3]$_DFF_P_.int_fwire_IQN (\__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[40]$_DFF_P_.CLK (\__mp_text_out[40]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[40]$_DFF_P_.QN (\__mp_text_out[40]$_DFF_P_.QN__gate ),
    .\__mp_text_out[40]$_DFF_P_.int_fwire_IQN (\__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[41]$_DFF_P_.CLK (\__mp_text_out[41]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[41]$_DFF_P_.QN (\__mp_text_out[41]$_DFF_P_.QN__gate ),
    .\__mp_text_out[41]$_DFF_P_.int_fwire_IQN (\__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[42]$_DFF_P_.CLK (\__mp_text_out[42]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[42]$_DFF_P_.QN (\__mp_text_out[42]$_DFF_P_.QN__gate ),
    .\__mp_text_out[42]$_DFF_P_.int_fwire_IQN (\__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[43]$_DFF_P_.CLK (\__mp_text_out[43]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[43]$_DFF_P_.QN (\__mp_text_out[43]$_DFF_P_.QN__gate ),
    .\__mp_text_out[43]$_DFF_P_.int_fwire_IQN (\__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[44]$_DFF_P_.CLK (\__mp_text_out[44]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[44]$_DFF_P_.QN (\__mp_text_out[44]$_DFF_P_.QN__gate ),
    .\__mp_text_out[44]$_DFF_P_.int_fwire_IQN (\__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[45]$_DFF_P_.CLK (\__mp_text_out[45]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[45]$_DFF_P_.QN (\__mp_text_out[45]$_DFF_P_.QN__gate ),
    .\__mp_text_out[45]$_DFF_P_.int_fwire_IQN (\__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[46]$_DFF_P_.CLK (\__mp_text_out[46]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[46]$_DFF_P_.QN (\__mp_text_out[46]$_DFF_P_.QN__gate ),
    .\__mp_text_out[46]$_DFF_P_.int_fwire_IQN (\__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[47]$_DFF_P_.CLK (\__mp_text_out[47]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[47]$_DFF_P_.QN (\__mp_text_out[47]$_DFF_P_.QN__gate ),
    .\__mp_text_out[47]$_DFF_P_.int_fwire_IQN (\__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[48]$_DFF_P_.CLK (\__mp_text_out[48]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[48]$_DFF_P_.QN (\__mp_text_out[48]$_DFF_P_.QN__gate ),
    .\__mp_text_out[48]$_DFF_P_.int_fwire_IQN (\__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[49]$_DFF_P_.CLK (\__mp_text_out[49]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[49]$_DFF_P_.QN (\__mp_text_out[49]$_DFF_P_.QN__gate ),
    .\__mp_text_out[49]$_DFF_P_.int_fwire_IQN (\__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[4]$_DFF_P_.CLK (\__mp_text_out[4]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[4]$_DFF_P_.QN (\__mp_text_out[4]$_DFF_P_.QN__gate ),
    .\__mp_text_out[4]$_DFF_P_.int_fwire_IQN (\__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[50]$_DFF_P_.CLK (\__mp_text_out[50]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[50]$_DFF_P_.QN (\__mp_text_out[50]$_DFF_P_.QN__gate ),
    .\__mp_text_out[50]$_DFF_P_.int_fwire_IQN (\__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[51]$_DFF_P_.CLK (\__mp_text_out[51]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[51]$_DFF_P_.QN (\__mp_text_out[51]$_DFF_P_.QN__gate ),
    .\__mp_text_out[51]$_DFF_P_.int_fwire_IQN (\__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[52]$_DFF_P_.CLK (\__mp_text_out[52]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[52]$_DFF_P_.QN (\__mp_text_out[52]$_DFF_P_.QN__gate ),
    .\__mp_text_out[52]$_DFF_P_.int_fwire_IQN (\__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[53]$_DFF_P_.CLK (\__mp_text_out[53]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[53]$_DFF_P_.QN (\__mp_text_out[53]$_DFF_P_.QN__gate ),
    .\__mp_text_out[53]$_DFF_P_.int_fwire_IQN (\__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[54]$_DFF_P_.CLK (\__mp_text_out[54]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[54]$_DFF_P_.QN (\__mp_text_out[54]$_DFF_P_.QN__gate ),
    .\__mp_text_out[54]$_DFF_P_.int_fwire_IQN (\__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[55]$_DFF_P_.CLK (\__mp_text_out[55]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[55]$_DFF_P_.QN (\__mp_text_out[55]$_DFF_P_.QN__gate ),
    .\__mp_text_out[55]$_DFF_P_.int_fwire_IQN (\__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[56]$_DFF_P_.CLK (\__mp_text_out[56]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[56]$_DFF_P_.QN (\__mp_text_out[56]$_DFF_P_.QN__gate ),
    .\__mp_text_out[56]$_DFF_P_.int_fwire_IQN (\__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[57]$_DFF_P_.CLK (\__mp_text_out[57]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[57]$_DFF_P_.QN (\__mp_text_out[57]$_DFF_P_.QN__gate ),
    .\__mp_text_out[57]$_DFF_P_.int_fwire_IQN (\__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[58]$_DFF_P_.CLK (\__mp_text_out[58]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[58]$_DFF_P_.QN (\__mp_text_out[58]$_DFF_P_.QN__gate ),
    .\__mp_text_out[58]$_DFF_P_.int_fwire_IQN (\__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[59]$_DFF_P_.CLK (\__mp_text_out[59]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[59]$_DFF_P_.QN (\__mp_text_out[59]$_DFF_P_.QN__gate ),
    .\__mp_text_out[59]$_DFF_P_.int_fwire_IQN (\__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[5]$_DFF_P_.CLK (\__mp_text_out[5]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[5]$_DFF_P_.QN (\__mp_text_out[5]$_DFF_P_.QN__gate ),
    .\__mp_text_out[5]$_DFF_P_.int_fwire_IQN (\__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[60]$_DFF_P_.CLK (\__mp_text_out[60]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[60]$_DFF_P_.QN (\__mp_text_out[60]$_DFF_P_.QN__gate ),
    .\__mp_text_out[60]$_DFF_P_.int_fwire_IQN (\__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[61]$_DFF_P_.CLK (\__mp_text_out[61]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[61]$_DFF_P_.QN (\__mp_text_out[61]$_DFF_P_.QN__gate ),
    .\__mp_text_out[61]$_DFF_P_.int_fwire_IQN (\__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[62]$_DFF_P_.CLK (\__mp_text_out[62]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[62]$_DFF_P_.QN (\__mp_text_out[62]$_DFF_P_.QN__gate ),
    .\__mp_text_out[62]$_DFF_P_.int_fwire_IQN (\__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[63]$_DFF_P_.CLK (\__mp_text_out[63]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[63]$_DFF_P_.QN (\__mp_text_out[63]$_DFF_P_.QN__gate ),
    .\__mp_text_out[63]$_DFF_P_.int_fwire_IQN (\__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[64]$_DFF_P_.CLK (\__mp_text_out[64]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[64]$_DFF_P_.QN (\__mp_text_out[64]$_DFF_P_.QN__gate ),
    .\__mp_text_out[64]$_DFF_P_.int_fwire_IQN (\__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[65]$_DFF_P_.CLK (\__mp_text_out[65]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[65]$_DFF_P_.QN (\__mp_text_out[65]$_DFF_P_.QN__gate ),
    .\__mp_text_out[65]$_DFF_P_.int_fwire_IQN (\__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[66]$_DFF_P_.CLK (\__mp_text_out[66]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[66]$_DFF_P_.QN (\__mp_text_out[66]$_DFF_P_.QN__gate ),
    .\__mp_text_out[66]$_DFF_P_.int_fwire_IQN (\__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[67]$_DFF_P_.CLK (\__mp_text_out[67]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[67]$_DFF_P_.QN (\__mp_text_out[67]$_DFF_P_.QN__gate ),
    .\__mp_text_out[67]$_DFF_P_.int_fwire_IQN (\__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[68]$_DFF_P_.CLK (\__mp_text_out[68]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[68]$_DFF_P_.QN (\__mp_text_out[68]$_DFF_P_.QN__gate ),
    .\__mp_text_out[68]$_DFF_P_.int_fwire_IQN (\__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[69]$_DFF_P_.CLK (\__mp_text_out[69]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[69]$_DFF_P_.QN (\__mp_text_out[69]$_DFF_P_.QN__gate ),
    .\__mp_text_out[69]$_DFF_P_.int_fwire_IQN (\__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[6]$_DFF_P_.CLK (\__mp_text_out[6]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[6]$_DFF_P_.QN (\__mp_text_out[6]$_DFF_P_.QN__gate ),
    .\__mp_text_out[6]$_DFF_P_.int_fwire_IQN (\__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[70]$_DFF_P_.CLK (\__mp_text_out[70]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[70]$_DFF_P_.QN (\__mp_text_out[70]$_DFF_P_.QN__gate ),
    .\__mp_text_out[70]$_DFF_P_.int_fwire_IQN (\__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[71]$_DFF_P_.CLK (\__mp_text_out[71]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[71]$_DFF_P_.QN (\__mp_text_out[71]$_DFF_P_.QN__gate ),
    .\__mp_text_out[71]$_DFF_P_.int_fwire_IQN (\__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[72]$_DFF_P_.CLK (\__mp_text_out[72]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[72]$_DFF_P_.QN (\__mp_text_out[72]$_DFF_P_.QN__gate ),
    .\__mp_text_out[72]$_DFF_P_.int_fwire_IQN (\__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[73]$_DFF_P_.CLK (\__mp_text_out[73]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[73]$_DFF_P_.QN (\__mp_text_out[73]$_DFF_P_.QN__gate ),
    .\__mp_text_out[73]$_DFF_P_.int_fwire_IQN (\__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[74]$_DFF_P_.CLK (\__mp_text_out[74]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[74]$_DFF_P_.QN (\__mp_text_out[74]$_DFF_P_.QN__gate ),
    .\__mp_text_out[74]$_DFF_P_.int_fwire_IQN (\__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[75]$_DFF_P_.CLK (\__mp_text_out[75]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[75]$_DFF_P_.QN (\__mp_text_out[75]$_DFF_P_.QN__gate ),
    .\__mp_text_out[75]$_DFF_P_.int_fwire_IQN (\__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[76]$_DFF_P_.CLK (\__mp_text_out[76]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[76]$_DFF_P_.QN (\__mp_text_out[76]$_DFF_P_.QN__gate ),
    .\__mp_text_out[76]$_DFF_P_.int_fwire_IQN (\__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[77]$_DFF_P_.CLK (\__mp_text_out[77]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[77]$_DFF_P_.QN (\__mp_text_out[77]$_DFF_P_.QN__gate ),
    .\__mp_text_out[77]$_DFF_P_.int_fwire_IQN (\__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[78]$_DFF_P_.CLK (\__mp_text_out[78]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[78]$_DFF_P_.QN (\__mp_text_out[78]$_DFF_P_.QN__gate ),
    .\__mp_text_out[78]$_DFF_P_.int_fwire_IQN (\__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[79]$_DFF_P_.CLK (\__mp_text_out[79]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[79]$_DFF_P_.QN (\__mp_text_out[79]$_DFF_P_.QN__gate ),
    .\__mp_text_out[79]$_DFF_P_.int_fwire_IQN (\__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[7]$_DFF_P_.CLK (\__mp_text_out[7]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[7]$_DFF_P_.QN (\__mp_text_out[7]$_DFF_P_.QN__gate ),
    .\__mp_text_out[7]$_DFF_P_.int_fwire_IQN (\__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[80]$_DFF_P_.CLK (\__mp_text_out[80]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[80]$_DFF_P_.QN (\__mp_text_out[80]$_DFF_P_.QN__gate ),
    .\__mp_text_out[80]$_DFF_P_.int_fwire_IQN (\__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[81]$_DFF_P_.CLK (\__mp_text_out[81]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[81]$_DFF_P_.QN (\__mp_text_out[81]$_DFF_P_.QN__gate ),
    .\__mp_text_out[81]$_DFF_P_.int_fwire_IQN (\__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[82]$_DFF_P_.CLK (\__mp_text_out[82]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[82]$_DFF_P_.QN (\__mp_text_out[82]$_DFF_P_.QN__gate ),
    .\__mp_text_out[82]$_DFF_P_.int_fwire_IQN (\__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[83]$_DFF_P_.CLK (\__mp_text_out[83]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[83]$_DFF_P_.QN (\__mp_text_out[83]$_DFF_P_.QN__gate ),
    .\__mp_text_out[83]$_DFF_P_.int_fwire_IQN (\__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[84]$_DFF_P_.CLK (\__mp_text_out[84]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[84]$_DFF_P_.QN (\__mp_text_out[84]$_DFF_P_.QN__gate ),
    .\__mp_text_out[84]$_DFF_P_.int_fwire_IQN (\__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[85]$_DFF_P_.CLK (\__mp_text_out[85]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[85]$_DFF_P_.QN (\__mp_text_out[85]$_DFF_P_.QN__gate ),
    .\__mp_text_out[85]$_DFF_P_.int_fwire_IQN (\__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[86]$_DFF_P_.CLK (\__mp_text_out[86]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[86]$_DFF_P_.QN (\__mp_text_out[86]$_DFF_P_.QN__gate ),
    .\__mp_text_out[86]$_DFF_P_.int_fwire_IQN (\__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[87]$_DFF_P_.CLK (\__mp_text_out[87]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[87]$_DFF_P_.QN (\__mp_text_out[87]$_DFF_P_.QN__gate ),
    .\__mp_text_out[87]$_DFF_P_.int_fwire_IQN (\__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[88]$_DFF_P_.CLK (\__mp_text_out[88]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[88]$_DFF_P_.QN (\__mp_text_out[88]$_DFF_P_.QN__gate ),
    .\__mp_text_out[88]$_DFF_P_.int_fwire_IQN (\__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[89]$_DFF_P_.CLK (\__mp_text_out[89]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[89]$_DFF_P_.QN (\__mp_text_out[89]$_DFF_P_.QN__gate ),
    .\__mp_text_out[89]$_DFF_P_.int_fwire_IQN (\__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[8]$_DFF_P_.CLK (\__mp_text_out[8]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[8]$_DFF_P_.QN (\__mp_text_out[8]$_DFF_P_.QN__gate ),
    .\__mp_text_out[8]$_DFF_P_.int_fwire_IQN (\__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[90]$_DFF_P_.CLK (\__mp_text_out[90]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[90]$_DFF_P_.QN (\__mp_text_out[90]$_DFF_P_.QN__gate ),
    .\__mp_text_out[90]$_DFF_P_.int_fwire_IQN (\__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[91]$_DFF_P_.CLK (\__mp_text_out[91]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[91]$_DFF_P_.QN (\__mp_text_out[91]$_DFF_P_.QN__gate ),
    .\__mp_text_out[91]$_DFF_P_.int_fwire_IQN (\__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[92]$_DFF_P_.CLK (\__mp_text_out[92]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[92]$_DFF_P_.QN (\__mp_text_out[92]$_DFF_P_.QN__gate ),
    .\__mp_text_out[92]$_DFF_P_.int_fwire_IQN (\__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[93]$_DFF_P_.CLK (\__mp_text_out[93]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[93]$_DFF_P_.QN (\__mp_text_out[93]$_DFF_P_.QN__gate ),
    .\__mp_text_out[93]$_DFF_P_.int_fwire_IQN (\__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[94]$_DFF_P_.CLK (\__mp_text_out[94]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[94]$_DFF_P_.QN (\__mp_text_out[94]$_DFF_P_.QN__gate ),
    .\__mp_text_out[94]$_DFF_P_.int_fwire_IQN (\__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[95]$_DFF_P_.CLK (\__mp_text_out[95]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[95]$_DFF_P_.QN (\__mp_text_out[95]$_DFF_P_.QN__gate ),
    .\__mp_text_out[95]$_DFF_P_.int_fwire_IQN (\__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[96]$_DFF_P_.CLK (\__mp_text_out[96]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[96]$_DFF_P_.QN (\__mp_text_out[96]$_DFF_P_.QN__gate ),
    .\__mp_text_out[96]$_DFF_P_.int_fwire_IQN (\__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[97]$_DFF_P_.CLK (\__mp_text_out[97]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[97]$_DFF_P_.QN (\__mp_text_out[97]$_DFF_P_.QN__gate ),
    .\__mp_text_out[97]$_DFF_P_.int_fwire_IQN (\__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[98]$_DFF_P_.CLK (\__mp_text_out[98]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[98]$_DFF_P_.QN (\__mp_text_out[98]$_DFF_P_.QN__gate ),
    .\__mp_text_out[98]$_DFF_P_.int_fwire_IQN (\__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[99]$_DFF_P_.CLK (\__mp_text_out[99]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[99]$_DFF_P_.QN (\__mp_text_out[99]$_DFF_P_.QN__gate ),
    .\__mp_text_out[99]$_DFF_P_.int_fwire_IQN (\__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_text_out[9]$_DFF_P_.CLK (\__mp_text_out[9]$_DFF_P_.CLK__gate ),
    .\__mp_text_out[9]$_DFF_P_.QN (\__mp_text_out[9]$_DFF_P_.QN__gate ),
    .\__mp_text_out[9]$_DFF_P_.int_fwire_IQN (\__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gate ),
    .\__mp_u0.r0.out[24]$_SDFF_PP1_.CLK (\__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gate ),
    .\__mp_u0.r0.out[25]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.out[26]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.out[27]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.out[28]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.out[29]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.out[30]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.out[31]$_SDFF_PP0_.CLK (\__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK (\__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gate ),
    .\__mp_u0.u0.d[0]$_DFF_P_.CLK (\__mp_u0.u0.d[0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u0.d[1]$_DFF_P_.CLK (\__mp_u0.u0.d[1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u0.d[2]$_DFF_P_.CLK (\__mp_u0.u0.d[2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u0.d[3]$_DFF_P_.CLK (\__mp_u0.u0.d[3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u0.d[4]$_DFF_P_.CLK (\__mp_u0.u0.d[4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u0.d[5]$_DFF_P_.CLK (\__mp_u0.u0.d[5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u0.d[6]$_DFF_P_.CLK (\__mp_u0.u0.d[6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u0.d[7]$_DFF_P_.CLK (\__mp_u0.u0.d[7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[0]$_DFF_P_.CLK (\__mp_u0.u1.d[0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[1]$_DFF_P_.CLK (\__mp_u0.u1.d[1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[2]$_DFF_P_.CLK (\__mp_u0.u1.d[2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[3]$_DFF_P_.CLK (\__mp_u0.u1.d[3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[4]$_DFF_P_.CLK (\__mp_u0.u1.d[4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[5]$_DFF_P_.CLK (\__mp_u0.u1.d[5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[6]$_DFF_P_.CLK (\__mp_u0.u1.d[6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u1.d[7]$_DFF_P_.CLK (\__mp_u0.u1.d[7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[0]$_DFF_P_.CLK (\__mp_u0.u2.d[0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[1]$_DFF_P_.CLK (\__mp_u0.u2.d[1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[2]$_DFF_P_.CLK (\__mp_u0.u2.d[2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[3]$_DFF_P_.CLK (\__mp_u0.u2.d[3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[4]$_DFF_P_.CLK (\__mp_u0.u2.d[4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[5]$_DFF_P_.CLK (\__mp_u0.u2.d[5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[6]$_DFF_P_.CLK (\__mp_u0.u2.d[6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u2.d[7]$_DFF_P_.CLK (\__mp_u0.u2.d[7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[0]$_DFF_P_.CLK (\__mp_u0.u3.d[0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[1]$_DFF_P_.CLK (\__mp_u0.u3.d[1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[2]$_DFF_P_.CLK (\__mp_u0.u3.d[2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[3]$_DFF_P_.CLK (\__mp_u0.u3.d[3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[4]$_DFF_P_.CLK (\__mp_u0.u3.d[4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[5]$_DFF_P_.CLK (\__mp_u0.u3.d[5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[6]$_DFF_P_.CLK (\__mp_u0.u3.d[6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.u3.d[7]$_DFF_P_.CLK (\__mp_u0.u3.d[7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][0]$_DFF_P_.CLK (\__mp_u0.w[0][0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][10]$_DFF_P_.CLK (\__mp_u0.w[0][10]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][11]$_DFF_P_.CLK (\__mp_u0.w[0][11]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][12]$_DFF_P_.CLK (\__mp_u0.w[0][12]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][13]$_DFF_P_.CLK (\__mp_u0.w[0][13]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][14]$_DFF_P_.CLK (\__mp_u0.w[0][14]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][15]$_DFF_P_.CLK (\__mp_u0.w[0][15]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][16]$_DFF_P_.CLK (\__mp_u0.w[0][16]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][17]$_DFF_P_.CLK (\__mp_u0.w[0][17]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][18]$_DFF_P_.CLK (\__mp_u0.w[0][18]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][19]$_DFF_P_.CLK (\__mp_u0.w[0][19]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][1]$_DFF_P_.CLK (\__mp_u0.w[0][1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][20]$_DFF_P_.CLK (\__mp_u0.w[0][20]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][21]$_DFF_P_.CLK (\__mp_u0.w[0][21]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][22]$_DFF_P_.CLK (\__mp_u0.w[0][22]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][23]$_DFF_P_.CLK (\__mp_u0.w[0][23]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][24]$_DFF_P_.CLK (\__mp_u0.w[0][24]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][25]$_DFF_P_.CLK (\__mp_u0.w[0][25]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][26]$_DFF_P_.CLK (\__mp_u0.w[0][26]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][27]$_DFF_P_.CLK (\__mp_u0.w[0][27]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][28]$_DFF_P_.CLK (\__mp_u0.w[0][28]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][29]$_DFF_P_.CLK (\__mp_u0.w[0][29]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][2]$_DFF_P_.CLK (\__mp_u0.w[0][2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][30]$_DFF_P_.CLK (\__mp_u0.w[0][30]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][31]$_DFF_P_.CLK (\__mp_u0.w[0][31]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][3]$_DFF_P_.CLK (\__mp_u0.w[0][3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][4]$_DFF_P_.CLK (\__mp_u0.w[0][4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][5]$_DFF_P_.CLK (\__mp_u0.w[0][5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][6]$_DFF_P_.CLK (\__mp_u0.w[0][6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][7]$_DFF_P_.CLK (\__mp_u0.w[0][7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][8]$_DFF_P_.CLK (\__mp_u0.w[0][8]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[0][9]$_DFF_P_.CLK (\__mp_u0.w[0][9]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][0]$_DFF_P_.CLK (\__mp_u0.w[1][0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][10]$_DFF_P_.CLK (\__mp_u0.w[1][10]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][11]$_DFF_P_.CLK (\__mp_u0.w[1][11]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][12]$_DFF_P_.CLK (\__mp_u0.w[1][12]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][13]$_DFF_P_.CLK (\__mp_u0.w[1][13]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][14]$_DFF_P_.CLK (\__mp_u0.w[1][14]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][15]$_DFF_P_.CLK (\__mp_u0.w[1][15]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][16]$_DFF_P_.CLK (\__mp_u0.w[1][16]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][17]$_DFF_P_.CLK (\__mp_u0.w[1][17]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][18]$_DFF_P_.CLK (\__mp_u0.w[1][18]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][19]$_DFF_P_.CLK (\__mp_u0.w[1][19]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][1]$_DFF_P_.CLK (\__mp_u0.w[1][1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][20]$_DFF_P_.CLK (\__mp_u0.w[1][20]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][21]$_DFF_P_.CLK (\__mp_u0.w[1][21]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][22]$_DFF_P_.CLK (\__mp_u0.w[1][22]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][23]$_DFF_P_.CLK (\__mp_u0.w[1][23]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][24]$_DFF_P_.CLK (\__mp_u0.w[1][24]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][25]$_DFF_P_.CLK (\__mp_u0.w[1][25]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][26]$_DFF_P_.CLK (\__mp_u0.w[1][26]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][27]$_DFF_P_.CLK (\__mp_u0.w[1][27]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][28]$_DFF_P_.CLK (\__mp_u0.w[1][28]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][29]$_DFF_P_.CLK (\__mp_u0.w[1][29]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][2]$_DFF_P_.CLK (\__mp_u0.w[1][2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][30]$_DFF_P_.CLK (\__mp_u0.w[1][30]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][31]$_DFF_P_.CLK (\__mp_u0.w[1][31]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][3]$_DFF_P_.CLK (\__mp_u0.w[1][3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][4]$_DFF_P_.CLK (\__mp_u0.w[1][4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][5]$_DFF_P_.CLK (\__mp_u0.w[1][5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][6]$_DFF_P_.CLK (\__mp_u0.w[1][6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][7]$_DFF_P_.CLK (\__mp_u0.w[1][7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][8]$_DFF_P_.CLK (\__mp_u0.w[1][8]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[1][9]$_DFF_P_.CLK (\__mp_u0.w[1][9]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][0]$_DFF_P_.CLK (\__mp_u0.w[2][0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][10]$_DFF_P_.CLK (\__mp_u0.w[2][10]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][11]$_DFF_P_.CLK (\__mp_u0.w[2][11]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][12]$_DFF_P_.CLK (\__mp_u0.w[2][12]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][13]$_DFF_P_.CLK (\__mp_u0.w[2][13]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][14]$_DFF_P_.CLK (\__mp_u0.w[2][14]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][15]$_DFF_P_.CLK (\__mp_u0.w[2][15]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][16]$_DFF_P_.CLK (\__mp_u0.w[2][16]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][17]$_DFF_P_.CLK (\__mp_u0.w[2][17]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][18]$_DFF_P_.CLK (\__mp_u0.w[2][18]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][19]$_DFF_P_.CLK (\__mp_u0.w[2][19]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][1]$_DFF_P_.CLK (\__mp_u0.w[2][1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][20]$_DFF_P_.CLK (\__mp_u0.w[2][20]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][21]$_DFF_P_.CLK (\__mp_u0.w[2][21]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][22]$_DFF_P_.CLK (\__mp_u0.w[2][22]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][23]$_DFF_P_.CLK (\__mp_u0.w[2][23]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][24]$_DFF_P_.CLK (\__mp_u0.w[2][24]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][25]$_DFF_P_.CLK (\__mp_u0.w[2][25]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][26]$_DFF_P_.CLK (\__mp_u0.w[2][26]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][27]$_DFF_P_.CLK (\__mp_u0.w[2][27]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][28]$_DFF_P_.CLK (\__mp_u0.w[2][28]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][29]$_DFF_P_.CLK (\__mp_u0.w[2][29]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][2]$_DFF_P_.CLK (\__mp_u0.w[2][2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][30]$_DFF_P_.CLK (\__mp_u0.w[2][30]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][31]$_DFF_P_.CLK (\__mp_u0.w[2][31]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][3]$_DFF_P_.CLK (\__mp_u0.w[2][3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][4]$_DFF_P_.CLK (\__mp_u0.w[2][4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][5]$_DFF_P_.CLK (\__mp_u0.w[2][5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][6]$_DFF_P_.CLK (\__mp_u0.w[2][6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][7]$_DFF_P_.CLK (\__mp_u0.w[2][7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][8]$_DFF_P_.CLK (\__mp_u0.w[2][8]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[2][9]$_DFF_P_.CLK (\__mp_u0.w[2][9]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][0]$_DFF_P_.CLK (\__mp_u0.w[3][0]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][10]$_DFF_P_.CLK (\__mp_u0.w[3][10]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][11]$_DFF_P_.CLK (\__mp_u0.w[3][11]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][12]$_DFF_P_.CLK (\__mp_u0.w[3][12]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][13]$_DFF_P_.CLK (\__mp_u0.w[3][13]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][14]$_DFF_P_.CLK (\__mp_u0.w[3][14]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][15]$_DFF_P_.CLK (\__mp_u0.w[3][15]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][16]$_DFF_P_.CLK (\__mp_u0.w[3][16]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][17]$_DFF_P_.CLK (\__mp_u0.w[3][17]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][18]$_DFF_P_.CLK (\__mp_u0.w[3][18]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][19]$_DFF_P_.CLK (\__mp_u0.w[3][19]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][1]$_DFF_P_.CLK (\__mp_u0.w[3][1]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][20]$_DFF_P_.CLK (\__mp_u0.w[3][20]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][21]$_DFF_P_.CLK (\__mp_u0.w[3][21]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][22]$_DFF_P_.CLK (\__mp_u0.w[3][22]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][23]$_DFF_P_.CLK (\__mp_u0.w[3][23]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][24]$_DFF_P_.CLK (\__mp_u0.w[3][24]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][25]$_DFF_P_.CLK (\__mp_u0.w[3][25]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][26]$_DFF_P_.CLK (\__mp_u0.w[3][26]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][27]$_DFF_P_.CLK (\__mp_u0.w[3][27]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][28]$_DFF_P_.CLK (\__mp_u0.w[3][28]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][29]$_DFF_P_.CLK (\__mp_u0.w[3][29]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][2]$_DFF_P_.CLK (\__mp_u0.w[3][2]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][30]$_DFF_P_.CLK (\__mp_u0.w[3][30]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][31]$_DFF_P_.CLK (\__mp_u0.w[3][31]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][3]$_DFF_P_.CLK (\__mp_u0.w[3][3]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][4]$_DFF_P_.CLK (\__mp_u0.w[3][4]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][5]$_DFF_P_.CLK (\__mp_u0.w[3][5]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][6]$_DFF_P_.CLK (\__mp_u0.w[3][6]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][7]$_DFF_P_.CLK (\__mp_u0.w[3][7]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][8]$_DFF_P_.CLK (\__mp_u0.w[3][8]$_DFF_P_.CLK__gate ),
    .\__mp_u0.w[3][9]$_DFF_P_.CLK (\__mp_u0.w[3][9]$_DFF_P_.CLK__gate ),
    .\__po_done (\__po_done__gate ),
    .\__po_text_out (\__po_text_out__gate )
  );
`ifdef ASSUME_DEFINED_INPUTS
  miter_def_prop #(1, "assume") \__pi_clk__assume (\__pi_clk );
  miter_def_prop #(128, "assume") \__pi_key__assume (\__pi_key );
  miter_def_prop #(1, "assume") \__pi_ld__assume (\__pi_ld );
  miter_def_prop #(1, "assume") \__pi_rst__assume (\__pi_rst );
  miter_def_prop #(128, "assume") \__pi_text_in__assume (\__pi_text_in );
`endif
`ifndef DIRECT_CROSS_POINTS
`endif
`ifdef CHECK_MATCH_POINTS
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_0_clk.A__assert (\__mp_clkbuf_0_clk.A__gold , \__mp_clkbuf_0_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_0_clk.Y__assert (\__mp_clkbuf_0_clk.Y__gold , \__mp_clkbuf_0_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_0_0_clk.A__assert (\__mp_clkbuf_2_0_0_clk.A__gold , \__mp_clkbuf_2_0_0_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_0_0_clk.Y__assert (\__mp_clkbuf_2_0_0_clk.Y__gold , \__mp_clkbuf_2_0_0_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_1_0_clk.A__assert (\__mp_clkbuf_2_1_0_clk.A__gold , \__mp_clkbuf_2_1_0_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_1_0_clk.Y__assert (\__mp_clkbuf_2_1_0_clk.Y__gold , \__mp_clkbuf_2_1_0_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_2_0_clk.A__assert (\__mp_clkbuf_2_2_0_clk.A__gold , \__mp_clkbuf_2_2_0_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_2_0_clk.Y__assert (\__mp_clkbuf_2_2_0_clk.Y__gold , \__mp_clkbuf_2_2_0_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_3_0_clk.A__assert (\__mp_clkbuf_2_3_0_clk.A__gold , \__mp_clkbuf_2_3_0_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_2_3_0_clk.Y__assert (\__mp_clkbuf_2_3_0_clk.Y__gold , \__mp_clkbuf_2_3_0_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_0_clk.A__assert (\__mp_clkbuf_leaf_0_clk.A__gold , \__mp_clkbuf_leaf_0_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_0_clk.Y__assert (\__mp_clkbuf_leaf_0_clk.Y__gold , \__mp_clkbuf_leaf_0_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_10_clk.A__assert (\__mp_clkbuf_leaf_10_clk.A__gold , \__mp_clkbuf_leaf_10_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_10_clk.Y__assert (\__mp_clkbuf_leaf_10_clk.Y__gold , \__mp_clkbuf_leaf_10_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_11_clk.A__assert (\__mp_clkbuf_leaf_11_clk.A__gold , \__mp_clkbuf_leaf_11_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_11_clk.Y__assert (\__mp_clkbuf_leaf_11_clk.Y__gold , \__mp_clkbuf_leaf_11_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_12_clk.A__assert (\__mp_clkbuf_leaf_12_clk.A__gold , \__mp_clkbuf_leaf_12_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_12_clk.Y__assert (\__mp_clkbuf_leaf_12_clk.Y__gold , \__mp_clkbuf_leaf_12_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_13_clk.A__assert (\__mp_clkbuf_leaf_13_clk.A__gold , \__mp_clkbuf_leaf_13_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_13_clk.Y__assert (\__mp_clkbuf_leaf_13_clk.Y__gold , \__mp_clkbuf_leaf_13_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_14_clk.A__assert (\__mp_clkbuf_leaf_14_clk.A__gold , \__mp_clkbuf_leaf_14_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_14_clk.Y__assert (\__mp_clkbuf_leaf_14_clk.Y__gold , \__mp_clkbuf_leaf_14_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_15_clk.A__assert (\__mp_clkbuf_leaf_15_clk.A__gold , \__mp_clkbuf_leaf_15_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_15_clk.Y__assert (\__mp_clkbuf_leaf_15_clk.Y__gold , \__mp_clkbuf_leaf_15_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_16_clk.A__assert (\__mp_clkbuf_leaf_16_clk.A__gold , \__mp_clkbuf_leaf_16_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_16_clk.Y__assert (\__mp_clkbuf_leaf_16_clk.Y__gold , \__mp_clkbuf_leaf_16_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_17_clk.A__assert (\__mp_clkbuf_leaf_17_clk.A__gold , \__mp_clkbuf_leaf_17_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_17_clk.Y__assert (\__mp_clkbuf_leaf_17_clk.Y__gold , \__mp_clkbuf_leaf_17_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_18_clk.A__assert (\__mp_clkbuf_leaf_18_clk.A__gold , \__mp_clkbuf_leaf_18_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_18_clk.Y__assert (\__mp_clkbuf_leaf_18_clk.Y__gold , \__mp_clkbuf_leaf_18_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_19_clk.A__assert (\__mp_clkbuf_leaf_19_clk.A__gold , \__mp_clkbuf_leaf_19_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_19_clk.Y__assert (\__mp_clkbuf_leaf_19_clk.Y__gold , \__mp_clkbuf_leaf_19_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_1_clk.A__assert (\__mp_clkbuf_leaf_1_clk.A__gold , \__mp_clkbuf_leaf_1_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_1_clk.Y__assert (\__mp_clkbuf_leaf_1_clk.Y__gold , \__mp_clkbuf_leaf_1_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_20_clk.A__assert (\__mp_clkbuf_leaf_20_clk.A__gold , \__mp_clkbuf_leaf_20_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_20_clk.Y__assert (\__mp_clkbuf_leaf_20_clk.Y__gold , \__mp_clkbuf_leaf_20_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_21_clk.A__assert (\__mp_clkbuf_leaf_21_clk.A__gold , \__mp_clkbuf_leaf_21_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_21_clk.Y__assert (\__mp_clkbuf_leaf_21_clk.Y__gold , \__mp_clkbuf_leaf_21_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_22_clk.A__assert (\__mp_clkbuf_leaf_22_clk.A__gold , \__mp_clkbuf_leaf_22_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_22_clk.Y__assert (\__mp_clkbuf_leaf_22_clk.Y__gold , \__mp_clkbuf_leaf_22_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_23_clk.A__assert (\__mp_clkbuf_leaf_23_clk.A__gold , \__mp_clkbuf_leaf_23_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_23_clk.Y__assert (\__mp_clkbuf_leaf_23_clk.Y__gold , \__mp_clkbuf_leaf_23_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_24_clk.A__assert (\__mp_clkbuf_leaf_24_clk.A__gold , \__mp_clkbuf_leaf_24_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_24_clk.Y__assert (\__mp_clkbuf_leaf_24_clk.Y__gold , \__mp_clkbuf_leaf_24_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_25_clk.A__assert (\__mp_clkbuf_leaf_25_clk.A__gold , \__mp_clkbuf_leaf_25_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_25_clk.Y__assert (\__mp_clkbuf_leaf_25_clk.Y__gold , \__mp_clkbuf_leaf_25_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_26_clk.A__assert (\__mp_clkbuf_leaf_26_clk.A__gold , \__mp_clkbuf_leaf_26_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_26_clk.Y__assert (\__mp_clkbuf_leaf_26_clk.Y__gold , \__mp_clkbuf_leaf_26_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_27_clk.A__assert (\__mp_clkbuf_leaf_27_clk.A__gold , \__mp_clkbuf_leaf_27_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_27_clk.Y__assert (\__mp_clkbuf_leaf_27_clk.Y__gold , \__mp_clkbuf_leaf_27_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_28_clk.A__assert (\__mp_clkbuf_leaf_28_clk.A__gold , \__mp_clkbuf_leaf_28_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_28_clk.Y__assert (\__mp_clkbuf_leaf_28_clk.Y__gold , \__mp_clkbuf_leaf_28_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_29_clk.A__assert (\__mp_clkbuf_leaf_29_clk.A__gold , \__mp_clkbuf_leaf_29_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_29_clk.Y__assert (\__mp_clkbuf_leaf_29_clk.Y__gold , \__mp_clkbuf_leaf_29_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_2_clk.A__assert (\__mp_clkbuf_leaf_2_clk.A__gold , \__mp_clkbuf_leaf_2_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_2_clk.Y__assert (\__mp_clkbuf_leaf_2_clk.Y__gold , \__mp_clkbuf_leaf_2_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_30_clk.A__assert (\__mp_clkbuf_leaf_30_clk.A__gold , \__mp_clkbuf_leaf_30_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_30_clk.Y__assert (\__mp_clkbuf_leaf_30_clk.Y__gold , \__mp_clkbuf_leaf_30_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_31_clk.A__assert (\__mp_clkbuf_leaf_31_clk.A__gold , \__mp_clkbuf_leaf_31_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_31_clk.Y__assert (\__mp_clkbuf_leaf_31_clk.Y__gold , \__mp_clkbuf_leaf_31_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_32_clk.A__assert (\__mp_clkbuf_leaf_32_clk.A__gold , \__mp_clkbuf_leaf_32_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_32_clk.Y__assert (\__mp_clkbuf_leaf_32_clk.Y__gold , \__mp_clkbuf_leaf_32_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_33_clk.A__assert (\__mp_clkbuf_leaf_33_clk.A__gold , \__mp_clkbuf_leaf_33_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_33_clk.Y__assert (\__mp_clkbuf_leaf_33_clk.Y__gold , \__mp_clkbuf_leaf_33_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_3_clk.A__assert (\__mp_clkbuf_leaf_3_clk.A__gold , \__mp_clkbuf_leaf_3_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_3_clk.Y__assert (\__mp_clkbuf_leaf_3_clk.Y__gold , \__mp_clkbuf_leaf_3_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_4_clk.A__assert (\__mp_clkbuf_leaf_4_clk.A__gold , \__mp_clkbuf_leaf_4_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_4_clk.Y__assert (\__mp_clkbuf_leaf_4_clk.Y__gold , \__mp_clkbuf_leaf_4_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_5_clk.A__assert (\__mp_clkbuf_leaf_5_clk.A__gold , \__mp_clkbuf_leaf_5_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_5_clk.Y__assert (\__mp_clkbuf_leaf_5_clk.Y__gold , \__mp_clkbuf_leaf_5_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_6_clk.A__assert (\__mp_clkbuf_leaf_6_clk.A__gold , \__mp_clkbuf_leaf_6_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_6_clk.Y__assert (\__mp_clkbuf_leaf_6_clk.Y__gold , \__mp_clkbuf_leaf_6_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_7_clk.A__assert (\__mp_clkbuf_leaf_7_clk.A__gold , \__mp_clkbuf_leaf_7_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_7_clk.Y__assert (\__mp_clkbuf_leaf_7_clk.Y__gold , \__mp_clkbuf_leaf_7_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_8_clk.A__assert (\__mp_clkbuf_leaf_8_clk.A__gold , \__mp_clkbuf_leaf_8_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_8_clk.Y__assert (\__mp_clkbuf_leaf_8_clk.Y__gold , \__mp_clkbuf_leaf_8_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_9_clk.A__assert (\__mp_clkbuf_leaf_9_clk.A__gold , \__mp_clkbuf_leaf_9_clk.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkbuf_leaf_9_clk.Y__assert (\__mp_clkbuf_leaf_9_clk.Y__gold , \__mp_clkbuf_leaf_9_clk.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload0.A__assert (\__mp_clkload0.A__gold , \__mp_clkload0.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload0.Y__assert (\__mp_clkload0.Y__gold , \__mp_clkload0.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload1.A__assert (\__mp_clkload1.A__gold , \__mp_clkload1.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload10.A__assert (\__mp_clkload10.A__gold , \__mp_clkload10.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload11.A__assert (\__mp_clkload11.A__gold , \__mp_clkload11.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload12.A__assert (\__mp_clkload12.A__gold , \__mp_clkload12.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload13.A__assert (\__mp_clkload13.A__gold , \__mp_clkload13.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload14.A__assert (\__mp_clkload14.A__gold , \__mp_clkload14.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload15.A__assert (\__mp_clkload15.A__gold , \__mp_clkload15.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload16.A__assert (\__mp_clkload16.A__gold , \__mp_clkload16.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload17.A__assert (\__mp_clkload17.A__gold , \__mp_clkload17.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload18.A__assert (\__mp_clkload18.A__gold , \__mp_clkload18.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload18.Y__assert (\__mp_clkload18.Y__gold , \__mp_clkload18.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload19.A__assert (\__mp_clkload19.A__gold , \__mp_clkload19.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload2.A__assert (\__mp_clkload2.A__gold , \__mp_clkload2.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload20.A__assert (\__mp_clkload20.A__gold , \__mp_clkload20.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload21.A__assert (\__mp_clkload21.A__gold , \__mp_clkload21.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload22.A__assert (\__mp_clkload22.A__gold , \__mp_clkload22.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload23.A__assert (\__mp_clkload23.A__gold , \__mp_clkload23.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload24.A__assert (\__mp_clkload24.A__gold , \__mp_clkload24.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload25.A__assert (\__mp_clkload25.A__gold , \__mp_clkload25.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload26.A__assert (\__mp_clkload26.A__gold , \__mp_clkload26.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload27.A__assert (\__mp_clkload27.A__gold , \__mp_clkload27.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload28.A__assert (\__mp_clkload28.A__gold , \__mp_clkload28.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload29.A__assert (\__mp_clkload29.A__gold , \__mp_clkload29.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload3.A__assert (\__mp_clkload3.A__gold , \__mp_clkload3.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload30.A__assert (\__mp_clkload30.A__gold , \__mp_clkload30.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload31.A__assert (\__mp_clkload31.A__gold , \__mp_clkload31.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload31.Y__assert (\__mp_clkload31.Y__gold , \__mp_clkload31.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload32.A__assert (\__mp_clkload32.A__gold , \__mp_clkload32.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload4.A__assert (\__mp_clkload4.A__gold , \__mp_clkload4.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload5.A__assert (\__mp_clkload5.A__gold , \__mp_clkload5.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload6.A__assert (\__mp_clkload6.A__gold , \__mp_clkload6.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload7.A__assert (\__mp_clkload7.A__gold , \__mp_clkload7.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload8.A__assert (\__mp_clkload8.A__gold , \__mp_clkload8.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clkload9.A__assert (\__mp_clkload9.A__gold , \__mp_clkload9.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_0_clk__assert (\__mp_clknet_0_clk__gold , \__mp_clknet_0_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_2_0_0_clk__assert (\__mp_clknet_2_0_0_clk__gold , \__mp_clknet_2_0_0_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_2_1_0_clk__assert (\__mp_clknet_2_1_0_clk__gold , \__mp_clknet_2_1_0_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_2_2_0_clk__assert (\__mp_clknet_2_2_0_clk__gold , \__mp_clknet_2_2_0_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_2_3_0_clk__assert (\__mp_clknet_2_3_0_clk__gold , \__mp_clknet_2_3_0_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_0_clk__assert (\__mp_clknet_leaf_0_clk__gold , \__mp_clknet_leaf_0_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_10_clk__assert (\__mp_clknet_leaf_10_clk__gold , \__mp_clknet_leaf_10_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_11_clk__assert (\__mp_clknet_leaf_11_clk__gold , \__mp_clknet_leaf_11_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_12_clk__assert (\__mp_clknet_leaf_12_clk__gold , \__mp_clknet_leaf_12_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_13_clk__assert (\__mp_clknet_leaf_13_clk__gold , \__mp_clknet_leaf_13_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_14_clk__assert (\__mp_clknet_leaf_14_clk__gold , \__mp_clknet_leaf_14_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_15_clk__assert (\__mp_clknet_leaf_15_clk__gold , \__mp_clknet_leaf_15_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_16_clk__assert (\__mp_clknet_leaf_16_clk__gold , \__mp_clknet_leaf_16_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_17_clk__assert (\__mp_clknet_leaf_17_clk__gold , \__mp_clknet_leaf_17_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_18_clk__assert (\__mp_clknet_leaf_18_clk__gold , \__mp_clknet_leaf_18_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_19_clk__assert (\__mp_clknet_leaf_19_clk__gold , \__mp_clknet_leaf_19_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_1_clk__assert (\__mp_clknet_leaf_1_clk__gold , \__mp_clknet_leaf_1_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_20_clk__assert (\__mp_clknet_leaf_20_clk__gold , \__mp_clknet_leaf_20_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_21_clk__assert (\__mp_clknet_leaf_21_clk__gold , \__mp_clknet_leaf_21_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_22_clk__assert (\__mp_clknet_leaf_22_clk__gold , \__mp_clknet_leaf_22_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_23_clk__assert (\__mp_clknet_leaf_23_clk__gold , \__mp_clknet_leaf_23_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_24_clk__assert (\__mp_clknet_leaf_24_clk__gold , \__mp_clknet_leaf_24_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_25_clk__assert (\__mp_clknet_leaf_25_clk__gold , \__mp_clknet_leaf_25_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_26_clk__assert (\__mp_clknet_leaf_26_clk__gold , \__mp_clknet_leaf_26_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_27_clk__assert (\__mp_clknet_leaf_27_clk__gold , \__mp_clknet_leaf_27_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_28_clk__assert (\__mp_clknet_leaf_28_clk__gold , \__mp_clknet_leaf_28_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_29_clk__assert (\__mp_clknet_leaf_29_clk__gold , \__mp_clknet_leaf_29_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_2_clk__assert (\__mp_clknet_leaf_2_clk__gold , \__mp_clknet_leaf_2_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_30_clk__assert (\__mp_clknet_leaf_30_clk__gold , \__mp_clknet_leaf_30_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_31_clk__assert (\__mp_clknet_leaf_31_clk__gold , \__mp_clknet_leaf_31_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_32_clk__assert (\__mp_clknet_leaf_32_clk__gold , \__mp_clknet_leaf_32_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_33_clk__assert (\__mp_clknet_leaf_33_clk__gold , \__mp_clknet_leaf_33_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_3_clk__assert (\__mp_clknet_leaf_3_clk__gold , \__mp_clknet_leaf_3_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_4_clk__assert (\__mp_clknet_leaf_4_clk__gold , \__mp_clknet_leaf_4_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_5_clk__assert (\__mp_clknet_leaf_5_clk__gold , \__mp_clknet_leaf_5_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_6_clk__assert (\__mp_clknet_leaf_6_clk__gold , \__mp_clknet_leaf_6_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_7_clk__assert (\__mp_clknet_leaf_7_clk__gold , \__mp_clknet_leaf_7_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_8_clk__assert (\__mp_clknet_leaf_8_clk__gold , \__mp_clknet_leaf_8_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_clknet_leaf_9_clk__assert (\__mp_clknet_leaf_9_clk__gold , \__mp_clknet_leaf_9_clk__gate );
  miter_cmp_prop #(1, "assert") \__mp_dcnt[0]$_SDFFE_PN0P_.CLK__assert (\__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gold , \__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_dcnt[1]$_SDFFE_PN0P_.CLK__assert (\__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gold , \__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_dcnt[2]$_SDFFE_PP0P_.CLK__assert (\__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gold , \__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_dcnt[3]$_SDFFE_PN0P_.CLK__assert (\__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gold , \__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_done$_DFF_P_.CLK__assert (\__mp_done$_DFF_P_.CLK__gold , \__mp_done$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_done$_DFF_P_.QN__assert (\__mp_done$_DFF_P_.QN__gold , \__mp_done$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_done$_DFF_P_.int_fwire_IQN__assert (\__mp_done$_DFF_P_.int_fwire_IQN__gold , \__mp_done$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_input1.A__assert (\__mp_input1.A__gold , \__mp_input1.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input1.Y__assert (\__mp_input1.Y__gold , \__mp_input1.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input10.A__assert (\__mp_input10.A__gold , \__mp_input10.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input10.Y__assert (\__mp_input10.Y__gold , \__mp_input10.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input100.A__assert (\__mp_input100.A__gold , \__mp_input100.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input100.Y__assert (\__mp_input100.Y__gold , \__mp_input100.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input101.A__assert (\__mp_input101.A__gold , \__mp_input101.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input101.Y__assert (\__mp_input101.Y__gold , \__mp_input101.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input102.A__assert (\__mp_input102.A__gold , \__mp_input102.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input102.Y__assert (\__mp_input102.Y__gold , \__mp_input102.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input103.A__assert (\__mp_input103.A__gold , \__mp_input103.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input103.Y__assert (\__mp_input103.Y__gold , \__mp_input103.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input104.A__assert (\__mp_input104.A__gold , \__mp_input104.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input104.Y__assert (\__mp_input104.Y__gold , \__mp_input104.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input105.A__assert (\__mp_input105.A__gold , \__mp_input105.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input105.Y__assert (\__mp_input105.Y__gold , \__mp_input105.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input106.A__assert (\__mp_input106.A__gold , \__mp_input106.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input106.Y__assert (\__mp_input106.Y__gold , \__mp_input106.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input107.A__assert (\__mp_input107.A__gold , \__mp_input107.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input107.Y__assert (\__mp_input107.Y__gold , \__mp_input107.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input108.A__assert (\__mp_input108.A__gold , \__mp_input108.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input108.Y__assert (\__mp_input108.Y__gold , \__mp_input108.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input109.A__assert (\__mp_input109.A__gold , \__mp_input109.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input109.Y__assert (\__mp_input109.Y__gold , \__mp_input109.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input11.A__assert (\__mp_input11.A__gold , \__mp_input11.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input11.Y__assert (\__mp_input11.Y__gold , \__mp_input11.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input110.A__assert (\__mp_input110.A__gold , \__mp_input110.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input110.Y__assert (\__mp_input110.Y__gold , \__mp_input110.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input111.A__assert (\__mp_input111.A__gold , \__mp_input111.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input111.Y__assert (\__mp_input111.Y__gold , \__mp_input111.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input112.A__assert (\__mp_input112.A__gold , \__mp_input112.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input112.Y__assert (\__mp_input112.Y__gold , \__mp_input112.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input113.A__assert (\__mp_input113.A__gold , \__mp_input113.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input113.Y__assert (\__mp_input113.Y__gold , \__mp_input113.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input114.A__assert (\__mp_input114.A__gold , \__mp_input114.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input114.Y__assert (\__mp_input114.Y__gold , \__mp_input114.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input115.A__assert (\__mp_input115.A__gold , \__mp_input115.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input115.Y__assert (\__mp_input115.Y__gold , \__mp_input115.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input116.A__assert (\__mp_input116.A__gold , \__mp_input116.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input116.Y__assert (\__mp_input116.Y__gold , \__mp_input116.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input117.A__assert (\__mp_input117.A__gold , \__mp_input117.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input117.Y__assert (\__mp_input117.Y__gold , \__mp_input117.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input118.A__assert (\__mp_input118.A__gold , \__mp_input118.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input118.Y__assert (\__mp_input118.Y__gold , \__mp_input118.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input119.A__assert (\__mp_input119.A__gold , \__mp_input119.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input119.Y__assert (\__mp_input119.Y__gold , \__mp_input119.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input12.A__assert (\__mp_input12.A__gold , \__mp_input12.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input12.Y__assert (\__mp_input12.Y__gold , \__mp_input12.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input120.A__assert (\__mp_input120.A__gold , \__mp_input120.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input120.Y__assert (\__mp_input120.Y__gold , \__mp_input120.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input121.A__assert (\__mp_input121.A__gold , \__mp_input121.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input121.Y__assert (\__mp_input121.Y__gold , \__mp_input121.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input122.A__assert (\__mp_input122.A__gold , \__mp_input122.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input122.Y__assert (\__mp_input122.Y__gold , \__mp_input122.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input123.A__assert (\__mp_input123.A__gold , \__mp_input123.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input123.Y__assert (\__mp_input123.Y__gold , \__mp_input123.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input124.A__assert (\__mp_input124.A__gold , \__mp_input124.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input124.Y__assert (\__mp_input124.Y__gold , \__mp_input124.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input125.A__assert (\__mp_input125.A__gold , \__mp_input125.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input125.Y__assert (\__mp_input125.Y__gold , \__mp_input125.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input126.A__assert (\__mp_input126.A__gold , \__mp_input126.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input126.Y__assert (\__mp_input126.Y__gold , \__mp_input126.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input127.A__assert (\__mp_input127.A__gold , \__mp_input127.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input127.Y__assert (\__mp_input127.Y__gold , \__mp_input127.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input128.A__assert (\__mp_input128.A__gold , \__mp_input128.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input128.Y__assert (\__mp_input128.Y__gold , \__mp_input128.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input129.A__assert (\__mp_input129.A__gold , \__mp_input129.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input129.Y__assert (\__mp_input129.Y__gold , \__mp_input129.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input13.A__assert (\__mp_input13.A__gold , \__mp_input13.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input13.Y__assert (\__mp_input13.Y__gold , \__mp_input13.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input130.A__assert (\__mp_input130.A__gold , \__mp_input130.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input130.Y__assert (\__mp_input130.Y__gold , \__mp_input130.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input131.A__assert (\__mp_input131.A__gold , \__mp_input131.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input131.Y__assert (\__mp_input131.Y__gold , \__mp_input131.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input132.A__assert (\__mp_input132.A__gold , \__mp_input132.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input132.Y__assert (\__mp_input132.Y__gold , \__mp_input132.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input133.A__assert (\__mp_input133.A__gold , \__mp_input133.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input133.Y__assert (\__mp_input133.Y__gold , \__mp_input133.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input134.A__assert (\__mp_input134.A__gold , \__mp_input134.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input134.Y__assert (\__mp_input134.Y__gold , \__mp_input134.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input135.A__assert (\__mp_input135.A__gold , \__mp_input135.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input135.Y__assert (\__mp_input135.Y__gold , \__mp_input135.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input136.A__assert (\__mp_input136.A__gold , \__mp_input136.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input136.Y__assert (\__mp_input136.Y__gold , \__mp_input136.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input137.A__assert (\__mp_input137.A__gold , \__mp_input137.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input137.Y__assert (\__mp_input137.Y__gold , \__mp_input137.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input138.A__assert (\__mp_input138.A__gold , \__mp_input138.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input138.Y__assert (\__mp_input138.Y__gold , \__mp_input138.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input139.A__assert (\__mp_input139.A__gold , \__mp_input139.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input139.Y__assert (\__mp_input139.Y__gold , \__mp_input139.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input14.A__assert (\__mp_input14.A__gold , \__mp_input14.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input14.Y__assert (\__mp_input14.Y__gold , \__mp_input14.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input140.A__assert (\__mp_input140.A__gold , \__mp_input140.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input140.Y__assert (\__mp_input140.Y__gold , \__mp_input140.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input141.A__assert (\__mp_input141.A__gold , \__mp_input141.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input141.Y__assert (\__mp_input141.Y__gold , \__mp_input141.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input142.A__assert (\__mp_input142.A__gold , \__mp_input142.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input142.Y__assert (\__mp_input142.Y__gold , \__mp_input142.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input143.A__assert (\__mp_input143.A__gold , \__mp_input143.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input143.Y__assert (\__mp_input143.Y__gold , \__mp_input143.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input144.A__assert (\__mp_input144.A__gold , \__mp_input144.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input144.Y__assert (\__mp_input144.Y__gold , \__mp_input144.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input145.A__assert (\__mp_input145.A__gold , \__mp_input145.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input145.Y__assert (\__mp_input145.Y__gold , \__mp_input145.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input146.A__assert (\__mp_input146.A__gold , \__mp_input146.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input146.Y__assert (\__mp_input146.Y__gold , \__mp_input146.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input147.A__assert (\__mp_input147.A__gold , \__mp_input147.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input147.Y__assert (\__mp_input147.Y__gold , \__mp_input147.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input148.A__assert (\__mp_input148.A__gold , \__mp_input148.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input148.Y__assert (\__mp_input148.Y__gold , \__mp_input148.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input149.A__assert (\__mp_input149.A__gold , \__mp_input149.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input149.Y__assert (\__mp_input149.Y__gold , \__mp_input149.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input15.A__assert (\__mp_input15.A__gold , \__mp_input15.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input15.Y__assert (\__mp_input15.Y__gold , \__mp_input15.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input150.A__assert (\__mp_input150.A__gold , \__mp_input150.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input150.Y__assert (\__mp_input150.Y__gold , \__mp_input150.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input151.A__assert (\__mp_input151.A__gold , \__mp_input151.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input151.Y__assert (\__mp_input151.Y__gold , \__mp_input151.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input152.A__assert (\__mp_input152.A__gold , \__mp_input152.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input152.Y__assert (\__mp_input152.Y__gold , \__mp_input152.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input153.A__assert (\__mp_input153.A__gold , \__mp_input153.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input153.Y__assert (\__mp_input153.Y__gold , \__mp_input153.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input154.A__assert (\__mp_input154.A__gold , \__mp_input154.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input154.Y__assert (\__mp_input154.Y__gold , \__mp_input154.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input155.A__assert (\__mp_input155.A__gold , \__mp_input155.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input155.Y__assert (\__mp_input155.Y__gold , \__mp_input155.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input156.A__assert (\__mp_input156.A__gold , \__mp_input156.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input156.Y__assert (\__mp_input156.Y__gold , \__mp_input156.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input157.A__assert (\__mp_input157.A__gold , \__mp_input157.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input157.Y__assert (\__mp_input157.Y__gold , \__mp_input157.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input158.A__assert (\__mp_input158.A__gold , \__mp_input158.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input158.Y__assert (\__mp_input158.Y__gold , \__mp_input158.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input159.A__assert (\__mp_input159.A__gold , \__mp_input159.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input159.Y__assert (\__mp_input159.Y__gold , \__mp_input159.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input16.A__assert (\__mp_input16.A__gold , \__mp_input16.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input16.Y__assert (\__mp_input16.Y__gold , \__mp_input16.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input160.A__assert (\__mp_input160.A__gold , \__mp_input160.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input160.Y__assert (\__mp_input160.Y__gold , \__mp_input160.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input161.A__assert (\__mp_input161.A__gold , \__mp_input161.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input161.Y__assert (\__mp_input161.Y__gold , \__mp_input161.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input162.A__assert (\__mp_input162.A__gold , \__mp_input162.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input162.Y__assert (\__mp_input162.Y__gold , \__mp_input162.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input163.A__assert (\__mp_input163.A__gold , \__mp_input163.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input163.Y__assert (\__mp_input163.Y__gold , \__mp_input163.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input164.A__assert (\__mp_input164.A__gold , \__mp_input164.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input164.Y__assert (\__mp_input164.Y__gold , \__mp_input164.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input165.A__assert (\__mp_input165.A__gold , \__mp_input165.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input165.Y__assert (\__mp_input165.Y__gold , \__mp_input165.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input166.A__assert (\__mp_input166.A__gold , \__mp_input166.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input166.Y__assert (\__mp_input166.Y__gold , \__mp_input166.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input167.A__assert (\__mp_input167.A__gold , \__mp_input167.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input167.Y__assert (\__mp_input167.Y__gold , \__mp_input167.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input168.A__assert (\__mp_input168.A__gold , \__mp_input168.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input168.Y__assert (\__mp_input168.Y__gold , \__mp_input168.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input169.A__assert (\__mp_input169.A__gold , \__mp_input169.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input169.Y__assert (\__mp_input169.Y__gold , \__mp_input169.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input17.A__assert (\__mp_input17.A__gold , \__mp_input17.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input17.Y__assert (\__mp_input17.Y__gold , \__mp_input17.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input170.A__assert (\__mp_input170.A__gold , \__mp_input170.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input170.Y__assert (\__mp_input170.Y__gold , \__mp_input170.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input171.A__assert (\__mp_input171.A__gold , \__mp_input171.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input171.Y__assert (\__mp_input171.Y__gold , \__mp_input171.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input172.A__assert (\__mp_input172.A__gold , \__mp_input172.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input172.Y__assert (\__mp_input172.Y__gold , \__mp_input172.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input173.A__assert (\__mp_input173.A__gold , \__mp_input173.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input173.Y__assert (\__mp_input173.Y__gold , \__mp_input173.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input174.A__assert (\__mp_input174.A__gold , \__mp_input174.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input174.Y__assert (\__mp_input174.Y__gold , \__mp_input174.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input175.A__assert (\__mp_input175.A__gold , \__mp_input175.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input175.Y__assert (\__mp_input175.Y__gold , \__mp_input175.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input176.A__assert (\__mp_input176.A__gold , \__mp_input176.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input176.Y__assert (\__mp_input176.Y__gold , \__mp_input176.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input177.A__assert (\__mp_input177.A__gold , \__mp_input177.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input177.Y__assert (\__mp_input177.Y__gold , \__mp_input177.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input178.A__assert (\__mp_input178.A__gold , \__mp_input178.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input178.Y__assert (\__mp_input178.Y__gold , \__mp_input178.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input179.A__assert (\__mp_input179.A__gold , \__mp_input179.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input179.Y__assert (\__mp_input179.Y__gold , \__mp_input179.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input18.A__assert (\__mp_input18.A__gold , \__mp_input18.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input18.Y__assert (\__mp_input18.Y__gold , \__mp_input18.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input180.A__assert (\__mp_input180.A__gold , \__mp_input180.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input180.Y__assert (\__mp_input180.Y__gold , \__mp_input180.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input181.A__assert (\__mp_input181.A__gold , \__mp_input181.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input181.Y__assert (\__mp_input181.Y__gold , \__mp_input181.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input182.A__assert (\__mp_input182.A__gold , \__mp_input182.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input182.Y__assert (\__mp_input182.Y__gold , \__mp_input182.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input183.A__assert (\__mp_input183.A__gold , \__mp_input183.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input183.Y__assert (\__mp_input183.Y__gold , \__mp_input183.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input184.A__assert (\__mp_input184.A__gold , \__mp_input184.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input184.Y__assert (\__mp_input184.Y__gold , \__mp_input184.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input185.A__assert (\__mp_input185.A__gold , \__mp_input185.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input185.Y__assert (\__mp_input185.Y__gold , \__mp_input185.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input186.A__assert (\__mp_input186.A__gold , \__mp_input186.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input186.Y__assert (\__mp_input186.Y__gold , \__mp_input186.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input187.A__assert (\__mp_input187.A__gold , \__mp_input187.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input187.Y__assert (\__mp_input187.Y__gold , \__mp_input187.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input188.A__assert (\__mp_input188.A__gold , \__mp_input188.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input188.Y__assert (\__mp_input188.Y__gold , \__mp_input188.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input189.A__assert (\__mp_input189.A__gold , \__mp_input189.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input189.Y__assert (\__mp_input189.Y__gold , \__mp_input189.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input19.A__assert (\__mp_input19.A__gold , \__mp_input19.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input19.Y__assert (\__mp_input19.Y__gold , \__mp_input19.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input190.A__assert (\__mp_input190.A__gold , \__mp_input190.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input190.Y__assert (\__mp_input190.Y__gold , \__mp_input190.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input191.A__assert (\__mp_input191.A__gold , \__mp_input191.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input191.Y__assert (\__mp_input191.Y__gold , \__mp_input191.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input192.A__assert (\__mp_input192.A__gold , \__mp_input192.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input192.Y__assert (\__mp_input192.Y__gold , \__mp_input192.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input193.A__assert (\__mp_input193.A__gold , \__mp_input193.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input193.Y__assert (\__mp_input193.Y__gold , \__mp_input193.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input194.A__assert (\__mp_input194.A__gold , \__mp_input194.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input194.Y__assert (\__mp_input194.Y__gold , \__mp_input194.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input195.A__assert (\__mp_input195.A__gold , \__mp_input195.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input195.Y__assert (\__mp_input195.Y__gold , \__mp_input195.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input196.A__assert (\__mp_input196.A__gold , \__mp_input196.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input196.Y__assert (\__mp_input196.Y__gold , \__mp_input196.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input197.A__assert (\__mp_input197.A__gold , \__mp_input197.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input197.Y__assert (\__mp_input197.Y__gold , \__mp_input197.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input198.A__assert (\__mp_input198.A__gold , \__mp_input198.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input198.Y__assert (\__mp_input198.Y__gold , \__mp_input198.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input199.A__assert (\__mp_input199.A__gold , \__mp_input199.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input199.Y__assert (\__mp_input199.Y__gold , \__mp_input199.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input2.A__assert (\__mp_input2.A__gold , \__mp_input2.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input2.Y__assert (\__mp_input2.Y__gold , \__mp_input2.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input20.A__assert (\__mp_input20.A__gold , \__mp_input20.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input20.Y__assert (\__mp_input20.Y__gold , \__mp_input20.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input200.A__assert (\__mp_input200.A__gold , \__mp_input200.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input200.Y__assert (\__mp_input200.Y__gold , \__mp_input200.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input201.A__assert (\__mp_input201.A__gold , \__mp_input201.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input201.Y__assert (\__mp_input201.Y__gold , \__mp_input201.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input202.A__assert (\__mp_input202.A__gold , \__mp_input202.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input202.Y__assert (\__mp_input202.Y__gold , \__mp_input202.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input203.A__assert (\__mp_input203.A__gold , \__mp_input203.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input203.Y__assert (\__mp_input203.Y__gold , \__mp_input203.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input204.A__assert (\__mp_input204.A__gold , \__mp_input204.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input204.Y__assert (\__mp_input204.Y__gold , \__mp_input204.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input205.A__assert (\__mp_input205.A__gold , \__mp_input205.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input205.Y__assert (\__mp_input205.Y__gold , \__mp_input205.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input206.A__assert (\__mp_input206.A__gold , \__mp_input206.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input206.Y__assert (\__mp_input206.Y__gold , \__mp_input206.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input207.A__assert (\__mp_input207.A__gold , \__mp_input207.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input207.Y__assert (\__mp_input207.Y__gold , \__mp_input207.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input208.A__assert (\__mp_input208.A__gold , \__mp_input208.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input208.Y__assert (\__mp_input208.Y__gold , \__mp_input208.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input209.A__assert (\__mp_input209.A__gold , \__mp_input209.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input209.Y__assert (\__mp_input209.Y__gold , \__mp_input209.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input21.A__assert (\__mp_input21.A__gold , \__mp_input21.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input21.Y__assert (\__mp_input21.Y__gold , \__mp_input21.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input210.A__assert (\__mp_input210.A__gold , \__mp_input210.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input210.Y__assert (\__mp_input210.Y__gold , \__mp_input210.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input211.A__assert (\__mp_input211.A__gold , \__mp_input211.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input211.Y__assert (\__mp_input211.Y__gold , \__mp_input211.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input212.A__assert (\__mp_input212.A__gold , \__mp_input212.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input212.Y__assert (\__mp_input212.Y__gold , \__mp_input212.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input213.A__assert (\__mp_input213.A__gold , \__mp_input213.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input213.Y__assert (\__mp_input213.Y__gold , \__mp_input213.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input214.A__assert (\__mp_input214.A__gold , \__mp_input214.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input214.Y__assert (\__mp_input214.Y__gold , \__mp_input214.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input215.A__assert (\__mp_input215.A__gold , \__mp_input215.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input215.Y__assert (\__mp_input215.Y__gold , \__mp_input215.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input216.A__assert (\__mp_input216.A__gold , \__mp_input216.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input216.Y__assert (\__mp_input216.Y__gold , \__mp_input216.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input217.A__assert (\__mp_input217.A__gold , \__mp_input217.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input217.Y__assert (\__mp_input217.Y__gold , \__mp_input217.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input218.A__assert (\__mp_input218.A__gold , \__mp_input218.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input218.Y__assert (\__mp_input218.Y__gold , \__mp_input218.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input219.A__assert (\__mp_input219.A__gold , \__mp_input219.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input219.Y__assert (\__mp_input219.Y__gold , \__mp_input219.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input22.A__assert (\__mp_input22.A__gold , \__mp_input22.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input22.Y__assert (\__mp_input22.Y__gold , \__mp_input22.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input220.A__assert (\__mp_input220.A__gold , \__mp_input220.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input220.Y__assert (\__mp_input220.Y__gold , \__mp_input220.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input221.A__assert (\__mp_input221.A__gold , \__mp_input221.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input221.Y__assert (\__mp_input221.Y__gold , \__mp_input221.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input222.A__assert (\__mp_input222.A__gold , \__mp_input222.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input222.Y__assert (\__mp_input222.Y__gold , \__mp_input222.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input223.A__assert (\__mp_input223.A__gold , \__mp_input223.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input223.Y__assert (\__mp_input223.Y__gold , \__mp_input223.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input224.A__assert (\__mp_input224.A__gold , \__mp_input224.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input224.Y__assert (\__mp_input224.Y__gold , \__mp_input224.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input225.A__assert (\__mp_input225.A__gold , \__mp_input225.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input225.Y__assert (\__mp_input225.Y__gold , \__mp_input225.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input226.A__assert (\__mp_input226.A__gold , \__mp_input226.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input226.Y__assert (\__mp_input226.Y__gold , \__mp_input226.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input227.A__assert (\__mp_input227.A__gold , \__mp_input227.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input227.Y__assert (\__mp_input227.Y__gold , \__mp_input227.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input228.A__assert (\__mp_input228.A__gold , \__mp_input228.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input228.Y__assert (\__mp_input228.Y__gold , \__mp_input228.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input229.A__assert (\__mp_input229.A__gold , \__mp_input229.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input229.Y__assert (\__mp_input229.Y__gold , \__mp_input229.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input23.A__assert (\__mp_input23.A__gold , \__mp_input23.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input23.Y__assert (\__mp_input23.Y__gold , \__mp_input23.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input230.A__assert (\__mp_input230.A__gold , \__mp_input230.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input230.Y__assert (\__mp_input230.Y__gold , \__mp_input230.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input231.A__assert (\__mp_input231.A__gold , \__mp_input231.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input231.Y__assert (\__mp_input231.Y__gold , \__mp_input231.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input232.A__assert (\__mp_input232.A__gold , \__mp_input232.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input232.Y__assert (\__mp_input232.Y__gold , \__mp_input232.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input233.A__assert (\__mp_input233.A__gold , \__mp_input233.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input233.Y__assert (\__mp_input233.Y__gold , \__mp_input233.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input234.A__assert (\__mp_input234.A__gold , \__mp_input234.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input234.Y__assert (\__mp_input234.Y__gold , \__mp_input234.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input235.A__assert (\__mp_input235.A__gold , \__mp_input235.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input235.Y__assert (\__mp_input235.Y__gold , \__mp_input235.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input236.A__assert (\__mp_input236.A__gold , \__mp_input236.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input236.Y__assert (\__mp_input236.Y__gold , \__mp_input236.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input237.A__assert (\__mp_input237.A__gold , \__mp_input237.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input237.Y__assert (\__mp_input237.Y__gold , \__mp_input237.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input238.A__assert (\__mp_input238.A__gold , \__mp_input238.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input238.Y__assert (\__mp_input238.Y__gold , \__mp_input238.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input239.A__assert (\__mp_input239.A__gold , \__mp_input239.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input239.Y__assert (\__mp_input239.Y__gold , \__mp_input239.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input24.A__assert (\__mp_input24.A__gold , \__mp_input24.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input24.Y__assert (\__mp_input24.Y__gold , \__mp_input24.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input240.A__assert (\__mp_input240.A__gold , \__mp_input240.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input240.Y__assert (\__mp_input240.Y__gold , \__mp_input240.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input241.A__assert (\__mp_input241.A__gold , \__mp_input241.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input241.Y__assert (\__mp_input241.Y__gold , \__mp_input241.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input242.A__assert (\__mp_input242.A__gold , \__mp_input242.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input242.Y__assert (\__mp_input242.Y__gold , \__mp_input242.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input243.A__assert (\__mp_input243.A__gold , \__mp_input243.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input243.Y__assert (\__mp_input243.Y__gold , \__mp_input243.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input244.A__assert (\__mp_input244.A__gold , \__mp_input244.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input244.Y__assert (\__mp_input244.Y__gold , \__mp_input244.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input245.A__assert (\__mp_input245.A__gold , \__mp_input245.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input245.Y__assert (\__mp_input245.Y__gold , \__mp_input245.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input246.A__assert (\__mp_input246.A__gold , \__mp_input246.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input246.Y__assert (\__mp_input246.Y__gold , \__mp_input246.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input247.A__assert (\__mp_input247.A__gold , \__mp_input247.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input247.Y__assert (\__mp_input247.Y__gold , \__mp_input247.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input248.A__assert (\__mp_input248.A__gold , \__mp_input248.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input248.Y__assert (\__mp_input248.Y__gold , \__mp_input248.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input249.A__assert (\__mp_input249.A__gold , \__mp_input249.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input249.Y__assert (\__mp_input249.Y__gold , \__mp_input249.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input25.A__assert (\__mp_input25.A__gold , \__mp_input25.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input25.Y__assert (\__mp_input25.Y__gold , \__mp_input25.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input250.A__assert (\__mp_input250.A__gold , \__mp_input250.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input250.Y__assert (\__mp_input250.Y__gold , \__mp_input250.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input251.A__assert (\__mp_input251.A__gold , \__mp_input251.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input251.Y__assert (\__mp_input251.Y__gold , \__mp_input251.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input252.A__assert (\__mp_input252.A__gold , \__mp_input252.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input252.Y__assert (\__mp_input252.Y__gold , \__mp_input252.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input253.A__assert (\__mp_input253.A__gold , \__mp_input253.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input253.Y__assert (\__mp_input253.Y__gold , \__mp_input253.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input254.A__assert (\__mp_input254.A__gold , \__mp_input254.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input254.Y__assert (\__mp_input254.Y__gold , \__mp_input254.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input255.A__assert (\__mp_input255.A__gold , \__mp_input255.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input255.Y__assert (\__mp_input255.Y__gold , \__mp_input255.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input256.A__assert (\__mp_input256.A__gold , \__mp_input256.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input256.Y__assert (\__mp_input256.Y__gold , \__mp_input256.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input257.A__assert (\__mp_input257.A__gold , \__mp_input257.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input257.Y__assert (\__mp_input257.Y__gold , \__mp_input257.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input258.A__assert (\__mp_input258.A__gold , \__mp_input258.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input258.Y__assert (\__mp_input258.Y__gold , \__mp_input258.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input26.A__assert (\__mp_input26.A__gold , \__mp_input26.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input26.Y__assert (\__mp_input26.Y__gold , \__mp_input26.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input27.A__assert (\__mp_input27.A__gold , \__mp_input27.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input27.Y__assert (\__mp_input27.Y__gold , \__mp_input27.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input28.A__assert (\__mp_input28.A__gold , \__mp_input28.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input28.Y__assert (\__mp_input28.Y__gold , \__mp_input28.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input29.A__assert (\__mp_input29.A__gold , \__mp_input29.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input29.Y__assert (\__mp_input29.Y__gold , \__mp_input29.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input3.A__assert (\__mp_input3.A__gold , \__mp_input3.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input3.Y__assert (\__mp_input3.Y__gold , \__mp_input3.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input30.A__assert (\__mp_input30.A__gold , \__mp_input30.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input30.Y__assert (\__mp_input30.Y__gold , \__mp_input30.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input31.A__assert (\__mp_input31.A__gold , \__mp_input31.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input31.Y__assert (\__mp_input31.Y__gold , \__mp_input31.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input32.A__assert (\__mp_input32.A__gold , \__mp_input32.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input32.Y__assert (\__mp_input32.Y__gold , \__mp_input32.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input33.A__assert (\__mp_input33.A__gold , \__mp_input33.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input33.Y__assert (\__mp_input33.Y__gold , \__mp_input33.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input34.A__assert (\__mp_input34.A__gold , \__mp_input34.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input34.Y__assert (\__mp_input34.Y__gold , \__mp_input34.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input35.A__assert (\__mp_input35.A__gold , \__mp_input35.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input35.Y__assert (\__mp_input35.Y__gold , \__mp_input35.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input36.A__assert (\__mp_input36.A__gold , \__mp_input36.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input36.Y__assert (\__mp_input36.Y__gold , \__mp_input36.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input37.A__assert (\__mp_input37.A__gold , \__mp_input37.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input37.Y__assert (\__mp_input37.Y__gold , \__mp_input37.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input38.A__assert (\__mp_input38.A__gold , \__mp_input38.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input38.Y__assert (\__mp_input38.Y__gold , \__mp_input38.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input39.A__assert (\__mp_input39.A__gold , \__mp_input39.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input39.Y__assert (\__mp_input39.Y__gold , \__mp_input39.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input4.A__assert (\__mp_input4.A__gold , \__mp_input4.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input4.Y__assert (\__mp_input4.Y__gold , \__mp_input4.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input40.A__assert (\__mp_input40.A__gold , \__mp_input40.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input40.Y__assert (\__mp_input40.Y__gold , \__mp_input40.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input41.A__assert (\__mp_input41.A__gold , \__mp_input41.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input41.Y__assert (\__mp_input41.Y__gold , \__mp_input41.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input42.A__assert (\__mp_input42.A__gold , \__mp_input42.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input42.Y__assert (\__mp_input42.Y__gold , \__mp_input42.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input43.A__assert (\__mp_input43.A__gold , \__mp_input43.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input43.Y__assert (\__mp_input43.Y__gold , \__mp_input43.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input44.A__assert (\__mp_input44.A__gold , \__mp_input44.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input44.Y__assert (\__mp_input44.Y__gold , \__mp_input44.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input45.A__assert (\__mp_input45.A__gold , \__mp_input45.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input45.Y__assert (\__mp_input45.Y__gold , \__mp_input45.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input46.A__assert (\__mp_input46.A__gold , \__mp_input46.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input46.Y__assert (\__mp_input46.Y__gold , \__mp_input46.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input47.A__assert (\__mp_input47.A__gold , \__mp_input47.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input47.Y__assert (\__mp_input47.Y__gold , \__mp_input47.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input48.A__assert (\__mp_input48.A__gold , \__mp_input48.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input48.Y__assert (\__mp_input48.Y__gold , \__mp_input48.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input49.A__assert (\__mp_input49.A__gold , \__mp_input49.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input49.Y__assert (\__mp_input49.Y__gold , \__mp_input49.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input5.A__assert (\__mp_input5.A__gold , \__mp_input5.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input5.Y__assert (\__mp_input5.Y__gold , \__mp_input5.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input50.A__assert (\__mp_input50.A__gold , \__mp_input50.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input50.Y__assert (\__mp_input50.Y__gold , \__mp_input50.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input51.A__assert (\__mp_input51.A__gold , \__mp_input51.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input51.Y__assert (\__mp_input51.Y__gold , \__mp_input51.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input52.A__assert (\__mp_input52.A__gold , \__mp_input52.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input52.Y__assert (\__mp_input52.Y__gold , \__mp_input52.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input53.A__assert (\__mp_input53.A__gold , \__mp_input53.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input53.Y__assert (\__mp_input53.Y__gold , \__mp_input53.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input54.A__assert (\__mp_input54.A__gold , \__mp_input54.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input54.Y__assert (\__mp_input54.Y__gold , \__mp_input54.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input55.A__assert (\__mp_input55.A__gold , \__mp_input55.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input55.Y__assert (\__mp_input55.Y__gold , \__mp_input55.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input56.A__assert (\__mp_input56.A__gold , \__mp_input56.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input56.Y__assert (\__mp_input56.Y__gold , \__mp_input56.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input57.A__assert (\__mp_input57.A__gold , \__mp_input57.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input57.Y__assert (\__mp_input57.Y__gold , \__mp_input57.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input58.A__assert (\__mp_input58.A__gold , \__mp_input58.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input58.Y__assert (\__mp_input58.Y__gold , \__mp_input58.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input59.A__assert (\__mp_input59.A__gold , \__mp_input59.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input59.Y__assert (\__mp_input59.Y__gold , \__mp_input59.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input6.A__assert (\__mp_input6.A__gold , \__mp_input6.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input6.Y__assert (\__mp_input6.Y__gold , \__mp_input6.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input60.A__assert (\__mp_input60.A__gold , \__mp_input60.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input60.Y__assert (\__mp_input60.Y__gold , \__mp_input60.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input61.A__assert (\__mp_input61.A__gold , \__mp_input61.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input61.Y__assert (\__mp_input61.Y__gold , \__mp_input61.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input62.A__assert (\__mp_input62.A__gold , \__mp_input62.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input62.Y__assert (\__mp_input62.Y__gold , \__mp_input62.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input63.A__assert (\__mp_input63.A__gold , \__mp_input63.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input63.Y__assert (\__mp_input63.Y__gold , \__mp_input63.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input64.A__assert (\__mp_input64.A__gold , \__mp_input64.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input64.Y__assert (\__mp_input64.Y__gold , \__mp_input64.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input65.A__assert (\__mp_input65.A__gold , \__mp_input65.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input65.Y__assert (\__mp_input65.Y__gold , \__mp_input65.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input66.A__assert (\__mp_input66.A__gold , \__mp_input66.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input66.Y__assert (\__mp_input66.Y__gold , \__mp_input66.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input67.A__assert (\__mp_input67.A__gold , \__mp_input67.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input67.Y__assert (\__mp_input67.Y__gold , \__mp_input67.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input68.A__assert (\__mp_input68.A__gold , \__mp_input68.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input68.Y__assert (\__mp_input68.Y__gold , \__mp_input68.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input69.A__assert (\__mp_input69.A__gold , \__mp_input69.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input69.Y__assert (\__mp_input69.Y__gold , \__mp_input69.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input7.A__assert (\__mp_input7.A__gold , \__mp_input7.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input7.Y__assert (\__mp_input7.Y__gold , \__mp_input7.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input70.A__assert (\__mp_input70.A__gold , \__mp_input70.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input70.Y__assert (\__mp_input70.Y__gold , \__mp_input70.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input71.A__assert (\__mp_input71.A__gold , \__mp_input71.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input71.Y__assert (\__mp_input71.Y__gold , \__mp_input71.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input72.A__assert (\__mp_input72.A__gold , \__mp_input72.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input72.Y__assert (\__mp_input72.Y__gold , \__mp_input72.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input73.A__assert (\__mp_input73.A__gold , \__mp_input73.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input73.Y__assert (\__mp_input73.Y__gold , \__mp_input73.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input74.A__assert (\__mp_input74.A__gold , \__mp_input74.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input74.Y__assert (\__mp_input74.Y__gold , \__mp_input74.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input75.A__assert (\__mp_input75.A__gold , \__mp_input75.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input75.Y__assert (\__mp_input75.Y__gold , \__mp_input75.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input76.A__assert (\__mp_input76.A__gold , \__mp_input76.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input76.Y__assert (\__mp_input76.Y__gold , \__mp_input76.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input77.A__assert (\__mp_input77.A__gold , \__mp_input77.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input77.Y__assert (\__mp_input77.Y__gold , \__mp_input77.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input78.A__assert (\__mp_input78.A__gold , \__mp_input78.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input78.Y__assert (\__mp_input78.Y__gold , \__mp_input78.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input79.A__assert (\__mp_input79.A__gold , \__mp_input79.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input79.Y__assert (\__mp_input79.Y__gold , \__mp_input79.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input8.A__assert (\__mp_input8.A__gold , \__mp_input8.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input8.Y__assert (\__mp_input8.Y__gold , \__mp_input8.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input80.A__assert (\__mp_input80.A__gold , \__mp_input80.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input80.Y__assert (\__mp_input80.Y__gold , \__mp_input80.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input81.A__assert (\__mp_input81.A__gold , \__mp_input81.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input81.Y__assert (\__mp_input81.Y__gold , \__mp_input81.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input82.A__assert (\__mp_input82.A__gold , \__mp_input82.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input82.Y__assert (\__mp_input82.Y__gold , \__mp_input82.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input83.A__assert (\__mp_input83.A__gold , \__mp_input83.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input83.Y__assert (\__mp_input83.Y__gold , \__mp_input83.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input84.A__assert (\__mp_input84.A__gold , \__mp_input84.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input84.Y__assert (\__mp_input84.Y__gold , \__mp_input84.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input85.A__assert (\__mp_input85.A__gold , \__mp_input85.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input85.Y__assert (\__mp_input85.Y__gold , \__mp_input85.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input86.A__assert (\__mp_input86.A__gold , \__mp_input86.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input86.Y__assert (\__mp_input86.Y__gold , \__mp_input86.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input87.A__assert (\__mp_input87.A__gold , \__mp_input87.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input87.Y__assert (\__mp_input87.Y__gold , \__mp_input87.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input88.A__assert (\__mp_input88.A__gold , \__mp_input88.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input88.Y__assert (\__mp_input88.Y__gold , \__mp_input88.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input89.A__assert (\__mp_input89.A__gold , \__mp_input89.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input89.Y__assert (\__mp_input89.Y__gold , \__mp_input89.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input9.A__assert (\__mp_input9.A__gold , \__mp_input9.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input9.Y__assert (\__mp_input9.Y__gold , \__mp_input9.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input90.A__assert (\__mp_input90.A__gold , \__mp_input90.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input90.Y__assert (\__mp_input90.Y__gold , \__mp_input90.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input91.A__assert (\__mp_input91.A__gold , \__mp_input91.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input91.Y__assert (\__mp_input91.Y__gold , \__mp_input91.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input92.A__assert (\__mp_input92.A__gold , \__mp_input92.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input92.Y__assert (\__mp_input92.Y__gold , \__mp_input92.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input93.A__assert (\__mp_input93.A__gold , \__mp_input93.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input93.Y__assert (\__mp_input93.Y__gold , \__mp_input93.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input94.A__assert (\__mp_input94.A__gold , \__mp_input94.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input94.Y__assert (\__mp_input94.Y__gold , \__mp_input94.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input95.A__assert (\__mp_input95.A__gold , \__mp_input95.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input95.Y__assert (\__mp_input95.Y__gold , \__mp_input95.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input96.A__assert (\__mp_input96.A__gold , \__mp_input96.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input96.Y__assert (\__mp_input96.Y__gold , \__mp_input96.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input97.A__assert (\__mp_input97.A__gold , \__mp_input97.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input97.Y__assert (\__mp_input97.Y__gold , \__mp_input97.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input98.A__assert (\__mp_input98.A__gold , \__mp_input98.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input98.Y__assert (\__mp_input98.Y__gold , \__mp_input98.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_input99.A__assert (\__mp_input99.A__gold , \__mp_input99.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_input99.Y__assert (\__mp_input99.Y__gold , \__mp_input99.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_ld_r$_DFF_P_.CLK__assert (\__mp_ld_r$_DFF_P_.CLK__gold , \__mp_ld_r$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_ld_r$_DFF_P_.D__assert (\__mp_ld_r$_DFF_P_.D__gold , \__mp_ld_r$_DFF_P_.D__gate );
  miter_cmp_prop #(1, "assert") \__mp_output259.A__assert (\__mp_output259.A__gold , \__mp_output259.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output259.Y__assert (\__mp_output259.Y__gold , \__mp_output259.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output260.A__assert (\__mp_output260.A__gold , \__mp_output260.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output260.Y__assert (\__mp_output260.Y__gold , \__mp_output260.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output261.A__assert (\__mp_output261.A__gold , \__mp_output261.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output261.Y__assert (\__mp_output261.Y__gold , \__mp_output261.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output262.A__assert (\__mp_output262.A__gold , \__mp_output262.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output262.Y__assert (\__mp_output262.Y__gold , \__mp_output262.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output263.A__assert (\__mp_output263.A__gold , \__mp_output263.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output263.Y__assert (\__mp_output263.Y__gold , \__mp_output263.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output264.A__assert (\__mp_output264.A__gold , \__mp_output264.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output264.Y__assert (\__mp_output264.Y__gold , \__mp_output264.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output265.A__assert (\__mp_output265.A__gold , \__mp_output265.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output265.Y__assert (\__mp_output265.Y__gold , \__mp_output265.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output266.A__assert (\__mp_output266.A__gold , \__mp_output266.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output266.Y__assert (\__mp_output266.Y__gold , \__mp_output266.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output267.A__assert (\__mp_output267.A__gold , \__mp_output267.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output267.Y__assert (\__mp_output267.Y__gold , \__mp_output267.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output268.A__assert (\__mp_output268.A__gold , \__mp_output268.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output268.Y__assert (\__mp_output268.Y__gold , \__mp_output268.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output269.A__assert (\__mp_output269.A__gold , \__mp_output269.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output269.Y__assert (\__mp_output269.Y__gold , \__mp_output269.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output270.A__assert (\__mp_output270.A__gold , \__mp_output270.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output270.Y__assert (\__mp_output270.Y__gold , \__mp_output270.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output271.A__assert (\__mp_output271.A__gold , \__mp_output271.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output271.Y__assert (\__mp_output271.Y__gold , \__mp_output271.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output272.A__assert (\__mp_output272.A__gold , \__mp_output272.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output272.Y__assert (\__mp_output272.Y__gold , \__mp_output272.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output273.A__assert (\__mp_output273.A__gold , \__mp_output273.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output273.Y__assert (\__mp_output273.Y__gold , \__mp_output273.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output274.A__assert (\__mp_output274.A__gold , \__mp_output274.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output274.Y__assert (\__mp_output274.Y__gold , \__mp_output274.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output275.A__assert (\__mp_output275.A__gold , \__mp_output275.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output275.Y__assert (\__mp_output275.Y__gold , \__mp_output275.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output276.A__assert (\__mp_output276.A__gold , \__mp_output276.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output276.Y__assert (\__mp_output276.Y__gold , \__mp_output276.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output277.A__assert (\__mp_output277.A__gold , \__mp_output277.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output277.Y__assert (\__mp_output277.Y__gold , \__mp_output277.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output278.A__assert (\__mp_output278.A__gold , \__mp_output278.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output278.Y__assert (\__mp_output278.Y__gold , \__mp_output278.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output279.A__assert (\__mp_output279.A__gold , \__mp_output279.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output279.Y__assert (\__mp_output279.Y__gold , \__mp_output279.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output280.A__assert (\__mp_output280.A__gold , \__mp_output280.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output280.Y__assert (\__mp_output280.Y__gold , \__mp_output280.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output281.A__assert (\__mp_output281.A__gold , \__mp_output281.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output281.Y__assert (\__mp_output281.Y__gold , \__mp_output281.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output282.A__assert (\__mp_output282.A__gold , \__mp_output282.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output282.Y__assert (\__mp_output282.Y__gold , \__mp_output282.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output283.A__assert (\__mp_output283.A__gold , \__mp_output283.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output283.Y__assert (\__mp_output283.Y__gold , \__mp_output283.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output284.A__assert (\__mp_output284.A__gold , \__mp_output284.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output284.Y__assert (\__mp_output284.Y__gold , \__mp_output284.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output285.A__assert (\__mp_output285.A__gold , \__mp_output285.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output285.Y__assert (\__mp_output285.Y__gold , \__mp_output285.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output286.A__assert (\__mp_output286.A__gold , \__mp_output286.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output286.Y__assert (\__mp_output286.Y__gold , \__mp_output286.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output287.A__assert (\__mp_output287.A__gold , \__mp_output287.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output287.Y__assert (\__mp_output287.Y__gold , \__mp_output287.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output288.A__assert (\__mp_output288.A__gold , \__mp_output288.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output288.Y__assert (\__mp_output288.Y__gold , \__mp_output288.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output289.A__assert (\__mp_output289.A__gold , \__mp_output289.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output289.Y__assert (\__mp_output289.Y__gold , \__mp_output289.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output290.A__assert (\__mp_output290.A__gold , \__mp_output290.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output290.Y__assert (\__mp_output290.Y__gold , \__mp_output290.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output291.A__assert (\__mp_output291.A__gold , \__mp_output291.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output291.Y__assert (\__mp_output291.Y__gold , \__mp_output291.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output292.A__assert (\__mp_output292.A__gold , \__mp_output292.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output292.Y__assert (\__mp_output292.Y__gold , \__mp_output292.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output293.A__assert (\__mp_output293.A__gold , \__mp_output293.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output293.Y__assert (\__mp_output293.Y__gold , \__mp_output293.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output294.A__assert (\__mp_output294.A__gold , \__mp_output294.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output294.Y__assert (\__mp_output294.Y__gold , \__mp_output294.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output295.A__assert (\__mp_output295.A__gold , \__mp_output295.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output295.Y__assert (\__mp_output295.Y__gold , \__mp_output295.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output296.A__assert (\__mp_output296.A__gold , \__mp_output296.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output296.Y__assert (\__mp_output296.Y__gold , \__mp_output296.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output297.A__assert (\__mp_output297.A__gold , \__mp_output297.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output297.Y__assert (\__mp_output297.Y__gold , \__mp_output297.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output298.A__assert (\__mp_output298.A__gold , \__mp_output298.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output298.Y__assert (\__mp_output298.Y__gold , \__mp_output298.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output299.A__assert (\__mp_output299.A__gold , \__mp_output299.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output299.Y__assert (\__mp_output299.Y__gold , \__mp_output299.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output300.A__assert (\__mp_output300.A__gold , \__mp_output300.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output300.Y__assert (\__mp_output300.Y__gold , \__mp_output300.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output301.A__assert (\__mp_output301.A__gold , \__mp_output301.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output301.Y__assert (\__mp_output301.Y__gold , \__mp_output301.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output302.A__assert (\__mp_output302.A__gold , \__mp_output302.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output302.Y__assert (\__mp_output302.Y__gold , \__mp_output302.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output303.A__assert (\__mp_output303.A__gold , \__mp_output303.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output303.Y__assert (\__mp_output303.Y__gold , \__mp_output303.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output304.A__assert (\__mp_output304.A__gold , \__mp_output304.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output304.Y__assert (\__mp_output304.Y__gold , \__mp_output304.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output305.A__assert (\__mp_output305.A__gold , \__mp_output305.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output305.Y__assert (\__mp_output305.Y__gold , \__mp_output305.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output306.A__assert (\__mp_output306.A__gold , \__mp_output306.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output306.Y__assert (\__mp_output306.Y__gold , \__mp_output306.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output307.A__assert (\__mp_output307.A__gold , \__mp_output307.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output307.Y__assert (\__mp_output307.Y__gold , \__mp_output307.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output308.A__assert (\__mp_output308.A__gold , \__mp_output308.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output308.Y__assert (\__mp_output308.Y__gold , \__mp_output308.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output309.A__assert (\__mp_output309.A__gold , \__mp_output309.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output309.Y__assert (\__mp_output309.Y__gold , \__mp_output309.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output310.A__assert (\__mp_output310.A__gold , \__mp_output310.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output310.Y__assert (\__mp_output310.Y__gold , \__mp_output310.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output311.A__assert (\__mp_output311.A__gold , \__mp_output311.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output311.Y__assert (\__mp_output311.Y__gold , \__mp_output311.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output312.A__assert (\__mp_output312.A__gold , \__mp_output312.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output312.Y__assert (\__mp_output312.Y__gold , \__mp_output312.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output313.A__assert (\__mp_output313.A__gold , \__mp_output313.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output313.Y__assert (\__mp_output313.Y__gold , \__mp_output313.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output314.A__assert (\__mp_output314.A__gold , \__mp_output314.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output314.Y__assert (\__mp_output314.Y__gold , \__mp_output314.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output315.A__assert (\__mp_output315.A__gold , \__mp_output315.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output315.Y__assert (\__mp_output315.Y__gold , \__mp_output315.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output316.A__assert (\__mp_output316.A__gold , \__mp_output316.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output316.Y__assert (\__mp_output316.Y__gold , \__mp_output316.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output317.A__assert (\__mp_output317.A__gold , \__mp_output317.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output317.Y__assert (\__mp_output317.Y__gold , \__mp_output317.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output318.A__assert (\__mp_output318.A__gold , \__mp_output318.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output318.Y__assert (\__mp_output318.Y__gold , \__mp_output318.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output319.A__assert (\__mp_output319.A__gold , \__mp_output319.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output319.Y__assert (\__mp_output319.Y__gold , \__mp_output319.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output320.A__assert (\__mp_output320.A__gold , \__mp_output320.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output320.Y__assert (\__mp_output320.Y__gold , \__mp_output320.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output321.A__assert (\__mp_output321.A__gold , \__mp_output321.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output321.Y__assert (\__mp_output321.Y__gold , \__mp_output321.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output322.A__assert (\__mp_output322.A__gold , \__mp_output322.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output322.Y__assert (\__mp_output322.Y__gold , \__mp_output322.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output323.A__assert (\__mp_output323.A__gold , \__mp_output323.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output323.Y__assert (\__mp_output323.Y__gold , \__mp_output323.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output324.A__assert (\__mp_output324.A__gold , \__mp_output324.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output324.Y__assert (\__mp_output324.Y__gold , \__mp_output324.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output325.A__assert (\__mp_output325.A__gold , \__mp_output325.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output325.Y__assert (\__mp_output325.Y__gold , \__mp_output325.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output326.A__assert (\__mp_output326.A__gold , \__mp_output326.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output326.Y__assert (\__mp_output326.Y__gold , \__mp_output326.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output327.A__assert (\__mp_output327.A__gold , \__mp_output327.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output327.Y__assert (\__mp_output327.Y__gold , \__mp_output327.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output328.A__assert (\__mp_output328.A__gold , \__mp_output328.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output328.Y__assert (\__mp_output328.Y__gold , \__mp_output328.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output329.A__assert (\__mp_output329.A__gold , \__mp_output329.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output329.Y__assert (\__mp_output329.Y__gold , \__mp_output329.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output330.A__assert (\__mp_output330.A__gold , \__mp_output330.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output330.Y__assert (\__mp_output330.Y__gold , \__mp_output330.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output331.A__assert (\__mp_output331.A__gold , \__mp_output331.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output331.Y__assert (\__mp_output331.Y__gold , \__mp_output331.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output332.A__assert (\__mp_output332.A__gold , \__mp_output332.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output332.Y__assert (\__mp_output332.Y__gold , \__mp_output332.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output333.A__assert (\__mp_output333.A__gold , \__mp_output333.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output333.Y__assert (\__mp_output333.Y__gold , \__mp_output333.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output334.A__assert (\__mp_output334.A__gold , \__mp_output334.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output334.Y__assert (\__mp_output334.Y__gold , \__mp_output334.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output335.A__assert (\__mp_output335.A__gold , \__mp_output335.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output335.Y__assert (\__mp_output335.Y__gold , \__mp_output335.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output336.A__assert (\__mp_output336.A__gold , \__mp_output336.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output336.Y__assert (\__mp_output336.Y__gold , \__mp_output336.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output337.A__assert (\__mp_output337.A__gold , \__mp_output337.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output337.Y__assert (\__mp_output337.Y__gold , \__mp_output337.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output338.A__assert (\__mp_output338.A__gold , \__mp_output338.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output338.Y__assert (\__mp_output338.Y__gold , \__mp_output338.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output339.A__assert (\__mp_output339.A__gold , \__mp_output339.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output339.Y__assert (\__mp_output339.Y__gold , \__mp_output339.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output340.A__assert (\__mp_output340.A__gold , \__mp_output340.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output340.Y__assert (\__mp_output340.Y__gold , \__mp_output340.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output341.A__assert (\__mp_output341.A__gold , \__mp_output341.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output341.Y__assert (\__mp_output341.Y__gold , \__mp_output341.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output342.A__assert (\__mp_output342.A__gold , \__mp_output342.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output342.Y__assert (\__mp_output342.Y__gold , \__mp_output342.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output343.A__assert (\__mp_output343.A__gold , \__mp_output343.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output343.Y__assert (\__mp_output343.Y__gold , \__mp_output343.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output344.A__assert (\__mp_output344.A__gold , \__mp_output344.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output344.Y__assert (\__mp_output344.Y__gold , \__mp_output344.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output345.A__assert (\__mp_output345.A__gold , \__mp_output345.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output345.Y__assert (\__mp_output345.Y__gold , \__mp_output345.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output346.A__assert (\__mp_output346.A__gold , \__mp_output346.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output346.Y__assert (\__mp_output346.Y__gold , \__mp_output346.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output347.A__assert (\__mp_output347.A__gold , \__mp_output347.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output347.Y__assert (\__mp_output347.Y__gold , \__mp_output347.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output348.A__assert (\__mp_output348.A__gold , \__mp_output348.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output348.Y__assert (\__mp_output348.Y__gold , \__mp_output348.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output349.A__assert (\__mp_output349.A__gold , \__mp_output349.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output349.Y__assert (\__mp_output349.Y__gold , \__mp_output349.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output350.A__assert (\__mp_output350.A__gold , \__mp_output350.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output350.Y__assert (\__mp_output350.Y__gold , \__mp_output350.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output351.A__assert (\__mp_output351.A__gold , \__mp_output351.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output351.Y__assert (\__mp_output351.Y__gold , \__mp_output351.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output352.A__assert (\__mp_output352.A__gold , \__mp_output352.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output352.Y__assert (\__mp_output352.Y__gold , \__mp_output352.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output353.A__assert (\__mp_output353.A__gold , \__mp_output353.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output353.Y__assert (\__mp_output353.Y__gold , \__mp_output353.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output354.A__assert (\__mp_output354.A__gold , \__mp_output354.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output354.Y__assert (\__mp_output354.Y__gold , \__mp_output354.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output355.A__assert (\__mp_output355.A__gold , \__mp_output355.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output355.Y__assert (\__mp_output355.Y__gold , \__mp_output355.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output356.A__assert (\__mp_output356.A__gold , \__mp_output356.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output356.Y__assert (\__mp_output356.Y__gold , \__mp_output356.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output357.A__assert (\__mp_output357.A__gold , \__mp_output357.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output357.Y__assert (\__mp_output357.Y__gold , \__mp_output357.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output358.A__assert (\__mp_output358.A__gold , \__mp_output358.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output358.Y__assert (\__mp_output358.Y__gold , \__mp_output358.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output359.A__assert (\__mp_output359.A__gold , \__mp_output359.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output359.Y__assert (\__mp_output359.Y__gold , \__mp_output359.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output360.A__assert (\__mp_output360.A__gold , \__mp_output360.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output360.Y__assert (\__mp_output360.Y__gold , \__mp_output360.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output361.A__assert (\__mp_output361.A__gold , \__mp_output361.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output361.Y__assert (\__mp_output361.Y__gold , \__mp_output361.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output362.A__assert (\__mp_output362.A__gold , \__mp_output362.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output362.Y__assert (\__mp_output362.Y__gold , \__mp_output362.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output363.A__assert (\__mp_output363.A__gold , \__mp_output363.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output363.Y__assert (\__mp_output363.Y__gold , \__mp_output363.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output364.A__assert (\__mp_output364.A__gold , \__mp_output364.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output364.Y__assert (\__mp_output364.Y__gold , \__mp_output364.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output365.A__assert (\__mp_output365.A__gold , \__mp_output365.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output365.Y__assert (\__mp_output365.Y__gold , \__mp_output365.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output366.A__assert (\__mp_output366.A__gold , \__mp_output366.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output366.Y__assert (\__mp_output366.Y__gold , \__mp_output366.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output367.A__assert (\__mp_output367.A__gold , \__mp_output367.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output367.Y__assert (\__mp_output367.Y__gold , \__mp_output367.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output368.A__assert (\__mp_output368.A__gold , \__mp_output368.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output368.Y__assert (\__mp_output368.Y__gold , \__mp_output368.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output369.A__assert (\__mp_output369.A__gold , \__mp_output369.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output369.Y__assert (\__mp_output369.Y__gold , \__mp_output369.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output370.A__assert (\__mp_output370.A__gold , \__mp_output370.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output370.Y__assert (\__mp_output370.Y__gold , \__mp_output370.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output371.A__assert (\__mp_output371.A__gold , \__mp_output371.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output371.Y__assert (\__mp_output371.Y__gold , \__mp_output371.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output372.A__assert (\__mp_output372.A__gold , \__mp_output372.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output372.Y__assert (\__mp_output372.Y__gold , \__mp_output372.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output373.A__assert (\__mp_output373.A__gold , \__mp_output373.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output373.Y__assert (\__mp_output373.Y__gold , \__mp_output373.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output374.A__assert (\__mp_output374.A__gold , \__mp_output374.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output374.Y__assert (\__mp_output374.Y__gold , \__mp_output374.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output375.A__assert (\__mp_output375.A__gold , \__mp_output375.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output375.Y__assert (\__mp_output375.Y__gold , \__mp_output375.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output376.A__assert (\__mp_output376.A__gold , \__mp_output376.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output376.Y__assert (\__mp_output376.Y__gold , \__mp_output376.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output377.A__assert (\__mp_output377.A__gold , \__mp_output377.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output377.Y__assert (\__mp_output377.Y__gold , \__mp_output377.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output378.A__assert (\__mp_output378.A__gold , \__mp_output378.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output378.Y__assert (\__mp_output378.Y__gold , \__mp_output378.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output379.A__assert (\__mp_output379.A__gold , \__mp_output379.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output379.Y__assert (\__mp_output379.Y__gold , \__mp_output379.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output380.A__assert (\__mp_output380.A__gold , \__mp_output380.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output380.Y__assert (\__mp_output380.Y__gold , \__mp_output380.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output381.A__assert (\__mp_output381.A__gold , \__mp_output381.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output381.Y__assert (\__mp_output381.Y__gold , \__mp_output381.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output382.A__assert (\__mp_output382.A__gold , \__mp_output382.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output382.Y__assert (\__mp_output382.Y__gold , \__mp_output382.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output383.A__assert (\__mp_output383.A__gold , \__mp_output383.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output383.Y__assert (\__mp_output383.Y__gold , \__mp_output383.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output384.A__assert (\__mp_output384.A__gold , \__mp_output384.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output384.Y__assert (\__mp_output384.Y__gold , \__mp_output384.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output385.A__assert (\__mp_output385.A__gold , \__mp_output385.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output385.Y__assert (\__mp_output385.Y__gold , \__mp_output385.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output386.A__assert (\__mp_output386.A__gold , \__mp_output386.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output386.Y__assert (\__mp_output386.Y__gold , \__mp_output386.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_output387.A__assert (\__mp_output387.A__gold , \__mp_output387.A__gate );
  miter_cmp_prop #(1, "assert") \__mp_output387.Y__assert (\__mp_output387.Y__gold , \__mp_output387.Y__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[0]$_DFF_P_.CLK__assert (\__mp_sa00_sr[0]$_DFF_P_.CLK__gold , \__mp_sa00_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[1]$_DFF_P_.CLK__assert (\__mp_sa00_sr[1]$_DFF_P_.CLK__gold , \__mp_sa00_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[2]$_DFF_P_.CLK__assert (\__mp_sa00_sr[2]$_DFF_P_.CLK__gold , \__mp_sa00_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[3]$_DFF_P_.CLK__assert (\__mp_sa00_sr[3]$_DFF_P_.CLK__gold , \__mp_sa00_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[4]$_DFF_P_.CLK__assert (\__mp_sa00_sr[4]$_DFF_P_.CLK__gold , \__mp_sa00_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[5]$_DFF_P_.CLK__assert (\__mp_sa00_sr[5]$_DFF_P_.CLK__gold , \__mp_sa00_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[6]$_DFF_P_.CLK__assert (\__mp_sa00_sr[6]$_DFF_P_.CLK__gold , \__mp_sa00_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa00_sr[7]$_DFF_P_.CLK__assert (\__mp_sa00_sr[7]$_DFF_P_.CLK__gold , \__mp_sa00_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[0]$_DFF_P_.CLK__assert (\__mp_sa01_sr[0]$_DFF_P_.CLK__gold , \__mp_sa01_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[1]$_DFF_P_.CLK__assert (\__mp_sa01_sr[1]$_DFF_P_.CLK__gold , \__mp_sa01_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[2]$_DFF_P_.CLK__assert (\__mp_sa01_sr[2]$_DFF_P_.CLK__gold , \__mp_sa01_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[3]$_DFF_P_.CLK__assert (\__mp_sa01_sr[3]$_DFF_P_.CLK__gold , \__mp_sa01_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[4]$_DFF_P_.CLK__assert (\__mp_sa01_sr[4]$_DFF_P_.CLK__gold , \__mp_sa01_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[5]$_DFF_P_.CLK__assert (\__mp_sa01_sr[5]$_DFF_P_.CLK__gold , \__mp_sa01_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[6]$_DFF_P_.CLK__assert (\__mp_sa01_sr[6]$_DFF_P_.CLK__gold , \__mp_sa01_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa01_sr[7]$_DFF_P_.CLK__assert (\__mp_sa01_sr[7]$_DFF_P_.CLK__gold , \__mp_sa01_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[0]$_DFF_P_.CLK__assert (\__mp_sa02_sr[0]$_DFF_P_.CLK__gold , \__mp_sa02_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[1]$_DFF_P_.CLK__assert (\__mp_sa02_sr[1]$_DFF_P_.CLK__gold , \__mp_sa02_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[2]$_DFF_P_.CLK__assert (\__mp_sa02_sr[2]$_DFF_P_.CLK__gold , \__mp_sa02_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[3]$_DFF_P_.CLK__assert (\__mp_sa02_sr[3]$_DFF_P_.CLK__gold , \__mp_sa02_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[4]$_DFF_P_.CLK__assert (\__mp_sa02_sr[4]$_DFF_P_.CLK__gold , \__mp_sa02_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[5]$_DFF_P_.CLK__assert (\__mp_sa02_sr[5]$_DFF_P_.CLK__gold , \__mp_sa02_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[6]$_DFF_P_.CLK__assert (\__mp_sa02_sr[6]$_DFF_P_.CLK__gold , \__mp_sa02_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa02_sr[7]$_DFF_P_.CLK__assert (\__mp_sa02_sr[7]$_DFF_P_.CLK__gold , \__mp_sa02_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[0]$_DFF_P_.CLK__assert (\__mp_sa03_sr[0]$_DFF_P_.CLK__gold , \__mp_sa03_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[1]$_DFF_P_.CLK__assert (\__mp_sa03_sr[1]$_DFF_P_.CLK__gold , \__mp_sa03_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[2]$_DFF_P_.CLK__assert (\__mp_sa03_sr[2]$_DFF_P_.CLK__gold , \__mp_sa03_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[3]$_DFF_P_.CLK__assert (\__mp_sa03_sr[3]$_DFF_P_.CLK__gold , \__mp_sa03_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[4]$_DFF_P_.CLK__assert (\__mp_sa03_sr[4]$_DFF_P_.CLK__gold , \__mp_sa03_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[5]$_DFF_P_.CLK__assert (\__mp_sa03_sr[5]$_DFF_P_.CLK__gold , \__mp_sa03_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[6]$_DFF_P_.CLK__assert (\__mp_sa03_sr[6]$_DFF_P_.CLK__gold , \__mp_sa03_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa03_sr[7]$_DFF_P_.CLK__assert (\__mp_sa03_sr[7]$_DFF_P_.CLK__gold , \__mp_sa03_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[0]$_DFF_P_.CLK__assert (\__mp_sa10_sr[0]$_DFF_P_.CLK__gold , \__mp_sa10_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[1]$_DFF_P_.CLK__assert (\__mp_sa10_sr[1]$_DFF_P_.CLK__gold , \__mp_sa10_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[2]$_DFF_P_.CLK__assert (\__mp_sa10_sr[2]$_DFF_P_.CLK__gold , \__mp_sa10_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[3]$_DFF_P_.CLK__assert (\__mp_sa10_sr[3]$_DFF_P_.CLK__gold , \__mp_sa10_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[4]$_DFF_P_.CLK__assert (\__mp_sa10_sr[4]$_DFF_P_.CLK__gold , \__mp_sa10_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[5]$_DFF_P_.CLK__assert (\__mp_sa10_sr[5]$_DFF_P_.CLK__gold , \__mp_sa10_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[6]$_DFF_P_.CLK__assert (\__mp_sa10_sr[6]$_DFF_P_.CLK__gold , \__mp_sa10_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa10_sr[7]$_DFF_P_.CLK__assert (\__mp_sa10_sr[7]$_DFF_P_.CLK__gold , \__mp_sa10_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[0]$_DFF_P_.CLK__assert (\__mp_sa11_sr[0]$_DFF_P_.CLK__gold , \__mp_sa11_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[1]$_DFF_P_.CLK__assert (\__mp_sa11_sr[1]$_DFF_P_.CLK__gold , \__mp_sa11_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[2]$_DFF_P_.CLK__assert (\__mp_sa11_sr[2]$_DFF_P_.CLK__gold , \__mp_sa11_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[3]$_DFF_P_.CLK__assert (\__mp_sa11_sr[3]$_DFF_P_.CLK__gold , \__mp_sa11_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[4]$_DFF_P_.CLK__assert (\__mp_sa11_sr[4]$_DFF_P_.CLK__gold , \__mp_sa11_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[5]$_DFF_P_.CLK__assert (\__mp_sa11_sr[5]$_DFF_P_.CLK__gold , \__mp_sa11_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[6]$_DFF_P_.CLK__assert (\__mp_sa11_sr[6]$_DFF_P_.CLK__gold , \__mp_sa11_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa11_sr[7]$_DFF_P_.CLK__assert (\__mp_sa11_sr[7]$_DFF_P_.CLK__gold , \__mp_sa11_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[0]$_DFF_P_.CLK__assert (\__mp_sa12_sr[0]$_DFF_P_.CLK__gold , \__mp_sa12_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[1]$_DFF_P_.CLK__assert (\__mp_sa12_sr[1]$_DFF_P_.CLK__gold , \__mp_sa12_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[2]$_DFF_P_.CLK__assert (\__mp_sa12_sr[2]$_DFF_P_.CLK__gold , \__mp_sa12_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[3]$_DFF_P_.CLK__assert (\__mp_sa12_sr[3]$_DFF_P_.CLK__gold , \__mp_sa12_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[4]$_DFF_P_.CLK__assert (\__mp_sa12_sr[4]$_DFF_P_.CLK__gold , \__mp_sa12_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[5]$_DFF_P_.CLK__assert (\__mp_sa12_sr[5]$_DFF_P_.CLK__gold , \__mp_sa12_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[6]$_DFF_P_.CLK__assert (\__mp_sa12_sr[6]$_DFF_P_.CLK__gold , \__mp_sa12_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa12_sr[7]$_DFF_P_.CLK__assert (\__mp_sa12_sr[7]$_DFF_P_.CLK__gold , \__mp_sa12_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[0]$_DFF_P_.CLK__assert (\__mp_sa13_sr[0]$_DFF_P_.CLK__gold , \__mp_sa13_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[1]$_DFF_P_.CLK__assert (\__mp_sa13_sr[1]$_DFF_P_.CLK__gold , \__mp_sa13_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[2]$_DFF_P_.CLK__assert (\__mp_sa13_sr[2]$_DFF_P_.CLK__gold , \__mp_sa13_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[3]$_DFF_P_.CLK__assert (\__mp_sa13_sr[3]$_DFF_P_.CLK__gold , \__mp_sa13_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[4]$_DFF_P_.CLK__assert (\__mp_sa13_sr[4]$_DFF_P_.CLK__gold , \__mp_sa13_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[5]$_DFF_P_.CLK__assert (\__mp_sa13_sr[5]$_DFF_P_.CLK__gold , \__mp_sa13_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[6]$_DFF_P_.CLK__assert (\__mp_sa13_sr[6]$_DFF_P_.CLK__gold , \__mp_sa13_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa13_sr[7]$_DFF_P_.CLK__assert (\__mp_sa13_sr[7]$_DFF_P_.CLK__gold , \__mp_sa13_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[0]$_DFF_P_.CLK__assert (\__mp_sa20_sr[0]$_DFF_P_.CLK__gold , \__mp_sa20_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[1]$_DFF_P_.CLK__assert (\__mp_sa20_sr[1]$_DFF_P_.CLK__gold , \__mp_sa20_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[2]$_DFF_P_.CLK__assert (\__mp_sa20_sr[2]$_DFF_P_.CLK__gold , \__mp_sa20_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[3]$_DFF_P_.CLK__assert (\__mp_sa20_sr[3]$_DFF_P_.CLK__gold , \__mp_sa20_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[4]$_DFF_P_.CLK__assert (\__mp_sa20_sr[4]$_DFF_P_.CLK__gold , \__mp_sa20_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[5]$_DFF_P_.CLK__assert (\__mp_sa20_sr[5]$_DFF_P_.CLK__gold , \__mp_sa20_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[6]$_DFF_P_.CLK__assert (\__mp_sa20_sr[6]$_DFF_P_.CLK__gold , \__mp_sa20_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa20_sr[7]$_DFF_P_.CLK__assert (\__mp_sa20_sr[7]$_DFF_P_.CLK__gold , \__mp_sa20_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[0]$_DFF_P_.CLK__assert (\__mp_sa21_sr[0]$_DFF_P_.CLK__gold , \__mp_sa21_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[1]$_DFF_P_.CLK__assert (\__mp_sa21_sr[1]$_DFF_P_.CLK__gold , \__mp_sa21_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[2]$_DFF_P_.CLK__assert (\__mp_sa21_sr[2]$_DFF_P_.CLK__gold , \__mp_sa21_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[3]$_DFF_P_.CLK__assert (\__mp_sa21_sr[3]$_DFF_P_.CLK__gold , \__mp_sa21_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[4]$_DFF_P_.CLK__assert (\__mp_sa21_sr[4]$_DFF_P_.CLK__gold , \__mp_sa21_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[5]$_DFF_P_.CLK__assert (\__mp_sa21_sr[5]$_DFF_P_.CLK__gold , \__mp_sa21_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[6]$_DFF_P_.CLK__assert (\__mp_sa21_sr[6]$_DFF_P_.CLK__gold , \__mp_sa21_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa21_sr[7]$_DFF_P_.CLK__assert (\__mp_sa21_sr[7]$_DFF_P_.CLK__gold , \__mp_sa21_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[0]$_DFF_P_.CLK__assert (\__mp_sa22_sr[0]$_DFF_P_.CLK__gold , \__mp_sa22_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[1]$_DFF_P_.CLK__assert (\__mp_sa22_sr[1]$_DFF_P_.CLK__gold , \__mp_sa22_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[2]$_DFF_P_.CLK__assert (\__mp_sa22_sr[2]$_DFF_P_.CLK__gold , \__mp_sa22_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[3]$_DFF_P_.CLK__assert (\__mp_sa22_sr[3]$_DFF_P_.CLK__gold , \__mp_sa22_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[4]$_DFF_P_.CLK__assert (\__mp_sa22_sr[4]$_DFF_P_.CLK__gold , \__mp_sa22_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[5]$_DFF_P_.CLK__assert (\__mp_sa22_sr[5]$_DFF_P_.CLK__gold , \__mp_sa22_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[6]$_DFF_P_.CLK__assert (\__mp_sa22_sr[6]$_DFF_P_.CLK__gold , \__mp_sa22_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa22_sr[7]$_DFF_P_.CLK__assert (\__mp_sa22_sr[7]$_DFF_P_.CLK__gold , \__mp_sa22_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[0]$_DFF_P_.CLK__assert (\__mp_sa23_sr[0]$_DFF_P_.CLK__gold , \__mp_sa23_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[1]$_DFF_P_.CLK__assert (\__mp_sa23_sr[1]$_DFF_P_.CLK__gold , \__mp_sa23_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[2]$_DFF_P_.CLK__assert (\__mp_sa23_sr[2]$_DFF_P_.CLK__gold , \__mp_sa23_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[3]$_DFF_P_.CLK__assert (\__mp_sa23_sr[3]$_DFF_P_.CLK__gold , \__mp_sa23_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[4]$_DFF_P_.CLK__assert (\__mp_sa23_sr[4]$_DFF_P_.CLK__gold , \__mp_sa23_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[5]$_DFF_P_.CLK__assert (\__mp_sa23_sr[5]$_DFF_P_.CLK__gold , \__mp_sa23_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[6]$_DFF_P_.CLK__assert (\__mp_sa23_sr[6]$_DFF_P_.CLK__gold , \__mp_sa23_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa23_sr[7]$_DFF_P_.CLK__assert (\__mp_sa23_sr[7]$_DFF_P_.CLK__gold , \__mp_sa23_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[0]$_DFF_P_.CLK__assert (\__mp_sa30_sr[0]$_DFF_P_.CLK__gold , \__mp_sa30_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[1]$_DFF_P_.CLK__assert (\__mp_sa30_sr[1]$_DFF_P_.CLK__gold , \__mp_sa30_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[2]$_DFF_P_.CLK__assert (\__mp_sa30_sr[2]$_DFF_P_.CLK__gold , \__mp_sa30_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[3]$_DFF_P_.CLK__assert (\__mp_sa30_sr[3]$_DFF_P_.CLK__gold , \__mp_sa30_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[4]$_DFF_P_.CLK__assert (\__mp_sa30_sr[4]$_DFF_P_.CLK__gold , \__mp_sa30_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[5]$_DFF_P_.CLK__assert (\__mp_sa30_sr[5]$_DFF_P_.CLK__gold , \__mp_sa30_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[6]$_DFF_P_.CLK__assert (\__mp_sa30_sr[6]$_DFF_P_.CLK__gold , \__mp_sa30_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa30_sr[7]$_DFF_P_.CLK__assert (\__mp_sa30_sr[7]$_DFF_P_.CLK__gold , \__mp_sa30_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[0]$_DFF_P_.CLK__assert (\__mp_sa31_sr[0]$_DFF_P_.CLK__gold , \__mp_sa31_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[1]$_DFF_P_.CLK__assert (\__mp_sa31_sr[1]$_DFF_P_.CLK__gold , \__mp_sa31_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[2]$_DFF_P_.CLK__assert (\__mp_sa31_sr[2]$_DFF_P_.CLK__gold , \__mp_sa31_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[3]$_DFF_P_.CLK__assert (\__mp_sa31_sr[3]$_DFF_P_.CLK__gold , \__mp_sa31_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[4]$_DFF_P_.CLK__assert (\__mp_sa31_sr[4]$_DFF_P_.CLK__gold , \__mp_sa31_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[5]$_DFF_P_.CLK__assert (\__mp_sa31_sr[5]$_DFF_P_.CLK__gold , \__mp_sa31_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[6]$_DFF_P_.CLK__assert (\__mp_sa31_sr[6]$_DFF_P_.CLK__gold , \__mp_sa31_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa31_sr[7]$_DFF_P_.CLK__assert (\__mp_sa31_sr[7]$_DFF_P_.CLK__gold , \__mp_sa31_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[0]$_DFF_P_.CLK__assert (\__mp_sa32_sr[0]$_DFF_P_.CLK__gold , \__mp_sa32_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[1]$_DFF_P_.CLK__assert (\__mp_sa32_sr[1]$_DFF_P_.CLK__gold , \__mp_sa32_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[2]$_DFF_P_.CLK__assert (\__mp_sa32_sr[2]$_DFF_P_.CLK__gold , \__mp_sa32_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[3]$_DFF_P_.CLK__assert (\__mp_sa32_sr[3]$_DFF_P_.CLK__gold , \__mp_sa32_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[4]$_DFF_P_.CLK__assert (\__mp_sa32_sr[4]$_DFF_P_.CLK__gold , \__mp_sa32_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[5]$_DFF_P_.CLK__assert (\__mp_sa32_sr[5]$_DFF_P_.CLK__gold , \__mp_sa32_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[6]$_DFF_P_.CLK__assert (\__mp_sa32_sr[6]$_DFF_P_.CLK__gold , \__mp_sa32_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa32_sr[7]$_DFF_P_.CLK__assert (\__mp_sa32_sr[7]$_DFF_P_.CLK__gold , \__mp_sa32_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[0]$_DFF_P_.CLK__assert (\__mp_sa33_sr[0]$_DFF_P_.CLK__gold , \__mp_sa33_sr[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[1]$_DFF_P_.CLK__assert (\__mp_sa33_sr[1]$_DFF_P_.CLK__gold , \__mp_sa33_sr[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[2]$_DFF_P_.CLK__assert (\__mp_sa33_sr[2]$_DFF_P_.CLK__gold , \__mp_sa33_sr[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[3]$_DFF_P_.CLK__assert (\__mp_sa33_sr[3]$_DFF_P_.CLK__gold , \__mp_sa33_sr[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[4]$_DFF_P_.CLK__assert (\__mp_sa33_sr[4]$_DFF_P_.CLK__gold , \__mp_sa33_sr[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[5]$_DFF_P_.CLK__assert (\__mp_sa33_sr[5]$_DFF_P_.CLK__gold , \__mp_sa33_sr[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[6]$_DFF_P_.CLK__assert (\__mp_sa33_sr[6]$_DFF_P_.CLK__gold , \__mp_sa33_sr[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_sa33_sr[7]$_DFF_P_.CLK__assert (\__mp_sa33_sr[7]$_DFF_P_.CLK__gold , \__mp_sa33_sr[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[0]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[0]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[0]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[100]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[100]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[100]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[101]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[101]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[101]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[102]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[102]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[102]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[103]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[103]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[103]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[104]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[104]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[104]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[105]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[105]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[105]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[106]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[106]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[106]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[107]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[107]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[107]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[108]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[108]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[108]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[109]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[109]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[109]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[10]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[10]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[10]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[110]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[110]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[110]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[111]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[111]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[111]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[112]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[112]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[112]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[113]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[113]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[113]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[114]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[114]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[114]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[115]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[115]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[115]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[116]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[116]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[116]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[117]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[117]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[117]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[118]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[118]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[118]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[119]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[119]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[119]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[11]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[11]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[11]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[120]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[120]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[120]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[121]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[121]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[121]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[122]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[122]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[122]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[123]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[123]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[123]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[124]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[124]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[124]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[125]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[125]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[125]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[126]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[126]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[126]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[127]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[127]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[127]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[12]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[12]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[12]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[13]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[13]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[13]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[14]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[14]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[14]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[15]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[15]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[15]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[16]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[16]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[16]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[17]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[17]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[17]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[18]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[18]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[18]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[19]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[19]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[19]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[1]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[1]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[1]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[20]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[20]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[20]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[21]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[21]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[21]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[22]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[22]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[22]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[23]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[23]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[23]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[24]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[24]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[24]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[25]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[25]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[25]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[26]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[26]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[26]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[27]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[27]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[27]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[28]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[28]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[28]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[29]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[29]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[29]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[2]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[2]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[2]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[30]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[30]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[30]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[31]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[31]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[31]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[32]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[32]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[32]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[33]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[33]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[33]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[34]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[34]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[34]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[35]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[35]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[35]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[36]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[36]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[36]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[37]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[37]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[37]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[38]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[38]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[38]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[39]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[39]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[39]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[3]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[3]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[3]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[40]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[40]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[40]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[41]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[41]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[41]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[42]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[42]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[42]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[43]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[43]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[43]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[44]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[44]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[44]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[45]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[45]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[45]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[46]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[46]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[46]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[47]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[47]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[47]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[48]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[48]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[48]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[49]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[49]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[49]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[4]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[4]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[4]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[50]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[50]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[50]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[51]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[51]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[51]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[52]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[52]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[52]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[53]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[53]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[53]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[54]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[54]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[54]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[55]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[55]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[55]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[56]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[56]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[56]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[57]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[57]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[57]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[58]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[58]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[58]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[59]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[59]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[59]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[5]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[5]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[5]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[60]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[60]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[60]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[61]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[61]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[61]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[62]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[62]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[62]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[63]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[63]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[63]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[64]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[64]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[64]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[65]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[65]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[65]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[66]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[66]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[66]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[67]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[67]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[67]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[68]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[68]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[68]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[69]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[69]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[69]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[6]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[6]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[6]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[70]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[70]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[70]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[71]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[71]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[71]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[72]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[72]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[72]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[73]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[73]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[73]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[74]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[74]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[74]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[75]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[75]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[75]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[76]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[76]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[76]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[77]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[77]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[77]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[78]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[78]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[78]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[79]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[79]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[79]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[7]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[7]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[7]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[80]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[80]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[80]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[81]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[81]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[81]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[82]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[82]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[82]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[83]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[83]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[83]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[84]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[84]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[84]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[85]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[85]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[85]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[86]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[86]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[86]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[87]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[87]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[87]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[88]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[88]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[88]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[89]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[89]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[89]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[8]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[8]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[8]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[90]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[90]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[90]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[91]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[91]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[91]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[92]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[92]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[92]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[93]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[93]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[93]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[94]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[94]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[94]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[95]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[95]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[95]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[96]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[96]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[96]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[97]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[97]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[97]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[98]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[98]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[98]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[99]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[99]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[99]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_in_r[9]$_DFFE_PP_.CLK__assert (\__mp_text_in_r[9]$_DFFE_PP_.CLK__gold , \__mp_text_in_r[9]$_DFFE_PP_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[0]$_DFF_P_.CLK__assert (\__mp_text_out[0]$_DFF_P_.CLK__gold , \__mp_text_out[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[0]$_DFF_P_.QN__assert (\__mp_text_out[0]$_DFF_P_.QN__gold , \__mp_text_out[0]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[0]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[100]$_DFF_P_.CLK__assert (\__mp_text_out[100]$_DFF_P_.CLK__gold , \__mp_text_out[100]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[100]$_DFF_P_.QN__assert (\__mp_text_out[100]$_DFF_P_.QN__gold , \__mp_text_out[100]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[100]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[101]$_DFF_P_.CLK__assert (\__mp_text_out[101]$_DFF_P_.CLK__gold , \__mp_text_out[101]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[101]$_DFF_P_.QN__assert (\__mp_text_out[101]$_DFF_P_.QN__gold , \__mp_text_out[101]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[101]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[102]$_DFF_P_.CLK__assert (\__mp_text_out[102]$_DFF_P_.CLK__gold , \__mp_text_out[102]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[102]$_DFF_P_.QN__assert (\__mp_text_out[102]$_DFF_P_.QN__gold , \__mp_text_out[102]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[102]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[103]$_DFF_P_.CLK__assert (\__mp_text_out[103]$_DFF_P_.CLK__gold , \__mp_text_out[103]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[103]$_DFF_P_.QN__assert (\__mp_text_out[103]$_DFF_P_.QN__gold , \__mp_text_out[103]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[103]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[104]$_DFF_P_.CLK__assert (\__mp_text_out[104]$_DFF_P_.CLK__gold , \__mp_text_out[104]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[104]$_DFF_P_.QN__assert (\__mp_text_out[104]$_DFF_P_.QN__gold , \__mp_text_out[104]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[104]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[105]$_DFF_P_.CLK__assert (\__mp_text_out[105]$_DFF_P_.CLK__gold , \__mp_text_out[105]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[105]$_DFF_P_.QN__assert (\__mp_text_out[105]$_DFF_P_.QN__gold , \__mp_text_out[105]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[105]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[106]$_DFF_P_.CLK__assert (\__mp_text_out[106]$_DFF_P_.CLK__gold , \__mp_text_out[106]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[106]$_DFF_P_.QN__assert (\__mp_text_out[106]$_DFF_P_.QN__gold , \__mp_text_out[106]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[106]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[107]$_DFF_P_.CLK__assert (\__mp_text_out[107]$_DFF_P_.CLK__gold , \__mp_text_out[107]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[107]$_DFF_P_.QN__assert (\__mp_text_out[107]$_DFF_P_.QN__gold , \__mp_text_out[107]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[107]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[108]$_DFF_P_.CLK__assert (\__mp_text_out[108]$_DFF_P_.CLK__gold , \__mp_text_out[108]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[108]$_DFF_P_.QN__assert (\__mp_text_out[108]$_DFF_P_.QN__gold , \__mp_text_out[108]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[108]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[109]$_DFF_P_.CLK__assert (\__mp_text_out[109]$_DFF_P_.CLK__gold , \__mp_text_out[109]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[109]$_DFF_P_.QN__assert (\__mp_text_out[109]$_DFF_P_.QN__gold , \__mp_text_out[109]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[109]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[10]$_DFF_P_.CLK__assert (\__mp_text_out[10]$_DFF_P_.CLK__gold , \__mp_text_out[10]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[10]$_DFF_P_.QN__assert (\__mp_text_out[10]$_DFF_P_.QN__gold , \__mp_text_out[10]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[10]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[110]$_DFF_P_.CLK__assert (\__mp_text_out[110]$_DFF_P_.CLK__gold , \__mp_text_out[110]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[110]$_DFF_P_.QN__assert (\__mp_text_out[110]$_DFF_P_.QN__gold , \__mp_text_out[110]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[110]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[111]$_DFF_P_.CLK__assert (\__mp_text_out[111]$_DFF_P_.CLK__gold , \__mp_text_out[111]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[111]$_DFF_P_.QN__assert (\__mp_text_out[111]$_DFF_P_.QN__gold , \__mp_text_out[111]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[111]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[112]$_DFF_P_.CLK__assert (\__mp_text_out[112]$_DFF_P_.CLK__gold , \__mp_text_out[112]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[112]$_DFF_P_.QN__assert (\__mp_text_out[112]$_DFF_P_.QN__gold , \__mp_text_out[112]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[112]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[113]$_DFF_P_.CLK__assert (\__mp_text_out[113]$_DFF_P_.CLK__gold , \__mp_text_out[113]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[113]$_DFF_P_.QN__assert (\__mp_text_out[113]$_DFF_P_.QN__gold , \__mp_text_out[113]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[113]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[114]$_DFF_P_.CLK__assert (\__mp_text_out[114]$_DFF_P_.CLK__gold , \__mp_text_out[114]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[114]$_DFF_P_.QN__assert (\__mp_text_out[114]$_DFF_P_.QN__gold , \__mp_text_out[114]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[114]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[115]$_DFF_P_.CLK__assert (\__mp_text_out[115]$_DFF_P_.CLK__gold , \__mp_text_out[115]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[115]$_DFF_P_.QN__assert (\__mp_text_out[115]$_DFF_P_.QN__gold , \__mp_text_out[115]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[115]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[116]$_DFF_P_.CLK__assert (\__mp_text_out[116]$_DFF_P_.CLK__gold , \__mp_text_out[116]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[116]$_DFF_P_.QN__assert (\__mp_text_out[116]$_DFF_P_.QN__gold , \__mp_text_out[116]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[116]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[117]$_DFF_P_.CLK__assert (\__mp_text_out[117]$_DFF_P_.CLK__gold , \__mp_text_out[117]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[117]$_DFF_P_.QN__assert (\__mp_text_out[117]$_DFF_P_.QN__gold , \__mp_text_out[117]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[117]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[118]$_DFF_P_.CLK__assert (\__mp_text_out[118]$_DFF_P_.CLK__gold , \__mp_text_out[118]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[118]$_DFF_P_.QN__assert (\__mp_text_out[118]$_DFF_P_.QN__gold , \__mp_text_out[118]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[118]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[119]$_DFF_P_.CLK__assert (\__mp_text_out[119]$_DFF_P_.CLK__gold , \__mp_text_out[119]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[119]$_DFF_P_.QN__assert (\__mp_text_out[119]$_DFF_P_.QN__gold , \__mp_text_out[119]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[119]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[11]$_DFF_P_.CLK__assert (\__mp_text_out[11]$_DFF_P_.CLK__gold , \__mp_text_out[11]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[11]$_DFF_P_.QN__assert (\__mp_text_out[11]$_DFF_P_.QN__gold , \__mp_text_out[11]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[11]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[120]$_DFF_P_.CLK__assert (\__mp_text_out[120]$_DFF_P_.CLK__gold , \__mp_text_out[120]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[120]$_DFF_P_.QN__assert (\__mp_text_out[120]$_DFF_P_.QN__gold , \__mp_text_out[120]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[120]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[121]$_DFF_P_.CLK__assert (\__mp_text_out[121]$_DFF_P_.CLK__gold , \__mp_text_out[121]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[121]$_DFF_P_.QN__assert (\__mp_text_out[121]$_DFF_P_.QN__gold , \__mp_text_out[121]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[121]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[122]$_DFF_P_.CLK__assert (\__mp_text_out[122]$_DFF_P_.CLK__gold , \__mp_text_out[122]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[122]$_DFF_P_.QN__assert (\__mp_text_out[122]$_DFF_P_.QN__gold , \__mp_text_out[122]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[122]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[123]$_DFF_P_.CLK__assert (\__mp_text_out[123]$_DFF_P_.CLK__gold , \__mp_text_out[123]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[123]$_DFF_P_.QN__assert (\__mp_text_out[123]$_DFF_P_.QN__gold , \__mp_text_out[123]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[123]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[124]$_DFF_P_.CLK__assert (\__mp_text_out[124]$_DFF_P_.CLK__gold , \__mp_text_out[124]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[124]$_DFF_P_.QN__assert (\__mp_text_out[124]$_DFF_P_.QN__gold , \__mp_text_out[124]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[124]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[125]$_DFF_P_.CLK__assert (\__mp_text_out[125]$_DFF_P_.CLK__gold , \__mp_text_out[125]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[125]$_DFF_P_.QN__assert (\__mp_text_out[125]$_DFF_P_.QN__gold , \__mp_text_out[125]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[125]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[126]$_DFF_P_.CLK__assert (\__mp_text_out[126]$_DFF_P_.CLK__gold , \__mp_text_out[126]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[126]$_DFF_P_.QN__assert (\__mp_text_out[126]$_DFF_P_.QN__gold , \__mp_text_out[126]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[126]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[127]$_DFF_P_.CLK__assert (\__mp_text_out[127]$_DFF_P_.CLK__gold , \__mp_text_out[127]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[127]$_DFF_P_.QN__assert (\__mp_text_out[127]$_DFF_P_.QN__gold , \__mp_text_out[127]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[127]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[12]$_DFF_P_.CLK__assert (\__mp_text_out[12]$_DFF_P_.CLK__gold , \__mp_text_out[12]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[12]$_DFF_P_.QN__assert (\__mp_text_out[12]$_DFF_P_.QN__gold , \__mp_text_out[12]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[12]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[13]$_DFF_P_.CLK__assert (\__mp_text_out[13]$_DFF_P_.CLK__gold , \__mp_text_out[13]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[13]$_DFF_P_.QN__assert (\__mp_text_out[13]$_DFF_P_.QN__gold , \__mp_text_out[13]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[13]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[14]$_DFF_P_.CLK__assert (\__mp_text_out[14]$_DFF_P_.CLK__gold , \__mp_text_out[14]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[14]$_DFF_P_.QN__assert (\__mp_text_out[14]$_DFF_P_.QN__gold , \__mp_text_out[14]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[14]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[15]$_DFF_P_.CLK__assert (\__mp_text_out[15]$_DFF_P_.CLK__gold , \__mp_text_out[15]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[15]$_DFF_P_.QN__assert (\__mp_text_out[15]$_DFF_P_.QN__gold , \__mp_text_out[15]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[15]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[16]$_DFF_P_.CLK__assert (\__mp_text_out[16]$_DFF_P_.CLK__gold , \__mp_text_out[16]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[16]$_DFF_P_.QN__assert (\__mp_text_out[16]$_DFF_P_.QN__gold , \__mp_text_out[16]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[16]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[17]$_DFF_P_.CLK__assert (\__mp_text_out[17]$_DFF_P_.CLK__gold , \__mp_text_out[17]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[17]$_DFF_P_.QN__assert (\__mp_text_out[17]$_DFF_P_.QN__gold , \__mp_text_out[17]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[17]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[18]$_DFF_P_.CLK__assert (\__mp_text_out[18]$_DFF_P_.CLK__gold , \__mp_text_out[18]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[18]$_DFF_P_.QN__assert (\__mp_text_out[18]$_DFF_P_.QN__gold , \__mp_text_out[18]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[18]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[19]$_DFF_P_.CLK__assert (\__mp_text_out[19]$_DFF_P_.CLK__gold , \__mp_text_out[19]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[19]$_DFF_P_.QN__assert (\__mp_text_out[19]$_DFF_P_.QN__gold , \__mp_text_out[19]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[19]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[1]$_DFF_P_.CLK__assert (\__mp_text_out[1]$_DFF_P_.CLK__gold , \__mp_text_out[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[1]$_DFF_P_.QN__assert (\__mp_text_out[1]$_DFF_P_.QN__gold , \__mp_text_out[1]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[1]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[20]$_DFF_P_.CLK__assert (\__mp_text_out[20]$_DFF_P_.CLK__gold , \__mp_text_out[20]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[20]$_DFF_P_.QN__assert (\__mp_text_out[20]$_DFF_P_.QN__gold , \__mp_text_out[20]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[20]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[21]$_DFF_P_.CLK__assert (\__mp_text_out[21]$_DFF_P_.CLK__gold , \__mp_text_out[21]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[21]$_DFF_P_.QN__assert (\__mp_text_out[21]$_DFF_P_.QN__gold , \__mp_text_out[21]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[21]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[22]$_DFF_P_.CLK__assert (\__mp_text_out[22]$_DFF_P_.CLK__gold , \__mp_text_out[22]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[22]$_DFF_P_.QN__assert (\__mp_text_out[22]$_DFF_P_.QN__gold , \__mp_text_out[22]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[22]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[23]$_DFF_P_.CLK__assert (\__mp_text_out[23]$_DFF_P_.CLK__gold , \__mp_text_out[23]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[23]$_DFF_P_.QN__assert (\__mp_text_out[23]$_DFF_P_.QN__gold , \__mp_text_out[23]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[23]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[24]$_DFF_P_.CLK__assert (\__mp_text_out[24]$_DFF_P_.CLK__gold , \__mp_text_out[24]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[24]$_DFF_P_.QN__assert (\__mp_text_out[24]$_DFF_P_.QN__gold , \__mp_text_out[24]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[24]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[25]$_DFF_P_.CLK__assert (\__mp_text_out[25]$_DFF_P_.CLK__gold , \__mp_text_out[25]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[25]$_DFF_P_.QN__assert (\__mp_text_out[25]$_DFF_P_.QN__gold , \__mp_text_out[25]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[25]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[26]$_DFF_P_.CLK__assert (\__mp_text_out[26]$_DFF_P_.CLK__gold , \__mp_text_out[26]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[26]$_DFF_P_.QN__assert (\__mp_text_out[26]$_DFF_P_.QN__gold , \__mp_text_out[26]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[26]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[27]$_DFF_P_.CLK__assert (\__mp_text_out[27]$_DFF_P_.CLK__gold , \__mp_text_out[27]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[27]$_DFF_P_.QN__assert (\__mp_text_out[27]$_DFF_P_.QN__gold , \__mp_text_out[27]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[27]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[28]$_DFF_P_.CLK__assert (\__mp_text_out[28]$_DFF_P_.CLK__gold , \__mp_text_out[28]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[28]$_DFF_P_.QN__assert (\__mp_text_out[28]$_DFF_P_.QN__gold , \__mp_text_out[28]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[28]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[29]$_DFF_P_.CLK__assert (\__mp_text_out[29]$_DFF_P_.CLK__gold , \__mp_text_out[29]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[29]$_DFF_P_.QN__assert (\__mp_text_out[29]$_DFF_P_.QN__gold , \__mp_text_out[29]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[29]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[2]$_DFF_P_.CLK__assert (\__mp_text_out[2]$_DFF_P_.CLK__gold , \__mp_text_out[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[2]$_DFF_P_.QN__assert (\__mp_text_out[2]$_DFF_P_.QN__gold , \__mp_text_out[2]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[2]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[30]$_DFF_P_.CLK__assert (\__mp_text_out[30]$_DFF_P_.CLK__gold , \__mp_text_out[30]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[30]$_DFF_P_.QN__assert (\__mp_text_out[30]$_DFF_P_.QN__gold , \__mp_text_out[30]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[30]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[31]$_DFF_P_.CLK__assert (\__mp_text_out[31]$_DFF_P_.CLK__gold , \__mp_text_out[31]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[31]$_DFF_P_.QN__assert (\__mp_text_out[31]$_DFF_P_.QN__gold , \__mp_text_out[31]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[31]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[32]$_DFF_P_.CLK__assert (\__mp_text_out[32]$_DFF_P_.CLK__gold , \__mp_text_out[32]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[32]$_DFF_P_.QN__assert (\__mp_text_out[32]$_DFF_P_.QN__gold , \__mp_text_out[32]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[32]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[33]$_DFF_P_.CLK__assert (\__mp_text_out[33]$_DFF_P_.CLK__gold , \__mp_text_out[33]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[33]$_DFF_P_.QN__assert (\__mp_text_out[33]$_DFF_P_.QN__gold , \__mp_text_out[33]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[33]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[34]$_DFF_P_.CLK__assert (\__mp_text_out[34]$_DFF_P_.CLK__gold , \__mp_text_out[34]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[34]$_DFF_P_.QN__assert (\__mp_text_out[34]$_DFF_P_.QN__gold , \__mp_text_out[34]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[34]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[35]$_DFF_P_.CLK__assert (\__mp_text_out[35]$_DFF_P_.CLK__gold , \__mp_text_out[35]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[35]$_DFF_P_.QN__assert (\__mp_text_out[35]$_DFF_P_.QN__gold , \__mp_text_out[35]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[35]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[36]$_DFF_P_.CLK__assert (\__mp_text_out[36]$_DFF_P_.CLK__gold , \__mp_text_out[36]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[36]$_DFF_P_.QN__assert (\__mp_text_out[36]$_DFF_P_.QN__gold , \__mp_text_out[36]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[36]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[37]$_DFF_P_.CLK__assert (\__mp_text_out[37]$_DFF_P_.CLK__gold , \__mp_text_out[37]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[37]$_DFF_P_.QN__assert (\__mp_text_out[37]$_DFF_P_.QN__gold , \__mp_text_out[37]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[37]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[38]$_DFF_P_.CLK__assert (\__mp_text_out[38]$_DFF_P_.CLK__gold , \__mp_text_out[38]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[38]$_DFF_P_.QN__assert (\__mp_text_out[38]$_DFF_P_.QN__gold , \__mp_text_out[38]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[38]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[39]$_DFF_P_.CLK__assert (\__mp_text_out[39]$_DFF_P_.CLK__gold , \__mp_text_out[39]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[39]$_DFF_P_.QN__assert (\__mp_text_out[39]$_DFF_P_.QN__gold , \__mp_text_out[39]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[39]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[3]$_DFF_P_.CLK__assert (\__mp_text_out[3]$_DFF_P_.CLK__gold , \__mp_text_out[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[3]$_DFF_P_.QN__assert (\__mp_text_out[3]$_DFF_P_.QN__gold , \__mp_text_out[3]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[3]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[40]$_DFF_P_.CLK__assert (\__mp_text_out[40]$_DFF_P_.CLK__gold , \__mp_text_out[40]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[40]$_DFF_P_.QN__assert (\__mp_text_out[40]$_DFF_P_.QN__gold , \__mp_text_out[40]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[40]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[41]$_DFF_P_.CLK__assert (\__mp_text_out[41]$_DFF_P_.CLK__gold , \__mp_text_out[41]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[41]$_DFF_P_.QN__assert (\__mp_text_out[41]$_DFF_P_.QN__gold , \__mp_text_out[41]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[41]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[42]$_DFF_P_.CLK__assert (\__mp_text_out[42]$_DFF_P_.CLK__gold , \__mp_text_out[42]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[42]$_DFF_P_.QN__assert (\__mp_text_out[42]$_DFF_P_.QN__gold , \__mp_text_out[42]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[42]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[43]$_DFF_P_.CLK__assert (\__mp_text_out[43]$_DFF_P_.CLK__gold , \__mp_text_out[43]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[43]$_DFF_P_.QN__assert (\__mp_text_out[43]$_DFF_P_.QN__gold , \__mp_text_out[43]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[43]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[44]$_DFF_P_.CLK__assert (\__mp_text_out[44]$_DFF_P_.CLK__gold , \__mp_text_out[44]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[44]$_DFF_P_.QN__assert (\__mp_text_out[44]$_DFF_P_.QN__gold , \__mp_text_out[44]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[44]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[45]$_DFF_P_.CLK__assert (\__mp_text_out[45]$_DFF_P_.CLK__gold , \__mp_text_out[45]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[45]$_DFF_P_.QN__assert (\__mp_text_out[45]$_DFF_P_.QN__gold , \__mp_text_out[45]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[45]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[46]$_DFF_P_.CLK__assert (\__mp_text_out[46]$_DFF_P_.CLK__gold , \__mp_text_out[46]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[46]$_DFF_P_.QN__assert (\__mp_text_out[46]$_DFF_P_.QN__gold , \__mp_text_out[46]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[46]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[47]$_DFF_P_.CLK__assert (\__mp_text_out[47]$_DFF_P_.CLK__gold , \__mp_text_out[47]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[47]$_DFF_P_.QN__assert (\__mp_text_out[47]$_DFF_P_.QN__gold , \__mp_text_out[47]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[47]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[48]$_DFF_P_.CLK__assert (\__mp_text_out[48]$_DFF_P_.CLK__gold , \__mp_text_out[48]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[48]$_DFF_P_.QN__assert (\__mp_text_out[48]$_DFF_P_.QN__gold , \__mp_text_out[48]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[48]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[49]$_DFF_P_.CLK__assert (\__mp_text_out[49]$_DFF_P_.CLK__gold , \__mp_text_out[49]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[49]$_DFF_P_.QN__assert (\__mp_text_out[49]$_DFF_P_.QN__gold , \__mp_text_out[49]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[49]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[4]$_DFF_P_.CLK__assert (\__mp_text_out[4]$_DFF_P_.CLK__gold , \__mp_text_out[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[4]$_DFF_P_.QN__assert (\__mp_text_out[4]$_DFF_P_.QN__gold , \__mp_text_out[4]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[4]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[50]$_DFF_P_.CLK__assert (\__mp_text_out[50]$_DFF_P_.CLK__gold , \__mp_text_out[50]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[50]$_DFF_P_.QN__assert (\__mp_text_out[50]$_DFF_P_.QN__gold , \__mp_text_out[50]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[50]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[51]$_DFF_P_.CLK__assert (\__mp_text_out[51]$_DFF_P_.CLK__gold , \__mp_text_out[51]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[51]$_DFF_P_.QN__assert (\__mp_text_out[51]$_DFF_P_.QN__gold , \__mp_text_out[51]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[51]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[52]$_DFF_P_.CLK__assert (\__mp_text_out[52]$_DFF_P_.CLK__gold , \__mp_text_out[52]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[52]$_DFF_P_.QN__assert (\__mp_text_out[52]$_DFF_P_.QN__gold , \__mp_text_out[52]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[52]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[53]$_DFF_P_.CLK__assert (\__mp_text_out[53]$_DFF_P_.CLK__gold , \__mp_text_out[53]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[53]$_DFF_P_.QN__assert (\__mp_text_out[53]$_DFF_P_.QN__gold , \__mp_text_out[53]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[53]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[54]$_DFF_P_.CLK__assert (\__mp_text_out[54]$_DFF_P_.CLK__gold , \__mp_text_out[54]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[54]$_DFF_P_.QN__assert (\__mp_text_out[54]$_DFF_P_.QN__gold , \__mp_text_out[54]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[54]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[55]$_DFF_P_.CLK__assert (\__mp_text_out[55]$_DFF_P_.CLK__gold , \__mp_text_out[55]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[55]$_DFF_P_.QN__assert (\__mp_text_out[55]$_DFF_P_.QN__gold , \__mp_text_out[55]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[55]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[56]$_DFF_P_.CLK__assert (\__mp_text_out[56]$_DFF_P_.CLK__gold , \__mp_text_out[56]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[56]$_DFF_P_.QN__assert (\__mp_text_out[56]$_DFF_P_.QN__gold , \__mp_text_out[56]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[56]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[57]$_DFF_P_.CLK__assert (\__mp_text_out[57]$_DFF_P_.CLK__gold , \__mp_text_out[57]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[57]$_DFF_P_.QN__assert (\__mp_text_out[57]$_DFF_P_.QN__gold , \__mp_text_out[57]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[57]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[58]$_DFF_P_.CLK__assert (\__mp_text_out[58]$_DFF_P_.CLK__gold , \__mp_text_out[58]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[58]$_DFF_P_.QN__assert (\__mp_text_out[58]$_DFF_P_.QN__gold , \__mp_text_out[58]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[58]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[59]$_DFF_P_.CLK__assert (\__mp_text_out[59]$_DFF_P_.CLK__gold , \__mp_text_out[59]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[59]$_DFF_P_.QN__assert (\__mp_text_out[59]$_DFF_P_.QN__gold , \__mp_text_out[59]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[59]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[5]$_DFF_P_.CLK__assert (\__mp_text_out[5]$_DFF_P_.CLK__gold , \__mp_text_out[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[5]$_DFF_P_.QN__assert (\__mp_text_out[5]$_DFF_P_.QN__gold , \__mp_text_out[5]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[5]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[60]$_DFF_P_.CLK__assert (\__mp_text_out[60]$_DFF_P_.CLK__gold , \__mp_text_out[60]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[60]$_DFF_P_.QN__assert (\__mp_text_out[60]$_DFF_P_.QN__gold , \__mp_text_out[60]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[60]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[61]$_DFF_P_.CLK__assert (\__mp_text_out[61]$_DFF_P_.CLK__gold , \__mp_text_out[61]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[61]$_DFF_P_.QN__assert (\__mp_text_out[61]$_DFF_P_.QN__gold , \__mp_text_out[61]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[61]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[62]$_DFF_P_.CLK__assert (\__mp_text_out[62]$_DFF_P_.CLK__gold , \__mp_text_out[62]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[62]$_DFF_P_.QN__assert (\__mp_text_out[62]$_DFF_P_.QN__gold , \__mp_text_out[62]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[62]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[63]$_DFF_P_.CLK__assert (\__mp_text_out[63]$_DFF_P_.CLK__gold , \__mp_text_out[63]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[63]$_DFF_P_.QN__assert (\__mp_text_out[63]$_DFF_P_.QN__gold , \__mp_text_out[63]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[63]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[64]$_DFF_P_.CLK__assert (\__mp_text_out[64]$_DFF_P_.CLK__gold , \__mp_text_out[64]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[64]$_DFF_P_.QN__assert (\__mp_text_out[64]$_DFF_P_.QN__gold , \__mp_text_out[64]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[64]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[65]$_DFF_P_.CLK__assert (\__mp_text_out[65]$_DFF_P_.CLK__gold , \__mp_text_out[65]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[65]$_DFF_P_.QN__assert (\__mp_text_out[65]$_DFF_P_.QN__gold , \__mp_text_out[65]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[65]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[66]$_DFF_P_.CLK__assert (\__mp_text_out[66]$_DFF_P_.CLK__gold , \__mp_text_out[66]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[66]$_DFF_P_.QN__assert (\__mp_text_out[66]$_DFF_P_.QN__gold , \__mp_text_out[66]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[66]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[67]$_DFF_P_.CLK__assert (\__mp_text_out[67]$_DFF_P_.CLK__gold , \__mp_text_out[67]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[67]$_DFF_P_.QN__assert (\__mp_text_out[67]$_DFF_P_.QN__gold , \__mp_text_out[67]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[67]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[68]$_DFF_P_.CLK__assert (\__mp_text_out[68]$_DFF_P_.CLK__gold , \__mp_text_out[68]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[68]$_DFF_P_.QN__assert (\__mp_text_out[68]$_DFF_P_.QN__gold , \__mp_text_out[68]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[68]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[69]$_DFF_P_.CLK__assert (\__mp_text_out[69]$_DFF_P_.CLK__gold , \__mp_text_out[69]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[69]$_DFF_P_.QN__assert (\__mp_text_out[69]$_DFF_P_.QN__gold , \__mp_text_out[69]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[69]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[6]$_DFF_P_.CLK__assert (\__mp_text_out[6]$_DFF_P_.CLK__gold , \__mp_text_out[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[6]$_DFF_P_.QN__assert (\__mp_text_out[6]$_DFF_P_.QN__gold , \__mp_text_out[6]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[6]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[70]$_DFF_P_.CLK__assert (\__mp_text_out[70]$_DFF_P_.CLK__gold , \__mp_text_out[70]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[70]$_DFF_P_.QN__assert (\__mp_text_out[70]$_DFF_P_.QN__gold , \__mp_text_out[70]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[70]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[71]$_DFF_P_.CLK__assert (\__mp_text_out[71]$_DFF_P_.CLK__gold , \__mp_text_out[71]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[71]$_DFF_P_.QN__assert (\__mp_text_out[71]$_DFF_P_.QN__gold , \__mp_text_out[71]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[71]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[72]$_DFF_P_.CLK__assert (\__mp_text_out[72]$_DFF_P_.CLK__gold , \__mp_text_out[72]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[72]$_DFF_P_.QN__assert (\__mp_text_out[72]$_DFF_P_.QN__gold , \__mp_text_out[72]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[72]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[73]$_DFF_P_.CLK__assert (\__mp_text_out[73]$_DFF_P_.CLK__gold , \__mp_text_out[73]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[73]$_DFF_P_.QN__assert (\__mp_text_out[73]$_DFF_P_.QN__gold , \__mp_text_out[73]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[73]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[74]$_DFF_P_.CLK__assert (\__mp_text_out[74]$_DFF_P_.CLK__gold , \__mp_text_out[74]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[74]$_DFF_P_.QN__assert (\__mp_text_out[74]$_DFF_P_.QN__gold , \__mp_text_out[74]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[74]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[75]$_DFF_P_.CLK__assert (\__mp_text_out[75]$_DFF_P_.CLK__gold , \__mp_text_out[75]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[75]$_DFF_P_.QN__assert (\__mp_text_out[75]$_DFF_P_.QN__gold , \__mp_text_out[75]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[75]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[76]$_DFF_P_.CLK__assert (\__mp_text_out[76]$_DFF_P_.CLK__gold , \__mp_text_out[76]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[76]$_DFF_P_.QN__assert (\__mp_text_out[76]$_DFF_P_.QN__gold , \__mp_text_out[76]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[76]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[77]$_DFF_P_.CLK__assert (\__mp_text_out[77]$_DFF_P_.CLK__gold , \__mp_text_out[77]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[77]$_DFF_P_.QN__assert (\__mp_text_out[77]$_DFF_P_.QN__gold , \__mp_text_out[77]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[77]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[78]$_DFF_P_.CLK__assert (\__mp_text_out[78]$_DFF_P_.CLK__gold , \__mp_text_out[78]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[78]$_DFF_P_.QN__assert (\__mp_text_out[78]$_DFF_P_.QN__gold , \__mp_text_out[78]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[78]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[79]$_DFF_P_.CLK__assert (\__mp_text_out[79]$_DFF_P_.CLK__gold , \__mp_text_out[79]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[79]$_DFF_P_.QN__assert (\__mp_text_out[79]$_DFF_P_.QN__gold , \__mp_text_out[79]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[79]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[7]$_DFF_P_.CLK__assert (\__mp_text_out[7]$_DFF_P_.CLK__gold , \__mp_text_out[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[7]$_DFF_P_.QN__assert (\__mp_text_out[7]$_DFF_P_.QN__gold , \__mp_text_out[7]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[7]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[80]$_DFF_P_.CLK__assert (\__mp_text_out[80]$_DFF_P_.CLK__gold , \__mp_text_out[80]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[80]$_DFF_P_.QN__assert (\__mp_text_out[80]$_DFF_P_.QN__gold , \__mp_text_out[80]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[80]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[81]$_DFF_P_.CLK__assert (\__mp_text_out[81]$_DFF_P_.CLK__gold , \__mp_text_out[81]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[81]$_DFF_P_.QN__assert (\__mp_text_out[81]$_DFF_P_.QN__gold , \__mp_text_out[81]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[81]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[82]$_DFF_P_.CLK__assert (\__mp_text_out[82]$_DFF_P_.CLK__gold , \__mp_text_out[82]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[82]$_DFF_P_.QN__assert (\__mp_text_out[82]$_DFF_P_.QN__gold , \__mp_text_out[82]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[82]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[83]$_DFF_P_.CLK__assert (\__mp_text_out[83]$_DFF_P_.CLK__gold , \__mp_text_out[83]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[83]$_DFF_P_.QN__assert (\__mp_text_out[83]$_DFF_P_.QN__gold , \__mp_text_out[83]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[83]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[84]$_DFF_P_.CLK__assert (\__mp_text_out[84]$_DFF_P_.CLK__gold , \__mp_text_out[84]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[84]$_DFF_P_.QN__assert (\__mp_text_out[84]$_DFF_P_.QN__gold , \__mp_text_out[84]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[84]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[85]$_DFF_P_.CLK__assert (\__mp_text_out[85]$_DFF_P_.CLK__gold , \__mp_text_out[85]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[85]$_DFF_P_.QN__assert (\__mp_text_out[85]$_DFF_P_.QN__gold , \__mp_text_out[85]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[85]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[86]$_DFF_P_.CLK__assert (\__mp_text_out[86]$_DFF_P_.CLK__gold , \__mp_text_out[86]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[86]$_DFF_P_.QN__assert (\__mp_text_out[86]$_DFF_P_.QN__gold , \__mp_text_out[86]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[86]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[87]$_DFF_P_.CLK__assert (\__mp_text_out[87]$_DFF_P_.CLK__gold , \__mp_text_out[87]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[87]$_DFF_P_.QN__assert (\__mp_text_out[87]$_DFF_P_.QN__gold , \__mp_text_out[87]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[87]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[88]$_DFF_P_.CLK__assert (\__mp_text_out[88]$_DFF_P_.CLK__gold , \__mp_text_out[88]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[88]$_DFF_P_.QN__assert (\__mp_text_out[88]$_DFF_P_.QN__gold , \__mp_text_out[88]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[88]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[89]$_DFF_P_.CLK__assert (\__mp_text_out[89]$_DFF_P_.CLK__gold , \__mp_text_out[89]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[89]$_DFF_P_.QN__assert (\__mp_text_out[89]$_DFF_P_.QN__gold , \__mp_text_out[89]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[89]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[8]$_DFF_P_.CLK__assert (\__mp_text_out[8]$_DFF_P_.CLK__gold , \__mp_text_out[8]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[8]$_DFF_P_.QN__assert (\__mp_text_out[8]$_DFF_P_.QN__gold , \__mp_text_out[8]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[8]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[90]$_DFF_P_.CLK__assert (\__mp_text_out[90]$_DFF_P_.CLK__gold , \__mp_text_out[90]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[90]$_DFF_P_.QN__assert (\__mp_text_out[90]$_DFF_P_.QN__gold , \__mp_text_out[90]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[90]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[91]$_DFF_P_.CLK__assert (\__mp_text_out[91]$_DFF_P_.CLK__gold , \__mp_text_out[91]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[91]$_DFF_P_.QN__assert (\__mp_text_out[91]$_DFF_P_.QN__gold , \__mp_text_out[91]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[91]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[92]$_DFF_P_.CLK__assert (\__mp_text_out[92]$_DFF_P_.CLK__gold , \__mp_text_out[92]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[92]$_DFF_P_.QN__assert (\__mp_text_out[92]$_DFF_P_.QN__gold , \__mp_text_out[92]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[92]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[93]$_DFF_P_.CLK__assert (\__mp_text_out[93]$_DFF_P_.CLK__gold , \__mp_text_out[93]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[93]$_DFF_P_.QN__assert (\__mp_text_out[93]$_DFF_P_.QN__gold , \__mp_text_out[93]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[93]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[94]$_DFF_P_.CLK__assert (\__mp_text_out[94]$_DFF_P_.CLK__gold , \__mp_text_out[94]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[94]$_DFF_P_.QN__assert (\__mp_text_out[94]$_DFF_P_.QN__gold , \__mp_text_out[94]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[94]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[95]$_DFF_P_.CLK__assert (\__mp_text_out[95]$_DFF_P_.CLK__gold , \__mp_text_out[95]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[95]$_DFF_P_.QN__assert (\__mp_text_out[95]$_DFF_P_.QN__gold , \__mp_text_out[95]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[95]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[96]$_DFF_P_.CLK__assert (\__mp_text_out[96]$_DFF_P_.CLK__gold , \__mp_text_out[96]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[96]$_DFF_P_.QN__assert (\__mp_text_out[96]$_DFF_P_.QN__gold , \__mp_text_out[96]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[96]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[97]$_DFF_P_.CLK__assert (\__mp_text_out[97]$_DFF_P_.CLK__gold , \__mp_text_out[97]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[97]$_DFF_P_.QN__assert (\__mp_text_out[97]$_DFF_P_.QN__gold , \__mp_text_out[97]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[97]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[98]$_DFF_P_.CLK__assert (\__mp_text_out[98]$_DFF_P_.CLK__gold , \__mp_text_out[98]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[98]$_DFF_P_.QN__assert (\__mp_text_out[98]$_DFF_P_.QN__gold , \__mp_text_out[98]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[98]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[99]$_DFF_P_.CLK__assert (\__mp_text_out[99]$_DFF_P_.CLK__gold , \__mp_text_out[99]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[99]$_DFF_P_.QN__assert (\__mp_text_out[99]$_DFF_P_.QN__gold , \__mp_text_out[99]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[99]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[9]$_DFF_P_.CLK__assert (\__mp_text_out[9]$_DFF_P_.CLK__gold , \__mp_text_out[9]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[9]$_DFF_P_.QN__assert (\__mp_text_out[9]$_DFF_P_.QN__gold , \__mp_text_out[9]$_DFF_P_.QN__gate );
  miter_cmp_prop #(1, "assert") \__mp_text_out[9]$_DFF_P_.int_fwire_IQN__assert (\__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gold , \__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__assert (\__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gold , \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__assert (\__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gold , \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[0]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[0]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[1]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[1]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[2]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[2]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[3]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[3]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[4]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[4]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[5]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[5]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[6]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[6]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u0.d[7]$_DFF_P_.CLK__assert (\__mp_u0.u0.d[7]$_DFF_P_.CLK__gold , \__mp_u0.u0.d[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[0]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[0]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[1]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[1]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[2]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[2]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[3]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[3]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[4]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[4]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[5]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[5]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[6]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[6]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u1.d[7]$_DFF_P_.CLK__assert (\__mp_u0.u1.d[7]$_DFF_P_.CLK__gold , \__mp_u0.u1.d[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[0]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[0]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[1]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[1]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[2]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[2]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[3]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[3]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[4]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[4]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[5]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[5]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[6]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[6]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u2.d[7]$_DFF_P_.CLK__assert (\__mp_u0.u2.d[7]$_DFF_P_.CLK__gold , \__mp_u0.u2.d[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[0]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[0]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[1]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[1]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[2]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[2]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[3]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[3]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[4]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[4]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[5]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[5]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[6]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[6]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.u3.d[7]$_DFF_P_.CLK__assert (\__mp_u0.u3.d[7]$_DFF_P_.CLK__gold , \__mp_u0.u3.d[7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][0]$_DFF_P_.CLK__assert (\__mp_u0.w[0][0]$_DFF_P_.CLK__gold , \__mp_u0.w[0][0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][10]$_DFF_P_.CLK__assert (\__mp_u0.w[0][10]$_DFF_P_.CLK__gold , \__mp_u0.w[0][10]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][11]$_DFF_P_.CLK__assert (\__mp_u0.w[0][11]$_DFF_P_.CLK__gold , \__mp_u0.w[0][11]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][12]$_DFF_P_.CLK__assert (\__mp_u0.w[0][12]$_DFF_P_.CLK__gold , \__mp_u0.w[0][12]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][13]$_DFF_P_.CLK__assert (\__mp_u0.w[0][13]$_DFF_P_.CLK__gold , \__mp_u0.w[0][13]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][14]$_DFF_P_.CLK__assert (\__mp_u0.w[0][14]$_DFF_P_.CLK__gold , \__mp_u0.w[0][14]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][15]$_DFF_P_.CLK__assert (\__mp_u0.w[0][15]$_DFF_P_.CLK__gold , \__mp_u0.w[0][15]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][16]$_DFF_P_.CLK__assert (\__mp_u0.w[0][16]$_DFF_P_.CLK__gold , \__mp_u0.w[0][16]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][17]$_DFF_P_.CLK__assert (\__mp_u0.w[0][17]$_DFF_P_.CLK__gold , \__mp_u0.w[0][17]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][18]$_DFF_P_.CLK__assert (\__mp_u0.w[0][18]$_DFF_P_.CLK__gold , \__mp_u0.w[0][18]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][19]$_DFF_P_.CLK__assert (\__mp_u0.w[0][19]$_DFF_P_.CLK__gold , \__mp_u0.w[0][19]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][1]$_DFF_P_.CLK__assert (\__mp_u0.w[0][1]$_DFF_P_.CLK__gold , \__mp_u0.w[0][1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][20]$_DFF_P_.CLK__assert (\__mp_u0.w[0][20]$_DFF_P_.CLK__gold , \__mp_u0.w[0][20]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][21]$_DFF_P_.CLK__assert (\__mp_u0.w[0][21]$_DFF_P_.CLK__gold , \__mp_u0.w[0][21]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][22]$_DFF_P_.CLK__assert (\__mp_u0.w[0][22]$_DFF_P_.CLK__gold , \__mp_u0.w[0][22]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][23]$_DFF_P_.CLK__assert (\__mp_u0.w[0][23]$_DFF_P_.CLK__gold , \__mp_u0.w[0][23]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][24]$_DFF_P_.CLK__assert (\__mp_u0.w[0][24]$_DFF_P_.CLK__gold , \__mp_u0.w[0][24]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][25]$_DFF_P_.CLK__assert (\__mp_u0.w[0][25]$_DFF_P_.CLK__gold , \__mp_u0.w[0][25]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][26]$_DFF_P_.CLK__assert (\__mp_u0.w[0][26]$_DFF_P_.CLK__gold , \__mp_u0.w[0][26]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][27]$_DFF_P_.CLK__assert (\__mp_u0.w[0][27]$_DFF_P_.CLK__gold , \__mp_u0.w[0][27]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][28]$_DFF_P_.CLK__assert (\__mp_u0.w[0][28]$_DFF_P_.CLK__gold , \__mp_u0.w[0][28]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][29]$_DFF_P_.CLK__assert (\__mp_u0.w[0][29]$_DFF_P_.CLK__gold , \__mp_u0.w[0][29]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][2]$_DFF_P_.CLK__assert (\__mp_u0.w[0][2]$_DFF_P_.CLK__gold , \__mp_u0.w[0][2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][30]$_DFF_P_.CLK__assert (\__mp_u0.w[0][30]$_DFF_P_.CLK__gold , \__mp_u0.w[0][30]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][31]$_DFF_P_.CLK__assert (\__mp_u0.w[0][31]$_DFF_P_.CLK__gold , \__mp_u0.w[0][31]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][3]$_DFF_P_.CLK__assert (\__mp_u0.w[0][3]$_DFF_P_.CLK__gold , \__mp_u0.w[0][3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][4]$_DFF_P_.CLK__assert (\__mp_u0.w[0][4]$_DFF_P_.CLK__gold , \__mp_u0.w[0][4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][5]$_DFF_P_.CLK__assert (\__mp_u0.w[0][5]$_DFF_P_.CLK__gold , \__mp_u0.w[0][5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][6]$_DFF_P_.CLK__assert (\__mp_u0.w[0][6]$_DFF_P_.CLK__gold , \__mp_u0.w[0][6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][7]$_DFF_P_.CLK__assert (\__mp_u0.w[0][7]$_DFF_P_.CLK__gold , \__mp_u0.w[0][7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][8]$_DFF_P_.CLK__assert (\__mp_u0.w[0][8]$_DFF_P_.CLK__gold , \__mp_u0.w[0][8]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[0][9]$_DFF_P_.CLK__assert (\__mp_u0.w[0][9]$_DFF_P_.CLK__gold , \__mp_u0.w[0][9]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][0]$_DFF_P_.CLK__assert (\__mp_u0.w[1][0]$_DFF_P_.CLK__gold , \__mp_u0.w[1][0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][10]$_DFF_P_.CLK__assert (\__mp_u0.w[1][10]$_DFF_P_.CLK__gold , \__mp_u0.w[1][10]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][11]$_DFF_P_.CLK__assert (\__mp_u0.w[1][11]$_DFF_P_.CLK__gold , \__mp_u0.w[1][11]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][12]$_DFF_P_.CLK__assert (\__mp_u0.w[1][12]$_DFF_P_.CLK__gold , \__mp_u0.w[1][12]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][13]$_DFF_P_.CLK__assert (\__mp_u0.w[1][13]$_DFF_P_.CLK__gold , \__mp_u0.w[1][13]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][14]$_DFF_P_.CLK__assert (\__mp_u0.w[1][14]$_DFF_P_.CLK__gold , \__mp_u0.w[1][14]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][15]$_DFF_P_.CLK__assert (\__mp_u0.w[1][15]$_DFF_P_.CLK__gold , \__mp_u0.w[1][15]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][16]$_DFF_P_.CLK__assert (\__mp_u0.w[1][16]$_DFF_P_.CLK__gold , \__mp_u0.w[1][16]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][17]$_DFF_P_.CLK__assert (\__mp_u0.w[1][17]$_DFF_P_.CLK__gold , \__mp_u0.w[1][17]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][18]$_DFF_P_.CLK__assert (\__mp_u0.w[1][18]$_DFF_P_.CLK__gold , \__mp_u0.w[1][18]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][19]$_DFF_P_.CLK__assert (\__mp_u0.w[1][19]$_DFF_P_.CLK__gold , \__mp_u0.w[1][19]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][1]$_DFF_P_.CLK__assert (\__mp_u0.w[1][1]$_DFF_P_.CLK__gold , \__mp_u0.w[1][1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][20]$_DFF_P_.CLK__assert (\__mp_u0.w[1][20]$_DFF_P_.CLK__gold , \__mp_u0.w[1][20]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][21]$_DFF_P_.CLK__assert (\__mp_u0.w[1][21]$_DFF_P_.CLK__gold , \__mp_u0.w[1][21]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][22]$_DFF_P_.CLK__assert (\__mp_u0.w[1][22]$_DFF_P_.CLK__gold , \__mp_u0.w[1][22]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][23]$_DFF_P_.CLK__assert (\__mp_u0.w[1][23]$_DFF_P_.CLK__gold , \__mp_u0.w[1][23]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][24]$_DFF_P_.CLK__assert (\__mp_u0.w[1][24]$_DFF_P_.CLK__gold , \__mp_u0.w[1][24]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][25]$_DFF_P_.CLK__assert (\__mp_u0.w[1][25]$_DFF_P_.CLK__gold , \__mp_u0.w[1][25]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][26]$_DFF_P_.CLK__assert (\__mp_u0.w[1][26]$_DFF_P_.CLK__gold , \__mp_u0.w[1][26]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][27]$_DFF_P_.CLK__assert (\__mp_u0.w[1][27]$_DFF_P_.CLK__gold , \__mp_u0.w[1][27]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][28]$_DFF_P_.CLK__assert (\__mp_u0.w[1][28]$_DFF_P_.CLK__gold , \__mp_u0.w[1][28]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][29]$_DFF_P_.CLK__assert (\__mp_u0.w[1][29]$_DFF_P_.CLK__gold , \__mp_u0.w[1][29]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][2]$_DFF_P_.CLK__assert (\__mp_u0.w[1][2]$_DFF_P_.CLK__gold , \__mp_u0.w[1][2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][30]$_DFF_P_.CLK__assert (\__mp_u0.w[1][30]$_DFF_P_.CLK__gold , \__mp_u0.w[1][30]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][31]$_DFF_P_.CLK__assert (\__mp_u0.w[1][31]$_DFF_P_.CLK__gold , \__mp_u0.w[1][31]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][3]$_DFF_P_.CLK__assert (\__mp_u0.w[1][3]$_DFF_P_.CLK__gold , \__mp_u0.w[1][3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][4]$_DFF_P_.CLK__assert (\__mp_u0.w[1][4]$_DFF_P_.CLK__gold , \__mp_u0.w[1][4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][5]$_DFF_P_.CLK__assert (\__mp_u0.w[1][5]$_DFF_P_.CLK__gold , \__mp_u0.w[1][5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][6]$_DFF_P_.CLK__assert (\__mp_u0.w[1][6]$_DFF_P_.CLK__gold , \__mp_u0.w[1][6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][7]$_DFF_P_.CLK__assert (\__mp_u0.w[1][7]$_DFF_P_.CLK__gold , \__mp_u0.w[1][7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][8]$_DFF_P_.CLK__assert (\__mp_u0.w[1][8]$_DFF_P_.CLK__gold , \__mp_u0.w[1][8]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[1][9]$_DFF_P_.CLK__assert (\__mp_u0.w[1][9]$_DFF_P_.CLK__gold , \__mp_u0.w[1][9]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][0]$_DFF_P_.CLK__assert (\__mp_u0.w[2][0]$_DFF_P_.CLK__gold , \__mp_u0.w[2][0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][10]$_DFF_P_.CLK__assert (\__mp_u0.w[2][10]$_DFF_P_.CLK__gold , \__mp_u0.w[2][10]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][11]$_DFF_P_.CLK__assert (\__mp_u0.w[2][11]$_DFF_P_.CLK__gold , \__mp_u0.w[2][11]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][12]$_DFF_P_.CLK__assert (\__mp_u0.w[2][12]$_DFF_P_.CLK__gold , \__mp_u0.w[2][12]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][13]$_DFF_P_.CLK__assert (\__mp_u0.w[2][13]$_DFF_P_.CLK__gold , \__mp_u0.w[2][13]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][14]$_DFF_P_.CLK__assert (\__mp_u0.w[2][14]$_DFF_P_.CLK__gold , \__mp_u0.w[2][14]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][15]$_DFF_P_.CLK__assert (\__mp_u0.w[2][15]$_DFF_P_.CLK__gold , \__mp_u0.w[2][15]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][16]$_DFF_P_.CLK__assert (\__mp_u0.w[2][16]$_DFF_P_.CLK__gold , \__mp_u0.w[2][16]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][17]$_DFF_P_.CLK__assert (\__mp_u0.w[2][17]$_DFF_P_.CLK__gold , \__mp_u0.w[2][17]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][18]$_DFF_P_.CLK__assert (\__mp_u0.w[2][18]$_DFF_P_.CLK__gold , \__mp_u0.w[2][18]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][19]$_DFF_P_.CLK__assert (\__mp_u0.w[2][19]$_DFF_P_.CLK__gold , \__mp_u0.w[2][19]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][1]$_DFF_P_.CLK__assert (\__mp_u0.w[2][1]$_DFF_P_.CLK__gold , \__mp_u0.w[2][1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][20]$_DFF_P_.CLK__assert (\__mp_u0.w[2][20]$_DFF_P_.CLK__gold , \__mp_u0.w[2][20]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][21]$_DFF_P_.CLK__assert (\__mp_u0.w[2][21]$_DFF_P_.CLK__gold , \__mp_u0.w[2][21]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][22]$_DFF_P_.CLK__assert (\__mp_u0.w[2][22]$_DFF_P_.CLK__gold , \__mp_u0.w[2][22]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][23]$_DFF_P_.CLK__assert (\__mp_u0.w[2][23]$_DFF_P_.CLK__gold , \__mp_u0.w[2][23]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][24]$_DFF_P_.CLK__assert (\__mp_u0.w[2][24]$_DFF_P_.CLK__gold , \__mp_u0.w[2][24]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][25]$_DFF_P_.CLK__assert (\__mp_u0.w[2][25]$_DFF_P_.CLK__gold , \__mp_u0.w[2][25]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][26]$_DFF_P_.CLK__assert (\__mp_u0.w[2][26]$_DFF_P_.CLK__gold , \__mp_u0.w[2][26]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][27]$_DFF_P_.CLK__assert (\__mp_u0.w[2][27]$_DFF_P_.CLK__gold , \__mp_u0.w[2][27]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][28]$_DFF_P_.CLK__assert (\__mp_u0.w[2][28]$_DFF_P_.CLK__gold , \__mp_u0.w[2][28]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][29]$_DFF_P_.CLK__assert (\__mp_u0.w[2][29]$_DFF_P_.CLK__gold , \__mp_u0.w[2][29]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][2]$_DFF_P_.CLK__assert (\__mp_u0.w[2][2]$_DFF_P_.CLK__gold , \__mp_u0.w[2][2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][30]$_DFF_P_.CLK__assert (\__mp_u0.w[2][30]$_DFF_P_.CLK__gold , \__mp_u0.w[2][30]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][31]$_DFF_P_.CLK__assert (\__mp_u0.w[2][31]$_DFF_P_.CLK__gold , \__mp_u0.w[2][31]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][3]$_DFF_P_.CLK__assert (\__mp_u0.w[2][3]$_DFF_P_.CLK__gold , \__mp_u0.w[2][3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][4]$_DFF_P_.CLK__assert (\__mp_u0.w[2][4]$_DFF_P_.CLK__gold , \__mp_u0.w[2][4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][5]$_DFF_P_.CLK__assert (\__mp_u0.w[2][5]$_DFF_P_.CLK__gold , \__mp_u0.w[2][5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][6]$_DFF_P_.CLK__assert (\__mp_u0.w[2][6]$_DFF_P_.CLK__gold , \__mp_u0.w[2][6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][7]$_DFF_P_.CLK__assert (\__mp_u0.w[2][7]$_DFF_P_.CLK__gold , \__mp_u0.w[2][7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][8]$_DFF_P_.CLK__assert (\__mp_u0.w[2][8]$_DFF_P_.CLK__gold , \__mp_u0.w[2][8]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[2][9]$_DFF_P_.CLK__assert (\__mp_u0.w[2][9]$_DFF_P_.CLK__gold , \__mp_u0.w[2][9]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][0]$_DFF_P_.CLK__assert (\__mp_u0.w[3][0]$_DFF_P_.CLK__gold , \__mp_u0.w[3][0]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][10]$_DFF_P_.CLK__assert (\__mp_u0.w[3][10]$_DFF_P_.CLK__gold , \__mp_u0.w[3][10]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][11]$_DFF_P_.CLK__assert (\__mp_u0.w[3][11]$_DFF_P_.CLK__gold , \__mp_u0.w[3][11]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][12]$_DFF_P_.CLK__assert (\__mp_u0.w[3][12]$_DFF_P_.CLK__gold , \__mp_u0.w[3][12]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][13]$_DFF_P_.CLK__assert (\__mp_u0.w[3][13]$_DFF_P_.CLK__gold , \__mp_u0.w[3][13]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][14]$_DFF_P_.CLK__assert (\__mp_u0.w[3][14]$_DFF_P_.CLK__gold , \__mp_u0.w[3][14]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][15]$_DFF_P_.CLK__assert (\__mp_u0.w[3][15]$_DFF_P_.CLK__gold , \__mp_u0.w[3][15]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][16]$_DFF_P_.CLK__assert (\__mp_u0.w[3][16]$_DFF_P_.CLK__gold , \__mp_u0.w[3][16]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][17]$_DFF_P_.CLK__assert (\__mp_u0.w[3][17]$_DFF_P_.CLK__gold , \__mp_u0.w[3][17]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][18]$_DFF_P_.CLK__assert (\__mp_u0.w[3][18]$_DFF_P_.CLK__gold , \__mp_u0.w[3][18]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][19]$_DFF_P_.CLK__assert (\__mp_u0.w[3][19]$_DFF_P_.CLK__gold , \__mp_u0.w[3][19]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][1]$_DFF_P_.CLK__assert (\__mp_u0.w[3][1]$_DFF_P_.CLK__gold , \__mp_u0.w[3][1]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][20]$_DFF_P_.CLK__assert (\__mp_u0.w[3][20]$_DFF_P_.CLK__gold , \__mp_u0.w[3][20]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][21]$_DFF_P_.CLK__assert (\__mp_u0.w[3][21]$_DFF_P_.CLK__gold , \__mp_u0.w[3][21]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][22]$_DFF_P_.CLK__assert (\__mp_u0.w[3][22]$_DFF_P_.CLK__gold , \__mp_u0.w[3][22]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][23]$_DFF_P_.CLK__assert (\__mp_u0.w[3][23]$_DFF_P_.CLK__gold , \__mp_u0.w[3][23]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][24]$_DFF_P_.CLK__assert (\__mp_u0.w[3][24]$_DFF_P_.CLK__gold , \__mp_u0.w[3][24]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][25]$_DFF_P_.CLK__assert (\__mp_u0.w[3][25]$_DFF_P_.CLK__gold , \__mp_u0.w[3][25]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][26]$_DFF_P_.CLK__assert (\__mp_u0.w[3][26]$_DFF_P_.CLK__gold , \__mp_u0.w[3][26]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][27]$_DFF_P_.CLK__assert (\__mp_u0.w[3][27]$_DFF_P_.CLK__gold , \__mp_u0.w[3][27]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][28]$_DFF_P_.CLK__assert (\__mp_u0.w[3][28]$_DFF_P_.CLK__gold , \__mp_u0.w[3][28]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][29]$_DFF_P_.CLK__assert (\__mp_u0.w[3][29]$_DFF_P_.CLK__gold , \__mp_u0.w[3][29]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][2]$_DFF_P_.CLK__assert (\__mp_u0.w[3][2]$_DFF_P_.CLK__gold , \__mp_u0.w[3][2]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][30]$_DFF_P_.CLK__assert (\__mp_u0.w[3][30]$_DFF_P_.CLK__gold , \__mp_u0.w[3][30]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][31]$_DFF_P_.CLK__assert (\__mp_u0.w[3][31]$_DFF_P_.CLK__gold , \__mp_u0.w[3][31]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][3]$_DFF_P_.CLK__assert (\__mp_u0.w[3][3]$_DFF_P_.CLK__gold , \__mp_u0.w[3][3]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][4]$_DFF_P_.CLK__assert (\__mp_u0.w[3][4]$_DFF_P_.CLK__gold , \__mp_u0.w[3][4]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][5]$_DFF_P_.CLK__assert (\__mp_u0.w[3][5]$_DFF_P_.CLK__gold , \__mp_u0.w[3][5]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][6]$_DFF_P_.CLK__assert (\__mp_u0.w[3][6]$_DFF_P_.CLK__gold , \__mp_u0.w[3][6]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][7]$_DFF_P_.CLK__assert (\__mp_u0.w[3][7]$_DFF_P_.CLK__gold , \__mp_u0.w[3][7]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][8]$_DFF_P_.CLK__assert (\__mp_u0.w[3][8]$_DFF_P_.CLK__gold , \__mp_u0.w[3][8]$_DFF_P_.CLK__gate );
  miter_cmp_prop #(1, "assert") \__mp_u0.w[3][9]$_DFF_P_.CLK__assert (\__mp_u0.w[3][9]$_DFF_P_.CLK__gold , \__mp_u0.w[3][9]$_DFF_P_.CLK__gate );
`endif
`ifdef CHECK_OUTPUTS
  miter_cmp_prop #(1, "assert") \__po_done__assert (\__po_done__gold , \__po_done__gate );
  miter_cmp_prop #(128, "assert") \__po_text_out__assert (\__po_text_out__gold , \__po_text_out__gate );
`endif
`ifdef COVER_DEF_CROSS_POINTS
  `ifdef DIRECT_CROSS_POINTS
  `else
  `endif
`endif
`ifdef COVER_DEF_GOLD_MATCH_POINTS
  miter_def_prop #(1, "cover") \__mp_clkbuf_0_clk.A__gold_cover (\__mp_clkbuf_0_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_0_clk.Y__gold_cover (\__mp_clkbuf_0_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_0_0_clk.A__gold_cover (\__mp_clkbuf_2_0_0_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_0_0_clk.Y__gold_cover (\__mp_clkbuf_2_0_0_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_1_0_clk.A__gold_cover (\__mp_clkbuf_2_1_0_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_1_0_clk.Y__gold_cover (\__mp_clkbuf_2_1_0_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_2_0_clk.A__gold_cover (\__mp_clkbuf_2_2_0_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_2_0_clk.Y__gold_cover (\__mp_clkbuf_2_2_0_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_3_0_clk.A__gold_cover (\__mp_clkbuf_2_3_0_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_3_0_clk.Y__gold_cover (\__mp_clkbuf_2_3_0_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_0_clk.A__gold_cover (\__mp_clkbuf_leaf_0_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_0_clk.Y__gold_cover (\__mp_clkbuf_leaf_0_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_10_clk.A__gold_cover (\__mp_clkbuf_leaf_10_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_10_clk.Y__gold_cover (\__mp_clkbuf_leaf_10_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_11_clk.A__gold_cover (\__mp_clkbuf_leaf_11_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_11_clk.Y__gold_cover (\__mp_clkbuf_leaf_11_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_12_clk.A__gold_cover (\__mp_clkbuf_leaf_12_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_12_clk.Y__gold_cover (\__mp_clkbuf_leaf_12_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_13_clk.A__gold_cover (\__mp_clkbuf_leaf_13_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_13_clk.Y__gold_cover (\__mp_clkbuf_leaf_13_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_14_clk.A__gold_cover (\__mp_clkbuf_leaf_14_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_14_clk.Y__gold_cover (\__mp_clkbuf_leaf_14_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_15_clk.A__gold_cover (\__mp_clkbuf_leaf_15_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_15_clk.Y__gold_cover (\__mp_clkbuf_leaf_15_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_16_clk.A__gold_cover (\__mp_clkbuf_leaf_16_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_16_clk.Y__gold_cover (\__mp_clkbuf_leaf_16_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_17_clk.A__gold_cover (\__mp_clkbuf_leaf_17_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_17_clk.Y__gold_cover (\__mp_clkbuf_leaf_17_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_18_clk.A__gold_cover (\__mp_clkbuf_leaf_18_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_18_clk.Y__gold_cover (\__mp_clkbuf_leaf_18_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_19_clk.A__gold_cover (\__mp_clkbuf_leaf_19_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_19_clk.Y__gold_cover (\__mp_clkbuf_leaf_19_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_1_clk.A__gold_cover (\__mp_clkbuf_leaf_1_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_1_clk.Y__gold_cover (\__mp_clkbuf_leaf_1_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_20_clk.A__gold_cover (\__mp_clkbuf_leaf_20_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_20_clk.Y__gold_cover (\__mp_clkbuf_leaf_20_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_21_clk.A__gold_cover (\__mp_clkbuf_leaf_21_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_21_clk.Y__gold_cover (\__mp_clkbuf_leaf_21_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_22_clk.A__gold_cover (\__mp_clkbuf_leaf_22_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_22_clk.Y__gold_cover (\__mp_clkbuf_leaf_22_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_23_clk.A__gold_cover (\__mp_clkbuf_leaf_23_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_23_clk.Y__gold_cover (\__mp_clkbuf_leaf_23_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_24_clk.A__gold_cover (\__mp_clkbuf_leaf_24_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_24_clk.Y__gold_cover (\__mp_clkbuf_leaf_24_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_25_clk.A__gold_cover (\__mp_clkbuf_leaf_25_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_25_clk.Y__gold_cover (\__mp_clkbuf_leaf_25_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_26_clk.A__gold_cover (\__mp_clkbuf_leaf_26_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_26_clk.Y__gold_cover (\__mp_clkbuf_leaf_26_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_27_clk.A__gold_cover (\__mp_clkbuf_leaf_27_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_27_clk.Y__gold_cover (\__mp_clkbuf_leaf_27_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_28_clk.A__gold_cover (\__mp_clkbuf_leaf_28_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_28_clk.Y__gold_cover (\__mp_clkbuf_leaf_28_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_29_clk.A__gold_cover (\__mp_clkbuf_leaf_29_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_29_clk.Y__gold_cover (\__mp_clkbuf_leaf_29_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_2_clk.A__gold_cover (\__mp_clkbuf_leaf_2_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_2_clk.Y__gold_cover (\__mp_clkbuf_leaf_2_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_30_clk.A__gold_cover (\__mp_clkbuf_leaf_30_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_30_clk.Y__gold_cover (\__mp_clkbuf_leaf_30_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_31_clk.A__gold_cover (\__mp_clkbuf_leaf_31_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_31_clk.Y__gold_cover (\__mp_clkbuf_leaf_31_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_32_clk.A__gold_cover (\__mp_clkbuf_leaf_32_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_32_clk.Y__gold_cover (\__mp_clkbuf_leaf_32_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_33_clk.A__gold_cover (\__mp_clkbuf_leaf_33_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_33_clk.Y__gold_cover (\__mp_clkbuf_leaf_33_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_3_clk.A__gold_cover (\__mp_clkbuf_leaf_3_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_3_clk.Y__gold_cover (\__mp_clkbuf_leaf_3_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_4_clk.A__gold_cover (\__mp_clkbuf_leaf_4_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_4_clk.Y__gold_cover (\__mp_clkbuf_leaf_4_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_5_clk.A__gold_cover (\__mp_clkbuf_leaf_5_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_5_clk.Y__gold_cover (\__mp_clkbuf_leaf_5_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_6_clk.A__gold_cover (\__mp_clkbuf_leaf_6_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_6_clk.Y__gold_cover (\__mp_clkbuf_leaf_6_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_7_clk.A__gold_cover (\__mp_clkbuf_leaf_7_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_7_clk.Y__gold_cover (\__mp_clkbuf_leaf_7_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_8_clk.A__gold_cover (\__mp_clkbuf_leaf_8_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_8_clk.Y__gold_cover (\__mp_clkbuf_leaf_8_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_9_clk.A__gold_cover (\__mp_clkbuf_leaf_9_clk.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_9_clk.Y__gold_cover (\__mp_clkbuf_leaf_9_clk.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkload0.A__gold_cover (\__mp_clkload0.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload0.Y__gold_cover (\__mp_clkload0.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkload1.A__gold_cover (\__mp_clkload1.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload10.A__gold_cover (\__mp_clkload10.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload11.A__gold_cover (\__mp_clkload11.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload12.A__gold_cover (\__mp_clkload12.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload13.A__gold_cover (\__mp_clkload13.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload14.A__gold_cover (\__mp_clkload14.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload15.A__gold_cover (\__mp_clkload15.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload16.A__gold_cover (\__mp_clkload16.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload17.A__gold_cover (\__mp_clkload17.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload18.A__gold_cover (\__mp_clkload18.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload18.Y__gold_cover (\__mp_clkload18.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkload19.A__gold_cover (\__mp_clkload19.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload2.A__gold_cover (\__mp_clkload2.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload20.A__gold_cover (\__mp_clkload20.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload21.A__gold_cover (\__mp_clkload21.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload22.A__gold_cover (\__mp_clkload22.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload23.A__gold_cover (\__mp_clkload23.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload24.A__gold_cover (\__mp_clkload24.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload25.A__gold_cover (\__mp_clkload25.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload26.A__gold_cover (\__mp_clkload26.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload27.A__gold_cover (\__mp_clkload27.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload28.A__gold_cover (\__mp_clkload28.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload29.A__gold_cover (\__mp_clkload29.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload3.A__gold_cover (\__mp_clkload3.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload30.A__gold_cover (\__mp_clkload30.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload31.A__gold_cover (\__mp_clkload31.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload31.Y__gold_cover (\__mp_clkload31.Y__gold );
  miter_def_prop #(1, "cover") \__mp_clkload32.A__gold_cover (\__mp_clkload32.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload4.A__gold_cover (\__mp_clkload4.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload5.A__gold_cover (\__mp_clkload5.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload6.A__gold_cover (\__mp_clkload6.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload7.A__gold_cover (\__mp_clkload7.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload8.A__gold_cover (\__mp_clkload8.A__gold );
  miter_def_prop #(1, "cover") \__mp_clkload9.A__gold_cover (\__mp_clkload9.A__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_0_clk__gold_cover (\__mp_clknet_0_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_2_0_0_clk__gold_cover (\__mp_clknet_2_0_0_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_2_1_0_clk__gold_cover (\__mp_clknet_2_1_0_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_2_2_0_clk__gold_cover (\__mp_clknet_2_2_0_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_2_3_0_clk__gold_cover (\__mp_clknet_2_3_0_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_0_clk__gold_cover (\__mp_clknet_leaf_0_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_10_clk__gold_cover (\__mp_clknet_leaf_10_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_11_clk__gold_cover (\__mp_clknet_leaf_11_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_12_clk__gold_cover (\__mp_clknet_leaf_12_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_13_clk__gold_cover (\__mp_clknet_leaf_13_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_14_clk__gold_cover (\__mp_clknet_leaf_14_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_15_clk__gold_cover (\__mp_clknet_leaf_15_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_16_clk__gold_cover (\__mp_clknet_leaf_16_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_17_clk__gold_cover (\__mp_clknet_leaf_17_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_18_clk__gold_cover (\__mp_clknet_leaf_18_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_19_clk__gold_cover (\__mp_clknet_leaf_19_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_1_clk__gold_cover (\__mp_clknet_leaf_1_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_20_clk__gold_cover (\__mp_clknet_leaf_20_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_21_clk__gold_cover (\__mp_clknet_leaf_21_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_22_clk__gold_cover (\__mp_clknet_leaf_22_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_23_clk__gold_cover (\__mp_clknet_leaf_23_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_24_clk__gold_cover (\__mp_clknet_leaf_24_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_25_clk__gold_cover (\__mp_clknet_leaf_25_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_26_clk__gold_cover (\__mp_clknet_leaf_26_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_27_clk__gold_cover (\__mp_clknet_leaf_27_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_28_clk__gold_cover (\__mp_clknet_leaf_28_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_29_clk__gold_cover (\__mp_clknet_leaf_29_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_2_clk__gold_cover (\__mp_clknet_leaf_2_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_30_clk__gold_cover (\__mp_clknet_leaf_30_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_31_clk__gold_cover (\__mp_clknet_leaf_31_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_32_clk__gold_cover (\__mp_clknet_leaf_32_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_33_clk__gold_cover (\__mp_clknet_leaf_33_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_3_clk__gold_cover (\__mp_clknet_leaf_3_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_4_clk__gold_cover (\__mp_clknet_leaf_4_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_5_clk__gold_cover (\__mp_clknet_leaf_5_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_6_clk__gold_cover (\__mp_clknet_leaf_6_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_7_clk__gold_cover (\__mp_clknet_leaf_7_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_8_clk__gold_cover (\__mp_clknet_leaf_8_clk__gold );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_9_clk__gold_cover (\__mp_clknet_leaf_9_clk__gold );
  miter_def_prop #(1, "cover") \__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gold_cover (\__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gold_cover (\__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gold_cover (\__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gold_cover (\__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_done$_DFF_P_.CLK__gold_cover (\__mp_done$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_done$_DFF_P_.QN__gold_cover (\__mp_done$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_done$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_done$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_input1.A__gold_cover (\__mp_input1.A__gold );
  miter_def_prop #(1, "cover") \__mp_input1.Y__gold_cover (\__mp_input1.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input10.A__gold_cover (\__mp_input10.A__gold );
  miter_def_prop #(1, "cover") \__mp_input10.Y__gold_cover (\__mp_input10.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input100.A__gold_cover (\__mp_input100.A__gold );
  miter_def_prop #(1, "cover") \__mp_input100.Y__gold_cover (\__mp_input100.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input101.A__gold_cover (\__mp_input101.A__gold );
  miter_def_prop #(1, "cover") \__mp_input101.Y__gold_cover (\__mp_input101.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input102.A__gold_cover (\__mp_input102.A__gold );
  miter_def_prop #(1, "cover") \__mp_input102.Y__gold_cover (\__mp_input102.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input103.A__gold_cover (\__mp_input103.A__gold );
  miter_def_prop #(1, "cover") \__mp_input103.Y__gold_cover (\__mp_input103.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input104.A__gold_cover (\__mp_input104.A__gold );
  miter_def_prop #(1, "cover") \__mp_input104.Y__gold_cover (\__mp_input104.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input105.A__gold_cover (\__mp_input105.A__gold );
  miter_def_prop #(1, "cover") \__mp_input105.Y__gold_cover (\__mp_input105.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input106.A__gold_cover (\__mp_input106.A__gold );
  miter_def_prop #(1, "cover") \__mp_input106.Y__gold_cover (\__mp_input106.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input107.A__gold_cover (\__mp_input107.A__gold );
  miter_def_prop #(1, "cover") \__mp_input107.Y__gold_cover (\__mp_input107.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input108.A__gold_cover (\__mp_input108.A__gold );
  miter_def_prop #(1, "cover") \__mp_input108.Y__gold_cover (\__mp_input108.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input109.A__gold_cover (\__mp_input109.A__gold );
  miter_def_prop #(1, "cover") \__mp_input109.Y__gold_cover (\__mp_input109.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input11.A__gold_cover (\__mp_input11.A__gold );
  miter_def_prop #(1, "cover") \__mp_input11.Y__gold_cover (\__mp_input11.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input110.A__gold_cover (\__mp_input110.A__gold );
  miter_def_prop #(1, "cover") \__mp_input110.Y__gold_cover (\__mp_input110.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input111.A__gold_cover (\__mp_input111.A__gold );
  miter_def_prop #(1, "cover") \__mp_input111.Y__gold_cover (\__mp_input111.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input112.A__gold_cover (\__mp_input112.A__gold );
  miter_def_prop #(1, "cover") \__mp_input112.Y__gold_cover (\__mp_input112.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input113.A__gold_cover (\__mp_input113.A__gold );
  miter_def_prop #(1, "cover") \__mp_input113.Y__gold_cover (\__mp_input113.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input114.A__gold_cover (\__mp_input114.A__gold );
  miter_def_prop #(1, "cover") \__mp_input114.Y__gold_cover (\__mp_input114.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input115.A__gold_cover (\__mp_input115.A__gold );
  miter_def_prop #(1, "cover") \__mp_input115.Y__gold_cover (\__mp_input115.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input116.A__gold_cover (\__mp_input116.A__gold );
  miter_def_prop #(1, "cover") \__mp_input116.Y__gold_cover (\__mp_input116.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input117.A__gold_cover (\__mp_input117.A__gold );
  miter_def_prop #(1, "cover") \__mp_input117.Y__gold_cover (\__mp_input117.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input118.A__gold_cover (\__mp_input118.A__gold );
  miter_def_prop #(1, "cover") \__mp_input118.Y__gold_cover (\__mp_input118.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input119.A__gold_cover (\__mp_input119.A__gold );
  miter_def_prop #(1, "cover") \__mp_input119.Y__gold_cover (\__mp_input119.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input12.A__gold_cover (\__mp_input12.A__gold );
  miter_def_prop #(1, "cover") \__mp_input12.Y__gold_cover (\__mp_input12.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input120.A__gold_cover (\__mp_input120.A__gold );
  miter_def_prop #(1, "cover") \__mp_input120.Y__gold_cover (\__mp_input120.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input121.A__gold_cover (\__mp_input121.A__gold );
  miter_def_prop #(1, "cover") \__mp_input121.Y__gold_cover (\__mp_input121.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input122.A__gold_cover (\__mp_input122.A__gold );
  miter_def_prop #(1, "cover") \__mp_input122.Y__gold_cover (\__mp_input122.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input123.A__gold_cover (\__mp_input123.A__gold );
  miter_def_prop #(1, "cover") \__mp_input123.Y__gold_cover (\__mp_input123.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input124.A__gold_cover (\__mp_input124.A__gold );
  miter_def_prop #(1, "cover") \__mp_input124.Y__gold_cover (\__mp_input124.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input125.A__gold_cover (\__mp_input125.A__gold );
  miter_def_prop #(1, "cover") \__mp_input125.Y__gold_cover (\__mp_input125.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input126.A__gold_cover (\__mp_input126.A__gold );
  miter_def_prop #(1, "cover") \__mp_input126.Y__gold_cover (\__mp_input126.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input127.A__gold_cover (\__mp_input127.A__gold );
  miter_def_prop #(1, "cover") \__mp_input127.Y__gold_cover (\__mp_input127.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input128.A__gold_cover (\__mp_input128.A__gold );
  miter_def_prop #(1, "cover") \__mp_input128.Y__gold_cover (\__mp_input128.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input129.A__gold_cover (\__mp_input129.A__gold );
  miter_def_prop #(1, "cover") \__mp_input129.Y__gold_cover (\__mp_input129.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input13.A__gold_cover (\__mp_input13.A__gold );
  miter_def_prop #(1, "cover") \__mp_input13.Y__gold_cover (\__mp_input13.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input130.A__gold_cover (\__mp_input130.A__gold );
  miter_def_prop #(1, "cover") \__mp_input130.Y__gold_cover (\__mp_input130.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input131.A__gold_cover (\__mp_input131.A__gold );
  miter_def_prop #(1, "cover") \__mp_input131.Y__gold_cover (\__mp_input131.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input132.A__gold_cover (\__mp_input132.A__gold );
  miter_def_prop #(1, "cover") \__mp_input132.Y__gold_cover (\__mp_input132.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input133.A__gold_cover (\__mp_input133.A__gold );
  miter_def_prop #(1, "cover") \__mp_input133.Y__gold_cover (\__mp_input133.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input134.A__gold_cover (\__mp_input134.A__gold );
  miter_def_prop #(1, "cover") \__mp_input134.Y__gold_cover (\__mp_input134.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input135.A__gold_cover (\__mp_input135.A__gold );
  miter_def_prop #(1, "cover") \__mp_input135.Y__gold_cover (\__mp_input135.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input136.A__gold_cover (\__mp_input136.A__gold );
  miter_def_prop #(1, "cover") \__mp_input136.Y__gold_cover (\__mp_input136.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input137.A__gold_cover (\__mp_input137.A__gold );
  miter_def_prop #(1, "cover") \__mp_input137.Y__gold_cover (\__mp_input137.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input138.A__gold_cover (\__mp_input138.A__gold );
  miter_def_prop #(1, "cover") \__mp_input138.Y__gold_cover (\__mp_input138.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input139.A__gold_cover (\__mp_input139.A__gold );
  miter_def_prop #(1, "cover") \__mp_input139.Y__gold_cover (\__mp_input139.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input14.A__gold_cover (\__mp_input14.A__gold );
  miter_def_prop #(1, "cover") \__mp_input14.Y__gold_cover (\__mp_input14.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input140.A__gold_cover (\__mp_input140.A__gold );
  miter_def_prop #(1, "cover") \__mp_input140.Y__gold_cover (\__mp_input140.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input141.A__gold_cover (\__mp_input141.A__gold );
  miter_def_prop #(1, "cover") \__mp_input141.Y__gold_cover (\__mp_input141.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input142.A__gold_cover (\__mp_input142.A__gold );
  miter_def_prop #(1, "cover") \__mp_input142.Y__gold_cover (\__mp_input142.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input143.A__gold_cover (\__mp_input143.A__gold );
  miter_def_prop #(1, "cover") \__mp_input143.Y__gold_cover (\__mp_input143.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input144.A__gold_cover (\__mp_input144.A__gold );
  miter_def_prop #(1, "cover") \__mp_input144.Y__gold_cover (\__mp_input144.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input145.A__gold_cover (\__mp_input145.A__gold );
  miter_def_prop #(1, "cover") \__mp_input145.Y__gold_cover (\__mp_input145.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input146.A__gold_cover (\__mp_input146.A__gold );
  miter_def_prop #(1, "cover") \__mp_input146.Y__gold_cover (\__mp_input146.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input147.A__gold_cover (\__mp_input147.A__gold );
  miter_def_prop #(1, "cover") \__mp_input147.Y__gold_cover (\__mp_input147.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input148.A__gold_cover (\__mp_input148.A__gold );
  miter_def_prop #(1, "cover") \__mp_input148.Y__gold_cover (\__mp_input148.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input149.A__gold_cover (\__mp_input149.A__gold );
  miter_def_prop #(1, "cover") \__mp_input149.Y__gold_cover (\__mp_input149.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input15.A__gold_cover (\__mp_input15.A__gold );
  miter_def_prop #(1, "cover") \__mp_input15.Y__gold_cover (\__mp_input15.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input150.A__gold_cover (\__mp_input150.A__gold );
  miter_def_prop #(1, "cover") \__mp_input150.Y__gold_cover (\__mp_input150.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input151.A__gold_cover (\__mp_input151.A__gold );
  miter_def_prop #(1, "cover") \__mp_input151.Y__gold_cover (\__mp_input151.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input152.A__gold_cover (\__mp_input152.A__gold );
  miter_def_prop #(1, "cover") \__mp_input152.Y__gold_cover (\__mp_input152.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input153.A__gold_cover (\__mp_input153.A__gold );
  miter_def_prop #(1, "cover") \__mp_input153.Y__gold_cover (\__mp_input153.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input154.A__gold_cover (\__mp_input154.A__gold );
  miter_def_prop #(1, "cover") \__mp_input154.Y__gold_cover (\__mp_input154.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input155.A__gold_cover (\__mp_input155.A__gold );
  miter_def_prop #(1, "cover") \__mp_input155.Y__gold_cover (\__mp_input155.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input156.A__gold_cover (\__mp_input156.A__gold );
  miter_def_prop #(1, "cover") \__mp_input156.Y__gold_cover (\__mp_input156.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input157.A__gold_cover (\__mp_input157.A__gold );
  miter_def_prop #(1, "cover") \__mp_input157.Y__gold_cover (\__mp_input157.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input158.A__gold_cover (\__mp_input158.A__gold );
  miter_def_prop #(1, "cover") \__mp_input158.Y__gold_cover (\__mp_input158.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input159.A__gold_cover (\__mp_input159.A__gold );
  miter_def_prop #(1, "cover") \__mp_input159.Y__gold_cover (\__mp_input159.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input16.A__gold_cover (\__mp_input16.A__gold );
  miter_def_prop #(1, "cover") \__mp_input16.Y__gold_cover (\__mp_input16.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input160.A__gold_cover (\__mp_input160.A__gold );
  miter_def_prop #(1, "cover") \__mp_input160.Y__gold_cover (\__mp_input160.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input161.A__gold_cover (\__mp_input161.A__gold );
  miter_def_prop #(1, "cover") \__mp_input161.Y__gold_cover (\__mp_input161.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input162.A__gold_cover (\__mp_input162.A__gold );
  miter_def_prop #(1, "cover") \__mp_input162.Y__gold_cover (\__mp_input162.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input163.A__gold_cover (\__mp_input163.A__gold );
  miter_def_prop #(1, "cover") \__mp_input163.Y__gold_cover (\__mp_input163.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input164.A__gold_cover (\__mp_input164.A__gold );
  miter_def_prop #(1, "cover") \__mp_input164.Y__gold_cover (\__mp_input164.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input165.A__gold_cover (\__mp_input165.A__gold );
  miter_def_prop #(1, "cover") \__mp_input165.Y__gold_cover (\__mp_input165.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input166.A__gold_cover (\__mp_input166.A__gold );
  miter_def_prop #(1, "cover") \__mp_input166.Y__gold_cover (\__mp_input166.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input167.A__gold_cover (\__mp_input167.A__gold );
  miter_def_prop #(1, "cover") \__mp_input167.Y__gold_cover (\__mp_input167.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input168.A__gold_cover (\__mp_input168.A__gold );
  miter_def_prop #(1, "cover") \__mp_input168.Y__gold_cover (\__mp_input168.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input169.A__gold_cover (\__mp_input169.A__gold );
  miter_def_prop #(1, "cover") \__mp_input169.Y__gold_cover (\__mp_input169.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input17.A__gold_cover (\__mp_input17.A__gold );
  miter_def_prop #(1, "cover") \__mp_input17.Y__gold_cover (\__mp_input17.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input170.A__gold_cover (\__mp_input170.A__gold );
  miter_def_prop #(1, "cover") \__mp_input170.Y__gold_cover (\__mp_input170.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input171.A__gold_cover (\__mp_input171.A__gold );
  miter_def_prop #(1, "cover") \__mp_input171.Y__gold_cover (\__mp_input171.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input172.A__gold_cover (\__mp_input172.A__gold );
  miter_def_prop #(1, "cover") \__mp_input172.Y__gold_cover (\__mp_input172.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input173.A__gold_cover (\__mp_input173.A__gold );
  miter_def_prop #(1, "cover") \__mp_input173.Y__gold_cover (\__mp_input173.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input174.A__gold_cover (\__mp_input174.A__gold );
  miter_def_prop #(1, "cover") \__mp_input174.Y__gold_cover (\__mp_input174.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input175.A__gold_cover (\__mp_input175.A__gold );
  miter_def_prop #(1, "cover") \__mp_input175.Y__gold_cover (\__mp_input175.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input176.A__gold_cover (\__mp_input176.A__gold );
  miter_def_prop #(1, "cover") \__mp_input176.Y__gold_cover (\__mp_input176.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input177.A__gold_cover (\__mp_input177.A__gold );
  miter_def_prop #(1, "cover") \__mp_input177.Y__gold_cover (\__mp_input177.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input178.A__gold_cover (\__mp_input178.A__gold );
  miter_def_prop #(1, "cover") \__mp_input178.Y__gold_cover (\__mp_input178.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input179.A__gold_cover (\__mp_input179.A__gold );
  miter_def_prop #(1, "cover") \__mp_input179.Y__gold_cover (\__mp_input179.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input18.A__gold_cover (\__mp_input18.A__gold );
  miter_def_prop #(1, "cover") \__mp_input18.Y__gold_cover (\__mp_input18.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input180.A__gold_cover (\__mp_input180.A__gold );
  miter_def_prop #(1, "cover") \__mp_input180.Y__gold_cover (\__mp_input180.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input181.A__gold_cover (\__mp_input181.A__gold );
  miter_def_prop #(1, "cover") \__mp_input181.Y__gold_cover (\__mp_input181.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input182.A__gold_cover (\__mp_input182.A__gold );
  miter_def_prop #(1, "cover") \__mp_input182.Y__gold_cover (\__mp_input182.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input183.A__gold_cover (\__mp_input183.A__gold );
  miter_def_prop #(1, "cover") \__mp_input183.Y__gold_cover (\__mp_input183.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input184.A__gold_cover (\__mp_input184.A__gold );
  miter_def_prop #(1, "cover") \__mp_input184.Y__gold_cover (\__mp_input184.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input185.A__gold_cover (\__mp_input185.A__gold );
  miter_def_prop #(1, "cover") \__mp_input185.Y__gold_cover (\__mp_input185.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input186.A__gold_cover (\__mp_input186.A__gold );
  miter_def_prop #(1, "cover") \__mp_input186.Y__gold_cover (\__mp_input186.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input187.A__gold_cover (\__mp_input187.A__gold );
  miter_def_prop #(1, "cover") \__mp_input187.Y__gold_cover (\__mp_input187.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input188.A__gold_cover (\__mp_input188.A__gold );
  miter_def_prop #(1, "cover") \__mp_input188.Y__gold_cover (\__mp_input188.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input189.A__gold_cover (\__mp_input189.A__gold );
  miter_def_prop #(1, "cover") \__mp_input189.Y__gold_cover (\__mp_input189.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input19.A__gold_cover (\__mp_input19.A__gold );
  miter_def_prop #(1, "cover") \__mp_input19.Y__gold_cover (\__mp_input19.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input190.A__gold_cover (\__mp_input190.A__gold );
  miter_def_prop #(1, "cover") \__mp_input190.Y__gold_cover (\__mp_input190.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input191.A__gold_cover (\__mp_input191.A__gold );
  miter_def_prop #(1, "cover") \__mp_input191.Y__gold_cover (\__mp_input191.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input192.A__gold_cover (\__mp_input192.A__gold );
  miter_def_prop #(1, "cover") \__mp_input192.Y__gold_cover (\__mp_input192.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input193.A__gold_cover (\__mp_input193.A__gold );
  miter_def_prop #(1, "cover") \__mp_input193.Y__gold_cover (\__mp_input193.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input194.A__gold_cover (\__mp_input194.A__gold );
  miter_def_prop #(1, "cover") \__mp_input194.Y__gold_cover (\__mp_input194.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input195.A__gold_cover (\__mp_input195.A__gold );
  miter_def_prop #(1, "cover") \__mp_input195.Y__gold_cover (\__mp_input195.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input196.A__gold_cover (\__mp_input196.A__gold );
  miter_def_prop #(1, "cover") \__mp_input196.Y__gold_cover (\__mp_input196.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input197.A__gold_cover (\__mp_input197.A__gold );
  miter_def_prop #(1, "cover") \__mp_input197.Y__gold_cover (\__mp_input197.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input198.A__gold_cover (\__mp_input198.A__gold );
  miter_def_prop #(1, "cover") \__mp_input198.Y__gold_cover (\__mp_input198.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input199.A__gold_cover (\__mp_input199.A__gold );
  miter_def_prop #(1, "cover") \__mp_input199.Y__gold_cover (\__mp_input199.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input2.A__gold_cover (\__mp_input2.A__gold );
  miter_def_prop #(1, "cover") \__mp_input2.Y__gold_cover (\__mp_input2.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input20.A__gold_cover (\__mp_input20.A__gold );
  miter_def_prop #(1, "cover") \__mp_input20.Y__gold_cover (\__mp_input20.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input200.A__gold_cover (\__mp_input200.A__gold );
  miter_def_prop #(1, "cover") \__mp_input200.Y__gold_cover (\__mp_input200.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input201.A__gold_cover (\__mp_input201.A__gold );
  miter_def_prop #(1, "cover") \__mp_input201.Y__gold_cover (\__mp_input201.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input202.A__gold_cover (\__mp_input202.A__gold );
  miter_def_prop #(1, "cover") \__mp_input202.Y__gold_cover (\__mp_input202.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input203.A__gold_cover (\__mp_input203.A__gold );
  miter_def_prop #(1, "cover") \__mp_input203.Y__gold_cover (\__mp_input203.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input204.A__gold_cover (\__mp_input204.A__gold );
  miter_def_prop #(1, "cover") \__mp_input204.Y__gold_cover (\__mp_input204.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input205.A__gold_cover (\__mp_input205.A__gold );
  miter_def_prop #(1, "cover") \__mp_input205.Y__gold_cover (\__mp_input205.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input206.A__gold_cover (\__mp_input206.A__gold );
  miter_def_prop #(1, "cover") \__mp_input206.Y__gold_cover (\__mp_input206.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input207.A__gold_cover (\__mp_input207.A__gold );
  miter_def_prop #(1, "cover") \__mp_input207.Y__gold_cover (\__mp_input207.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input208.A__gold_cover (\__mp_input208.A__gold );
  miter_def_prop #(1, "cover") \__mp_input208.Y__gold_cover (\__mp_input208.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input209.A__gold_cover (\__mp_input209.A__gold );
  miter_def_prop #(1, "cover") \__mp_input209.Y__gold_cover (\__mp_input209.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input21.A__gold_cover (\__mp_input21.A__gold );
  miter_def_prop #(1, "cover") \__mp_input21.Y__gold_cover (\__mp_input21.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input210.A__gold_cover (\__mp_input210.A__gold );
  miter_def_prop #(1, "cover") \__mp_input210.Y__gold_cover (\__mp_input210.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input211.A__gold_cover (\__mp_input211.A__gold );
  miter_def_prop #(1, "cover") \__mp_input211.Y__gold_cover (\__mp_input211.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input212.A__gold_cover (\__mp_input212.A__gold );
  miter_def_prop #(1, "cover") \__mp_input212.Y__gold_cover (\__mp_input212.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input213.A__gold_cover (\__mp_input213.A__gold );
  miter_def_prop #(1, "cover") \__mp_input213.Y__gold_cover (\__mp_input213.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input214.A__gold_cover (\__mp_input214.A__gold );
  miter_def_prop #(1, "cover") \__mp_input214.Y__gold_cover (\__mp_input214.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input215.A__gold_cover (\__mp_input215.A__gold );
  miter_def_prop #(1, "cover") \__mp_input215.Y__gold_cover (\__mp_input215.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input216.A__gold_cover (\__mp_input216.A__gold );
  miter_def_prop #(1, "cover") \__mp_input216.Y__gold_cover (\__mp_input216.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input217.A__gold_cover (\__mp_input217.A__gold );
  miter_def_prop #(1, "cover") \__mp_input217.Y__gold_cover (\__mp_input217.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input218.A__gold_cover (\__mp_input218.A__gold );
  miter_def_prop #(1, "cover") \__mp_input218.Y__gold_cover (\__mp_input218.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input219.A__gold_cover (\__mp_input219.A__gold );
  miter_def_prop #(1, "cover") \__mp_input219.Y__gold_cover (\__mp_input219.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input22.A__gold_cover (\__mp_input22.A__gold );
  miter_def_prop #(1, "cover") \__mp_input22.Y__gold_cover (\__mp_input22.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input220.A__gold_cover (\__mp_input220.A__gold );
  miter_def_prop #(1, "cover") \__mp_input220.Y__gold_cover (\__mp_input220.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input221.A__gold_cover (\__mp_input221.A__gold );
  miter_def_prop #(1, "cover") \__mp_input221.Y__gold_cover (\__mp_input221.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input222.A__gold_cover (\__mp_input222.A__gold );
  miter_def_prop #(1, "cover") \__mp_input222.Y__gold_cover (\__mp_input222.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input223.A__gold_cover (\__mp_input223.A__gold );
  miter_def_prop #(1, "cover") \__mp_input223.Y__gold_cover (\__mp_input223.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input224.A__gold_cover (\__mp_input224.A__gold );
  miter_def_prop #(1, "cover") \__mp_input224.Y__gold_cover (\__mp_input224.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input225.A__gold_cover (\__mp_input225.A__gold );
  miter_def_prop #(1, "cover") \__mp_input225.Y__gold_cover (\__mp_input225.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input226.A__gold_cover (\__mp_input226.A__gold );
  miter_def_prop #(1, "cover") \__mp_input226.Y__gold_cover (\__mp_input226.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input227.A__gold_cover (\__mp_input227.A__gold );
  miter_def_prop #(1, "cover") \__mp_input227.Y__gold_cover (\__mp_input227.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input228.A__gold_cover (\__mp_input228.A__gold );
  miter_def_prop #(1, "cover") \__mp_input228.Y__gold_cover (\__mp_input228.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input229.A__gold_cover (\__mp_input229.A__gold );
  miter_def_prop #(1, "cover") \__mp_input229.Y__gold_cover (\__mp_input229.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input23.A__gold_cover (\__mp_input23.A__gold );
  miter_def_prop #(1, "cover") \__mp_input23.Y__gold_cover (\__mp_input23.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input230.A__gold_cover (\__mp_input230.A__gold );
  miter_def_prop #(1, "cover") \__mp_input230.Y__gold_cover (\__mp_input230.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input231.A__gold_cover (\__mp_input231.A__gold );
  miter_def_prop #(1, "cover") \__mp_input231.Y__gold_cover (\__mp_input231.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input232.A__gold_cover (\__mp_input232.A__gold );
  miter_def_prop #(1, "cover") \__mp_input232.Y__gold_cover (\__mp_input232.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input233.A__gold_cover (\__mp_input233.A__gold );
  miter_def_prop #(1, "cover") \__mp_input233.Y__gold_cover (\__mp_input233.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input234.A__gold_cover (\__mp_input234.A__gold );
  miter_def_prop #(1, "cover") \__mp_input234.Y__gold_cover (\__mp_input234.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input235.A__gold_cover (\__mp_input235.A__gold );
  miter_def_prop #(1, "cover") \__mp_input235.Y__gold_cover (\__mp_input235.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input236.A__gold_cover (\__mp_input236.A__gold );
  miter_def_prop #(1, "cover") \__mp_input236.Y__gold_cover (\__mp_input236.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input237.A__gold_cover (\__mp_input237.A__gold );
  miter_def_prop #(1, "cover") \__mp_input237.Y__gold_cover (\__mp_input237.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input238.A__gold_cover (\__mp_input238.A__gold );
  miter_def_prop #(1, "cover") \__mp_input238.Y__gold_cover (\__mp_input238.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input239.A__gold_cover (\__mp_input239.A__gold );
  miter_def_prop #(1, "cover") \__mp_input239.Y__gold_cover (\__mp_input239.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input24.A__gold_cover (\__mp_input24.A__gold );
  miter_def_prop #(1, "cover") \__mp_input24.Y__gold_cover (\__mp_input24.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input240.A__gold_cover (\__mp_input240.A__gold );
  miter_def_prop #(1, "cover") \__mp_input240.Y__gold_cover (\__mp_input240.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input241.A__gold_cover (\__mp_input241.A__gold );
  miter_def_prop #(1, "cover") \__mp_input241.Y__gold_cover (\__mp_input241.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input242.A__gold_cover (\__mp_input242.A__gold );
  miter_def_prop #(1, "cover") \__mp_input242.Y__gold_cover (\__mp_input242.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input243.A__gold_cover (\__mp_input243.A__gold );
  miter_def_prop #(1, "cover") \__mp_input243.Y__gold_cover (\__mp_input243.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input244.A__gold_cover (\__mp_input244.A__gold );
  miter_def_prop #(1, "cover") \__mp_input244.Y__gold_cover (\__mp_input244.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input245.A__gold_cover (\__mp_input245.A__gold );
  miter_def_prop #(1, "cover") \__mp_input245.Y__gold_cover (\__mp_input245.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input246.A__gold_cover (\__mp_input246.A__gold );
  miter_def_prop #(1, "cover") \__mp_input246.Y__gold_cover (\__mp_input246.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input247.A__gold_cover (\__mp_input247.A__gold );
  miter_def_prop #(1, "cover") \__mp_input247.Y__gold_cover (\__mp_input247.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input248.A__gold_cover (\__mp_input248.A__gold );
  miter_def_prop #(1, "cover") \__mp_input248.Y__gold_cover (\__mp_input248.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input249.A__gold_cover (\__mp_input249.A__gold );
  miter_def_prop #(1, "cover") \__mp_input249.Y__gold_cover (\__mp_input249.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input25.A__gold_cover (\__mp_input25.A__gold );
  miter_def_prop #(1, "cover") \__mp_input25.Y__gold_cover (\__mp_input25.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input250.A__gold_cover (\__mp_input250.A__gold );
  miter_def_prop #(1, "cover") \__mp_input250.Y__gold_cover (\__mp_input250.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input251.A__gold_cover (\__mp_input251.A__gold );
  miter_def_prop #(1, "cover") \__mp_input251.Y__gold_cover (\__mp_input251.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input252.A__gold_cover (\__mp_input252.A__gold );
  miter_def_prop #(1, "cover") \__mp_input252.Y__gold_cover (\__mp_input252.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input253.A__gold_cover (\__mp_input253.A__gold );
  miter_def_prop #(1, "cover") \__mp_input253.Y__gold_cover (\__mp_input253.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input254.A__gold_cover (\__mp_input254.A__gold );
  miter_def_prop #(1, "cover") \__mp_input254.Y__gold_cover (\__mp_input254.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input255.A__gold_cover (\__mp_input255.A__gold );
  miter_def_prop #(1, "cover") \__mp_input255.Y__gold_cover (\__mp_input255.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input256.A__gold_cover (\__mp_input256.A__gold );
  miter_def_prop #(1, "cover") \__mp_input256.Y__gold_cover (\__mp_input256.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input257.A__gold_cover (\__mp_input257.A__gold );
  miter_def_prop #(1, "cover") \__mp_input257.Y__gold_cover (\__mp_input257.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input258.A__gold_cover (\__mp_input258.A__gold );
  miter_def_prop #(1, "cover") \__mp_input258.Y__gold_cover (\__mp_input258.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input26.A__gold_cover (\__mp_input26.A__gold );
  miter_def_prop #(1, "cover") \__mp_input26.Y__gold_cover (\__mp_input26.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input27.A__gold_cover (\__mp_input27.A__gold );
  miter_def_prop #(1, "cover") \__mp_input27.Y__gold_cover (\__mp_input27.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input28.A__gold_cover (\__mp_input28.A__gold );
  miter_def_prop #(1, "cover") \__mp_input28.Y__gold_cover (\__mp_input28.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input29.A__gold_cover (\__mp_input29.A__gold );
  miter_def_prop #(1, "cover") \__mp_input29.Y__gold_cover (\__mp_input29.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input3.A__gold_cover (\__mp_input3.A__gold );
  miter_def_prop #(1, "cover") \__mp_input3.Y__gold_cover (\__mp_input3.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input30.A__gold_cover (\__mp_input30.A__gold );
  miter_def_prop #(1, "cover") \__mp_input30.Y__gold_cover (\__mp_input30.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input31.A__gold_cover (\__mp_input31.A__gold );
  miter_def_prop #(1, "cover") \__mp_input31.Y__gold_cover (\__mp_input31.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input32.A__gold_cover (\__mp_input32.A__gold );
  miter_def_prop #(1, "cover") \__mp_input32.Y__gold_cover (\__mp_input32.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input33.A__gold_cover (\__mp_input33.A__gold );
  miter_def_prop #(1, "cover") \__mp_input33.Y__gold_cover (\__mp_input33.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input34.A__gold_cover (\__mp_input34.A__gold );
  miter_def_prop #(1, "cover") \__mp_input34.Y__gold_cover (\__mp_input34.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input35.A__gold_cover (\__mp_input35.A__gold );
  miter_def_prop #(1, "cover") \__mp_input35.Y__gold_cover (\__mp_input35.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input36.A__gold_cover (\__mp_input36.A__gold );
  miter_def_prop #(1, "cover") \__mp_input36.Y__gold_cover (\__mp_input36.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input37.A__gold_cover (\__mp_input37.A__gold );
  miter_def_prop #(1, "cover") \__mp_input37.Y__gold_cover (\__mp_input37.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input38.A__gold_cover (\__mp_input38.A__gold );
  miter_def_prop #(1, "cover") \__mp_input38.Y__gold_cover (\__mp_input38.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input39.A__gold_cover (\__mp_input39.A__gold );
  miter_def_prop #(1, "cover") \__mp_input39.Y__gold_cover (\__mp_input39.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input4.A__gold_cover (\__mp_input4.A__gold );
  miter_def_prop #(1, "cover") \__mp_input4.Y__gold_cover (\__mp_input4.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input40.A__gold_cover (\__mp_input40.A__gold );
  miter_def_prop #(1, "cover") \__mp_input40.Y__gold_cover (\__mp_input40.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input41.A__gold_cover (\__mp_input41.A__gold );
  miter_def_prop #(1, "cover") \__mp_input41.Y__gold_cover (\__mp_input41.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input42.A__gold_cover (\__mp_input42.A__gold );
  miter_def_prop #(1, "cover") \__mp_input42.Y__gold_cover (\__mp_input42.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input43.A__gold_cover (\__mp_input43.A__gold );
  miter_def_prop #(1, "cover") \__mp_input43.Y__gold_cover (\__mp_input43.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input44.A__gold_cover (\__mp_input44.A__gold );
  miter_def_prop #(1, "cover") \__mp_input44.Y__gold_cover (\__mp_input44.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input45.A__gold_cover (\__mp_input45.A__gold );
  miter_def_prop #(1, "cover") \__mp_input45.Y__gold_cover (\__mp_input45.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input46.A__gold_cover (\__mp_input46.A__gold );
  miter_def_prop #(1, "cover") \__mp_input46.Y__gold_cover (\__mp_input46.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input47.A__gold_cover (\__mp_input47.A__gold );
  miter_def_prop #(1, "cover") \__mp_input47.Y__gold_cover (\__mp_input47.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input48.A__gold_cover (\__mp_input48.A__gold );
  miter_def_prop #(1, "cover") \__mp_input48.Y__gold_cover (\__mp_input48.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input49.A__gold_cover (\__mp_input49.A__gold );
  miter_def_prop #(1, "cover") \__mp_input49.Y__gold_cover (\__mp_input49.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input5.A__gold_cover (\__mp_input5.A__gold );
  miter_def_prop #(1, "cover") \__mp_input5.Y__gold_cover (\__mp_input5.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input50.A__gold_cover (\__mp_input50.A__gold );
  miter_def_prop #(1, "cover") \__mp_input50.Y__gold_cover (\__mp_input50.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input51.A__gold_cover (\__mp_input51.A__gold );
  miter_def_prop #(1, "cover") \__mp_input51.Y__gold_cover (\__mp_input51.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input52.A__gold_cover (\__mp_input52.A__gold );
  miter_def_prop #(1, "cover") \__mp_input52.Y__gold_cover (\__mp_input52.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input53.A__gold_cover (\__mp_input53.A__gold );
  miter_def_prop #(1, "cover") \__mp_input53.Y__gold_cover (\__mp_input53.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input54.A__gold_cover (\__mp_input54.A__gold );
  miter_def_prop #(1, "cover") \__mp_input54.Y__gold_cover (\__mp_input54.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input55.A__gold_cover (\__mp_input55.A__gold );
  miter_def_prop #(1, "cover") \__mp_input55.Y__gold_cover (\__mp_input55.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input56.A__gold_cover (\__mp_input56.A__gold );
  miter_def_prop #(1, "cover") \__mp_input56.Y__gold_cover (\__mp_input56.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input57.A__gold_cover (\__mp_input57.A__gold );
  miter_def_prop #(1, "cover") \__mp_input57.Y__gold_cover (\__mp_input57.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input58.A__gold_cover (\__mp_input58.A__gold );
  miter_def_prop #(1, "cover") \__mp_input58.Y__gold_cover (\__mp_input58.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input59.A__gold_cover (\__mp_input59.A__gold );
  miter_def_prop #(1, "cover") \__mp_input59.Y__gold_cover (\__mp_input59.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input6.A__gold_cover (\__mp_input6.A__gold );
  miter_def_prop #(1, "cover") \__mp_input6.Y__gold_cover (\__mp_input6.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input60.A__gold_cover (\__mp_input60.A__gold );
  miter_def_prop #(1, "cover") \__mp_input60.Y__gold_cover (\__mp_input60.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input61.A__gold_cover (\__mp_input61.A__gold );
  miter_def_prop #(1, "cover") \__mp_input61.Y__gold_cover (\__mp_input61.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input62.A__gold_cover (\__mp_input62.A__gold );
  miter_def_prop #(1, "cover") \__mp_input62.Y__gold_cover (\__mp_input62.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input63.A__gold_cover (\__mp_input63.A__gold );
  miter_def_prop #(1, "cover") \__mp_input63.Y__gold_cover (\__mp_input63.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input64.A__gold_cover (\__mp_input64.A__gold );
  miter_def_prop #(1, "cover") \__mp_input64.Y__gold_cover (\__mp_input64.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input65.A__gold_cover (\__mp_input65.A__gold );
  miter_def_prop #(1, "cover") \__mp_input65.Y__gold_cover (\__mp_input65.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input66.A__gold_cover (\__mp_input66.A__gold );
  miter_def_prop #(1, "cover") \__mp_input66.Y__gold_cover (\__mp_input66.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input67.A__gold_cover (\__mp_input67.A__gold );
  miter_def_prop #(1, "cover") \__mp_input67.Y__gold_cover (\__mp_input67.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input68.A__gold_cover (\__mp_input68.A__gold );
  miter_def_prop #(1, "cover") \__mp_input68.Y__gold_cover (\__mp_input68.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input69.A__gold_cover (\__mp_input69.A__gold );
  miter_def_prop #(1, "cover") \__mp_input69.Y__gold_cover (\__mp_input69.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input7.A__gold_cover (\__mp_input7.A__gold );
  miter_def_prop #(1, "cover") \__mp_input7.Y__gold_cover (\__mp_input7.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input70.A__gold_cover (\__mp_input70.A__gold );
  miter_def_prop #(1, "cover") \__mp_input70.Y__gold_cover (\__mp_input70.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input71.A__gold_cover (\__mp_input71.A__gold );
  miter_def_prop #(1, "cover") \__mp_input71.Y__gold_cover (\__mp_input71.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input72.A__gold_cover (\__mp_input72.A__gold );
  miter_def_prop #(1, "cover") \__mp_input72.Y__gold_cover (\__mp_input72.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input73.A__gold_cover (\__mp_input73.A__gold );
  miter_def_prop #(1, "cover") \__mp_input73.Y__gold_cover (\__mp_input73.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input74.A__gold_cover (\__mp_input74.A__gold );
  miter_def_prop #(1, "cover") \__mp_input74.Y__gold_cover (\__mp_input74.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input75.A__gold_cover (\__mp_input75.A__gold );
  miter_def_prop #(1, "cover") \__mp_input75.Y__gold_cover (\__mp_input75.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input76.A__gold_cover (\__mp_input76.A__gold );
  miter_def_prop #(1, "cover") \__mp_input76.Y__gold_cover (\__mp_input76.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input77.A__gold_cover (\__mp_input77.A__gold );
  miter_def_prop #(1, "cover") \__mp_input77.Y__gold_cover (\__mp_input77.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input78.A__gold_cover (\__mp_input78.A__gold );
  miter_def_prop #(1, "cover") \__mp_input78.Y__gold_cover (\__mp_input78.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input79.A__gold_cover (\__mp_input79.A__gold );
  miter_def_prop #(1, "cover") \__mp_input79.Y__gold_cover (\__mp_input79.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input8.A__gold_cover (\__mp_input8.A__gold );
  miter_def_prop #(1, "cover") \__mp_input8.Y__gold_cover (\__mp_input8.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input80.A__gold_cover (\__mp_input80.A__gold );
  miter_def_prop #(1, "cover") \__mp_input80.Y__gold_cover (\__mp_input80.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input81.A__gold_cover (\__mp_input81.A__gold );
  miter_def_prop #(1, "cover") \__mp_input81.Y__gold_cover (\__mp_input81.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input82.A__gold_cover (\__mp_input82.A__gold );
  miter_def_prop #(1, "cover") \__mp_input82.Y__gold_cover (\__mp_input82.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input83.A__gold_cover (\__mp_input83.A__gold );
  miter_def_prop #(1, "cover") \__mp_input83.Y__gold_cover (\__mp_input83.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input84.A__gold_cover (\__mp_input84.A__gold );
  miter_def_prop #(1, "cover") \__mp_input84.Y__gold_cover (\__mp_input84.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input85.A__gold_cover (\__mp_input85.A__gold );
  miter_def_prop #(1, "cover") \__mp_input85.Y__gold_cover (\__mp_input85.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input86.A__gold_cover (\__mp_input86.A__gold );
  miter_def_prop #(1, "cover") \__mp_input86.Y__gold_cover (\__mp_input86.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input87.A__gold_cover (\__mp_input87.A__gold );
  miter_def_prop #(1, "cover") \__mp_input87.Y__gold_cover (\__mp_input87.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input88.A__gold_cover (\__mp_input88.A__gold );
  miter_def_prop #(1, "cover") \__mp_input88.Y__gold_cover (\__mp_input88.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input89.A__gold_cover (\__mp_input89.A__gold );
  miter_def_prop #(1, "cover") \__mp_input89.Y__gold_cover (\__mp_input89.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input9.A__gold_cover (\__mp_input9.A__gold );
  miter_def_prop #(1, "cover") \__mp_input9.Y__gold_cover (\__mp_input9.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input90.A__gold_cover (\__mp_input90.A__gold );
  miter_def_prop #(1, "cover") \__mp_input90.Y__gold_cover (\__mp_input90.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input91.A__gold_cover (\__mp_input91.A__gold );
  miter_def_prop #(1, "cover") \__mp_input91.Y__gold_cover (\__mp_input91.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input92.A__gold_cover (\__mp_input92.A__gold );
  miter_def_prop #(1, "cover") \__mp_input92.Y__gold_cover (\__mp_input92.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input93.A__gold_cover (\__mp_input93.A__gold );
  miter_def_prop #(1, "cover") \__mp_input93.Y__gold_cover (\__mp_input93.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input94.A__gold_cover (\__mp_input94.A__gold );
  miter_def_prop #(1, "cover") \__mp_input94.Y__gold_cover (\__mp_input94.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input95.A__gold_cover (\__mp_input95.A__gold );
  miter_def_prop #(1, "cover") \__mp_input95.Y__gold_cover (\__mp_input95.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input96.A__gold_cover (\__mp_input96.A__gold );
  miter_def_prop #(1, "cover") \__mp_input96.Y__gold_cover (\__mp_input96.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input97.A__gold_cover (\__mp_input97.A__gold );
  miter_def_prop #(1, "cover") \__mp_input97.Y__gold_cover (\__mp_input97.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input98.A__gold_cover (\__mp_input98.A__gold );
  miter_def_prop #(1, "cover") \__mp_input98.Y__gold_cover (\__mp_input98.Y__gold );
  miter_def_prop #(1, "cover") \__mp_input99.A__gold_cover (\__mp_input99.A__gold );
  miter_def_prop #(1, "cover") \__mp_input99.Y__gold_cover (\__mp_input99.Y__gold );
  miter_def_prop #(1, "cover") \__mp_ld_r$_DFF_P_.CLK__gold_cover (\__mp_ld_r$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_ld_r$_DFF_P_.D__gold_cover (\__mp_ld_r$_DFF_P_.D__gold );
  miter_def_prop #(1, "cover") \__mp_output259.A__gold_cover (\__mp_output259.A__gold );
  miter_def_prop #(1, "cover") \__mp_output259.Y__gold_cover (\__mp_output259.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output260.A__gold_cover (\__mp_output260.A__gold );
  miter_def_prop #(1, "cover") \__mp_output260.Y__gold_cover (\__mp_output260.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output261.A__gold_cover (\__mp_output261.A__gold );
  miter_def_prop #(1, "cover") \__mp_output261.Y__gold_cover (\__mp_output261.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output262.A__gold_cover (\__mp_output262.A__gold );
  miter_def_prop #(1, "cover") \__mp_output262.Y__gold_cover (\__mp_output262.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output263.A__gold_cover (\__mp_output263.A__gold );
  miter_def_prop #(1, "cover") \__mp_output263.Y__gold_cover (\__mp_output263.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output264.A__gold_cover (\__mp_output264.A__gold );
  miter_def_prop #(1, "cover") \__mp_output264.Y__gold_cover (\__mp_output264.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output265.A__gold_cover (\__mp_output265.A__gold );
  miter_def_prop #(1, "cover") \__mp_output265.Y__gold_cover (\__mp_output265.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output266.A__gold_cover (\__mp_output266.A__gold );
  miter_def_prop #(1, "cover") \__mp_output266.Y__gold_cover (\__mp_output266.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output267.A__gold_cover (\__mp_output267.A__gold );
  miter_def_prop #(1, "cover") \__mp_output267.Y__gold_cover (\__mp_output267.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output268.A__gold_cover (\__mp_output268.A__gold );
  miter_def_prop #(1, "cover") \__mp_output268.Y__gold_cover (\__mp_output268.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output269.A__gold_cover (\__mp_output269.A__gold );
  miter_def_prop #(1, "cover") \__mp_output269.Y__gold_cover (\__mp_output269.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output270.A__gold_cover (\__mp_output270.A__gold );
  miter_def_prop #(1, "cover") \__mp_output270.Y__gold_cover (\__mp_output270.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output271.A__gold_cover (\__mp_output271.A__gold );
  miter_def_prop #(1, "cover") \__mp_output271.Y__gold_cover (\__mp_output271.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output272.A__gold_cover (\__mp_output272.A__gold );
  miter_def_prop #(1, "cover") \__mp_output272.Y__gold_cover (\__mp_output272.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output273.A__gold_cover (\__mp_output273.A__gold );
  miter_def_prop #(1, "cover") \__mp_output273.Y__gold_cover (\__mp_output273.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output274.A__gold_cover (\__mp_output274.A__gold );
  miter_def_prop #(1, "cover") \__mp_output274.Y__gold_cover (\__mp_output274.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output275.A__gold_cover (\__mp_output275.A__gold );
  miter_def_prop #(1, "cover") \__mp_output275.Y__gold_cover (\__mp_output275.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output276.A__gold_cover (\__mp_output276.A__gold );
  miter_def_prop #(1, "cover") \__mp_output276.Y__gold_cover (\__mp_output276.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output277.A__gold_cover (\__mp_output277.A__gold );
  miter_def_prop #(1, "cover") \__mp_output277.Y__gold_cover (\__mp_output277.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output278.A__gold_cover (\__mp_output278.A__gold );
  miter_def_prop #(1, "cover") \__mp_output278.Y__gold_cover (\__mp_output278.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output279.A__gold_cover (\__mp_output279.A__gold );
  miter_def_prop #(1, "cover") \__mp_output279.Y__gold_cover (\__mp_output279.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output280.A__gold_cover (\__mp_output280.A__gold );
  miter_def_prop #(1, "cover") \__mp_output280.Y__gold_cover (\__mp_output280.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output281.A__gold_cover (\__mp_output281.A__gold );
  miter_def_prop #(1, "cover") \__mp_output281.Y__gold_cover (\__mp_output281.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output282.A__gold_cover (\__mp_output282.A__gold );
  miter_def_prop #(1, "cover") \__mp_output282.Y__gold_cover (\__mp_output282.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output283.A__gold_cover (\__mp_output283.A__gold );
  miter_def_prop #(1, "cover") \__mp_output283.Y__gold_cover (\__mp_output283.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output284.A__gold_cover (\__mp_output284.A__gold );
  miter_def_prop #(1, "cover") \__mp_output284.Y__gold_cover (\__mp_output284.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output285.A__gold_cover (\__mp_output285.A__gold );
  miter_def_prop #(1, "cover") \__mp_output285.Y__gold_cover (\__mp_output285.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output286.A__gold_cover (\__mp_output286.A__gold );
  miter_def_prop #(1, "cover") \__mp_output286.Y__gold_cover (\__mp_output286.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output287.A__gold_cover (\__mp_output287.A__gold );
  miter_def_prop #(1, "cover") \__mp_output287.Y__gold_cover (\__mp_output287.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output288.A__gold_cover (\__mp_output288.A__gold );
  miter_def_prop #(1, "cover") \__mp_output288.Y__gold_cover (\__mp_output288.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output289.A__gold_cover (\__mp_output289.A__gold );
  miter_def_prop #(1, "cover") \__mp_output289.Y__gold_cover (\__mp_output289.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output290.A__gold_cover (\__mp_output290.A__gold );
  miter_def_prop #(1, "cover") \__mp_output290.Y__gold_cover (\__mp_output290.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output291.A__gold_cover (\__mp_output291.A__gold );
  miter_def_prop #(1, "cover") \__mp_output291.Y__gold_cover (\__mp_output291.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output292.A__gold_cover (\__mp_output292.A__gold );
  miter_def_prop #(1, "cover") \__mp_output292.Y__gold_cover (\__mp_output292.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output293.A__gold_cover (\__mp_output293.A__gold );
  miter_def_prop #(1, "cover") \__mp_output293.Y__gold_cover (\__mp_output293.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output294.A__gold_cover (\__mp_output294.A__gold );
  miter_def_prop #(1, "cover") \__mp_output294.Y__gold_cover (\__mp_output294.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output295.A__gold_cover (\__mp_output295.A__gold );
  miter_def_prop #(1, "cover") \__mp_output295.Y__gold_cover (\__mp_output295.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output296.A__gold_cover (\__mp_output296.A__gold );
  miter_def_prop #(1, "cover") \__mp_output296.Y__gold_cover (\__mp_output296.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output297.A__gold_cover (\__mp_output297.A__gold );
  miter_def_prop #(1, "cover") \__mp_output297.Y__gold_cover (\__mp_output297.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output298.A__gold_cover (\__mp_output298.A__gold );
  miter_def_prop #(1, "cover") \__mp_output298.Y__gold_cover (\__mp_output298.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output299.A__gold_cover (\__mp_output299.A__gold );
  miter_def_prop #(1, "cover") \__mp_output299.Y__gold_cover (\__mp_output299.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output300.A__gold_cover (\__mp_output300.A__gold );
  miter_def_prop #(1, "cover") \__mp_output300.Y__gold_cover (\__mp_output300.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output301.A__gold_cover (\__mp_output301.A__gold );
  miter_def_prop #(1, "cover") \__mp_output301.Y__gold_cover (\__mp_output301.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output302.A__gold_cover (\__mp_output302.A__gold );
  miter_def_prop #(1, "cover") \__mp_output302.Y__gold_cover (\__mp_output302.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output303.A__gold_cover (\__mp_output303.A__gold );
  miter_def_prop #(1, "cover") \__mp_output303.Y__gold_cover (\__mp_output303.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output304.A__gold_cover (\__mp_output304.A__gold );
  miter_def_prop #(1, "cover") \__mp_output304.Y__gold_cover (\__mp_output304.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output305.A__gold_cover (\__mp_output305.A__gold );
  miter_def_prop #(1, "cover") \__mp_output305.Y__gold_cover (\__mp_output305.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output306.A__gold_cover (\__mp_output306.A__gold );
  miter_def_prop #(1, "cover") \__mp_output306.Y__gold_cover (\__mp_output306.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output307.A__gold_cover (\__mp_output307.A__gold );
  miter_def_prop #(1, "cover") \__mp_output307.Y__gold_cover (\__mp_output307.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output308.A__gold_cover (\__mp_output308.A__gold );
  miter_def_prop #(1, "cover") \__mp_output308.Y__gold_cover (\__mp_output308.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output309.A__gold_cover (\__mp_output309.A__gold );
  miter_def_prop #(1, "cover") \__mp_output309.Y__gold_cover (\__mp_output309.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output310.A__gold_cover (\__mp_output310.A__gold );
  miter_def_prop #(1, "cover") \__mp_output310.Y__gold_cover (\__mp_output310.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output311.A__gold_cover (\__mp_output311.A__gold );
  miter_def_prop #(1, "cover") \__mp_output311.Y__gold_cover (\__mp_output311.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output312.A__gold_cover (\__mp_output312.A__gold );
  miter_def_prop #(1, "cover") \__mp_output312.Y__gold_cover (\__mp_output312.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output313.A__gold_cover (\__mp_output313.A__gold );
  miter_def_prop #(1, "cover") \__mp_output313.Y__gold_cover (\__mp_output313.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output314.A__gold_cover (\__mp_output314.A__gold );
  miter_def_prop #(1, "cover") \__mp_output314.Y__gold_cover (\__mp_output314.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output315.A__gold_cover (\__mp_output315.A__gold );
  miter_def_prop #(1, "cover") \__mp_output315.Y__gold_cover (\__mp_output315.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output316.A__gold_cover (\__mp_output316.A__gold );
  miter_def_prop #(1, "cover") \__mp_output316.Y__gold_cover (\__mp_output316.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output317.A__gold_cover (\__mp_output317.A__gold );
  miter_def_prop #(1, "cover") \__mp_output317.Y__gold_cover (\__mp_output317.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output318.A__gold_cover (\__mp_output318.A__gold );
  miter_def_prop #(1, "cover") \__mp_output318.Y__gold_cover (\__mp_output318.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output319.A__gold_cover (\__mp_output319.A__gold );
  miter_def_prop #(1, "cover") \__mp_output319.Y__gold_cover (\__mp_output319.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output320.A__gold_cover (\__mp_output320.A__gold );
  miter_def_prop #(1, "cover") \__mp_output320.Y__gold_cover (\__mp_output320.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output321.A__gold_cover (\__mp_output321.A__gold );
  miter_def_prop #(1, "cover") \__mp_output321.Y__gold_cover (\__mp_output321.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output322.A__gold_cover (\__mp_output322.A__gold );
  miter_def_prop #(1, "cover") \__mp_output322.Y__gold_cover (\__mp_output322.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output323.A__gold_cover (\__mp_output323.A__gold );
  miter_def_prop #(1, "cover") \__mp_output323.Y__gold_cover (\__mp_output323.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output324.A__gold_cover (\__mp_output324.A__gold );
  miter_def_prop #(1, "cover") \__mp_output324.Y__gold_cover (\__mp_output324.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output325.A__gold_cover (\__mp_output325.A__gold );
  miter_def_prop #(1, "cover") \__mp_output325.Y__gold_cover (\__mp_output325.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output326.A__gold_cover (\__mp_output326.A__gold );
  miter_def_prop #(1, "cover") \__mp_output326.Y__gold_cover (\__mp_output326.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output327.A__gold_cover (\__mp_output327.A__gold );
  miter_def_prop #(1, "cover") \__mp_output327.Y__gold_cover (\__mp_output327.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output328.A__gold_cover (\__mp_output328.A__gold );
  miter_def_prop #(1, "cover") \__mp_output328.Y__gold_cover (\__mp_output328.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output329.A__gold_cover (\__mp_output329.A__gold );
  miter_def_prop #(1, "cover") \__mp_output329.Y__gold_cover (\__mp_output329.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output330.A__gold_cover (\__mp_output330.A__gold );
  miter_def_prop #(1, "cover") \__mp_output330.Y__gold_cover (\__mp_output330.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output331.A__gold_cover (\__mp_output331.A__gold );
  miter_def_prop #(1, "cover") \__mp_output331.Y__gold_cover (\__mp_output331.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output332.A__gold_cover (\__mp_output332.A__gold );
  miter_def_prop #(1, "cover") \__mp_output332.Y__gold_cover (\__mp_output332.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output333.A__gold_cover (\__mp_output333.A__gold );
  miter_def_prop #(1, "cover") \__mp_output333.Y__gold_cover (\__mp_output333.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output334.A__gold_cover (\__mp_output334.A__gold );
  miter_def_prop #(1, "cover") \__mp_output334.Y__gold_cover (\__mp_output334.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output335.A__gold_cover (\__mp_output335.A__gold );
  miter_def_prop #(1, "cover") \__mp_output335.Y__gold_cover (\__mp_output335.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output336.A__gold_cover (\__mp_output336.A__gold );
  miter_def_prop #(1, "cover") \__mp_output336.Y__gold_cover (\__mp_output336.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output337.A__gold_cover (\__mp_output337.A__gold );
  miter_def_prop #(1, "cover") \__mp_output337.Y__gold_cover (\__mp_output337.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output338.A__gold_cover (\__mp_output338.A__gold );
  miter_def_prop #(1, "cover") \__mp_output338.Y__gold_cover (\__mp_output338.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output339.A__gold_cover (\__mp_output339.A__gold );
  miter_def_prop #(1, "cover") \__mp_output339.Y__gold_cover (\__mp_output339.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output340.A__gold_cover (\__mp_output340.A__gold );
  miter_def_prop #(1, "cover") \__mp_output340.Y__gold_cover (\__mp_output340.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output341.A__gold_cover (\__mp_output341.A__gold );
  miter_def_prop #(1, "cover") \__mp_output341.Y__gold_cover (\__mp_output341.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output342.A__gold_cover (\__mp_output342.A__gold );
  miter_def_prop #(1, "cover") \__mp_output342.Y__gold_cover (\__mp_output342.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output343.A__gold_cover (\__mp_output343.A__gold );
  miter_def_prop #(1, "cover") \__mp_output343.Y__gold_cover (\__mp_output343.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output344.A__gold_cover (\__mp_output344.A__gold );
  miter_def_prop #(1, "cover") \__mp_output344.Y__gold_cover (\__mp_output344.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output345.A__gold_cover (\__mp_output345.A__gold );
  miter_def_prop #(1, "cover") \__mp_output345.Y__gold_cover (\__mp_output345.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output346.A__gold_cover (\__mp_output346.A__gold );
  miter_def_prop #(1, "cover") \__mp_output346.Y__gold_cover (\__mp_output346.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output347.A__gold_cover (\__mp_output347.A__gold );
  miter_def_prop #(1, "cover") \__mp_output347.Y__gold_cover (\__mp_output347.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output348.A__gold_cover (\__mp_output348.A__gold );
  miter_def_prop #(1, "cover") \__mp_output348.Y__gold_cover (\__mp_output348.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output349.A__gold_cover (\__mp_output349.A__gold );
  miter_def_prop #(1, "cover") \__mp_output349.Y__gold_cover (\__mp_output349.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output350.A__gold_cover (\__mp_output350.A__gold );
  miter_def_prop #(1, "cover") \__mp_output350.Y__gold_cover (\__mp_output350.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output351.A__gold_cover (\__mp_output351.A__gold );
  miter_def_prop #(1, "cover") \__mp_output351.Y__gold_cover (\__mp_output351.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output352.A__gold_cover (\__mp_output352.A__gold );
  miter_def_prop #(1, "cover") \__mp_output352.Y__gold_cover (\__mp_output352.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output353.A__gold_cover (\__mp_output353.A__gold );
  miter_def_prop #(1, "cover") \__mp_output353.Y__gold_cover (\__mp_output353.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output354.A__gold_cover (\__mp_output354.A__gold );
  miter_def_prop #(1, "cover") \__mp_output354.Y__gold_cover (\__mp_output354.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output355.A__gold_cover (\__mp_output355.A__gold );
  miter_def_prop #(1, "cover") \__mp_output355.Y__gold_cover (\__mp_output355.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output356.A__gold_cover (\__mp_output356.A__gold );
  miter_def_prop #(1, "cover") \__mp_output356.Y__gold_cover (\__mp_output356.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output357.A__gold_cover (\__mp_output357.A__gold );
  miter_def_prop #(1, "cover") \__mp_output357.Y__gold_cover (\__mp_output357.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output358.A__gold_cover (\__mp_output358.A__gold );
  miter_def_prop #(1, "cover") \__mp_output358.Y__gold_cover (\__mp_output358.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output359.A__gold_cover (\__mp_output359.A__gold );
  miter_def_prop #(1, "cover") \__mp_output359.Y__gold_cover (\__mp_output359.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output360.A__gold_cover (\__mp_output360.A__gold );
  miter_def_prop #(1, "cover") \__mp_output360.Y__gold_cover (\__mp_output360.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output361.A__gold_cover (\__mp_output361.A__gold );
  miter_def_prop #(1, "cover") \__mp_output361.Y__gold_cover (\__mp_output361.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output362.A__gold_cover (\__mp_output362.A__gold );
  miter_def_prop #(1, "cover") \__mp_output362.Y__gold_cover (\__mp_output362.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output363.A__gold_cover (\__mp_output363.A__gold );
  miter_def_prop #(1, "cover") \__mp_output363.Y__gold_cover (\__mp_output363.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output364.A__gold_cover (\__mp_output364.A__gold );
  miter_def_prop #(1, "cover") \__mp_output364.Y__gold_cover (\__mp_output364.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output365.A__gold_cover (\__mp_output365.A__gold );
  miter_def_prop #(1, "cover") \__mp_output365.Y__gold_cover (\__mp_output365.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output366.A__gold_cover (\__mp_output366.A__gold );
  miter_def_prop #(1, "cover") \__mp_output366.Y__gold_cover (\__mp_output366.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output367.A__gold_cover (\__mp_output367.A__gold );
  miter_def_prop #(1, "cover") \__mp_output367.Y__gold_cover (\__mp_output367.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output368.A__gold_cover (\__mp_output368.A__gold );
  miter_def_prop #(1, "cover") \__mp_output368.Y__gold_cover (\__mp_output368.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output369.A__gold_cover (\__mp_output369.A__gold );
  miter_def_prop #(1, "cover") \__mp_output369.Y__gold_cover (\__mp_output369.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output370.A__gold_cover (\__mp_output370.A__gold );
  miter_def_prop #(1, "cover") \__mp_output370.Y__gold_cover (\__mp_output370.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output371.A__gold_cover (\__mp_output371.A__gold );
  miter_def_prop #(1, "cover") \__mp_output371.Y__gold_cover (\__mp_output371.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output372.A__gold_cover (\__mp_output372.A__gold );
  miter_def_prop #(1, "cover") \__mp_output372.Y__gold_cover (\__mp_output372.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output373.A__gold_cover (\__mp_output373.A__gold );
  miter_def_prop #(1, "cover") \__mp_output373.Y__gold_cover (\__mp_output373.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output374.A__gold_cover (\__mp_output374.A__gold );
  miter_def_prop #(1, "cover") \__mp_output374.Y__gold_cover (\__mp_output374.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output375.A__gold_cover (\__mp_output375.A__gold );
  miter_def_prop #(1, "cover") \__mp_output375.Y__gold_cover (\__mp_output375.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output376.A__gold_cover (\__mp_output376.A__gold );
  miter_def_prop #(1, "cover") \__mp_output376.Y__gold_cover (\__mp_output376.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output377.A__gold_cover (\__mp_output377.A__gold );
  miter_def_prop #(1, "cover") \__mp_output377.Y__gold_cover (\__mp_output377.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output378.A__gold_cover (\__mp_output378.A__gold );
  miter_def_prop #(1, "cover") \__mp_output378.Y__gold_cover (\__mp_output378.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output379.A__gold_cover (\__mp_output379.A__gold );
  miter_def_prop #(1, "cover") \__mp_output379.Y__gold_cover (\__mp_output379.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output380.A__gold_cover (\__mp_output380.A__gold );
  miter_def_prop #(1, "cover") \__mp_output380.Y__gold_cover (\__mp_output380.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output381.A__gold_cover (\__mp_output381.A__gold );
  miter_def_prop #(1, "cover") \__mp_output381.Y__gold_cover (\__mp_output381.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output382.A__gold_cover (\__mp_output382.A__gold );
  miter_def_prop #(1, "cover") \__mp_output382.Y__gold_cover (\__mp_output382.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output383.A__gold_cover (\__mp_output383.A__gold );
  miter_def_prop #(1, "cover") \__mp_output383.Y__gold_cover (\__mp_output383.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output384.A__gold_cover (\__mp_output384.A__gold );
  miter_def_prop #(1, "cover") \__mp_output384.Y__gold_cover (\__mp_output384.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output385.A__gold_cover (\__mp_output385.A__gold );
  miter_def_prop #(1, "cover") \__mp_output385.Y__gold_cover (\__mp_output385.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output386.A__gold_cover (\__mp_output386.A__gold );
  miter_def_prop #(1, "cover") \__mp_output386.Y__gold_cover (\__mp_output386.Y__gold );
  miter_def_prop #(1, "cover") \__mp_output387.A__gold_cover (\__mp_output387.A__gold );
  miter_def_prop #(1, "cover") \__mp_output387.Y__gold_cover (\__mp_output387.Y__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa00_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa01_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa02_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa03_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa10_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa11_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa12_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa13_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa20_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa21_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa22_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa23_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa30_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa31_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa32_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[0]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[1]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[2]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[3]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[4]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[5]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[6]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[7]$_DFF_P_.CLK__gold_cover (\__mp_sa33_sr[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[0]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[0]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[100]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[100]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[101]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[101]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[102]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[102]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[103]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[103]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[104]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[104]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[105]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[105]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[106]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[106]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[107]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[107]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[108]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[108]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[109]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[109]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[10]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[10]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[110]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[110]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[111]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[111]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[112]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[112]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[113]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[113]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[114]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[114]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[115]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[115]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[116]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[116]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[117]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[117]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[118]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[118]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[119]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[119]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[11]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[11]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[120]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[120]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[121]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[121]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[122]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[122]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[123]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[123]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[124]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[124]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[125]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[125]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[126]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[126]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[127]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[127]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[12]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[12]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[13]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[13]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[14]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[14]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[15]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[15]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[16]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[16]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[17]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[17]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[18]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[18]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[19]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[19]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[1]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[1]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[20]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[20]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[21]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[21]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[22]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[22]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[23]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[23]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[24]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[24]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[25]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[25]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[26]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[26]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[27]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[27]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[28]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[28]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[29]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[29]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[2]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[2]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[30]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[30]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[31]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[31]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[32]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[32]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[33]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[33]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[34]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[34]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[35]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[35]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[36]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[36]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[37]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[37]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[38]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[38]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[39]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[39]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[3]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[3]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[40]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[40]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[41]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[41]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[42]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[42]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[43]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[43]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[44]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[44]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[45]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[45]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[46]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[46]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[47]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[47]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[48]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[48]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[49]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[49]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[4]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[4]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[50]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[50]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[51]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[51]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[52]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[52]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[53]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[53]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[54]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[54]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[55]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[55]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[56]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[56]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[57]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[57]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[58]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[58]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[59]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[59]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[5]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[5]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[60]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[60]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[61]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[61]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[62]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[62]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[63]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[63]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[64]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[64]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[65]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[65]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[66]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[66]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[67]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[67]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[68]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[68]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[69]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[69]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[6]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[6]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[70]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[70]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[71]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[71]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[72]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[72]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[73]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[73]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[74]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[74]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[75]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[75]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[76]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[76]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[77]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[77]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[78]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[78]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[79]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[79]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[7]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[7]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[80]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[80]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[81]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[81]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[82]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[82]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[83]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[83]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[84]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[84]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[85]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[85]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[86]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[86]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[87]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[87]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[88]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[88]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[89]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[89]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[8]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[8]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[90]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[90]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[91]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[91]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[92]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[92]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[93]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[93]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[94]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[94]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[95]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[95]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[96]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[96]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[97]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[97]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[98]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[98]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[99]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[99]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_in_r[9]$_DFFE_PP_.CLK__gold_cover (\__mp_text_in_r[9]$_DFFE_PP_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[0]$_DFF_P_.CLK__gold_cover (\__mp_text_out[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[0]$_DFF_P_.QN__gold_cover (\__mp_text_out[0]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[100]$_DFF_P_.CLK__gold_cover (\__mp_text_out[100]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[100]$_DFF_P_.QN__gold_cover (\__mp_text_out[100]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[101]$_DFF_P_.CLK__gold_cover (\__mp_text_out[101]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[101]$_DFF_P_.QN__gold_cover (\__mp_text_out[101]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[102]$_DFF_P_.CLK__gold_cover (\__mp_text_out[102]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[102]$_DFF_P_.QN__gold_cover (\__mp_text_out[102]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[103]$_DFF_P_.CLK__gold_cover (\__mp_text_out[103]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[103]$_DFF_P_.QN__gold_cover (\__mp_text_out[103]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[104]$_DFF_P_.CLK__gold_cover (\__mp_text_out[104]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[104]$_DFF_P_.QN__gold_cover (\__mp_text_out[104]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[105]$_DFF_P_.CLK__gold_cover (\__mp_text_out[105]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[105]$_DFF_P_.QN__gold_cover (\__mp_text_out[105]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[106]$_DFF_P_.CLK__gold_cover (\__mp_text_out[106]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[106]$_DFF_P_.QN__gold_cover (\__mp_text_out[106]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[107]$_DFF_P_.CLK__gold_cover (\__mp_text_out[107]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[107]$_DFF_P_.QN__gold_cover (\__mp_text_out[107]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[108]$_DFF_P_.CLK__gold_cover (\__mp_text_out[108]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[108]$_DFF_P_.QN__gold_cover (\__mp_text_out[108]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[109]$_DFF_P_.CLK__gold_cover (\__mp_text_out[109]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[109]$_DFF_P_.QN__gold_cover (\__mp_text_out[109]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[10]$_DFF_P_.CLK__gold_cover (\__mp_text_out[10]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[10]$_DFF_P_.QN__gold_cover (\__mp_text_out[10]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[110]$_DFF_P_.CLK__gold_cover (\__mp_text_out[110]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[110]$_DFF_P_.QN__gold_cover (\__mp_text_out[110]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[111]$_DFF_P_.CLK__gold_cover (\__mp_text_out[111]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[111]$_DFF_P_.QN__gold_cover (\__mp_text_out[111]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[112]$_DFF_P_.CLK__gold_cover (\__mp_text_out[112]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[112]$_DFF_P_.QN__gold_cover (\__mp_text_out[112]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[113]$_DFF_P_.CLK__gold_cover (\__mp_text_out[113]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[113]$_DFF_P_.QN__gold_cover (\__mp_text_out[113]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[114]$_DFF_P_.CLK__gold_cover (\__mp_text_out[114]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[114]$_DFF_P_.QN__gold_cover (\__mp_text_out[114]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[115]$_DFF_P_.CLK__gold_cover (\__mp_text_out[115]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[115]$_DFF_P_.QN__gold_cover (\__mp_text_out[115]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[116]$_DFF_P_.CLK__gold_cover (\__mp_text_out[116]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[116]$_DFF_P_.QN__gold_cover (\__mp_text_out[116]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[117]$_DFF_P_.CLK__gold_cover (\__mp_text_out[117]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[117]$_DFF_P_.QN__gold_cover (\__mp_text_out[117]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[118]$_DFF_P_.CLK__gold_cover (\__mp_text_out[118]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[118]$_DFF_P_.QN__gold_cover (\__mp_text_out[118]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[119]$_DFF_P_.CLK__gold_cover (\__mp_text_out[119]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[119]$_DFF_P_.QN__gold_cover (\__mp_text_out[119]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[11]$_DFF_P_.CLK__gold_cover (\__mp_text_out[11]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[11]$_DFF_P_.QN__gold_cover (\__mp_text_out[11]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[120]$_DFF_P_.CLK__gold_cover (\__mp_text_out[120]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[120]$_DFF_P_.QN__gold_cover (\__mp_text_out[120]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[121]$_DFF_P_.CLK__gold_cover (\__mp_text_out[121]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[121]$_DFF_P_.QN__gold_cover (\__mp_text_out[121]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[122]$_DFF_P_.CLK__gold_cover (\__mp_text_out[122]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[122]$_DFF_P_.QN__gold_cover (\__mp_text_out[122]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[123]$_DFF_P_.CLK__gold_cover (\__mp_text_out[123]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[123]$_DFF_P_.QN__gold_cover (\__mp_text_out[123]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[124]$_DFF_P_.CLK__gold_cover (\__mp_text_out[124]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[124]$_DFF_P_.QN__gold_cover (\__mp_text_out[124]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[125]$_DFF_P_.CLK__gold_cover (\__mp_text_out[125]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[125]$_DFF_P_.QN__gold_cover (\__mp_text_out[125]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[126]$_DFF_P_.CLK__gold_cover (\__mp_text_out[126]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[126]$_DFF_P_.QN__gold_cover (\__mp_text_out[126]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[127]$_DFF_P_.CLK__gold_cover (\__mp_text_out[127]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[127]$_DFF_P_.QN__gold_cover (\__mp_text_out[127]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[12]$_DFF_P_.CLK__gold_cover (\__mp_text_out[12]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[12]$_DFF_P_.QN__gold_cover (\__mp_text_out[12]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[13]$_DFF_P_.CLK__gold_cover (\__mp_text_out[13]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[13]$_DFF_P_.QN__gold_cover (\__mp_text_out[13]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[14]$_DFF_P_.CLK__gold_cover (\__mp_text_out[14]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[14]$_DFF_P_.QN__gold_cover (\__mp_text_out[14]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[15]$_DFF_P_.CLK__gold_cover (\__mp_text_out[15]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[15]$_DFF_P_.QN__gold_cover (\__mp_text_out[15]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[16]$_DFF_P_.CLK__gold_cover (\__mp_text_out[16]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[16]$_DFF_P_.QN__gold_cover (\__mp_text_out[16]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[17]$_DFF_P_.CLK__gold_cover (\__mp_text_out[17]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[17]$_DFF_P_.QN__gold_cover (\__mp_text_out[17]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[18]$_DFF_P_.CLK__gold_cover (\__mp_text_out[18]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[18]$_DFF_P_.QN__gold_cover (\__mp_text_out[18]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[19]$_DFF_P_.CLK__gold_cover (\__mp_text_out[19]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[19]$_DFF_P_.QN__gold_cover (\__mp_text_out[19]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[1]$_DFF_P_.CLK__gold_cover (\__mp_text_out[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[1]$_DFF_P_.QN__gold_cover (\__mp_text_out[1]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[20]$_DFF_P_.CLK__gold_cover (\__mp_text_out[20]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[20]$_DFF_P_.QN__gold_cover (\__mp_text_out[20]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[21]$_DFF_P_.CLK__gold_cover (\__mp_text_out[21]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[21]$_DFF_P_.QN__gold_cover (\__mp_text_out[21]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[22]$_DFF_P_.CLK__gold_cover (\__mp_text_out[22]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[22]$_DFF_P_.QN__gold_cover (\__mp_text_out[22]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[23]$_DFF_P_.CLK__gold_cover (\__mp_text_out[23]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[23]$_DFF_P_.QN__gold_cover (\__mp_text_out[23]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[24]$_DFF_P_.CLK__gold_cover (\__mp_text_out[24]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[24]$_DFF_P_.QN__gold_cover (\__mp_text_out[24]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[25]$_DFF_P_.CLK__gold_cover (\__mp_text_out[25]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[25]$_DFF_P_.QN__gold_cover (\__mp_text_out[25]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[26]$_DFF_P_.CLK__gold_cover (\__mp_text_out[26]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[26]$_DFF_P_.QN__gold_cover (\__mp_text_out[26]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[27]$_DFF_P_.CLK__gold_cover (\__mp_text_out[27]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[27]$_DFF_P_.QN__gold_cover (\__mp_text_out[27]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[28]$_DFF_P_.CLK__gold_cover (\__mp_text_out[28]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[28]$_DFF_P_.QN__gold_cover (\__mp_text_out[28]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[29]$_DFF_P_.CLK__gold_cover (\__mp_text_out[29]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[29]$_DFF_P_.QN__gold_cover (\__mp_text_out[29]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[2]$_DFF_P_.CLK__gold_cover (\__mp_text_out[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[2]$_DFF_P_.QN__gold_cover (\__mp_text_out[2]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[30]$_DFF_P_.CLK__gold_cover (\__mp_text_out[30]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[30]$_DFF_P_.QN__gold_cover (\__mp_text_out[30]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[31]$_DFF_P_.CLK__gold_cover (\__mp_text_out[31]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[31]$_DFF_P_.QN__gold_cover (\__mp_text_out[31]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[32]$_DFF_P_.CLK__gold_cover (\__mp_text_out[32]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[32]$_DFF_P_.QN__gold_cover (\__mp_text_out[32]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[33]$_DFF_P_.CLK__gold_cover (\__mp_text_out[33]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[33]$_DFF_P_.QN__gold_cover (\__mp_text_out[33]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[34]$_DFF_P_.CLK__gold_cover (\__mp_text_out[34]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[34]$_DFF_P_.QN__gold_cover (\__mp_text_out[34]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[35]$_DFF_P_.CLK__gold_cover (\__mp_text_out[35]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[35]$_DFF_P_.QN__gold_cover (\__mp_text_out[35]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[36]$_DFF_P_.CLK__gold_cover (\__mp_text_out[36]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[36]$_DFF_P_.QN__gold_cover (\__mp_text_out[36]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[37]$_DFF_P_.CLK__gold_cover (\__mp_text_out[37]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[37]$_DFF_P_.QN__gold_cover (\__mp_text_out[37]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[38]$_DFF_P_.CLK__gold_cover (\__mp_text_out[38]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[38]$_DFF_P_.QN__gold_cover (\__mp_text_out[38]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[39]$_DFF_P_.CLK__gold_cover (\__mp_text_out[39]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[39]$_DFF_P_.QN__gold_cover (\__mp_text_out[39]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[3]$_DFF_P_.CLK__gold_cover (\__mp_text_out[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[3]$_DFF_P_.QN__gold_cover (\__mp_text_out[3]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[40]$_DFF_P_.CLK__gold_cover (\__mp_text_out[40]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[40]$_DFF_P_.QN__gold_cover (\__mp_text_out[40]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[41]$_DFF_P_.CLK__gold_cover (\__mp_text_out[41]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[41]$_DFF_P_.QN__gold_cover (\__mp_text_out[41]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[42]$_DFF_P_.CLK__gold_cover (\__mp_text_out[42]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[42]$_DFF_P_.QN__gold_cover (\__mp_text_out[42]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[43]$_DFF_P_.CLK__gold_cover (\__mp_text_out[43]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[43]$_DFF_P_.QN__gold_cover (\__mp_text_out[43]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[44]$_DFF_P_.CLK__gold_cover (\__mp_text_out[44]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[44]$_DFF_P_.QN__gold_cover (\__mp_text_out[44]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[45]$_DFF_P_.CLK__gold_cover (\__mp_text_out[45]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[45]$_DFF_P_.QN__gold_cover (\__mp_text_out[45]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[46]$_DFF_P_.CLK__gold_cover (\__mp_text_out[46]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[46]$_DFF_P_.QN__gold_cover (\__mp_text_out[46]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[47]$_DFF_P_.CLK__gold_cover (\__mp_text_out[47]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[47]$_DFF_P_.QN__gold_cover (\__mp_text_out[47]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[48]$_DFF_P_.CLK__gold_cover (\__mp_text_out[48]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[48]$_DFF_P_.QN__gold_cover (\__mp_text_out[48]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[49]$_DFF_P_.CLK__gold_cover (\__mp_text_out[49]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[49]$_DFF_P_.QN__gold_cover (\__mp_text_out[49]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[4]$_DFF_P_.CLK__gold_cover (\__mp_text_out[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[4]$_DFF_P_.QN__gold_cover (\__mp_text_out[4]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[50]$_DFF_P_.CLK__gold_cover (\__mp_text_out[50]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[50]$_DFF_P_.QN__gold_cover (\__mp_text_out[50]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[51]$_DFF_P_.CLK__gold_cover (\__mp_text_out[51]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[51]$_DFF_P_.QN__gold_cover (\__mp_text_out[51]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[52]$_DFF_P_.CLK__gold_cover (\__mp_text_out[52]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[52]$_DFF_P_.QN__gold_cover (\__mp_text_out[52]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[53]$_DFF_P_.CLK__gold_cover (\__mp_text_out[53]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[53]$_DFF_P_.QN__gold_cover (\__mp_text_out[53]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[54]$_DFF_P_.CLK__gold_cover (\__mp_text_out[54]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[54]$_DFF_P_.QN__gold_cover (\__mp_text_out[54]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[55]$_DFF_P_.CLK__gold_cover (\__mp_text_out[55]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[55]$_DFF_P_.QN__gold_cover (\__mp_text_out[55]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[56]$_DFF_P_.CLK__gold_cover (\__mp_text_out[56]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[56]$_DFF_P_.QN__gold_cover (\__mp_text_out[56]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[57]$_DFF_P_.CLK__gold_cover (\__mp_text_out[57]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[57]$_DFF_P_.QN__gold_cover (\__mp_text_out[57]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[58]$_DFF_P_.CLK__gold_cover (\__mp_text_out[58]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[58]$_DFF_P_.QN__gold_cover (\__mp_text_out[58]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[59]$_DFF_P_.CLK__gold_cover (\__mp_text_out[59]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[59]$_DFF_P_.QN__gold_cover (\__mp_text_out[59]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[5]$_DFF_P_.CLK__gold_cover (\__mp_text_out[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[5]$_DFF_P_.QN__gold_cover (\__mp_text_out[5]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[60]$_DFF_P_.CLK__gold_cover (\__mp_text_out[60]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[60]$_DFF_P_.QN__gold_cover (\__mp_text_out[60]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[61]$_DFF_P_.CLK__gold_cover (\__mp_text_out[61]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[61]$_DFF_P_.QN__gold_cover (\__mp_text_out[61]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[62]$_DFF_P_.CLK__gold_cover (\__mp_text_out[62]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[62]$_DFF_P_.QN__gold_cover (\__mp_text_out[62]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[63]$_DFF_P_.CLK__gold_cover (\__mp_text_out[63]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[63]$_DFF_P_.QN__gold_cover (\__mp_text_out[63]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[64]$_DFF_P_.CLK__gold_cover (\__mp_text_out[64]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[64]$_DFF_P_.QN__gold_cover (\__mp_text_out[64]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[65]$_DFF_P_.CLK__gold_cover (\__mp_text_out[65]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[65]$_DFF_P_.QN__gold_cover (\__mp_text_out[65]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[66]$_DFF_P_.CLK__gold_cover (\__mp_text_out[66]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[66]$_DFF_P_.QN__gold_cover (\__mp_text_out[66]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[67]$_DFF_P_.CLK__gold_cover (\__mp_text_out[67]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[67]$_DFF_P_.QN__gold_cover (\__mp_text_out[67]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[68]$_DFF_P_.CLK__gold_cover (\__mp_text_out[68]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[68]$_DFF_P_.QN__gold_cover (\__mp_text_out[68]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[69]$_DFF_P_.CLK__gold_cover (\__mp_text_out[69]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[69]$_DFF_P_.QN__gold_cover (\__mp_text_out[69]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[6]$_DFF_P_.CLK__gold_cover (\__mp_text_out[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[6]$_DFF_P_.QN__gold_cover (\__mp_text_out[6]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[70]$_DFF_P_.CLK__gold_cover (\__mp_text_out[70]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[70]$_DFF_P_.QN__gold_cover (\__mp_text_out[70]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[71]$_DFF_P_.CLK__gold_cover (\__mp_text_out[71]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[71]$_DFF_P_.QN__gold_cover (\__mp_text_out[71]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[72]$_DFF_P_.CLK__gold_cover (\__mp_text_out[72]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[72]$_DFF_P_.QN__gold_cover (\__mp_text_out[72]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[73]$_DFF_P_.CLK__gold_cover (\__mp_text_out[73]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[73]$_DFF_P_.QN__gold_cover (\__mp_text_out[73]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[74]$_DFF_P_.CLK__gold_cover (\__mp_text_out[74]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[74]$_DFF_P_.QN__gold_cover (\__mp_text_out[74]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[75]$_DFF_P_.CLK__gold_cover (\__mp_text_out[75]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[75]$_DFF_P_.QN__gold_cover (\__mp_text_out[75]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[76]$_DFF_P_.CLK__gold_cover (\__mp_text_out[76]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[76]$_DFF_P_.QN__gold_cover (\__mp_text_out[76]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[77]$_DFF_P_.CLK__gold_cover (\__mp_text_out[77]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[77]$_DFF_P_.QN__gold_cover (\__mp_text_out[77]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[78]$_DFF_P_.CLK__gold_cover (\__mp_text_out[78]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[78]$_DFF_P_.QN__gold_cover (\__mp_text_out[78]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[79]$_DFF_P_.CLK__gold_cover (\__mp_text_out[79]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[79]$_DFF_P_.QN__gold_cover (\__mp_text_out[79]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[7]$_DFF_P_.CLK__gold_cover (\__mp_text_out[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[7]$_DFF_P_.QN__gold_cover (\__mp_text_out[7]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[80]$_DFF_P_.CLK__gold_cover (\__mp_text_out[80]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[80]$_DFF_P_.QN__gold_cover (\__mp_text_out[80]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[81]$_DFF_P_.CLK__gold_cover (\__mp_text_out[81]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[81]$_DFF_P_.QN__gold_cover (\__mp_text_out[81]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[82]$_DFF_P_.CLK__gold_cover (\__mp_text_out[82]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[82]$_DFF_P_.QN__gold_cover (\__mp_text_out[82]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[83]$_DFF_P_.CLK__gold_cover (\__mp_text_out[83]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[83]$_DFF_P_.QN__gold_cover (\__mp_text_out[83]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[84]$_DFF_P_.CLK__gold_cover (\__mp_text_out[84]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[84]$_DFF_P_.QN__gold_cover (\__mp_text_out[84]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[85]$_DFF_P_.CLK__gold_cover (\__mp_text_out[85]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[85]$_DFF_P_.QN__gold_cover (\__mp_text_out[85]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[86]$_DFF_P_.CLK__gold_cover (\__mp_text_out[86]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[86]$_DFF_P_.QN__gold_cover (\__mp_text_out[86]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[87]$_DFF_P_.CLK__gold_cover (\__mp_text_out[87]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[87]$_DFF_P_.QN__gold_cover (\__mp_text_out[87]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[88]$_DFF_P_.CLK__gold_cover (\__mp_text_out[88]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[88]$_DFF_P_.QN__gold_cover (\__mp_text_out[88]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[89]$_DFF_P_.CLK__gold_cover (\__mp_text_out[89]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[89]$_DFF_P_.QN__gold_cover (\__mp_text_out[89]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[8]$_DFF_P_.CLK__gold_cover (\__mp_text_out[8]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[8]$_DFF_P_.QN__gold_cover (\__mp_text_out[8]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[90]$_DFF_P_.CLK__gold_cover (\__mp_text_out[90]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[90]$_DFF_P_.QN__gold_cover (\__mp_text_out[90]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[91]$_DFF_P_.CLK__gold_cover (\__mp_text_out[91]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[91]$_DFF_P_.QN__gold_cover (\__mp_text_out[91]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[92]$_DFF_P_.CLK__gold_cover (\__mp_text_out[92]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[92]$_DFF_P_.QN__gold_cover (\__mp_text_out[92]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[93]$_DFF_P_.CLK__gold_cover (\__mp_text_out[93]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[93]$_DFF_P_.QN__gold_cover (\__mp_text_out[93]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[94]$_DFF_P_.CLK__gold_cover (\__mp_text_out[94]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[94]$_DFF_P_.QN__gold_cover (\__mp_text_out[94]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[95]$_DFF_P_.CLK__gold_cover (\__mp_text_out[95]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[95]$_DFF_P_.QN__gold_cover (\__mp_text_out[95]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[96]$_DFF_P_.CLK__gold_cover (\__mp_text_out[96]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[96]$_DFF_P_.QN__gold_cover (\__mp_text_out[96]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[97]$_DFF_P_.CLK__gold_cover (\__mp_text_out[97]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[97]$_DFF_P_.QN__gold_cover (\__mp_text_out[97]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[98]$_DFF_P_.CLK__gold_cover (\__mp_text_out[98]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[98]$_DFF_P_.QN__gold_cover (\__mp_text_out[98]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[99]$_DFF_P_.CLK__gold_cover (\__mp_text_out[99]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[99]$_DFF_P_.QN__gold_cover (\__mp_text_out[99]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[9]$_DFF_P_.CLK__gold_cover (\__mp_text_out[9]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[9]$_DFF_P_.QN__gold_cover (\__mp_text_out[9]$_DFF_P_.QN__gold );
  miter_def_prop #(1, "cover") \__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gold_cover (\__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gold_cover (\__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gold_cover (\__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[0]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[1]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[2]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[3]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[4]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[5]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[6]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[7]$_DFF_P_.CLK__gold_cover (\__mp_u0.u0.d[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[0]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[1]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[2]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[3]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[4]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[5]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[6]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[7]$_DFF_P_.CLK__gold_cover (\__mp_u0.u1.d[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[0]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[1]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[2]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[3]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[4]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[5]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[6]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[7]$_DFF_P_.CLK__gold_cover (\__mp_u0.u2.d[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[0]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[1]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[2]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[3]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[4]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[5]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[6]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[7]$_DFF_P_.CLK__gold_cover (\__mp_u0.u3.d[7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][0]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][10]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][10]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][11]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][11]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][12]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][12]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][13]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][13]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][14]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][14]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][15]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][15]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][16]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][16]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][17]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][17]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][18]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][18]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][19]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][19]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][1]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][20]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][20]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][21]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][21]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][22]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][22]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][23]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][23]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][24]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][24]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][25]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][25]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][26]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][26]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][27]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][27]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][28]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][28]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][29]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][29]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][2]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][30]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][30]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][31]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][31]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][3]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][4]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][5]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][6]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][7]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][8]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][8]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][9]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[0][9]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][0]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][10]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][10]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][11]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][11]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][12]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][12]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][13]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][13]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][14]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][14]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][15]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][15]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][16]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][16]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][17]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][17]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][18]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][18]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][19]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][19]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][1]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][20]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][20]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][21]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][21]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][22]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][22]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][23]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][23]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][24]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][24]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][25]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][25]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][26]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][26]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][27]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][27]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][28]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][28]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][29]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][29]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][2]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][30]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][30]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][31]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][31]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][3]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][4]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][5]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][6]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][7]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][8]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][8]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][9]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[1][9]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][0]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][10]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][10]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][11]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][11]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][12]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][12]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][13]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][13]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][14]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][14]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][15]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][15]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][16]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][16]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][17]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][17]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][18]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][18]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][19]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][19]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][1]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][20]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][20]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][21]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][21]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][22]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][22]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][23]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][23]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][24]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][24]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][25]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][25]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][26]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][26]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][27]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][27]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][28]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][28]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][29]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][29]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][2]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][30]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][30]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][31]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][31]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][3]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][4]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][5]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][6]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][7]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][8]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][8]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][9]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[2][9]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][0]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][0]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][10]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][10]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][11]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][11]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][12]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][12]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][13]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][13]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][14]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][14]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][15]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][15]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][16]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][16]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][17]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][17]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][18]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][18]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][19]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][19]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][1]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][1]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][20]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][20]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][21]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][21]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][22]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][22]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][23]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][23]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][24]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][24]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][25]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][25]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][26]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][26]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][27]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][27]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][28]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][28]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][29]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][29]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][2]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][2]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][30]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][30]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][31]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][31]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][3]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][3]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][4]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][4]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][5]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][5]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][6]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][6]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][7]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][7]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][8]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][8]$_DFF_P_.CLK__gold );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][9]$_DFF_P_.CLK__gold_cover (\__mp_u0.w[3][9]$_DFF_P_.CLK__gold );
`endif
`ifdef COVER_DEF_GATE_MATCH_POINTS
  miter_def_prop #(1, "cover") \__mp_clkbuf_0_clk.A__gate_cover (\__mp_clkbuf_0_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_0_clk.Y__gate_cover (\__mp_clkbuf_0_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_0_0_clk.A__gate_cover (\__mp_clkbuf_2_0_0_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_0_0_clk.Y__gate_cover (\__mp_clkbuf_2_0_0_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_1_0_clk.A__gate_cover (\__mp_clkbuf_2_1_0_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_1_0_clk.Y__gate_cover (\__mp_clkbuf_2_1_0_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_2_0_clk.A__gate_cover (\__mp_clkbuf_2_2_0_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_2_0_clk.Y__gate_cover (\__mp_clkbuf_2_2_0_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_3_0_clk.A__gate_cover (\__mp_clkbuf_2_3_0_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_2_3_0_clk.Y__gate_cover (\__mp_clkbuf_2_3_0_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_0_clk.A__gate_cover (\__mp_clkbuf_leaf_0_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_0_clk.Y__gate_cover (\__mp_clkbuf_leaf_0_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_10_clk.A__gate_cover (\__mp_clkbuf_leaf_10_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_10_clk.Y__gate_cover (\__mp_clkbuf_leaf_10_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_11_clk.A__gate_cover (\__mp_clkbuf_leaf_11_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_11_clk.Y__gate_cover (\__mp_clkbuf_leaf_11_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_12_clk.A__gate_cover (\__mp_clkbuf_leaf_12_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_12_clk.Y__gate_cover (\__mp_clkbuf_leaf_12_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_13_clk.A__gate_cover (\__mp_clkbuf_leaf_13_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_13_clk.Y__gate_cover (\__mp_clkbuf_leaf_13_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_14_clk.A__gate_cover (\__mp_clkbuf_leaf_14_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_14_clk.Y__gate_cover (\__mp_clkbuf_leaf_14_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_15_clk.A__gate_cover (\__mp_clkbuf_leaf_15_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_15_clk.Y__gate_cover (\__mp_clkbuf_leaf_15_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_16_clk.A__gate_cover (\__mp_clkbuf_leaf_16_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_16_clk.Y__gate_cover (\__mp_clkbuf_leaf_16_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_17_clk.A__gate_cover (\__mp_clkbuf_leaf_17_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_17_clk.Y__gate_cover (\__mp_clkbuf_leaf_17_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_18_clk.A__gate_cover (\__mp_clkbuf_leaf_18_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_18_clk.Y__gate_cover (\__mp_clkbuf_leaf_18_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_19_clk.A__gate_cover (\__mp_clkbuf_leaf_19_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_19_clk.Y__gate_cover (\__mp_clkbuf_leaf_19_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_1_clk.A__gate_cover (\__mp_clkbuf_leaf_1_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_1_clk.Y__gate_cover (\__mp_clkbuf_leaf_1_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_20_clk.A__gate_cover (\__mp_clkbuf_leaf_20_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_20_clk.Y__gate_cover (\__mp_clkbuf_leaf_20_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_21_clk.A__gate_cover (\__mp_clkbuf_leaf_21_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_21_clk.Y__gate_cover (\__mp_clkbuf_leaf_21_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_22_clk.A__gate_cover (\__mp_clkbuf_leaf_22_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_22_clk.Y__gate_cover (\__mp_clkbuf_leaf_22_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_23_clk.A__gate_cover (\__mp_clkbuf_leaf_23_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_23_clk.Y__gate_cover (\__mp_clkbuf_leaf_23_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_24_clk.A__gate_cover (\__mp_clkbuf_leaf_24_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_24_clk.Y__gate_cover (\__mp_clkbuf_leaf_24_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_25_clk.A__gate_cover (\__mp_clkbuf_leaf_25_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_25_clk.Y__gate_cover (\__mp_clkbuf_leaf_25_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_26_clk.A__gate_cover (\__mp_clkbuf_leaf_26_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_26_clk.Y__gate_cover (\__mp_clkbuf_leaf_26_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_27_clk.A__gate_cover (\__mp_clkbuf_leaf_27_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_27_clk.Y__gate_cover (\__mp_clkbuf_leaf_27_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_28_clk.A__gate_cover (\__mp_clkbuf_leaf_28_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_28_clk.Y__gate_cover (\__mp_clkbuf_leaf_28_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_29_clk.A__gate_cover (\__mp_clkbuf_leaf_29_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_29_clk.Y__gate_cover (\__mp_clkbuf_leaf_29_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_2_clk.A__gate_cover (\__mp_clkbuf_leaf_2_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_2_clk.Y__gate_cover (\__mp_clkbuf_leaf_2_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_30_clk.A__gate_cover (\__mp_clkbuf_leaf_30_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_30_clk.Y__gate_cover (\__mp_clkbuf_leaf_30_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_31_clk.A__gate_cover (\__mp_clkbuf_leaf_31_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_31_clk.Y__gate_cover (\__mp_clkbuf_leaf_31_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_32_clk.A__gate_cover (\__mp_clkbuf_leaf_32_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_32_clk.Y__gate_cover (\__mp_clkbuf_leaf_32_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_33_clk.A__gate_cover (\__mp_clkbuf_leaf_33_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_33_clk.Y__gate_cover (\__mp_clkbuf_leaf_33_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_3_clk.A__gate_cover (\__mp_clkbuf_leaf_3_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_3_clk.Y__gate_cover (\__mp_clkbuf_leaf_3_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_4_clk.A__gate_cover (\__mp_clkbuf_leaf_4_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_4_clk.Y__gate_cover (\__mp_clkbuf_leaf_4_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_5_clk.A__gate_cover (\__mp_clkbuf_leaf_5_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_5_clk.Y__gate_cover (\__mp_clkbuf_leaf_5_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_6_clk.A__gate_cover (\__mp_clkbuf_leaf_6_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_6_clk.Y__gate_cover (\__mp_clkbuf_leaf_6_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_7_clk.A__gate_cover (\__mp_clkbuf_leaf_7_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_7_clk.Y__gate_cover (\__mp_clkbuf_leaf_7_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_8_clk.A__gate_cover (\__mp_clkbuf_leaf_8_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_8_clk.Y__gate_cover (\__mp_clkbuf_leaf_8_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_9_clk.A__gate_cover (\__mp_clkbuf_leaf_9_clk.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkbuf_leaf_9_clk.Y__gate_cover (\__mp_clkbuf_leaf_9_clk.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkload0.A__gate_cover (\__mp_clkload0.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload0.Y__gate_cover (\__mp_clkload0.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkload1.A__gate_cover (\__mp_clkload1.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload10.A__gate_cover (\__mp_clkload10.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload11.A__gate_cover (\__mp_clkload11.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload12.A__gate_cover (\__mp_clkload12.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload13.A__gate_cover (\__mp_clkload13.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload14.A__gate_cover (\__mp_clkload14.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload15.A__gate_cover (\__mp_clkload15.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload16.A__gate_cover (\__mp_clkload16.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload17.A__gate_cover (\__mp_clkload17.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload18.A__gate_cover (\__mp_clkload18.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload18.Y__gate_cover (\__mp_clkload18.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkload19.A__gate_cover (\__mp_clkload19.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload2.A__gate_cover (\__mp_clkload2.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload20.A__gate_cover (\__mp_clkload20.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload21.A__gate_cover (\__mp_clkload21.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload22.A__gate_cover (\__mp_clkload22.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload23.A__gate_cover (\__mp_clkload23.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload24.A__gate_cover (\__mp_clkload24.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload25.A__gate_cover (\__mp_clkload25.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload26.A__gate_cover (\__mp_clkload26.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload27.A__gate_cover (\__mp_clkload27.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload28.A__gate_cover (\__mp_clkload28.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload29.A__gate_cover (\__mp_clkload29.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload3.A__gate_cover (\__mp_clkload3.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload30.A__gate_cover (\__mp_clkload30.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload31.A__gate_cover (\__mp_clkload31.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload31.Y__gate_cover (\__mp_clkload31.Y__gate );
  miter_def_prop #(1, "cover") \__mp_clkload32.A__gate_cover (\__mp_clkload32.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload4.A__gate_cover (\__mp_clkload4.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload5.A__gate_cover (\__mp_clkload5.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload6.A__gate_cover (\__mp_clkload6.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload7.A__gate_cover (\__mp_clkload7.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload8.A__gate_cover (\__mp_clkload8.A__gate );
  miter_def_prop #(1, "cover") \__mp_clkload9.A__gate_cover (\__mp_clkload9.A__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_0_clk__gate_cover (\__mp_clknet_0_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_2_0_0_clk__gate_cover (\__mp_clknet_2_0_0_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_2_1_0_clk__gate_cover (\__mp_clknet_2_1_0_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_2_2_0_clk__gate_cover (\__mp_clknet_2_2_0_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_2_3_0_clk__gate_cover (\__mp_clknet_2_3_0_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_0_clk__gate_cover (\__mp_clknet_leaf_0_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_10_clk__gate_cover (\__mp_clknet_leaf_10_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_11_clk__gate_cover (\__mp_clknet_leaf_11_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_12_clk__gate_cover (\__mp_clknet_leaf_12_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_13_clk__gate_cover (\__mp_clknet_leaf_13_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_14_clk__gate_cover (\__mp_clknet_leaf_14_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_15_clk__gate_cover (\__mp_clknet_leaf_15_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_16_clk__gate_cover (\__mp_clknet_leaf_16_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_17_clk__gate_cover (\__mp_clknet_leaf_17_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_18_clk__gate_cover (\__mp_clknet_leaf_18_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_19_clk__gate_cover (\__mp_clknet_leaf_19_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_1_clk__gate_cover (\__mp_clknet_leaf_1_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_20_clk__gate_cover (\__mp_clknet_leaf_20_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_21_clk__gate_cover (\__mp_clknet_leaf_21_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_22_clk__gate_cover (\__mp_clknet_leaf_22_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_23_clk__gate_cover (\__mp_clknet_leaf_23_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_24_clk__gate_cover (\__mp_clknet_leaf_24_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_25_clk__gate_cover (\__mp_clknet_leaf_25_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_26_clk__gate_cover (\__mp_clknet_leaf_26_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_27_clk__gate_cover (\__mp_clknet_leaf_27_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_28_clk__gate_cover (\__mp_clknet_leaf_28_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_29_clk__gate_cover (\__mp_clknet_leaf_29_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_2_clk__gate_cover (\__mp_clknet_leaf_2_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_30_clk__gate_cover (\__mp_clknet_leaf_30_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_31_clk__gate_cover (\__mp_clknet_leaf_31_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_32_clk__gate_cover (\__mp_clknet_leaf_32_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_33_clk__gate_cover (\__mp_clknet_leaf_33_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_3_clk__gate_cover (\__mp_clknet_leaf_3_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_4_clk__gate_cover (\__mp_clknet_leaf_4_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_5_clk__gate_cover (\__mp_clknet_leaf_5_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_6_clk__gate_cover (\__mp_clknet_leaf_6_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_7_clk__gate_cover (\__mp_clknet_leaf_7_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_8_clk__gate_cover (\__mp_clknet_leaf_8_clk__gate );
  miter_def_prop #(1, "cover") \__mp_clknet_leaf_9_clk__gate_cover (\__mp_clknet_leaf_9_clk__gate );
  miter_def_prop #(1, "cover") \__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gate_cover (\__mp_dcnt[0]$_SDFFE_PN0P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gate_cover (\__mp_dcnt[1]$_SDFFE_PN0P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gate_cover (\__mp_dcnt[2]$_SDFFE_PP0P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gate_cover (\__mp_dcnt[3]$_SDFFE_PN0P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_done$_DFF_P_.CLK__gate_cover (\__mp_done$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_done$_DFF_P_.QN__gate_cover (\__mp_done$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_done$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_done$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_input1.A__gate_cover (\__mp_input1.A__gate );
  miter_def_prop #(1, "cover") \__mp_input1.Y__gate_cover (\__mp_input1.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input10.A__gate_cover (\__mp_input10.A__gate );
  miter_def_prop #(1, "cover") \__mp_input10.Y__gate_cover (\__mp_input10.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input100.A__gate_cover (\__mp_input100.A__gate );
  miter_def_prop #(1, "cover") \__mp_input100.Y__gate_cover (\__mp_input100.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input101.A__gate_cover (\__mp_input101.A__gate );
  miter_def_prop #(1, "cover") \__mp_input101.Y__gate_cover (\__mp_input101.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input102.A__gate_cover (\__mp_input102.A__gate );
  miter_def_prop #(1, "cover") \__mp_input102.Y__gate_cover (\__mp_input102.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input103.A__gate_cover (\__mp_input103.A__gate );
  miter_def_prop #(1, "cover") \__mp_input103.Y__gate_cover (\__mp_input103.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input104.A__gate_cover (\__mp_input104.A__gate );
  miter_def_prop #(1, "cover") \__mp_input104.Y__gate_cover (\__mp_input104.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input105.A__gate_cover (\__mp_input105.A__gate );
  miter_def_prop #(1, "cover") \__mp_input105.Y__gate_cover (\__mp_input105.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input106.A__gate_cover (\__mp_input106.A__gate );
  miter_def_prop #(1, "cover") \__mp_input106.Y__gate_cover (\__mp_input106.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input107.A__gate_cover (\__mp_input107.A__gate );
  miter_def_prop #(1, "cover") \__mp_input107.Y__gate_cover (\__mp_input107.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input108.A__gate_cover (\__mp_input108.A__gate );
  miter_def_prop #(1, "cover") \__mp_input108.Y__gate_cover (\__mp_input108.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input109.A__gate_cover (\__mp_input109.A__gate );
  miter_def_prop #(1, "cover") \__mp_input109.Y__gate_cover (\__mp_input109.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input11.A__gate_cover (\__mp_input11.A__gate );
  miter_def_prop #(1, "cover") \__mp_input11.Y__gate_cover (\__mp_input11.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input110.A__gate_cover (\__mp_input110.A__gate );
  miter_def_prop #(1, "cover") \__mp_input110.Y__gate_cover (\__mp_input110.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input111.A__gate_cover (\__mp_input111.A__gate );
  miter_def_prop #(1, "cover") \__mp_input111.Y__gate_cover (\__mp_input111.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input112.A__gate_cover (\__mp_input112.A__gate );
  miter_def_prop #(1, "cover") \__mp_input112.Y__gate_cover (\__mp_input112.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input113.A__gate_cover (\__mp_input113.A__gate );
  miter_def_prop #(1, "cover") \__mp_input113.Y__gate_cover (\__mp_input113.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input114.A__gate_cover (\__mp_input114.A__gate );
  miter_def_prop #(1, "cover") \__mp_input114.Y__gate_cover (\__mp_input114.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input115.A__gate_cover (\__mp_input115.A__gate );
  miter_def_prop #(1, "cover") \__mp_input115.Y__gate_cover (\__mp_input115.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input116.A__gate_cover (\__mp_input116.A__gate );
  miter_def_prop #(1, "cover") \__mp_input116.Y__gate_cover (\__mp_input116.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input117.A__gate_cover (\__mp_input117.A__gate );
  miter_def_prop #(1, "cover") \__mp_input117.Y__gate_cover (\__mp_input117.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input118.A__gate_cover (\__mp_input118.A__gate );
  miter_def_prop #(1, "cover") \__mp_input118.Y__gate_cover (\__mp_input118.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input119.A__gate_cover (\__mp_input119.A__gate );
  miter_def_prop #(1, "cover") \__mp_input119.Y__gate_cover (\__mp_input119.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input12.A__gate_cover (\__mp_input12.A__gate );
  miter_def_prop #(1, "cover") \__mp_input12.Y__gate_cover (\__mp_input12.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input120.A__gate_cover (\__mp_input120.A__gate );
  miter_def_prop #(1, "cover") \__mp_input120.Y__gate_cover (\__mp_input120.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input121.A__gate_cover (\__mp_input121.A__gate );
  miter_def_prop #(1, "cover") \__mp_input121.Y__gate_cover (\__mp_input121.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input122.A__gate_cover (\__mp_input122.A__gate );
  miter_def_prop #(1, "cover") \__mp_input122.Y__gate_cover (\__mp_input122.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input123.A__gate_cover (\__mp_input123.A__gate );
  miter_def_prop #(1, "cover") \__mp_input123.Y__gate_cover (\__mp_input123.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input124.A__gate_cover (\__mp_input124.A__gate );
  miter_def_prop #(1, "cover") \__mp_input124.Y__gate_cover (\__mp_input124.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input125.A__gate_cover (\__mp_input125.A__gate );
  miter_def_prop #(1, "cover") \__mp_input125.Y__gate_cover (\__mp_input125.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input126.A__gate_cover (\__mp_input126.A__gate );
  miter_def_prop #(1, "cover") \__mp_input126.Y__gate_cover (\__mp_input126.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input127.A__gate_cover (\__mp_input127.A__gate );
  miter_def_prop #(1, "cover") \__mp_input127.Y__gate_cover (\__mp_input127.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input128.A__gate_cover (\__mp_input128.A__gate );
  miter_def_prop #(1, "cover") \__mp_input128.Y__gate_cover (\__mp_input128.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input129.A__gate_cover (\__mp_input129.A__gate );
  miter_def_prop #(1, "cover") \__mp_input129.Y__gate_cover (\__mp_input129.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input13.A__gate_cover (\__mp_input13.A__gate );
  miter_def_prop #(1, "cover") \__mp_input13.Y__gate_cover (\__mp_input13.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input130.A__gate_cover (\__mp_input130.A__gate );
  miter_def_prop #(1, "cover") \__mp_input130.Y__gate_cover (\__mp_input130.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input131.A__gate_cover (\__mp_input131.A__gate );
  miter_def_prop #(1, "cover") \__mp_input131.Y__gate_cover (\__mp_input131.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input132.A__gate_cover (\__mp_input132.A__gate );
  miter_def_prop #(1, "cover") \__mp_input132.Y__gate_cover (\__mp_input132.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input133.A__gate_cover (\__mp_input133.A__gate );
  miter_def_prop #(1, "cover") \__mp_input133.Y__gate_cover (\__mp_input133.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input134.A__gate_cover (\__mp_input134.A__gate );
  miter_def_prop #(1, "cover") \__mp_input134.Y__gate_cover (\__mp_input134.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input135.A__gate_cover (\__mp_input135.A__gate );
  miter_def_prop #(1, "cover") \__mp_input135.Y__gate_cover (\__mp_input135.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input136.A__gate_cover (\__mp_input136.A__gate );
  miter_def_prop #(1, "cover") \__mp_input136.Y__gate_cover (\__mp_input136.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input137.A__gate_cover (\__mp_input137.A__gate );
  miter_def_prop #(1, "cover") \__mp_input137.Y__gate_cover (\__mp_input137.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input138.A__gate_cover (\__mp_input138.A__gate );
  miter_def_prop #(1, "cover") \__mp_input138.Y__gate_cover (\__mp_input138.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input139.A__gate_cover (\__mp_input139.A__gate );
  miter_def_prop #(1, "cover") \__mp_input139.Y__gate_cover (\__mp_input139.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input14.A__gate_cover (\__mp_input14.A__gate );
  miter_def_prop #(1, "cover") \__mp_input14.Y__gate_cover (\__mp_input14.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input140.A__gate_cover (\__mp_input140.A__gate );
  miter_def_prop #(1, "cover") \__mp_input140.Y__gate_cover (\__mp_input140.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input141.A__gate_cover (\__mp_input141.A__gate );
  miter_def_prop #(1, "cover") \__mp_input141.Y__gate_cover (\__mp_input141.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input142.A__gate_cover (\__mp_input142.A__gate );
  miter_def_prop #(1, "cover") \__mp_input142.Y__gate_cover (\__mp_input142.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input143.A__gate_cover (\__mp_input143.A__gate );
  miter_def_prop #(1, "cover") \__mp_input143.Y__gate_cover (\__mp_input143.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input144.A__gate_cover (\__mp_input144.A__gate );
  miter_def_prop #(1, "cover") \__mp_input144.Y__gate_cover (\__mp_input144.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input145.A__gate_cover (\__mp_input145.A__gate );
  miter_def_prop #(1, "cover") \__mp_input145.Y__gate_cover (\__mp_input145.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input146.A__gate_cover (\__mp_input146.A__gate );
  miter_def_prop #(1, "cover") \__mp_input146.Y__gate_cover (\__mp_input146.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input147.A__gate_cover (\__mp_input147.A__gate );
  miter_def_prop #(1, "cover") \__mp_input147.Y__gate_cover (\__mp_input147.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input148.A__gate_cover (\__mp_input148.A__gate );
  miter_def_prop #(1, "cover") \__mp_input148.Y__gate_cover (\__mp_input148.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input149.A__gate_cover (\__mp_input149.A__gate );
  miter_def_prop #(1, "cover") \__mp_input149.Y__gate_cover (\__mp_input149.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input15.A__gate_cover (\__mp_input15.A__gate );
  miter_def_prop #(1, "cover") \__mp_input15.Y__gate_cover (\__mp_input15.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input150.A__gate_cover (\__mp_input150.A__gate );
  miter_def_prop #(1, "cover") \__mp_input150.Y__gate_cover (\__mp_input150.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input151.A__gate_cover (\__mp_input151.A__gate );
  miter_def_prop #(1, "cover") \__mp_input151.Y__gate_cover (\__mp_input151.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input152.A__gate_cover (\__mp_input152.A__gate );
  miter_def_prop #(1, "cover") \__mp_input152.Y__gate_cover (\__mp_input152.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input153.A__gate_cover (\__mp_input153.A__gate );
  miter_def_prop #(1, "cover") \__mp_input153.Y__gate_cover (\__mp_input153.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input154.A__gate_cover (\__mp_input154.A__gate );
  miter_def_prop #(1, "cover") \__mp_input154.Y__gate_cover (\__mp_input154.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input155.A__gate_cover (\__mp_input155.A__gate );
  miter_def_prop #(1, "cover") \__mp_input155.Y__gate_cover (\__mp_input155.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input156.A__gate_cover (\__mp_input156.A__gate );
  miter_def_prop #(1, "cover") \__mp_input156.Y__gate_cover (\__mp_input156.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input157.A__gate_cover (\__mp_input157.A__gate );
  miter_def_prop #(1, "cover") \__mp_input157.Y__gate_cover (\__mp_input157.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input158.A__gate_cover (\__mp_input158.A__gate );
  miter_def_prop #(1, "cover") \__mp_input158.Y__gate_cover (\__mp_input158.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input159.A__gate_cover (\__mp_input159.A__gate );
  miter_def_prop #(1, "cover") \__mp_input159.Y__gate_cover (\__mp_input159.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input16.A__gate_cover (\__mp_input16.A__gate );
  miter_def_prop #(1, "cover") \__mp_input16.Y__gate_cover (\__mp_input16.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input160.A__gate_cover (\__mp_input160.A__gate );
  miter_def_prop #(1, "cover") \__mp_input160.Y__gate_cover (\__mp_input160.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input161.A__gate_cover (\__mp_input161.A__gate );
  miter_def_prop #(1, "cover") \__mp_input161.Y__gate_cover (\__mp_input161.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input162.A__gate_cover (\__mp_input162.A__gate );
  miter_def_prop #(1, "cover") \__mp_input162.Y__gate_cover (\__mp_input162.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input163.A__gate_cover (\__mp_input163.A__gate );
  miter_def_prop #(1, "cover") \__mp_input163.Y__gate_cover (\__mp_input163.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input164.A__gate_cover (\__mp_input164.A__gate );
  miter_def_prop #(1, "cover") \__mp_input164.Y__gate_cover (\__mp_input164.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input165.A__gate_cover (\__mp_input165.A__gate );
  miter_def_prop #(1, "cover") \__mp_input165.Y__gate_cover (\__mp_input165.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input166.A__gate_cover (\__mp_input166.A__gate );
  miter_def_prop #(1, "cover") \__mp_input166.Y__gate_cover (\__mp_input166.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input167.A__gate_cover (\__mp_input167.A__gate );
  miter_def_prop #(1, "cover") \__mp_input167.Y__gate_cover (\__mp_input167.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input168.A__gate_cover (\__mp_input168.A__gate );
  miter_def_prop #(1, "cover") \__mp_input168.Y__gate_cover (\__mp_input168.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input169.A__gate_cover (\__mp_input169.A__gate );
  miter_def_prop #(1, "cover") \__mp_input169.Y__gate_cover (\__mp_input169.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input17.A__gate_cover (\__mp_input17.A__gate );
  miter_def_prop #(1, "cover") \__mp_input17.Y__gate_cover (\__mp_input17.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input170.A__gate_cover (\__mp_input170.A__gate );
  miter_def_prop #(1, "cover") \__mp_input170.Y__gate_cover (\__mp_input170.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input171.A__gate_cover (\__mp_input171.A__gate );
  miter_def_prop #(1, "cover") \__mp_input171.Y__gate_cover (\__mp_input171.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input172.A__gate_cover (\__mp_input172.A__gate );
  miter_def_prop #(1, "cover") \__mp_input172.Y__gate_cover (\__mp_input172.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input173.A__gate_cover (\__mp_input173.A__gate );
  miter_def_prop #(1, "cover") \__mp_input173.Y__gate_cover (\__mp_input173.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input174.A__gate_cover (\__mp_input174.A__gate );
  miter_def_prop #(1, "cover") \__mp_input174.Y__gate_cover (\__mp_input174.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input175.A__gate_cover (\__mp_input175.A__gate );
  miter_def_prop #(1, "cover") \__mp_input175.Y__gate_cover (\__mp_input175.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input176.A__gate_cover (\__mp_input176.A__gate );
  miter_def_prop #(1, "cover") \__mp_input176.Y__gate_cover (\__mp_input176.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input177.A__gate_cover (\__mp_input177.A__gate );
  miter_def_prop #(1, "cover") \__mp_input177.Y__gate_cover (\__mp_input177.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input178.A__gate_cover (\__mp_input178.A__gate );
  miter_def_prop #(1, "cover") \__mp_input178.Y__gate_cover (\__mp_input178.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input179.A__gate_cover (\__mp_input179.A__gate );
  miter_def_prop #(1, "cover") \__mp_input179.Y__gate_cover (\__mp_input179.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input18.A__gate_cover (\__mp_input18.A__gate );
  miter_def_prop #(1, "cover") \__mp_input18.Y__gate_cover (\__mp_input18.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input180.A__gate_cover (\__mp_input180.A__gate );
  miter_def_prop #(1, "cover") \__mp_input180.Y__gate_cover (\__mp_input180.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input181.A__gate_cover (\__mp_input181.A__gate );
  miter_def_prop #(1, "cover") \__mp_input181.Y__gate_cover (\__mp_input181.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input182.A__gate_cover (\__mp_input182.A__gate );
  miter_def_prop #(1, "cover") \__mp_input182.Y__gate_cover (\__mp_input182.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input183.A__gate_cover (\__mp_input183.A__gate );
  miter_def_prop #(1, "cover") \__mp_input183.Y__gate_cover (\__mp_input183.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input184.A__gate_cover (\__mp_input184.A__gate );
  miter_def_prop #(1, "cover") \__mp_input184.Y__gate_cover (\__mp_input184.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input185.A__gate_cover (\__mp_input185.A__gate );
  miter_def_prop #(1, "cover") \__mp_input185.Y__gate_cover (\__mp_input185.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input186.A__gate_cover (\__mp_input186.A__gate );
  miter_def_prop #(1, "cover") \__mp_input186.Y__gate_cover (\__mp_input186.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input187.A__gate_cover (\__mp_input187.A__gate );
  miter_def_prop #(1, "cover") \__mp_input187.Y__gate_cover (\__mp_input187.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input188.A__gate_cover (\__mp_input188.A__gate );
  miter_def_prop #(1, "cover") \__mp_input188.Y__gate_cover (\__mp_input188.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input189.A__gate_cover (\__mp_input189.A__gate );
  miter_def_prop #(1, "cover") \__mp_input189.Y__gate_cover (\__mp_input189.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input19.A__gate_cover (\__mp_input19.A__gate );
  miter_def_prop #(1, "cover") \__mp_input19.Y__gate_cover (\__mp_input19.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input190.A__gate_cover (\__mp_input190.A__gate );
  miter_def_prop #(1, "cover") \__mp_input190.Y__gate_cover (\__mp_input190.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input191.A__gate_cover (\__mp_input191.A__gate );
  miter_def_prop #(1, "cover") \__mp_input191.Y__gate_cover (\__mp_input191.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input192.A__gate_cover (\__mp_input192.A__gate );
  miter_def_prop #(1, "cover") \__mp_input192.Y__gate_cover (\__mp_input192.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input193.A__gate_cover (\__mp_input193.A__gate );
  miter_def_prop #(1, "cover") \__mp_input193.Y__gate_cover (\__mp_input193.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input194.A__gate_cover (\__mp_input194.A__gate );
  miter_def_prop #(1, "cover") \__mp_input194.Y__gate_cover (\__mp_input194.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input195.A__gate_cover (\__mp_input195.A__gate );
  miter_def_prop #(1, "cover") \__mp_input195.Y__gate_cover (\__mp_input195.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input196.A__gate_cover (\__mp_input196.A__gate );
  miter_def_prop #(1, "cover") \__mp_input196.Y__gate_cover (\__mp_input196.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input197.A__gate_cover (\__mp_input197.A__gate );
  miter_def_prop #(1, "cover") \__mp_input197.Y__gate_cover (\__mp_input197.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input198.A__gate_cover (\__mp_input198.A__gate );
  miter_def_prop #(1, "cover") \__mp_input198.Y__gate_cover (\__mp_input198.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input199.A__gate_cover (\__mp_input199.A__gate );
  miter_def_prop #(1, "cover") \__mp_input199.Y__gate_cover (\__mp_input199.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input2.A__gate_cover (\__mp_input2.A__gate );
  miter_def_prop #(1, "cover") \__mp_input2.Y__gate_cover (\__mp_input2.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input20.A__gate_cover (\__mp_input20.A__gate );
  miter_def_prop #(1, "cover") \__mp_input20.Y__gate_cover (\__mp_input20.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input200.A__gate_cover (\__mp_input200.A__gate );
  miter_def_prop #(1, "cover") \__mp_input200.Y__gate_cover (\__mp_input200.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input201.A__gate_cover (\__mp_input201.A__gate );
  miter_def_prop #(1, "cover") \__mp_input201.Y__gate_cover (\__mp_input201.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input202.A__gate_cover (\__mp_input202.A__gate );
  miter_def_prop #(1, "cover") \__mp_input202.Y__gate_cover (\__mp_input202.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input203.A__gate_cover (\__mp_input203.A__gate );
  miter_def_prop #(1, "cover") \__mp_input203.Y__gate_cover (\__mp_input203.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input204.A__gate_cover (\__mp_input204.A__gate );
  miter_def_prop #(1, "cover") \__mp_input204.Y__gate_cover (\__mp_input204.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input205.A__gate_cover (\__mp_input205.A__gate );
  miter_def_prop #(1, "cover") \__mp_input205.Y__gate_cover (\__mp_input205.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input206.A__gate_cover (\__mp_input206.A__gate );
  miter_def_prop #(1, "cover") \__mp_input206.Y__gate_cover (\__mp_input206.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input207.A__gate_cover (\__mp_input207.A__gate );
  miter_def_prop #(1, "cover") \__mp_input207.Y__gate_cover (\__mp_input207.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input208.A__gate_cover (\__mp_input208.A__gate );
  miter_def_prop #(1, "cover") \__mp_input208.Y__gate_cover (\__mp_input208.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input209.A__gate_cover (\__mp_input209.A__gate );
  miter_def_prop #(1, "cover") \__mp_input209.Y__gate_cover (\__mp_input209.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input21.A__gate_cover (\__mp_input21.A__gate );
  miter_def_prop #(1, "cover") \__mp_input21.Y__gate_cover (\__mp_input21.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input210.A__gate_cover (\__mp_input210.A__gate );
  miter_def_prop #(1, "cover") \__mp_input210.Y__gate_cover (\__mp_input210.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input211.A__gate_cover (\__mp_input211.A__gate );
  miter_def_prop #(1, "cover") \__mp_input211.Y__gate_cover (\__mp_input211.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input212.A__gate_cover (\__mp_input212.A__gate );
  miter_def_prop #(1, "cover") \__mp_input212.Y__gate_cover (\__mp_input212.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input213.A__gate_cover (\__mp_input213.A__gate );
  miter_def_prop #(1, "cover") \__mp_input213.Y__gate_cover (\__mp_input213.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input214.A__gate_cover (\__mp_input214.A__gate );
  miter_def_prop #(1, "cover") \__mp_input214.Y__gate_cover (\__mp_input214.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input215.A__gate_cover (\__mp_input215.A__gate );
  miter_def_prop #(1, "cover") \__mp_input215.Y__gate_cover (\__mp_input215.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input216.A__gate_cover (\__mp_input216.A__gate );
  miter_def_prop #(1, "cover") \__mp_input216.Y__gate_cover (\__mp_input216.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input217.A__gate_cover (\__mp_input217.A__gate );
  miter_def_prop #(1, "cover") \__mp_input217.Y__gate_cover (\__mp_input217.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input218.A__gate_cover (\__mp_input218.A__gate );
  miter_def_prop #(1, "cover") \__mp_input218.Y__gate_cover (\__mp_input218.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input219.A__gate_cover (\__mp_input219.A__gate );
  miter_def_prop #(1, "cover") \__mp_input219.Y__gate_cover (\__mp_input219.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input22.A__gate_cover (\__mp_input22.A__gate );
  miter_def_prop #(1, "cover") \__mp_input22.Y__gate_cover (\__mp_input22.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input220.A__gate_cover (\__mp_input220.A__gate );
  miter_def_prop #(1, "cover") \__mp_input220.Y__gate_cover (\__mp_input220.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input221.A__gate_cover (\__mp_input221.A__gate );
  miter_def_prop #(1, "cover") \__mp_input221.Y__gate_cover (\__mp_input221.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input222.A__gate_cover (\__mp_input222.A__gate );
  miter_def_prop #(1, "cover") \__mp_input222.Y__gate_cover (\__mp_input222.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input223.A__gate_cover (\__mp_input223.A__gate );
  miter_def_prop #(1, "cover") \__mp_input223.Y__gate_cover (\__mp_input223.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input224.A__gate_cover (\__mp_input224.A__gate );
  miter_def_prop #(1, "cover") \__mp_input224.Y__gate_cover (\__mp_input224.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input225.A__gate_cover (\__mp_input225.A__gate );
  miter_def_prop #(1, "cover") \__mp_input225.Y__gate_cover (\__mp_input225.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input226.A__gate_cover (\__mp_input226.A__gate );
  miter_def_prop #(1, "cover") \__mp_input226.Y__gate_cover (\__mp_input226.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input227.A__gate_cover (\__mp_input227.A__gate );
  miter_def_prop #(1, "cover") \__mp_input227.Y__gate_cover (\__mp_input227.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input228.A__gate_cover (\__mp_input228.A__gate );
  miter_def_prop #(1, "cover") \__mp_input228.Y__gate_cover (\__mp_input228.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input229.A__gate_cover (\__mp_input229.A__gate );
  miter_def_prop #(1, "cover") \__mp_input229.Y__gate_cover (\__mp_input229.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input23.A__gate_cover (\__mp_input23.A__gate );
  miter_def_prop #(1, "cover") \__mp_input23.Y__gate_cover (\__mp_input23.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input230.A__gate_cover (\__mp_input230.A__gate );
  miter_def_prop #(1, "cover") \__mp_input230.Y__gate_cover (\__mp_input230.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input231.A__gate_cover (\__mp_input231.A__gate );
  miter_def_prop #(1, "cover") \__mp_input231.Y__gate_cover (\__mp_input231.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input232.A__gate_cover (\__mp_input232.A__gate );
  miter_def_prop #(1, "cover") \__mp_input232.Y__gate_cover (\__mp_input232.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input233.A__gate_cover (\__mp_input233.A__gate );
  miter_def_prop #(1, "cover") \__mp_input233.Y__gate_cover (\__mp_input233.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input234.A__gate_cover (\__mp_input234.A__gate );
  miter_def_prop #(1, "cover") \__mp_input234.Y__gate_cover (\__mp_input234.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input235.A__gate_cover (\__mp_input235.A__gate );
  miter_def_prop #(1, "cover") \__mp_input235.Y__gate_cover (\__mp_input235.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input236.A__gate_cover (\__mp_input236.A__gate );
  miter_def_prop #(1, "cover") \__mp_input236.Y__gate_cover (\__mp_input236.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input237.A__gate_cover (\__mp_input237.A__gate );
  miter_def_prop #(1, "cover") \__mp_input237.Y__gate_cover (\__mp_input237.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input238.A__gate_cover (\__mp_input238.A__gate );
  miter_def_prop #(1, "cover") \__mp_input238.Y__gate_cover (\__mp_input238.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input239.A__gate_cover (\__mp_input239.A__gate );
  miter_def_prop #(1, "cover") \__mp_input239.Y__gate_cover (\__mp_input239.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input24.A__gate_cover (\__mp_input24.A__gate );
  miter_def_prop #(1, "cover") \__mp_input24.Y__gate_cover (\__mp_input24.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input240.A__gate_cover (\__mp_input240.A__gate );
  miter_def_prop #(1, "cover") \__mp_input240.Y__gate_cover (\__mp_input240.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input241.A__gate_cover (\__mp_input241.A__gate );
  miter_def_prop #(1, "cover") \__mp_input241.Y__gate_cover (\__mp_input241.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input242.A__gate_cover (\__mp_input242.A__gate );
  miter_def_prop #(1, "cover") \__mp_input242.Y__gate_cover (\__mp_input242.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input243.A__gate_cover (\__mp_input243.A__gate );
  miter_def_prop #(1, "cover") \__mp_input243.Y__gate_cover (\__mp_input243.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input244.A__gate_cover (\__mp_input244.A__gate );
  miter_def_prop #(1, "cover") \__mp_input244.Y__gate_cover (\__mp_input244.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input245.A__gate_cover (\__mp_input245.A__gate );
  miter_def_prop #(1, "cover") \__mp_input245.Y__gate_cover (\__mp_input245.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input246.A__gate_cover (\__mp_input246.A__gate );
  miter_def_prop #(1, "cover") \__mp_input246.Y__gate_cover (\__mp_input246.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input247.A__gate_cover (\__mp_input247.A__gate );
  miter_def_prop #(1, "cover") \__mp_input247.Y__gate_cover (\__mp_input247.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input248.A__gate_cover (\__mp_input248.A__gate );
  miter_def_prop #(1, "cover") \__mp_input248.Y__gate_cover (\__mp_input248.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input249.A__gate_cover (\__mp_input249.A__gate );
  miter_def_prop #(1, "cover") \__mp_input249.Y__gate_cover (\__mp_input249.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input25.A__gate_cover (\__mp_input25.A__gate );
  miter_def_prop #(1, "cover") \__mp_input25.Y__gate_cover (\__mp_input25.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input250.A__gate_cover (\__mp_input250.A__gate );
  miter_def_prop #(1, "cover") \__mp_input250.Y__gate_cover (\__mp_input250.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input251.A__gate_cover (\__mp_input251.A__gate );
  miter_def_prop #(1, "cover") \__mp_input251.Y__gate_cover (\__mp_input251.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input252.A__gate_cover (\__mp_input252.A__gate );
  miter_def_prop #(1, "cover") \__mp_input252.Y__gate_cover (\__mp_input252.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input253.A__gate_cover (\__mp_input253.A__gate );
  miter_def_prop #(1, "cover") \__mp_input253.Y__gate_cover (\__mp_input253.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input254.A__gate_cover (\__mp_input254.A__gate );
  miter_def_prop #(1, "cover") \__mp_input254.Y__gate_cover (\__mp_input254.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input255.A__gate_cover (\__mp_input255.A__gate );
  miter_def_prop #(1, "cover") \__mp_input255.Y__gate_cover (\__mp_input255.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input256.A__gate_cover (\__mp_input256.A__gate );
  miter_def_prop #(1, "cover") \__mp_input256.Y__gate_cover (\__mp_input256.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input257.A__gate_cover (\__mp_input257.A__gate );
  miter_def_prop #(1, "cover") \__mp_input257.Y__gate_cover (\__mp_input257.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input258.A__gate_cover (\__mp_input258.A__gate );
  miter_def_prop #(1, "cover") \__mp_input258.Y__gate_cover (\__mp_input258.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input26.A__gate_cover (\__mp_input26.A__gate );
  miter_def_prop #(1, "cover") \__mp_input26.Y__gate_cover (\__mp_input26.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input27.A__gate_cover (\__mp_input27.A__gate );
  miter_def_prop #(1, "cover") \__mp_input27.Y__gate_cover (\__mp_input27.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input28.A__gate_cover (\__mp_input28.A__gate );
  miter_def_prop #(1, "cover") \__mp_input28.Y__gate_cover (\__mp_input28.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input29.A__gate_cover (\__mp_input29.A__gate );
  miter_def_prop #(1, "cover") \__mp_input29.Y__gate_cover (\__mp_input29.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input3.A__gate_cover (\__mp_input3.A__gate );
  miter_def_prop #(1, "cover") \__mp_input3.Y__gate_cover (\__mp_input3.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input30.A__gate_cover (\__mp_input30.A__gate );
  miter_def_prop #(1, "cover") \__mp_input30.Y__gate_cover (\__mp_input30.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input31.A__gate_cover (\__mp_input31.A__gate );
  miter_def_prop #(1, "cover") \__mp_input31.Y__gate_cover (\__mp_input31.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input32.A__gate_cover (\__mp_input32.A__gate );
  miter_def_prop #(1, "cover") \__mp_input32.Y__gate_cover (\__mp_input32.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input33.A__gate_cover (\__mp_input33.A__gate );
  miter_def_prop #(1, "cover") \__mp_input33.Y__gate_cover (\__mp_input33.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input34.A__gate_cover (\__mp_input34.A__gate );
  miter_def_prop #(1, "cover") \__mp_input34.Y__gate_cover (\__mp_input34.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input35.A__gate_cover (\__mp_input35.A__gate );
  miter_def_prop #(1, "cover") \__mp_input35.Y__gate_cover (\__mp_input35.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input36.A__gate_cover (\__mp_input36.A__gate );
  miter_def_prop #(1, "cover") \__mp_input36.Y__gate_cover (\__mp_input36.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input37.A__gate_cover (\__mp_input37.A__gate );
  miter_def_prop #(1, "cover") \__mp_input37.Y__gate_cover (\__mp_input37.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input38.A__gate_cover (\__mp_input38.A__gate );
  miter_def_prop #(1, "cover") \__mp_input38.Y__gate_cover (\__mp_input38.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input39.A__gate_cover (\__mp_input39.A__gate );
  miter_def_prop #(1, "cover") \__mp_input39.Y__gate_cover (\__mp_input39.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input4.A__gate_cover (\__mp_input4.A__gate );
  miter_def_prop #(1, "cover") \__mp_input4.Y__gate_cover (\__mp_input4.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input40.A__gate_cover (\__mp_input40.A__gate );
  miter_def_prop #(1, "cover") \__mp_input40.Y__gate_cover (\__mp_input40.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input41.A__gate_cover (\__mp_input41.A__gate );
  miter_def_prop #(1, "cover") \__mp_input41.Y__gate_cover (\__mp_input41.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input42.A__gate_cover (\__mp_input42.A__gate );
  miter_def_prop #(1, "cover") \__mp_input42.Y__gate_cover (\__mp_input42.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input43.A__gate_cover (\__mp_input43.A__gate );
  miter_def_prop #(1, "cover") \__mp_input43.Y__gate_cover (\__mp_input43.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input44.A__gate_cover (\__mp_input44.A__gate );
  miter_def_prop #(1, "cover") \__mp_input44.Y__gate_cover (\__mp_input44.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input45.A__gate_cover (\__mp_input45.A__gate );
  miter_def_prop #(1, "cover") \__mp_input45.Y__gate_cover (\__mp_input45.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input46.A__gate_cover (\__mp_input46.A__gate );
  miter_def_prop #(1, "cover") \__mp_input46.Y__gate_cover (\__mp_input46.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input47.A__gate_cover (\__mp_input47.A__gate );
  miter_def_prop #(1, "cover") \__mp_input47.Y__gate_cover (\__mp_input47.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input48.A__gate_cover (\__mp_input48.A__gate );
  miter_def_prop #(1, "cover") \__mp_input48.Y__gate_cover (\__mp_input48.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input49.A__gate_cover (\__mp_input49.A__gate );
  miter_def_prop #(1, "cover") \__mp_input49.Y__gate_cover (\__mp_input49.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input5.A__gate_cover (\__mp_input5.A__gate );
  miter_def_prop #(1, "cover") \__mp_input5.Y__gate_cover (\__mp_input5.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input50.A__gate_cover (\__mp_input50.A__gate );
  miter_def_prop #(1, "cover") \__mp_input50.Y__gate_cover (\__mp_input50.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input51.A__gate_cover (\__mp_input51.A__gate );
  miter_def_prop #(1, "cover") \__mp_input51.Y__gate_cover (\__mp_input51.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input52.A__gate_cover (\__mp_input52.A__gate );
  miter_def_prop #(1, "cover") \__mp_input52.Y__gate_cover (\__mp_input52.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input53.A__gate_cover (\__mp_input53.A__gate );
  miter_def_prop #(1, "cover") \__mp_input53.Y__gate_cover (\__mp_input53.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input54.A__gate_cover (\__mp_input54.A__gate );
  miter_def_prop #(1, "cover") \__mp_input54.Y__gate_cover (\__mp_input54.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input55.A__gate_cover (\__mp_input55.A__gate );
  miter_def_prop #(1, "cover") \__mp_input55.Y__gate_cover (\__mp_input55.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input56.A__gate_cover (\__mp_input56.A__gate );
  miter_def_prop #(1, "cover") \__mp_input56.Y__gate_cover (\__mp_input56.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input57.A__gate_cover (\__mp_input57.A__gate );
  miter_def_prop #(1, "cover") \__mp_input57.Y__gate_cover (\__mp_input57.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input58.A__gate_cover (\__mp_input58.A__gate );
  miter_def_prop #(1, "cover") \__mp_input58.Y__gate_cover (\__mp_input58.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input59.A__gate_cover (\__mp_input59.A__gate );
  miter_def_prop #(1, "cover") \__mp_input59.Y__gate_cover (\__mp_input59.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input6.A__gate_cover (\__mp_input6.A__gate );
  miter_def_prop #(1, "cover") \__mp_input6.Y__gate_cover (\__mp_input6.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input60.A__gate_cover (\__mp_input60.A__gate );
  miter_def_prop #(1, "cover") \__mp_input60.Y__gate_cover (\__mp_input60.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input61.A__gate_cover (\__mp_input61.A__gate );
  miter_def_prop #(1, "cover") \__mp_input61.Y__gate_cover (\__mp_input61.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input62.A__gate_cover (\__mp_input62.A__gate );
  miter_def_prop #(1, "cover") \__mp_input62.Y__gate_cover (\__mp_input62.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input63.A__gate_cover (\__mp_input63.A__gate );
  miter_def_prop #(1, "cover") \__mp_input63.Y__gate_cover (\__mp_input63.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input64.A__gate_cover (\__mp_input64.A__gate );
  miter_def_prop #(1, "cover") \__mp_input64.Y__gate_cover (\__mp_input64.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input65.A__gate_cover (\__mp_input65.A__gate );
  miter_def_prop #(1, "cover") \__mp_input65.Y__gate_cover (\__mp_input65.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input66.A__gate_cover (\__mp_input66.A__gate );
  miter_def_prop #(1, "cover") \__mp_input66.Y__gate_cover (\__mp_input66.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input67.A__gate_cover (\__mp_input67.A__gate );
  miter_def_prop #(1, "cover") \__mp_input67.Y__gate_cover (\__mp_input67.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input68.A__gate_cover (\__mp_input68.A__gate );
  miter_def_prop #(1, "cover") \__mp_input68.Y__gate_cover (\__mp_input68.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input69.A__gate_cover (\__mp_input69.A__gate );
  miter_def_prop #(1, "cover") \__mp_input69.Y__gate_cover (\__mp_input69.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input7.A__gate_cover (\__mp_input7.A__gate );
  miter_def_prop #(1, "cover") \__mp_input7.Y__gate_cover (\__mp_input7.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input70.A__gate_cover (\__mp_input70.A__gate );
  miter_def_prop #(1, "cover") \__mp_input70.Y__gate_cover (\__mp_input70.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input71.A__gate_cover (\__mp_input71.A__gate );
  miter_def_prop #(1, "cover") \__mp_input71.Y__gate_cover (\__mp_input71.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input72.A__gate_cover (\__mp_input72.A__gate );
  miter_def_prop #(1, "cover") \__mp_input72.Y__gate_cover (\__mp_input72.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input73.A__gate_cover (\__mp_input73.A__gate );
  miter_def_prop #(1, "cover") \__mp_input73.Y__gate_cover (\__mp_input73.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input74.A__gate_cover (\__mp_input74.A__gate );
  miter_def_prop #(1, "cover") \__mp_input74.Y__gate_cover (\__mp_input74.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input75.A__gate_cover (\__mp_input75.A__gate );
  miter_def_prop #(1, "cover") \__mp_input75.Y__gate_cover (\__mp_input75.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input76.A__gate_cover (\__mp_input76.A__gate );
  miter_def_prop #(1, "cover") \__mp_input76.Y__gate_cover (\__mp_input76.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input77.A__gate_cover (\__mp_input77.A__gate );
  miter_def_prop #(1, "cover") \__mp_input77.Y__gate_cover (\__mp_input77.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input78.A__gate_cover (\__mp_input78.A__gate );
  miter_def_prop #(1, "cover") \__mp_input78.Y__gate_cover (\__mp_input78.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input79.A__gate_cover (\__mp_input79.A__gate );
  miter_def_prop #(1, "cover") \__mp_input79.Y__gate_cover (\__mp_input79.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input8.A__gate_cover (\__mp_input8.A__gate );
  miter_def_prop #(1, "cover") \__mp_input8.Y__gate_cover (\__mp_input8.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input80.A__gate_cover (\__mp_input80.A__gate );
  miter_def_prop #(1, "cover") \__mp_input80.Y__gate_cover (\__mp_input80.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input81.A__gate_cover (\__mp_input81.A__gate );
  miter_def_prop #(1, "cover") \__mp_input81.Y__gate_cover (\__mp_input81.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input82.A__gate_cover (\__mp_input82.A__gate );
  miter_def_prop #(1, "cover") \__mp_input82.Y__gate_cover (\__mp_input82.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input83.A__gate_cover (\__mp_input83.A__gate );
  miter_def_prop #(1, "cover") \__mp_input83.Y__gate_cover (\__mp_input83.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input84.A__gate_cover (\__mp_input84.A__gate );
  miter_def_prop #(1, "cover") \__mp_input84.Y__gate_cover (\__mp_input84.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input85.A__gate_cover (\__mp_input85.A__gate );
  miter_def_prop #(1, "cover") \__mp_input85.Y__gate_cover (\__mp_input85.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input86.A__gate_cover (\__mp_input86.A__gate );
  miter_def_prop #(1, "cover") \__mp_input86.Y__gate_cover (\__mp_input86.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input87.A__gate_cover (\__mp_input87.A__gate );
  miter_def_prop #(1, "cover") \__mp_input87.Y__gate_cover (\__mp_input87.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input88.A__gate_cover (\__mp_input88.A__gate );
  miter_def_prop #(1, "cover") \__mp_input88.Y__gate_cover (\__mp_input88.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input89.A__gate_cover (\__mp_input89.A__gate );
  miter_def_prop #(1, "cover") \__mp_input89.Y__gate_cover (\__mp_input89.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input9.A__gate_cover (\__mp_input9.A__gate );
  miter_def_prop #(1, "cover") \__mp_input9.Y__gate_cover (\__mp_input9.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input90.A__gate_cover (\__mp_input90.A__gate );
  miter_def_prop #(1, "cover") \__mp_input90.Y__gate_cover (\__mp_input90.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input91.A__gate_cover (\__mp_input91.A__gate );
  miter_def_prop #(1, "cover") \__mp_input91.Y__gate_cover (\__mp_input91.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input92.A__gate_cover (\__mp_input92.A__gate );
  miter_def_prop #(1, "cover") \__mp_input92.Y__gate_cover (\__mp_input92.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input93.A__gate_cover (\__mp_input93.A__gate );
  miter_def_prop #(1, "cover") \__mp_input93.Y__gate_cover (\__mp_input93.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input94.A__gate_cover (\__mp_input94.A__gate );
  miter_def_prop #(1, "cover") \__mp_input94.Y__gate_cover (\__mp_input94.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input95.A__gate_cover (\__mp_input95.A__gate );
  miter_def_prop #(1, "cover") \__mp_input95.Y__gate_cover (\__mp_input95.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input96.A__gate_cover (\__mp_input96.A__gate );
  miter_def_prop #(1, "cover") \__mp_input96.Y__gate_cover (\__mp_input96.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input97.A__gate_cover (\__mp_input97.A__gate );
  miter_def_prop #(1, "cover") \__mp_input97.Y__gate_cover (\__mp_input97.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input98.A__gate_cover (\__mp_input98.A__gate );
  miter_def_prop #(1, "cover") \__mp_input98.Y__gate_cover (\__mp_input98.Y__gate );
  miter_def_prop #(1, "cover") \__mp_input99.A__gate_cover (\__mp_input99.A__gate );
  miter_def_prop #(1, "cover") \__mp_input99.Y__gate_cover (\__mp_input99.Y__gate );
  miter_def_prop #(1, "cover") \__mp_ld_r$_DFF_P_.CLK__gate_cover (\__mp_ld_r$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_ld_r$_DFF_P_.D__gate_cover (\__mp_ld_r$_DFF_P_.D__gate );
  miter_def_prop #(1, "cover") \__mp_output259.A__gate_cover (\__mp_output259.A__gate );
  miter_def_prop #(1, "cover") \__mp_output259.Y__gate_cover (\__mp_output259.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output260.A__gate_cover (\__mp_output260.A__gate );
  miter_def_prop #(1, "cover") \__mp_output260.Y__gate_cover (\__mp_output260.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output261.A__gate_cover (\__mp_output261.A__gate );
  miter_def_prop #(1, "cover") \__mp_output261.Y__gate_cover (\__mp_output261.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output262.A__gate_cover (\__mp_output262.A__gate );
  miter_def_prop #(1, "cover") \__mp_output262.Y__gate_cover (\__mp_output262.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output263.A__gate_cover (\__mp_output263.A__gate );
  miter_def_prop #(1, "cover") \__mp_output263.Y__gate_cover (\__mp_output263.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output264.A__gate_cover (\__mp_output264.A__gate );
  miter_def_prop #(1, "cover") \__mp_output264.Y__gate_cover (\__mp_output264.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output265.A__gate_cover (\__mp_output265.A__gate );
  miter_def_prop #(1, "cover") \__mp_output265.Y__gate_cover (\__mp_output265.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output266.A__gate_cover (\__mp_output266.A__gate );
  miter_def_prop #(1, "cover") \__mp_output266.Y__gate_cover (\__mp_output266.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output267.A__gate_cover (\__mp_output267.A__gate );
  miter_def_prop #(1, "cover") \__mp_output267.Y__gate_cover (\__mp_output267.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output268.A__gate_cover (\__mp_output268.A__gate );
  miter_def_prop #(1, "cover") \__mp_output268.Y__gate_cover (\__mp_output268.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output269.A__gate_cover (\__mp_output269.A__gate );
  miter_def_prop #(1, "cover") \__mp_output269.Y__gate_cover (\__mp_output269.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output270.A__gate_cover (\__mp_output270.A__gate );
  miter_def_prop #(1, "cover") \__mp_output270.Y__gate_cover (\__mp_output270.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output271.A__gate_cover (\__mp_output271.A__gate );
  miter_def_prop #(1, "cover") \__mp_output271.Y__gate_cover (\__mp_output271.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output272.A__gate_cover (\__mp_output272.A__gate );
  miter_def_prop #(1, "cover") \__mp_output272.Y__gate_cover (\__mp_output272.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output273.A__gate_cover (\__mp_output273.A__gate );
  miter_def_prop #(1, "cover") \__mp_output273.Y__gate_cover (\__mp_output273.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output274.A__gate_cover (\__mp_output274.A__gate );
  miter_def_prop #(1, "cover") \__mp_output274.Y__gate_cover (\__mp_output274.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output275.A__gate_cover (\__mp_output275.A__gate );
  miter_def_prop #(1, "cover") \__mp_output275.Y__gate_cover (\__mp_output275.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output276.A__gate_cover (\__mp_output276.A__gate );
  miter_def_prop #(1, "cover") \__mp_output276.Y__gate_cover (\__mp_output276.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output277.A__gate_cover (\__mp_output277.A__gate );
  miter_def_prop #(1, "cover") \__mp_output277.Y__gate_cover (\__mp_output277.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output278.A__gate_cover (\__mp_output278.A__gate );
  miter_def_prop #(1, "cover") \__mp_output278.Y__gate_cover (\__mp_output278.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output279.A__gate_cover (\__mp_output279.A__gate );
  miter_def_prop #(1, "cover") \__mp_output279.Y__gate_cover (\__mp_output279.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output280.A__gate_cover (\__mp_output280.A__gate );
  miter_def_prop #(1, "cover") \__mp_output280.Y__gate_cover (\__mp_output280.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output281.A__gate_cover (\__mp_output281.A__gate );
  miter_def_prop #(1, "cover") \__mp_output281.Y__gate_cover (\__mp_output281.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output282.A__gate_cover (\__mp_output282.A__gate );
  miter_def_prop #(1, "cover") \__mp_output282.Y__gate_cover (\__mp_output282.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output283.A__gate_cover (\__mp_output283.A__gate );
  miter_def_prop #(1, "cover") \__mp_output283.Y__gate_cover (\__mp_output283.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output284.A__gate_cover (\__mp_output284.A__gate );
  miter_def_prop #(1, "cover") \__mp_output284.Y__gate_cover (\__mp_output284.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output285.A__gate_cover (\__mp_output285.A__gate );
  miter_def_prop #(1, "cover") \__mp_output285.Y__gate_cover (\__mp_output285.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output286.A__gate_cover (\__mp_output286.A__gate );
  miter_def_prop #(1, "cover") \__mp_output286.Y__gate_cover (\__mp_output286.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output287.A__gate_cover (\__mp_output287.A__gate );
  miter_def_prop #(1, "cover") \__mp_output287.Y__gate_cover (\__mp_output287.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output288.A__gate_cover (\__mp_output288.A__gate );
  miter_def_prop #(1, "cover") \__mp_output288.Y__gate_cover (\__mp_output288.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output289.A__gate_cover (\__mp_output289.A__gate );
  miter_def_prop #(1, "cover") \__mp_output289.Y__gate_cover (\__mp_output289.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output290.A__gate_cover (\__mp_output290.A__gate );
  miter_def_prop #(1, "cover") \__mp_output290.Y__gate_cover (\__mp_output290.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output291.A__gate_cover (\__mp_output291.A__gate );
  miter_def_prop #(1, "cover") \__mp_output291.Y__gate_cover (\__mp_output291.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output292.A__gate_cover (\__mp_output292.A__gate );
  miter_def_prop #(1, "cover") \__mp_output292.Y__gate_cover (\__mp_output292.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output293.A__gate_cover (\__mp_output293.A__gate );
  miter_def_prop #(1, "cover") \__mp_output293.Y__gate_cover (\__mp_output293.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output294.A__gate_cover (\__mp_output294.A__gate );
  miter_def_prop #(1, "cover") \__mp_output294.Y__gate_cover (\__mp_output294.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output295.A__gate_cover (\__mp_output295.A__gate );
  miter_def_prop #(1, "cover") \__mp_output295.Y__gate_cover (\__mp_output295.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output296.A__gate_cover (\__mp_output296.A__gate );
  miter_def_prop #(1, "cover") \__mp_output296.Y__gate_cover (\__mp_output296.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output297.A__gate_cover (\__mp_output297.A__gate );
  miter_def_prop #(1, "cover") \__mp_output297.Y__gate_cover (\__mp_output297.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output298.A__gate_cover (\__mp_output298.A__gate );
  miter_def_prop #(1, "cover") \__mp_output298.Y__gate_cover (\__mp_output298.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output299.A__gate_cover (\__mp_output299.A__gate );
  miter_def_prop #(1, "cover") \__mp_output299.Y__gate_cover (\__mp_output299.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output300.A__gate_cover (\__mp_output300.A__gate );
  miter_def_prop #(1, "cover") \__mp_output300.Y__gate_cover (\__mp_output300.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output301.A__gate_cover (\__mp_output301.A__gate );
  miter_def_prop #(1, "cover") \__mp_output301.Y__gate_cover (\__mp_output301.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output302.A__gate_cover (\__mp_output302.A__gate );
  miter_def_prop #(1, "cover") \__mp_output302.Y__gate_cover (\__mp_output302.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output303.A__gate_cover (\__mp_output303.A__gate );
  miter_def_prop #(1, "cover") \__mp_output303.Y__gate_cover (\__mp_output303.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output304.A__gate_cover (\__mp_output304.A__gate );
  miter_def_prop #(1, "cover") \__mp_output304.Y__gate_cover (\__mp_output304.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output305.A__gate_cover (\__mp_output305.A__gate );
  miter_def_prop #(1, "cover") \__mp_output305.Y__gate_cover (\__mp_output305.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output306.A__gate_cover (\__mp_output306.A__gate );
  miter_def_prop #(1, "cover") \__mp_output306.Y__gate_cover (\__mp_output306.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output307.A__gate_cover (\__mp_output307.A__gate );
  miter_def_prop #(1, "cover") \__mp_output307.Y__gate_cover (\__mp_output307.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output308.A__gate_cover (\__mp_output308.A__gate );
  miter_def_prop #(1, "cover") \__mp_output308.Y__gate_cover (\__mp_output308.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output309.A__gate_cover (\__mp_output309.A__gate );
  miter_def_prop #(1, "cover") \__mp_output309.Y__gate_cover (\__mp_output309.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output310.A__gate_cover (\__mp_output310.A__gate );
  miter_def_prop #(1, "cover") \__mp_output310.Y__gate_cover (\__mp_output310.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output311.A__gate_cover (\__mp_output311.A__gate );
  miter_def_prop #(1, "cover") \__mp_output311.Y__gate_cover (\__mp_output311.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output312.A__gate_cover (\__mp_output312.A__gate );
  miter_def_prop #(1, "cover") \__mp_output312.Y__gate_cover (\__mp_output312.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output313.A__gate_cover (\__mp_output313.A__gate );
  miter_def_prop #(1, "cover") \__mp_output313.Y__gate_cover (\__mp_output313.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output314.A__gate_cover (\__mp_output314.A__gate );
  miter_def_prop #(1, "cover") \__mp_output314.Y__gate_cover (\__mp_output314.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output315.A__gate_cover (\__mp_output315.A__gate );
  miter_def_prop #(1, "cover") \__mp_output315.Y__gate_cover (\__mp_output315.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output316.A__gate_cover (\__mp_output316.A__gate );
  miter_def_prop #(1, "cover") \__mp_output316.Y__gate_cover (\__mp_output316.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output317.A__gate_cover (\__mp_output317.A__gate );
  miter_def_prop #(1, "cover") \__mp_output317.Y__gate_cover (\__mp_output317.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output318.A__gate_cover (\__mp_output318.A__gate );
  miter_def_prop #(1, "cover") \__mp_output318.Y__gate_cover (\__mp_output318.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output319.A__gate_cover (\__mp_output319.A__gate );
  miter_def_prop #(1, "cover") \__mp_output319.Y__gate_cover (\__mp_output319.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output320.A__gate_cover (\__mp_output320.A__gate );
  miter_def_prop #(1, "cover") \__mp_output320.Y__gate_cover (\__mp_output320.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output321.A__gate_cover (\__mp_output321.A__gate );
  miter_def_prop #(1, "cover") \__mp_output321.Y__gate_cover (\__mp_output321.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output322.A__gate_cover (\__mp_output322.A__gate );
  miter_def_prop #(1, "cover") \__mp_output322.Y__gate_cover (\__mp_output322.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output323.A__gate_cover (\__mp_output323.A__gate );
  miter_def_prop #(1, "cover") \__mp_output323.Y__gate_cover (\__mp_output323.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output324.A__gate_cover (\__mp_output324.A__gate );
  miter_def_prop #(1, "cover") \__mp_output324.Y__gate_cover (\__mp_output324.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output325.A__gate_cover (\__mp_output325.A__gate );
  miter_def_prop #(1, "cover") \__mp_output325.Y__gate_cover (\__mp_output325.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output326.A__gate_cover (\__mp_output326.A__gate );
  miter_def_prop #(1, "cover") \__mp_output326.Y__gate_cover (\__mp_output326.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output327.A__gate_cover (\__mp_output327.A__gate );
  miter_def_prop #(1, "cover") \__mp_output327.Y__gate_cover (\__mp_output327.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output328.A__gate_cover (\__mp_output328.A__gate );
  miter_def_prop #(1, "cover") \__mp_output328.Y__gate_cover (\__mp_output328.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output329.A__gate_cover (\__mp_output329.A__gate );
  miter_def_prop #(1, "cover") \__mp_output329.Y__gate_cover (\__mp_output329.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output330.A__gate_cover (\__mp_output330.A__gate );
  miter_def_prop #(1, "cover") \__mp_output330.Y__gate_cover (\__mp_output330.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output331.A__gate_cover (\__mp_output331.A__gate );
  miter_def_prop #(1, "cover") \__mp_output331.Y__gate_cover (\__mp_output331.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output332.A__gate_cover (\__mp_output332.A__gate );
  miter_def_prop #(1, "cover") \__mp_output332.Y__gate_cover (\__mp_output332.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output333.A__gate_cover (\__mp_output333.A__gate );
  miter_def_prop #(1, "cover") \__mp_output333.Y__gate_cover (\__mp_output333.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output334.A__gate_cover (\__mp_output334.A__gate );
  miter_def_prop #(1, "cover") \__mp_output334.Y__gate_cover (\__mp_output334.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output335.A__gate_cover (\__mp_output335.A__gate );
  miter_def_prop #(1, "cover") \__mp_output335.Y__gate_cover (\__mp_output335.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output336.A__gate_cover (\__mp_output336.A__gate );
  miter_def_prop #(1, "cover") \__mp_output336.Y__gate_cover (\__mp_output336.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output337.A__gate_cover (\__mp_output337.A__gate );
  miter_def_prop #(1, "cover") \__mp_output337.Y__gate_cover (\__mp_output337.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output338.A__gate_cover (\__mp_output338.A__gate );
  miter_def_prop #(1, "cover") \__mp_output338.Y__gate_cover (\__mp_output338.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output339.A__gate_cover (\__mp_output339.A__gate );
  miter_def_prop #(1, "cover") \__mp_output339.Y__gate_cover (\__mp_output339.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output340.A__gate_cover (\__mp_output340.A__gate );
  miter_def_prop #(1, "cover") \__mp_output340.Y__gate_cover (\__mp_output340.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output341.A__gate_cover (\__mp_output341.A__gate );
  miter_def_prop #(1, "cover") \__mp_output341.Y__gate_cover (\__mp_output341.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output342.A__gate_cover (\__mp_output342.A__gate );
  miter_def_prop #(1, "cover") \__mp_output342.Y__gate_cover (\__mp_output342.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output343.A__gate_cover (\__mp_output343.A__gate );
  miter_def_prop #(1, "cover") \__mp_output343.Y__gate_cover (\__mp_output343.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output344.A__gate_cover (\__mp_output344.A__gate );
  miter_def_prop #(1, "cover") \__mp_output344.Y__gate_cover (\__mp_output344.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output345.A__gate_cover (\__mp_output345.A__gate );
  miter_def_prop #(1, "cover") \__mp_output345.Y__gate_cover (\__mp_output345.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output346.A__gate_cover (\__mp_output346.A__gate );
  miter_def_prop #(1, "cover") \__mp_output346.Y__gate_cover (\__mp_output346.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output347.A__gate_cover (\__mp_output347.A__gate );
  miter_def_prop #(1, "cover") \__mp_output347.Y__gate_cover (\__mp_output347.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output348.A__gate_cover (\__mp_output348.A__gate );
  miter_def_prop #(1, "cover") \__mp_output348.Y__gate_cover (\__mp_output348.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output349.A__gate_cover (\__mp_output349.A__gate );
  miter_def_prop #(1, "cover") \__mp_output349.Y__gate_cover (\__mp_output349.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output350.A__gate_cover (\__mp_output350.A__gate );
  miter_def_prop #(1, "cover") \__mp_output350.Y__gate_cover (\__mp_output350.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output351.A__gate_cover (\__mp_output351.A__gate );
  miter_def_prop #(1, "cover") \__mp_output351.Y__gate_cover (\__mp_output351.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output352.A__gate_cover (\__mp_output352.A__gate );
  miter_def_prop #(1, "cover") \__mp_output352.Y__gate_cover (\__mp_output352.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output353.A__gate_cover (\__mp_output353.A__gate );
  miter_def_prop #(1, "cover") \__mp_output353.Y__gate_cover (\__mp_output353.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output354.A__gate_cover (\__mp_output354.A__gate );
  miter_def_prop #(1, "cover") \__mp_output354.Y__gate_cover (\__mp_output354.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output355.A__gate_cover (\__mp_output355.A__gate );
  miter_def_prop #(1, "cover") \__mp_output355.Y__gate_cover (\__mp_output355.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output356.A__gate_cover (\__mp_output356.A__gate );
  miter_def_prop #(1, "cover") \__mp_output356.Y__gate_cover (\__mp_output356.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output357.A__gate_cover (\__mp_output357.A__gate );
  miter_def_prop #(1, "cover") \__mp_output357.Y__gate_cover (\__mp_output357.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output358.A__gate_cover (\__mp_output358.A__gate );
  miter_def_prop #(1, "cover") \__mp_output358.Y__gate_cover (\__mp_output358.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output359.A__gate_cover (\__mp_output359.A__gate );
  miter_def_prop #(1, "cover") \__mp_output359.Y__gate_cover (\__mp_output359.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output360.A__gate_cover (\__mp_output360.A__gate );
  miter_def_prop #(1, "cover") \__mp_output360.Y__gate_cover (\__mp_output360.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output361.A__gate_cover (\__mp_output361.A__gate );
  miter_def_prop #(1, "cover") \__mp_output361.Y__gate_cover (\__mp_output361.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output362.A__gate_cover (\__mp_output362.A__gate );
  miter_def_prop #(1, "cover") \__mp_output362.Y__gate_cover (\__mp_output362.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output363.A__gate_cover (\__mp_output363.A__gate );
  miter_def_prop #(1, "cover") \__mp_output363.Y__gate_cover (\__mp_output363.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output364.A__gate_cover (\__mp_output364.A__gate );
  miter_def_prop #(1, "cover") \__mp_output364.Y__gate_cover (\__mp_output364.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output365.A__gate_cover (\__mp_output365.A__gate );
  miter_def_prop #(1, "cover") \__mp_output365.Y__gate_cover (\__mp_output365.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output366.A__gate_cover (\__mp_output366.A__gate );
  miter_def_prop #(1, "cover") \__mp_output366.Y__gate_cover (\__mp_output366.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output367.A__gate_cover (\__mp_output367.A__gate );
  miter_def_prop #(1, "cover") \__mp_output367.Y__gate_cover (\__mp_output367.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output368.A__gate_cover (\__mp_output368.A__gate );
  miter_def_prop #(1, "cover") \__mp_output368.Y__gate_cover (\__mp_output368.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output369.A__gate_cover (\__mp_output369.A__gate );
  miter_def_prop #(1, "cover") \__mp_output369.Y__gate_cover (\__mp_output369.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output370.A__gate_cover (\__mp_output370.A__gate );
  miter_def_prop #(1, "cover") \__mp_output370.Y__gate_cover (\__mp_output370.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output371.A__gate_cover (\__mp_output371.A__gate );
  miter_def_prop #(1, "cover") \__mp_output371.Y__gate_cover (\__mp_output371.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output372.A__gate_cover (\__mp_output372.A__gate );
  miter_def_prop #(1, "cover") \__mp_output372.Y__gate_cover (\__mp_output372.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output373.A__gate_cover (\__mp_output373.A__gate );
  miter_def_prop #(1, "cover") \__mp_output373.Y__gate_cover (\__mp_output373.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output374.A__gate_cover (\__mp_output374.A__gate );
  miter_def_prop #(1, "cover") \__mp_output374.Y__gate_cover (\__mp_output374.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output375.A__gate_cover (\__mp_output375.A__gate );
  miter_def_prop #(1, "cover") \__mp_output375.Y__gate_cover (\__mp_output375.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output376.A__gate_cover (\__mp_output376.A__gate );
  miter_def_prop #(1, "cover") \__mp_output376.Y__gate_cover (\__mp_output376.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output377.A__gate_cover (\__mp_output377.A__gate );
  miter_def_prop #(1, "cover") \__mp_output377.Y__gate_cover (\__mp_output377.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output378.A__gate_cover (\__mp_output378.A__gate );
  miter_def_prop #(1, "cover") \__mp_output378.Y__gate_cover (\__mp_output378.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output379.A__gate_cover (\__mp_output379.A__gate );
  miter_def_prop #(1, "cover") \__mp_output379.Y__gate_cover (\__mp_output379.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output380.A__gate_cover (\__mp_output380.A__gate );
  miter_def_prop #(1, "cover") \__mp_output380.Y__gate_cover (\__mp_output380.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output381.A__gate_cover (\__mp_output381.A__gate );
  miter_def_prop #(1, "cover") \__mp_output381.Y__gate_cover (\__mp_output381.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output382.A__gate_cover (\__mp_output382.A__gate );
  miter_def_prop #(1, "cover") \__mp_output382.Y__gate_cover (\__mp_output382.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output383.A__gate_cover (\__mp_output383.A__gate );
  miter_def_prop #(1, "cover") \__mp_output383.Y__gate_cover (\__mp_output383.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output384.A__gate_cover (\__mp_output384.A__gate );
  miter_def_prop #(1, "cover") \__mp_output384.Y__gate_cover (\__mp_output384.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output385.A__gate_cover (\__mp_output385.A__gate );
  miter_def_prop #(1, "cover") \__mp_output385.Y__gate_cover (\__mp_output385.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output386.A__gate_cover (\__mp_output386.A__gate );
  miter_def_prop #(1, "cover") \__mp_output386.Y__gate_cover (\__mp_output386.Y__gate );
  miter_def_prop #(1, "cover") \__mp_output387.A__gate_cover (\__mp_output387.A__gate );
  miter_def_prop #(1, "cover") \__mp_output387.Y__gate_cover (\__mp_output387.Y__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa00_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa00_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa01_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa01_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa02_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa02_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa03_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa03_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa10_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa10_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa11_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa11_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa12_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa12_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa13_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa13_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa20_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa20_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa21_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa21_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa22_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa22_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa23_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa23_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa30_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa30_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa31_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa31_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa32_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa32_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[0]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[1]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[2]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[3]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[4]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[5]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[6]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_sa33_sr[7]$_DFF_P_.CLK__gate_cover (\__mp_sa33_sr[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[0]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[0]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[100]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[100]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[101]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[101]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[102]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[102]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[103]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[103]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[104]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[104]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[105]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[105]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[106]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[106]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[107]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[107]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[108]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[108]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[109]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[109]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[10]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[10]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[110]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[110]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[111]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[111]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[112]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[112]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[113]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[113]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[114]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[114]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[115]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[115]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[116]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[116]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[117]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[117]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[118]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[118]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[119]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[119]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[11]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[11]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[120]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[120]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[121]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[121]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[122]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[122]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[123]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[123]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[124]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[124]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[125]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[125]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[126]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[126]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[127]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[127]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[12]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[12]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[13]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[13]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[14]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[14]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[15]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[15]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[16]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[16]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[17]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[17]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[18]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[18]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[19]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[19]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[1]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[1]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[20]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[20]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[21]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[21]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[22]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[22]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[23]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[23]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[24]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[24]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[25]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[25]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[26]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[26]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[27]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[27]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[28]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[28]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[29]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[29]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[2]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[2]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[30]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[30]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[31]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[31]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[32]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[32]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[33]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[33]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[34]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[34]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[35]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[35]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[36]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[36]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[37]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[37]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[38]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[38]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[39]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[39]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[3]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[3]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[40]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[40]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[41]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[41]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[42]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[42]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[43]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[43]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[44]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[44]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[45]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[45]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[46]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[46]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[47]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[47]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[48]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[48]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[49]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[49]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[4]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[4]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[50]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[50]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[51]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[51]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[52]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[52]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[53]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[53]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[54]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[54]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[55]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[55]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[56]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[56]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[57]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[57]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[58]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[58]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[59]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[59]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[5]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[5]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[60]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[60]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[61]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[61]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[62]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[62]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[63]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[63]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[64]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[64]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[65]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[65]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[66]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[66]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[67]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[67]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[68]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[68]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[69]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[69]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[6]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[6]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[70]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[70]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[71]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[71]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[72]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[72]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[73]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[73]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[74]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[74]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[75]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[75]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[76]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[76]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[77]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[77]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[78]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[78]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[79]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[79]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[7]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[7]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[80]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[80]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[81]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[81]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[82]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[82]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[83]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[83]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[84]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[84]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[85]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[85]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[86]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[86]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[87]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[87]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[88]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[88]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[89]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[89]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[8]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[8]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[90]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[90]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[91]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[91]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[92]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[92]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[93]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[93]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[94]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[94]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[95]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[95]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[96]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[96]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[97]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[97]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[98]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[98]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[99]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[99]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_in_r[9]$_DFFE_PP_.CLK__gate_cover (\__mp_text_in_r[9]$_DFFE_PP_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[0]$_DFF_P_.CLK__gate_cover (\__mp_text_out[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[0]$_DFF_P_.QN__gate_cover (\__mp_text_out[0]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[0]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[100]$_DFF_P_.CLK__gate_cover (\__mp_text_out[100]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[100]$_DFF_P_.QN__gate_cover (\__mp_text_out[100]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[100]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[101]$_DFF_P_.CLK__gate_cover (\__mp_text_out[101]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[101]$_DFF_P_.QN__gate_cover (\__mp_text_out[101]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[101]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[102]$_DFF_P_.CLK__gate_cover (\__mp_text_out[102]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[102]$_DFF_P_.QN__gate_cover (\__mp_text_out[102]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[102]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[103]$_DFF_P_.CLK__gate_cover (\__mp_text_out[103]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[103]$_DFF_P_.QN__gate_cover (\__mp_text_out[103]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[103]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[104]$_DFF_P_.CLK__gate_cover (\__mp_text_out[104]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[104]$_DFF_P_.QN__gate_cover (\__mp_text_out[104]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[104]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[105]$_DFF_P_.CLK__gate_cover (\__mp_text_out[105]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[105]$_DFF_P_.QN__gate_cover (\__mp_text_out[105]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[105]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[106]$_DFF_P_.CLK__gate_cover (\__mp_text_out[106]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[106]$_DFF_P_.QN__gate_cover (\__mp_text_out[106]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[106]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[107]$_DFF_P_.CLK__gate_cover (\__mp_text_out[107]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[107]$_DFF_P_.QN__gate_cover (\__mp_text_out[107]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[107]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[108]$_DFF_P_.CLK__gate_cover (\__mp_text_out[108]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[108]$_DFF_P_.QN__gate_cover (\__mp_text_out[108]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[108]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[109]$_DFF_P_.CLK__gate_cover (\__mp_text_out[109]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[109]$_DFF_P_.QN__gate_cover (\__mp_text_out[109]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[109]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[10]$_DFF_P_.CLK__gate_cover (\__mp_text_out[10]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[10]$_DFF_P_.QN__gate_cover (\__mp_text_out[10]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[10]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[110]$_DFF_P_.CLK__gate_cover (\__mp_text_out[110]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[110]$_DFF_P_.QN__gate_cover (\__mp_text_out[110]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[110]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[111]$_DFF_P_.CLK__gate_cover (\__mp_text_out[111]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[111]$_DFF_P_.QN__gate_cover (\__mp_text_out[111]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[111]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[112]$_DFF_P_.CLK__gate_cover (\__mp_text_out[112]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[112]$_DFF_P_.QN__gate_cover (\__mp_text_out[112]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[112]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[113]$_DFF_P_.CLK__gate_cover (\__mp_text_out[113]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[113]$_DFF_P_.QN__gate_cover (\__mp_text_out[113]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[113]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[114]$_DFF_P_.CLK__gate_cover (\__mp_text_out[114]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[114]$_DFF_P_.QN__gate_cover (\__mp_text_out[114]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[114]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[115]$_DFF_P_.CLK__gate_cover (\__mp_text_out[115]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[115]$_DFF_P_.QN__gate_cover (\__mp_text_out[115]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[115]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[116]$_DFF_P_.CLK__gate_cover (\__mp_text_out[116]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[116]$_DFF_P_.QN__gate_cover (\__mp_text_out[116]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[116]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[117]$_DFF_P_.CLK__gate_cover (\__mp_text_out[117]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[117]$_DFF_P_.QN__gate_cover (\__mp_text_out[117]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[117]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[118]$_DFF_P_.CLK__gate_cover (\__mp_text_out[118]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[118]$_DFF_P_.QN__gate_cover (\__mp_text_out[118]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[118]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[119]$_DFF_P_.CLK__gate_cover (\__mp_text_out[119]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[119]$_DFF_P_.QN__gate_cover (\__mp_text_out[119]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[119]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[11]$_DFF_P_.CLK__gate_cover (\__mp_text_out[11]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[11]$_DFF_P_.QN__gate_cover (\__mp_text_out[11]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[11]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[120]$_DFF_P_.CLK__gate_cover (\__mp_text_out[120]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[120]$_DFF_P_.QN__gate_cover (\__mp_text_out[120]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[120]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[121]$_DFF_P_.CLK__gate_cover (\__mp_text_out[121]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[121]$_DFF_P_.QN__gate_cover (\__mp_text_out[121]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[121]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[122]$_DFF_P_.CLK__gate_cover (\__mp_text_out[122]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[122]$_DFF_P_.QN__gate_cover (\__mp_text_out[122]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[122]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[123]$_DFF_P_.CLK__gate_cover (\__mp_text_out[123]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[123]$_DFF_P_.QN__gate_cover (\__mp_text_out[123]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[123]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[124]$_DFF_P_.CLK__gate_cover (\__mp_text_out[124]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[124]$_DFF_P_.QN__gate_cover (\__mp_text_out[124]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[124]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[125]$_DFF_P_.CLK__gate_cover (\__mp_text_out[125]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[125]$_DFF_P_.QN__gate_cover (\__mp_text_out[125]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[125]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[126]$_DFF_P_.CLK__gate_cover (\__mp_text_out[126]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[126]$_DFF_P_.QN__gate_cover (\__mp_text_out[126]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[126]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[127]$_DFF_P_.CLK__gate_cover (\__mp_text_out[127]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[127]$_DFF_P_.QN__gate_cover (\__mp_text_out[127]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[127]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[12]$_DFF_P_.CLK__gate_cover (\__mp_text_out[12]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[12]$_DFF_P_.QN__gate_cover (\__mp_text_out[12]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[12]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[13]$_DFF_P_.CLK__gate_cover (\__mp_text_out[13]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[13]$_DFF_P_.QN__gate_cover (\__mp_text_out[13]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[13]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[14]$_DFF_P_.CLK__gate_cover (\__mp_text_out[14]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[14]$_DFF_P_.QN__gate_cover (\__mp_text_out[14]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[14]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[15]$_DFF_P_.CLK__gate_cover (\__mp_text_out[15]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[15]$_DFF_P_.QN__gate_cover (\__mp_text_out[15]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[15]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[16]$_DFF_P_.CLK__gate_cover (\__mp_text_out[16]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[16]$_DFF_P_.QN__gate_cover (\__mp_text_out[16]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[16]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[17]$_DFF_P_.CLK__gate_cover (\__mp_text_out[17]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[17]$_DFF_P_.QN__gate_cover (\__mp_text_out[17]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[17]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[18]$_DFF_P_.CLK__gate_cover (\__mp_text_out[18]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[18]$_DFF_P_.QN__gate_cover (\__mp_text_out[18]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[18]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[19]$_DFF_P_.CLK__gate_cover (\__mp_text_out[19]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[19]$_DFF_P_.QN__gate_cover (\__mp_text_out[19]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[19]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[1]$_DFF_P_.CLK__gate_cover (\__mp_text_out[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[1]$_DFF_P_.QN__gate_cover (\__mp_text_out[1]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[1]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[20]$_DFF_P_.CLK__gate_cover (\__mp_text_out[20]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[20]$_DFF_P_.QN__gate_cover (\__mp_text_out[20]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[20]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[21]$_DFF_P_.CLK__gate_cover (\__mp_text_out[21]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[21]$_DFF_P_.QN__gate_cover (\__mp_text_out[21]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[21]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[22]$_DFF_P_.CLK__gate_cover (\__mp_text_out[22]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[22]$_DFF_P_.QN__gate_cover (\__mp_text_out[22]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[22]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[23]$_DFF_P_.CLK__gate_cover (\__mp_text_out[23]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[23]$_DFF_P_.QN__gate_cover (\__mp_text_out[23]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[23]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[24]$_DFF_P_.CLK__gate_cover (\__mp_text_out[24]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[24]$_DFF_P_.QN__gate_cover (\__mp_text_out[24]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[24]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[25]$_DFF_P_.CLK__gate_cover (\__mp_text_out[25]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[25]$_DFF_P_.QN__gate_cover (\__mp_text_out[25]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[25]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[26]$_DFF_P_.CLK__gate_cover (\__mp_text_out[26]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[26]$_DFF_P_.QN__gate_cover (\__mp_text_out[26]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[26]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[27]$_DFF_P_.CLK__gate_cover (\__mp_text_out[27]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[27]$_DFF_P_.QN__gate_cover (\__mp_text_out[27]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[27]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[28]$_DFF_P_.CLK__gate_cover (\__mp_text_out[28]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[28]$_DFF_P_.QN__gate_cover (\__mp_text_out[28]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[28]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[29]$_DFF_P_.CLK__gate_cover (\__mp_text_out[29]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[29]$_DFF_P_.QN__gate_cover (\__mp_text_out[29]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[29]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[2]$_DFF_P_.CLK__gate_cover (\__mp_text_out[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[2]$_DFF_P_.QN__gate_cover (\__mp_text_out[2]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[2]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[30]$_DFF_P_.CLK__gate_cover (\__mp_text_out[30]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[30]$_DFF_P_.QN__gate_cover (\__mp_text_out[30]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[30]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[31]$_DFF_P_.CLK__gate_cover (\__mp_text_out[31]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[31]$_DFF_P_.QN__gate_cover (\__mp_text_out[31]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[31]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[32]$_DFF_P_.CLK__gate_cover (\__mp_text_out[32]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[32]$_DFF_P_.QN__gate_cover (\__mp_text_out[32]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[32]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[33]$_DFF_P_.CLK__gate_cover (\__mp_text_out[33]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[33]$_DFF_P_.QN__gate_cover (\__mp_text_out[33]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[33]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[34]$_DFF_P_.CLK__gate_cover (\__mp_text_out[34]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[34]$_DFF_P_.QN__gate_cover (\__mp_text_out[34]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[34]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[35]$_DFF_P_.CLK__gate_cover (\__mp_text_out[35]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[35]$_DFF_P_.QN__gate_cover (\__mp_text_out[35]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[35]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[36]$_DFF_P_.CLK__gate_cover (\__mp_text_out[36]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[36]$_DFF_P_.QN__gate_cover (\__mp_text_out[36]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[36]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[37]$_DFF_P_.CLK__gate_cover (\__mp_text_out[37]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[37]$_DFF_P_.QN__gate_cover (\__mp_text_out[37]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[37]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[38]$_DFF_P_.CLK__gate_cover (\__mp_text_out[38]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[38]$_DFF_P_.QN__gate_cover (\__mp_text_out[38]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[38]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[39]$_DFF_P_.CLK__gate_cover (\__mp_text_out[39]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[39]$_DFF_P_.QN__gate_cover (\__mp_text_out[39]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[39]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[3]$_DFF_P_.CLK__gate_cover (\__mp_text_out[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[3]$_DFF_P_.QN__gate_cover (\__mp_text_out[3]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[3]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[40]$_DFF_P_.CLK__gate_cover (\__mp_text_out[40]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[40]$_DFF_P_.QN__gate_cover (\__mp_text_out[40]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[40]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[41]$_DFF_P_.CLK__gate_cover (\__mp_text_out[41]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[41]$_DFF_P_.QN__gate_cover (\__mp_text_out[41]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[41]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[42]$_DFF_P_.CLK__gate_cover (\__mp_text_out[42]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[42]$_DFF_P_.QN__gate_cover (\__mp_text_out[42]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[42]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[43]$_DFF_P_.CLK__gate_cover (\__mp_text_out[43]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[43]$_DFF_P_.QN__gate_cover (\__mp_text_out[43]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[43]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[44]$_DFF_P_.CLK__gate_cover (\__mp_text_out[44]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[44]$_DFF_P_.QN__gate_cover (\__mp_text_out[44]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[44]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[45]$_DFF_P_.CLK__gate_cover (\__mp_text_out[45]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[45]$_DFF_P_.QN__gate_cover (\__mp_text_out[45]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[45]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[46]$_DFF_P_.CLK__gate_cover (\__mp_text_out[46]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[46]$_DFF_P_.QN__gate_cover (\__mp_text_out[46]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[46]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[47]$_DFF_P_.CLK__gate_cover (\__mp_text_out[47]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[47]$_DFF_P_.QN__gate_cover (\__mp_text_out[47]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[47]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[48]$_DFF_P_.CLK__gate_cover (\__mp_text_out[48]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[48]$_DFF_P_.QN__gate_cover (\__mp_text_out[48]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[48]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[49]$_DFF_P_.CLK__gate_cover (\__mp_text_out[49]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[49]$_DFF_P_.QN__gate_cover (\__mp_text_out[49]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[49]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[4]$_DFF_P_.CLK__gate_cover (\__mp_text_out[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[4]$_DFF_P_.QN__gate_cover (\__mp_text_out[4]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[4]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[50]$_DFF_P_.CLK__gate_cover (\__mp_text_out[50]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[50]$_DFF_P_.QN__gate_cover (\__mp_text_out[50]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[50]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[51]$_DFF_P_.CLK__gate_cover (\__mp_text_out[51]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[51]$_DFF_P_.QN__gate_cover (\__mp_text_out[51]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[51]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[52]$_DFF_P_.CLK__gate_cover (\__mp_text_out[52]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[52]$_DFF_P_.QN__gate_cover (\__mp_text_out[52]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[52]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[53]$_DFF_P_.CLK__gate_cover (\__mp_text_out[53]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[53]$_DFF_P_.QN__gate_cover (\__mp_text_out[53]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[53]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[54]$_DFF_P_.CLK__gate_cover (\__mp_text_out[54]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[54]$_DFF_P_.QN__gate_cover (\__mp_text_out[54]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[54]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[55]$_DFF_P_.CLK__gate_cover (\__mp_text_out[55]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[55]$_DFF_P_.QN__gate_cover (\__mp_text_out[55]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[55]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[56]$_DFF_P_.CLK__gate_cover (\__mp_text_out[56]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[56]$_DFF_P_.QN__gate_cover (\__mp_text_out[56]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[56]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[57]$_DFF_P_.CLK__gate_cover (\__mp_text_out[57]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[57]$_DFF_P_.QN__gate_cover (\__mp_text_out[57]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[57]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[58]$_DFF_P_.CLK__gate_cover (\__mp_text_out[58]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[58]$_DFF_P_.QN__gate_cover (\__mp_text_out[58]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[58]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[59]$_DFF_P_.CLK__gate_cover (\__mp_text_out[59]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[59]$_DFF_P_.QN__gate_cover (\__mp_text_out[59]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[59]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[5]$_DFF_P_.CLK__gate_cover (\__mp_text_out[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[5]$_DFF_P_.QN__gate_cover (\__mp_text_out[5]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[5]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[60]$_DFF_P_.CLK__gate_cover (\__mp_text_out[60]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[60]$_DFF_P_.QN__gate_cover (\__mp_text_out[60]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[60]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[61]$_DFF_P_.CLK__gate_cover (\__mp_text_out[61]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[61]$_DFF_P_.QN__gate_cover (\__mp_text_out[61]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[61]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[62]$_DFF_P_.CLK__gate_cover (\__mp_text_out[62]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[62]$_DFF_P_.QN__gate_cover (\__mp_text_out[62]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[62]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[63]$_DFF_P_.CLK__gate_cover (\__mp_text_out[63]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[63]$_DFF_P_.QN__gate_cover (\__mp_text_out[63]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[63]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[64]$_DFF_P_.CLK__gate_cover (\__mp_text_out[64]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[64]$_DFF_P_.QN__gate_cover (\__mp_text_out[64]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[64]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[65]$_DFF_P_.CLK__gate_cover (\__mp_text_out[65]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[65]$_DFF_P_.QN__gate_cover (\__mp_text_out[65]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[65]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[66]$_DFF_P_.CLK__gate_cover (\__mp_text_out[66]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[66]$_DFF_P_.QN__gate_cover (\__mp_text_out[66]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[66]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[67]$_DFF_P_.CLK__gate_cover (\__mp_text_out[67]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[67]$_DFF_P_.QN__gate_cover (\__mp_text_out[67]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[67]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[68]$_DFF_P_.CLK__gate_cover (\__mp_text_out[68]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[68]$_DFF_P_.QN__gate_cover (\__mp_text_out[68]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[68]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[69]$_DFF_P_.CLK__gate_cover (\__mp_text_out[69]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[69]$_DFF_P_.QN__gate_cover (\__mp_text_out[69]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[69]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[6]$_DFF_P_.CLK__gate_cover (\__mp_text_out[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[6]$_DFF_P_.QN__gate_cover (\__mp_text_out[6]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[6]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[70]$_DFF_P_.CLK__gate_cover (\__mp_text_out[70]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[70]$_DFF_P_.QN__gate_cover (\__mp_text_out[70]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[70]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[71]$_DFF_P_.CLK__gate_cover (\__mp_text_out[71]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[71]$_DFF_P_.QN__gate_cover (\__mp_text_out[71]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[71]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[72]$_DFF_P_.CLK__gate_cover (\__mp_text_out[72]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[72]$_DFF_P_.QN__gate_cover (\__mp_text_out[72]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[72]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[73]$_DFF_P_.CLK__gate_cover (\__mp_text_out[73]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[73]$_DFF_P_.QN__gate_cover (\__mp_text_out[73]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[73]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[74]$_DFF_P_.CLK__gate_cover (\__mp_text_out[74]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[74]$_DFF_P_.QN__gate_cover (\__mp_text_out[74]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[74]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[75]$_DFF_P_.CLK__gate_cover (\__mp_text_out[75]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[75]$_DFF_P_.QN__gate_cover (\__mp_text_out[75]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[75]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[76]$_DFF_P_.CLK__gate_cover (\__mp_text_out[76]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[76]$_DFF_P_.QN__gate_cover (\__mp_text_out[76]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[76]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[77]$_DFF_P_.CLK__gate_cover (\__mp_text_out[77]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[77]$_DFF_P_.QN__gate_cover (\__mp_text_out[77]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[77]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[78]$_DFF_P_.CLK__gate_cover (\__mp_text_out[78]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[78]$_DFF_P_.QN__gate_cover (\__mp_text_out[78]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[78]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[79]$_DFF_P_.CLK__gate_cover (\__mp_text_out[79]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[79]$_DFF_P_.QN__gate_cover (\__mp_text_out[79]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[79]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[7]$_DFF_P_.CLK__gate_cover (\__mp_text_out[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[7]$_DFF_P_.QN__gate_cover (\__mp_text_out[7]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[7]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[80]$_DFF_P_.CLK__gate_cover (\__mp_text_out[80]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[80]$_DFF_P_.QN__gate_cover (\__mp_text_out[80]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[80]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[81]$_DFF_P_.CLK__gate_cover (\__mp_text_out[81]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[81]$_DFF_P_.QN__gate_cover (\__mp_text_out[81]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[81]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[82]$_DFF_P_.CLK__gate_cover (\__mp_text_out[82]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[82]$_DFF_P_.QN__gate_cover (\__mp_text_out[82]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[82]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[83]$_DFF_P_.CLK__gate_cover (\__mp_text_out[83]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[83]$_DFF_P_.QN__gate_cover (\__mp_text_out[83]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[83]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[84]$_DFF_P_.CLK__gate_cover (\__mp_text_out[84]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[84]$_DFF_P_.QN__gate_cover (\__mp_text_out[84]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[84]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[85]$_DFF_P_.CLK__gate_cover (\__mp_text_out[85]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[85]$_DFF_P_.QN__gate_cover (\__mp_text_out[85]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[85]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[86]$_DFF_P_.CLK__gate_cover (\__mp_text_out[86]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[86]$_DFF_P_.QN__gate_cover (\__mp_text_out[86]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[86]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[87]$_DFF_P_.CLK__gate_cover (\__mp_text_out[87]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[87]$_DFF_P_.QN__gate_cover (\__mp_text_out[87]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[87]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[88]$_DFF_P_.CLK__gate_cover (\__mp_text_out[88]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[88]$_DFF_P_.QN__gate_cover (\__mp_text_out[88]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[88]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[89]$_DFF_P_.CLK__gate_cover (\__mp_text_out[89]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[89]$_DFF_P_.QN__gate_cover (\__mp_text_out[89]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[89]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[8]$_DFF_P_.CLK__gate_cover (\__mp_text_out[8]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[8]$_DFF_P_.QN__gate_cover (\__mp_text_out[8]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[8]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[90]$_DFF_P_.CLK__gate_cover (\__mp_text_out[90]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[90]$_DFF_P_.QN__gate_cover (\__mp_text_out[90]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[90]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[91]$_DFF_P_.CLK__gate_cover (\__mp_text_out[91]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[91]$_DFF_P_.QN__gate_cover (\__mp_text_out[91]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[91]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[92]$_DFF_P_.CLK__gate_cover (\__mp_text_out[92]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[92]$_DFF_P_.QN__gate_cover (\__mp_text_out[92]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[92]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[93]$_DFF_P_.CLK__gate_cover (\__mp_text_out[93]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[93]$_DFF_P_.QN__gate_cover (\__mp_text_out[93]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[93]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[94]$_DFF_P_.CLK__gate_cover (\__mp_text_out[94]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[94]$_DFF_P_.QN__gate_cover (\__mp_text_out[94]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[94]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[95]$_DFF_P_.CLK__gate_cover (\__mp_text_out[95]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[95]$_DFF_P_.QN__gate_cover (\__mp_text_out[95]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[95]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[96]$_DFF_P_.CLK__gate_cover (\__mp_text_out[96]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[96]$_DFF_P_.QN__gate_cover (\__mp_text_out[96]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[96]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[97]$_DFF_P_.CLK__gate_cover (\__mp_text_out[97]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[97]$_DFF_P_.QN__gate_cover (\__mp_text_out[97]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[97]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[98]$_DFF_P_.CLK__gate_cover (\__mp_text_out[98]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[98]$_DFF_P_.QN__gate_cover (\__mp_text_out[98]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[98]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[99]$_DFF_P_.CLK__gate_cover (\__mp_text_out[99]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[99]$_DFF_P_.QN__gate_cover (\__mp_text_out[99]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[99]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[9]$_DFF_P_.CLK__gate_cover (\__mp_text_out[9]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[9]$_DFF_P_.QN__gate_cover (\__mp_text_out[9]$_DFF_P_.QN__gate );
  miter_def_prop #(1, "cover") \__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gate_cover (\__mp_text_out[9]$_DFF_P_.int_fwire_IQN__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gate_cover (\__mp_u0.r0.out[24]$_SDFF_PP1_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.out[25]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.out[26]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.out[27]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.out[28]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.out[29]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.out[30]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.out[31]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gate_cover (\__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[0]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[1]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[2]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[3]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[4]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[5]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[6]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u0.d[7]$_DFF_P_.CLK__gate_cover (\__mp_u0.u0.d[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[0]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[1]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[2]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[3]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[4]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[5]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[6]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u1.d[7]$_DFF_P_.CLK__gate_cover (\__mp_u0.u1.d[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[0]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[1]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[2]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[3]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[4]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[5]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[6]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u2.d[7]$_DFF_P_.CLK__gate_cover (\__mp_u0.u2.d[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[0]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[1]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[2]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[3]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[4]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[5]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[6]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.u3.d[7]$_DFF_P_.CLK__gate_cover (\__mp_u0.u3.d[7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][0]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][10]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][10]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][11]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][11]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][12]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][12]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][13]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][13]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][14]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][14]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][15]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][15]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][16]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][16]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][17]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][17]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][18]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][18]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][19]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][19]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][1]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][20]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][20]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][21]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][21]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][22]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][22]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][23]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][23]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][24]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][24]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][25]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][25]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][26]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][26]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][27]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][27]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][28]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][28]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][29]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][29]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][2]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][30]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][30]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][31]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][31]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][3]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][4]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][5]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][6]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][7]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][8]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][8]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[0][9]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[0][9]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][0]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][10]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][10]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][11]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][11]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][12]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][12]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][13]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][13]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][14]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][14]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][15]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][15]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][16]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][16]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][17]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][17]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][18]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][18]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][19]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][19]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][1]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][20]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][20]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][21]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][21]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][22]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][22]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][23]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][23]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][24]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][24]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][25]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][25]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][26]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][26]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][27]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][27]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][28]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][28]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][29]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][29]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][2]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][30]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][30]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][31]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][31]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][3]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][4]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][5]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][6]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][7]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][8]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][8]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[1][9]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[1][9]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][0]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][10]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][10]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][11]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][11]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][12]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][12]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][13]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][13]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][14]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][14]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][15]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][15]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][16]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][16]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][17]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][17]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][18]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][18]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][19]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][19]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][1]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][20]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][20]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][21]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][21]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][22]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][22]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][23]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][23]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][24]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][24]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][25]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][25]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][26]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][26]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][27]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][27]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][28]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][28]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][29]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][29]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][2]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][30]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][30]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][31]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][31]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][3]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][4]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][5]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][6]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][7]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][8]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][8]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[2][9]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[2][9]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][0]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][0]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][10]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][10]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][11]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][11]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][12]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][12]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][13]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][13]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][14]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][14]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][15]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][15]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][16]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][16]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][17]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][17]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][18]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][18]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][19]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][19]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][1]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][1]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][20]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][20]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][21]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][21]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][22]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][22]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][23]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][23]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][24]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][24]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][25]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][25]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][26]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][26]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][27]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][27]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][28]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][28]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][29]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][29]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][2]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][2]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][30]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][30]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][31]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][31]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][3]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][3]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][4]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][4]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][5]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][5]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][6]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][6]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][7]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][7]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][8]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][8]$_DFF_P_.CLK__gate );
  miter_def_prop #(1, "cover") \__mp_u0.w[3][9]$_DFF_P_.CLK__gate_cover (\__mp_u0.w[3][9]$_DFF_P_.CLK__gate );
`endif
`ifdef COVER_DEF_GOLD_OUTPUTS
  miter_def_prop #(1, "cover") \__po_done__gold_cover (\__po_done__gold );
  miter_def_prop #(128, "cover") \__po_text_out__gold_cover (\__po_text_out__gold );
`endif
`ifdef COVER_DEF_GATE_OUTPUTS
  miter_def_prop #(1, "cover") \__po_done__gate_cover (\__po_done__gate );
  miter_def_prop #(128, "cover") \__po_text_out__gate_cover (\__po_text_out__gate );
`endif
endmodule
module miter_cmp_prop #(parameter WIDTH=1, parameter TYPE="assert") (input [WIDTH-1:0] in_gold, in_gate);
  reg okay;
  integer i;
  always @* begin
    okay = 1;
    for (i = 0; i < WIDTH; i = i+1)
      okay = okay && (in_gold[i] === 1'bx || in_gold[i] === in_gate[i]);
  end
  generate
    if (TYPE == "assert") always @* assert(okay);
    if (TYPE == "assume") always @* assume(okay);
    if (TYPE == "cover")  always @* cover(okay);
  endgenerate
endmodule
module miter_def_prop #(parameter WIDTH=1, parameter TYPE="assert") (input [WIDTH-1:0] in);
  wire okay = ^in !== 1'bx;
  generate
    if (TYPE == "assert") always @* assert(okay);
    if (TYPE == "assume") always @* assume(okay);
    if (TYPE == "cover")  always @* cover(okay);
  endgenerate
endmodule
module \gold.aes_cipher_top (
  input  [  0:0] \__pi_clk ,
  input  [127:0] \__pi_key ,
  input  [  0:0] \__pi_ld ,
  input  [  0:0] \__pi_rst ,
  input  [127:0] \__pi_text_in ,
  output [  0:0] \__mp_clkbuf_0_clk.A ,
  output [  0:0] \__mp_clkbuf_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.Y ,
  output [  0:0] \__mp_clkload0.A ,
  output [  0:0] \__mp_clkload0.Y ,
  output [  0:0] \__mp_clkload1.A ,
  output [  0:0] \__mp_clkload10.A ,
  output [  0:0] \__mp_clkload11.A ,
  output [  0:0] \__mp_clkload12.A ,
  output [  0:0] \__mp_clkload13.A ,
  output [  0:0] \__mp_clkload14.A ,
  output [  0:0] \__mp_clkload15.A ,
  output [  0:0] \__mp_clkload16.A ,
  output [  0:0] \__mp_clkload17.A ,
  output [  0:0] \__mp_clkload18.A ,
  output [  0:0] \__mp_clkload18.Y ,
  output [  0:0] \__mp_clkload19.A ,
  output [  0:0] \__mp_clkload2.A ,
  output [  0:0] \__mp_clkload20.A ,
  output [  0:0] \__mp_clkload21.A ,
  output [  0:0] \__mp_clkload22.A ,
  output [  0:0] \__mp_clkload23.A ,
  output [  0:0] \__mp_clkload24.A ,
  output [  0:0] \__mp_clkload25.A ,
  output [  0:0] \__mp_clkload26.A ,
  output [  0:0] \__mp_clkload27.A ,
  output [  0:0] \__mp_clkload28.A ,
  output [  0:0] \__mp_clkload29.A ,
  output [  0:0] \__mp_clkload3.A ,
  output [  0:0] \__mp_clkload30.A ,
  output [  0:0] \__mp_clkload31.A ,
  output [  0:0] \__mp_clkload31.Y ,
  output [  0:0] \__mp_clkload32.A ,
  output [  0:0] \__mp_clkload4.A ,
  output [  0:0] \__mp_clkload5.A ,
  output [  0:0] \__mp_clkload6.A ,
  output [  0:0] \__mp_clkload7.A ,
  output [  0:0] \__mp_clkload8.A ,
  output [  0:0] \__mp_clkload9.A ,
  output [  0:0] \__mp_clknet_0_clk ,
  output [  0:0] \__mp_clknet_2_0_0_clk ,
  output [  0:0] \__mp_clknet_2_1_0_clk ,
  output [  0:0] \__mp_clknet_2_2_0_clk ,
  output [  0:0] \__mp_clknet_2_3_0_clk ,
  output [  0:0] \__mp_clknet_leaf_0_clk ,
  output [  0:0] \__mp_clknet_leaf_10_clk ,
  output [  0:0] \__mp_clknet_leaf_11_clk ,
  output [  0:0] \__mp_clknet_leaf_12_clk ,
  output [  0:0] \__mp_clknet_leaf_13_clk ,
  output [  0:0] \__mp_clknet_leaf_14_clk ,
  output [  0:0] \__mp_clknet_leaf_15_clk ,
  output [  0:0] \__mp_clknet_leaf_16_clk ,
  output [  0:0] \__mp_clknet_leaf_17_clk ,
  output [  0:0] \__mp_clknet_leaf_18_clk ,
  output [  0:0] \__mp_clknet_leaf_19_clk ,
  output [  0:0] \__mp_clknet_leaf_1_clk ,
  output [  0:0] \__mp_clknet_leaf_20_clk ,
  output [  0:0] \__mp_clknet_leaf_21_clk ,
  output [  0:0] \__mp_clknet_leaf_22_clk ,
  output [  0:0] \__mp_clknet_leaf_23_clk ,
  output [  0:0] \__mp_clknet_leaf_24_clk ,
  output [  0:0] \__mp_clknet_leaf_25_clk ,
  output [  0:0] \__mp_clknet_leaf_26_clk ,
  output [  0:0] \__mp_clknet_leaf_27_clk ,
  output [  0:0] \__mp_clknet_leaf_28_clk ,
  output [  0:0] \__mp_clknet_leaf_29_clk ,
  output [  0:0] \__mp_clknet_leaf_2_clk ,
  output [  0:0] \__mp_clknet_leaf_30_clk ,
  output [  0:0] \__mp_clknet_leaf_31_clk ,
  output [  0:0] \__mp_clknet_leaf_32_clk ,
  output [  0:0] \__mp_clknet_leaf_33_clk ,
  output [  0:0] \__mp_clknet_leaf_3_clk ,
  output [  0:0] \__mp_clknet_leaf_4_clk ,
  output [  0:0] \__mp_clknet_leaf_5_clk ,
  output [  0:0] \__mp_clknet_leaf_6_clk ,
  output [  0:0] \__mp_clknet_leaf_7_clk ,
  output [  0:0] \__mp_clknet_leaf_8_clk ,
  output [  0:0] \__mp_clknet_leaf_9_clk ,
  output [  0:0] \__mp_dcnt[0]$_SDFFE_PN0P_.CLK ,
  output [  0:0] \__mp_dcnt[1]$_SDFFE_PN0P_.CLK ,
  output [  0:0] \__mp_dcnt[2]$_SDFFE_PP0P_.CLK ,
  output [  0:0] \__mp_dcnt[3]$_SDFFE_PN0P_.CLK ,
  output [  0:0] \__mp_done$_DFF_P_.CLK ,
  output [  0:0] \__mp_done$_DFF_P_.QN ,
  output [  0:0] \__mp_done$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_input1.A ,
  output [  0:0] \__mp_input1.Y ,
  output [  0:0] \__mp_input10.A ,
  output [  0:0] \__mp_input10.Y ,
  output [  0:0] \__mp_input100.A ,
  output [  0:0] \__mp_input100.Y ,
  output [  0:0] \__mp_input101.A ,
  output [  0:0] \__mp_input101.Y ,
  output [  0:0] \__mp_input102.A ,
  output [  0:0] \__mp_input102.Y ,
  output [  0:0] \__mp_input103.A ,
  output [  0:0] \__mp_input103.Y ,
  output [  0:0] \__mp_input104.A ,
  output [  0:0] \__mp_input104.Y ,
  output [  0:0] \__mp_input105.A ,
  output [  0:0] \__mp_input105.Y ,
  output [  0:0] \__mp_input106.A ,
  output [  0:0] \__mp_input106.Y ,
  output [  0:0] \__mp_input107.A ,
  output [  0:0] \__mp_input107.Y ,
  output [  0:0] \__mp_input108.A ,
  output [  0:0] \__mp_input108.Y ,
  output [  0:0] \__mp_input109.A ,
  output [  0:0] \__mp_input109.Y ,
  output [  0:0] \__mp_input11.A ,
  output [  0:0] \__mp_input11.Y ,
  output [  0:0] \__mp_input110.A ,
  output [  0:0] \__mp_input110.Y ,
  output [  0:0] \__mp_input111.A ,
  output [  0:0] \__mp_input111.Y ,
  output [  0:0] \__mp_input112.A ,
  output [  0:0] \__mp_input112.Y ,
  output [  0:0] \__mp_input113.A ,
  output [  0:0] \__mp_input113.Y ,
  output [  0:0] \__mp_input114.A ,
  output [  0:0] \__mp_input114.Y ,
  output [  0:0] \__mp_input115.A ,
  output [  0:0] \__mp_input115.Y ,
  output [  0:0] \__mp_input116.A ,
  output [  0:0] \__mp_input116.Y ,
  output [  0:0] \__mp_input117.A ,
  output [  0:0] \__mp_input117.Y ,
  output [  0:0] \__mp_input118.A ,
  output [  0:0] \__mp_input118.Y ,
  output [  0:0] \__mp_input119.A ,
  output [  0:0] \__mp_input119.Y ,
  output [  0:0] \__mp_input12.A ,
  output [  0:0] \__mp_input12.Y ,
  output [  0:0] \__mp_input120.A ,
  output [  0:0] \__mp_input120.Y ,
  output [  0:0] \__mp_input121.A ,
  output [  0:0] \__mp_input121.Y ,
  output [  0:0] \__mp_input122.A ,
  output [  0:0] \__mp_input122.Y ,
  output [  0:0] \__mp_input123.A ,
  output [  0:0] \__mp_input123.Y ,
  output [  0:0] \__mp_input124.A ,
  output [  0:0] \__mp_input124.Y ,
  output [  0:0] \__mp_input125.A ,
  output [  0:0] \__mp_input125.Y ,
  output [  0:0] \__mp_input126.A ,
  output [  0:0] \__mp_input126.Y ,
  output [  0:0] \__mp_input127.A ,
  output [  0:0] \__mp_input127.Y ,
  output [  0:0] \__mp_input128.A ,
  output [  0:0] \__mp_input128.Y ,
  output [  0:0] \__mp_input129.A ,
  output [  0:0] \__mp_input129.Y ,
  output [  0:0] \__mp_input13.A ,
  output [  0:0] \__mp_input13.Y ,
  output [  0:0] \__mp_input130.A ,
  output [  0:0] \__mp_input130.Y ,
  output [  0:0] \__mp_input131.A ,
  output [  0:0] \__mp_input131.Y ,
  output [  0:0] \__mp_input132.A ,
  output [  0:0] \__mp_input132.Y ,
  output [  0:0] \__mp_input133.A ,
  output [  0:0] \__mp_input133.Y ,
  output [  0:0] \__mp_input134.A ,
  output [  0:0] \__mp_input134.Y ,
  output [  0:0] \__mp_input135.A ,
  output [  0:0] \__mp_input135.Y ,
  output [  0:0] \__mp_input136.A ,
  output [  0:0] \__mp_input136.Y ,
  output [  0:0] \__mp_input137.A ,
  output [  0:0] \__mp_input137.Y ,
  output [  0:0] \__mp_input138.A ,
  output [  0:0] \__mp_input138.Y ,
  output [  0:0] \__mp_input139.A ,
  output [  0:0] \__mp_input139.Y ,
  output [  0:0] \__mp_input14.A ,
  output [  0:0] \__mp_input14.Y ,
  output [  0:0] \__mp_input140.A ,
  output [  0:0] \__mp_input140.Y ,
  output [  0:0] \__mp_input141.A ,
  output [  0:0] \__mp_input141.Y ,
  output [  0:0] \__mp_input142.A ,
  output [  0:0] \__mp_input142.Y ,
  output [  0:0] \__mp_input143.A ,
  output [  0:0] \__mp_input143.Y ,
  output [  0:0] \__mp_input144.A ,
  output [  0:0] \__mp_input144.Y ,
  output [  0:0] \__mp_input145.A ,
  output [  0:0] \__mp_input145.Y ,
  output [  0:0] \__mp_input146.A ,
  output [  0:0] \__mp_input146.Y ,
  output [  0:0] \__mp_input147.A ,
  output [  0:0] \__mp_input147.Y ,
  output [  0:0] \__mp_input148.A ,
  output [  0:0] \__mp_input148.Y ,
  output [  0:0] \__mp_input149.A ,
  output [  0:0] \__mp_input149.Y ,
  output [  0:0] \__mp_input15.A ,
  output [  0:0] \__mp_input15.Y ,
  output [  0:0] \__mp_input150.A ,
  output [  0:0] \__mp_input150.Y ,
  output [  0:0] \__mp_input151.A ,
  output [  0:0] \__mp_input151.Y ,
  output [  0:0] \__mp_input152.A ,
  output [  0:0] \__mp_input152.Y ,
  output [  0:0] \__mp_input153.A ,
  output [  0:0] \__mp_input153.Y ,
  output [  0:0] \__mp_input154.A ,
  output [  0:0] \__mp_input154.Y ,
  output [  0:0] \__mp_input155.A ,
  output [  0:0] \__mp_input155.Y ,
  output [  0:0] \__mp_input156.A ,
  output [  0:0] \__mp_input156.Y ,
  output [  0:0] \__mp_input157.A ,
  output [  0:0] \__mp_input157.Y ,
  output [  0:0] \__mp_input158.A ,
  output [  0:0] \__mp_input158.Y ,
  output [  0:0] \__mp_input159.A ,
  output [  0:0] \__mp_input159.Y ,
  output [  0:0] \__mp_input16.A ,
  output [  0:0] \__mp_input16.Y ,
  output [  0:0] \__mp_input160.A ,
  output [  0:0] \__mp_input160.Y ,
  output [  0:0] \__mp_input161.A ,
  output [  0:0] \__mp_input161.Y ,
  output [  0:0] \__mp_input162.A ,
  output [  0:0] \__mp_input162.Y ,
  output [  0:0] \__mp_input163.A ,
  output [  0:0] \__mp_input163.Y ,
  output [  0:0] \__mp_input164.A ,
  output [  0:0] \__mp_input164.Y ,
  output [  0:0] \__mp_input165.A ,
  output [  0:0] \__mp_input165.Y ,
  output [  0:0] \__mp_input166.A ,
  output [  0:0] \__mp_input166.Y ,
  output [  0:0] \__mp_input167.A ,
  output [  0:0] \__mp_input167.Y ,
  output [  0:0] \__mp_input168.A ,
  output [  0:0] \__mp_input168.Y ,
  output [  0:0] \__mp_input169.A ,
  output [  0:0] \__mp_input169.Y ,
  output [  0:0] \__mp_input17.A ,
  output [  0:0] \__mp_input17.Y ,
  output [  0:0] \__mp_input170.A ,
  output [  0:0] \__mp_input170.Y ,
  output [  0:0] \__mp_input171.A ,
  output [  0:0] \__mp_input171.Y ,
  output [  0:0] \__mp_input172.A ,
  output [  0:0] \__mp_input172.Y ,
  output [  0:0] \__mp_input173.A ,
  output [  0:0] \__mp_input173.Y ,
  output [  0:0] \__mp_input174.A ,
  output [  0:0] \__mp_input174.Y ,
  output [  0:0] \__mp_input175.A ,
  output [  0:0] \__mp_input175.Y ,
  output [  0:0] \__mp_input176.A ,
  output [  0:0] \__mp_input176.Y ,
  output [  0:0] \__mp_input177.A ,
  output [  0:0] \__mp_input177.Y ,
  output [  0:0] \__mp_input178.A ,
  output [  0:0] \__mp_input178.Y ,
  output [  0:0] \__mp_input179.A ,
  output [  0:0] \__mp_input179.Y ,
  output [  0:0] \__mp_input18.A ,
  output [  0:0] \__mp_input18.Y ,
  output [  0:0] \__mp_input180.A ,
  output [  0:0] \__mp_input180.Y ,
  output [  0:0] \__mp_input181.A ,
  output [  0:0] \__mp_input181.Y ,
  output [  0:0] \__mp_input182.A ,
  output [  0:0] \__mp_input182.Y ,
  output [  0:0] \__mp_input183.A ,
  output [  0:0] \__mp_input183.Y ,
  output [  0:0] \__mp_input184.A ,
  output [  0:0] \__mp_input184.Y ,
  output [  0:0] \__mp_input185.A ,
  output [  0:0] \__mp_input185.Y ,
  output [  0:0] \__mp_input186.A ,
  output [  0:0] \__mp_input186.Y ,
  output [  0:0] \__mp_input187.A ,
  output [  0:0] \__mp_input187.Y ,
  output [  0:0] \__mp_input188.A ,
  output [  0:0] \__mp_input188.Y ,
  output [  0:0] \__mp_input189.A ,
  output [  0:0] \__mp_input189.Y ,
  output [  0:0] \__mp_input19.A ,
  output [  0:0] \__mp_input19.Y ,
  output [  0:0] \__mp_input190.A ,
  output [  0:0] \__mp_input190.Y ,
  output [  0:0] \__mp_input191.A ,
  output [  0:0] \__mp_input191.Y ,
  output [  0:0] \__mp_input192.A ,
  output [  0:0] \__mp_input192.Y ,
  output [  0:0] \__mp_input193.A ,
  output [  0:0] \__mp_input193.Y ,
  output [  0:0] \__mp_input194.A ,
  output [  0:0] \__mp_input194.Y ,
  output [  0:0] \__mp_input195.A ,
  output [  0:0] \__mp_input195.Y ,
  output [  0:0] \__mp_input196.A ,
  output [  0:0] \__mp_input196.Y ,
  output [  0:0] \__mp_input197.A ,
  output [  0:0] \__mp_input197.Y ,
  output [  0:0] \__mp_input198.A ,
  output [  0:0] \__mp_input198.Y ,
  output [  0:0] \__mp_input199.A ,
  output [  0:0] \__mp_input199.Y ,
  output [  0:0] \__mp_input2.A ,
  output [  0:0] \__mp_input2.Y ,
  output [  0:0] \__mp_input20.A ,
  output [  0:0] \__mp_input20.Y ,
  output [  0:0] \__mp_input200.A ,
  output [  0:0] \__mp_input200.Y ,
  output [  0:0] \__mp_input201.A ,
  output [  0:0] \__mp_input201.Y ,
  output [  0:0] \__mp_input202.A ,
  output [  0:0] \__mp_input202.Y ,
  output [  0:0] \__mp_input203.A ,
  output [  0:0] \__mp_input203.Y ,
  output [  0:0] \__mp_input204.A ,
  output [  0:0] \__mp_input204.Y ,
  output [  0:0] \__mp_input205.A ,
  output [  0:0] \__mp_input205.Y ,
  output [  0:0] \__mp_input206.A ,
  output [  0:0] \__mp_input206.Y ,
  output [  0:0] \__mp_input207.A ,
  output [  0:0] \__mp_input207.Y ,
  output [  0:0] \__mp_input208.A ,
  output [  0:0] \__mp_input208.Y ,
  output [  0:0] \__mp_input209.A ,
  output [  0:0] \__mp_input209.Y ,
  output [  0:0] \__mp_input21.A ,
  output [  0:0] \__mp_input21.Y ,
  output [  0:0] \__mp_input210.A ,
  output [  0:0] \__mp_input210.Y ,
  output [  0:0] \__mp_input211.A ,
  output [  0:0] \__mp_input211.Y ,
  output [  0:0] \__mp_input212.A ,
  output [  0:0] \__mp_input212.Y ,
  output [  0:0] \__mp_input213.A ,
  output [  0:0] \__mp_input213.Y ,
  output [  0:0] \__mp_input214.A ,
  output [  0:0] \__mp_input214.Y ,
  output [  0:0] \__mp_input215.A ,
  output [  0:0] \__mp_input215.Y ,
  output [  0:0] \__mp_input216.A ,
  output [  0:0] \__mp_input216.Y ,
  output [  0:0] \__mp_input217.A ,
  output [  0:0] \__mp_input217.Y ,
  output [  0:0] \__mp_input218.A ,
  output [  0:0] \__mp_input218.Y ,
  output [  0:0] \__mp_input219.A ,
  output [  0:0] \__mp_input219.Y ,
  output [  0:0] \__mp_input22.A ,
  output [  0:0] \__mp_input22.Y ,
  output [  0:0] \__mp_input220.A ,
  output [  0:0] \__mp_input220.Y ,
  output [  0:0] \__mp_input221.A ,
  output [  0:0] \__mp_input221.Y ,
  output [  0:0] \__mp_input222.A ,
  output [  0:0] \__mp_input222.Y ,
  output [  0:0] \__mp_input223.A ,
  output [  0:0] \__mp_input223.Y ,
  output [  0:0] \__mp_input224.A ,
  output [  0:0] \__mp_input224.Y ,
  output [  0:0] \__mp_input225.A ,
  output [  0:0] \__mp_input225.Y ,
  output [  0:0] \__mp_input226.A ,
  output [  0:0] \__mp_input226.Y ,
  output [  0:0] \__mp_input227.A ,
  output [  0:0] \__mp_input227.Y ,
  output [  0:0] \__mp_input228.A ,
  output [  0:0] \__mp_input228.Y ,
  output [  0:0] \__mp_input229.A ,
  output [  0:0] \__mp_input229.Y ,
  output [  0:0] \__mp_input23.A ,
  output [  0:0] \__mp_input23.Y ,
  output [  0:0] \__mp_input230.A ,
  output [  0:0] \__mp_input230.Y ,
  output [  0:0] \__mp_input231.A ,
  output [  0:0] \__mp_input231.Y ,
  output [  0:0] \__mp_input232.A ,
  output [  0:0] \__mp_input232.Y ,
  output [  0:0] \__mp_input233.A ,
  output [  0:0] \__mp_input233.Y ,
  output [  0:0] \__mp_input234.A ,
  output [  0:0] \__mp_input234.Y ,
  output [  0:0] \__mp_input235.A ,
  output [  0:0] \__mp_input235.Y ,
  output [  0:0] \__mp_input236.A ,
  output [  0:0] \__mp_input236.Y ,
  output [  0:0] \__mp_input237.A ,
  output [  0:0] \__mp_input237.Y ,
  output [  0:0] \__mp_input238.A ,
  output [  0:0] \__mp_input238.Y ,
  output [  0:0] \__mp_input239.A ,
  output [  0:0] \__mp_input239.Y ,
  output [  0:0] \__mp_input24.A ,
  output [  0:0] \__mp_input24.Y ,
  output [  0:0] \__mp_input240.A ,
  output [  0:0] \__mp_input240.Y ,
  output [  0:0] \__mp_input241.A ,
  output [  0:0] \__mp_input241.Y ,
  output [  0:0] \__mp_input242.A ,
  output [  0:0] \__mp_input242.Y ,
  output [  0:0] \__mp_input243.A ,
  output [  0:0] \__mp_input243.Y ,
  output [  0:0] \__mp_input244.A ,
  output [  0:0] \__mp_input244.Y ,
  output [  0:0] \__mp_input245.A ,
  output [  0:0] \__mp_input245.Y ,
  output [  0:0] \__mp_input246.A ,
  output [  0:0] \__mp_input246.Y ,
  output [  0:0] \__mp_input247.A ,
  output [  0:0] \__mp_input247.Y ,
  output [  0:0] \__mp_input248.A ,
  output [  0:0] \__mp_input248.Y ,
  output [  0:0] \__mp_input249.A ,
  output [  0:0] \__mp_input249.Y ,
  output [  0:0] \__mp_input25.A ,
  output [  0:0] \__mp_input25.Y ,
  output [  0:0] \__mp_input250.A ,
  output [  0:0] \__mp_input250.Y ,
  output [  0:0] \__mp_input251.A ,
  output [  0:0] \__mp_input251.Y ,
  output [  0:0] \__mp_input252.A ,
  output [  0:0] \__mp_input252.Y ,
  output [  0:0] \__mp_input253.A ,
  output [  0:0] \__mp_input253.Y ,
  output [  0:0] \__mp_input254.A ,
  output [  0:0] \__mp_input254.Y ,
  output [  0:0] \__mp_input255.A ,
  output [  0:0] \__mp_input255.Y ,
  output [  0:0] \__mp_input256.A ,
  output [  0:0] \__mp_input256.Y ,
  output [  0:0] \__mp_input257.A ,
  output [  0:0] \__mp_input257.Y ,
  output [  0:0] \__mp_input258.A ,
  output [  0:0] \__mp_input258.Y ,
  output [  0:0] \__mp_input26.A ,
  output [  0:0] \__mp_input26.Y ,
  output [  0:0] \__mp_input27.A ,
  output [  0:0] \__mp_input27.Y ,
  output [  0:0] \__mp_input28.A ,
  output [  0:0] \__mp_input28.Y ,
  output [  0:0] \__mp_input29.A ,
  output [  0:0] \__mp_input29.Y ,
  output [  0:0] \__mp_input3.A ,
  output [  0:0] \__mp_input3.Y ,
  output [  0:0] \__mp_input30.A ,
  output [  0:0] \__mp_input30.Y ,
  output [  0:0] \__mp_input31.A ,
  output [  0:0] \__mp_input31.Y ,
  output [  0:0] \__mp_input32.A ,
  output [  0:0] \__mp_input32.Y ,
  output [  0:0] \__mp_input33.A ,
  output [  0:0] \__mp_input33.Y ,
  output [  0:0] \__mp_input34.A ,
  output [  0:0] \__mp_input34.Y ,
  output [  0:0] \__mp_input35.A ,
  output [  0:0] \__mp_input35.Y ,
  output [  0:0] \__mp_input36.A ,
  output [  0:0] \__mp_input36.Y ,
  output [  0:0] \__mp_input37.A ,
  output [  0:0] \__mp_input37.Y ,
  output [  0:0] \__mp_input38.A ,
  output [  0:0] \__mp_input38.Y ,
  output [  0:0] \__mp_input39.A ,
  output [  0:0] \__mp_input39.Y ,
  output [  0:0] \__mp_input4.A ,
  output [  0:0] \__mp_input4.Y ,
  output [  0:0] \__mp_input40.A ,
  output [  0:0] \__mp_input40.Y ,
  output [  0:0] \__mp_input41.A ,
  output [  0:0] \__mp_input41.Y ,
  output [  0:0] \__mp_input42.A ,
  output [  0:0] \__mp_input42.Y ,
  output [  0:0] \__mp_input43.A ,
  output [  0:0] \__mp_input43.Y ,
  output [  0:0] \__mp_input44.A ,
  output [  0:0] \__mp_input44.Y ,
  output [  0:0] \__mp_input45.A ,
  output [  0:0] \__mp_input45.Y ,
  output [  0:0] \__mp_input46.A ,
  output [  0:0] \__mp_input46.Y ,
  output [  0:0] \__mp_input47.A ,
  output [  0:0] \__mp_input47.Y ,
  output [  0:0] \__mp_input48.A ,
  output [  0:0] \__mp_input48.Y ,
  output [  0:0] \__mp_input49.A ,
  output [  0:0] \__mp_input49.Y ,
  output [  0:0] \__mp_input5.A ,
  output [  0:0] \__mp_input5.Y ,
  output [  0:0] \__mp_input50.A ,
  output [  0:0] \__mp_input50.Y ,
  output [  0:0] \__mp_input51.A ,
  output [  0:0] \__mp_input51.Y ,
  output [  0:0] \__mp_input52.A ,
  output [  0:0] \__mp_input52.Y ,
  output [  0:0] \__mp_input53.A ,
  output [  0:0] \__mp_input53.Y ,
  output [  0:0] \__mp_input54.A ,
  output [  0:0] \__mp_input54.Y ,
  output [  0:0] \__mp_input55.A ,
  output [  0:0] \__mp_input55.Y ,
  output [  0:0] \__mp_input56.A ,
  output [  0:0] \__mp_input56.Y ,
  output [  0:0] \__mp_input57.A ,
  output [  0:0] \__mp_input57.Y ,
  output [  0:0] \__mp_input58.A ,
  output [  0:0] \__mp_input58.Y ,
  output [  0:0] \__mp_input59.A ,
  output [  0:0] \__mp_input59.Y ,
  output [  0:0] \__mp_input6.A ,
  output [  0:0] \__mp_input6.Y ,
  output [  0:0] \__mp_input60.A ,
  output [  0:0] \__mp_input60.Y ,
  output [  0:0] \__mp_input61.A ,
  output [  0:0] \__mp_input61.Y ,
  output [  0:0] \__mp_input62.A ,
  output [  0:0] \__mp_input62.Y ,
  output [  0:0] \__mp_input63.A ,
  output [  0:0] \__mp_input63.Y ,
  output [  0:0] \__mp_input64.A ,
  output [  0:0] \__mp_input64.Y ,
  output [  0:0] \__mp_input65.A ,
  output [  0:0] \__mp_input65.Y ,
  output [  0:0] \__mp_input66.A ,
  output [  0:0] \__mp_input66.Y ,
  output [  0:0] \__mp_input67.A ,
  output [  0:0] \__mp_input67.Y ,
  output [  0:0] \__mp_input68.A ,
  output [  0:0] \__mp_input68.Y ,
  output [  0:0] \__mp_input69.A ,
  output [  0:0] \__mp_input69.Y ,
  output [  0:0] \__mp_input7.A ,
  output [  0:0] \__mp_input7.Y ,
  output [  0:0] \__mp_input70.A ,
  output [  0:0] \__mp_input70.Y ,
  output [  0:0] \__mp_input71.A ,
  output [  0:0] \__mp_input71.Y ,
  output [  0:0] \__mp_input72.A ,
  output [  0:0] \__mp_input72.Y ,
  output [  0:0] \__mp_input73.A ,
  output [  0:0] \__mp_input73.Y ,
  output [  0:0] \__mp_input74.A ,
  output [  0:0] \__mp_input74.Y ,
  output [  0:0] \__mp_input75.A ,
  output [  0:0] \__mp_input75.Y ,
  output [  0:0] \__mp_input76.A ,
  output [  0:0] \__mp_input76.Y ,
  output [  0:0] \__mp_input77.A ,
  output [  0:0] \__mp_input77.Y ,
  output [  0:0] \__mp_input78.A ,
  output [  0:0] \__mp_input78.Y ,
  output [  0:0] \__mp_input79.A ,
  output [  0:0] \__mp_input79.Y ,
  output [  0:0] \__mp_input8.A ,
  output [  0:0] \__mp_input8.Y ,
  output [  0:0] \__mp_input80.A ,
  output [  0:0] \__mp_input80.Y ,
  output [  0:0] \__mp_input81.A ,
  output [  0:0] \__mp_input81.Y ,
  output [  0:0] \__mp_input82.A ,
  output [  0:0] \__mp_input82.Y ,
  output [  0:0] \__mp_input83.A ,
  output [  0:0] \__mp_input83.Y ,
  output [  0:0] \__mp_input84.A ,
  output [  0:0] \__mp_input84.Y ,
  output [  0:0] \__mp_input85.A ,
  output [  0:0] \__mp_input85.Y ,
  output [  0:0] \__mp_input86.A ,
  output [  0:0] \__mp_input86.Y ,
  output [  0:0] \__mp_input87.A ,
  output [  0:0] \__mp_input87.Y ,
  output [  0:0] \__mp_input88.A ,
  output [  0:0] \__mp_input88.Y ,
  output [  0:0] \__mp_input89.A ,
  output [  0:0] \__mp_input89.Y ,
  output [  0:0] \__mp_input9.A ,
  output [  0:0] \__mp_input9.Y ,
  output [  0:0] \__mp_input90.A ,
  output [  0:0] \__mp_input90.Y ,
  output [  0:0] \__mp_input91.A ,
  output [  0:0] \__mp_input91.Y ,
  output [  0:0] \__mp_input92.A ,
  output [  0:0] \__mp_input92.Y ,
  output [  0:0] \__mp_input93.A ,
  output [  0:0] \__mp_input93.Y ,
  output [  0:0] \__mp_input94.A ,
  output [  0:0] \__mp_input94.Y ,
  output [  0:0] \__mp_input95.A ,
  output [  0:0] \__mp_input95.Y ,
  output [  0:0] \__mp_input96.A ,
  output [  0:0] \__mp_input96.Y ,
  output [  0:0] \__mp_input97.A ,
  output [  0:0] \__mp_input97.Y ,
  output [  0:0] \__mp_input98.A ,
  output [  0:0] \__mp_input98.Y ,
  output [  0:0] \__mp_input99.A ,
  output [  0:0] \__mp_input99.Y ,
  output [  0:0] \__mp_ld_r$_DFF_P_.CLK ,
  output [  0:0] \__mp_ld_r$_DFF_P_.D ,
  output [  0:0] \__mp_output259.A ,
  output [  0:0] \__mp_output259.Y ,
  output [  0:0] \__mp_output260.A ,
  output [  0:0] \__mp_output260.Y ,
  output [  0:0] \__mp_output261.A ,
  output [  0:0] \__mp_output261.Y ,
  output [  0:0] \__mp_output262.A ,
  output [  0:0] \__mp_output262.Y ,
  output [  0:0] \__mp_output263.A ,
  output [  0:0] \__mp_output263.Y ,
  output [  0:0] \__mp_output264.A ,
  output [  0:0] \__mp_output264.Y ,
  output [  0:0] \__mp_output265.A ,
  output [  0:0] \__mp_output265.Y ,
  output [  0:0] \__mp_output266.A ,
  output [  0:0] \__mp_output266.Y ,
  output [  0:0] \__mp_output267.A ,
  output [  0:0] \__mp_output267.Y ,
  output [  0:0] \__mp_output268.A ,
  output [  0:0] \__mp_output268.Y ,
  output [  0:0] \__mp_output269.A ,
  output [  0:0] \__mp_output269.Y ,
  output [  0:0] \__mp_output270.A ,
  output [  0:0] \__mp_output270.Y ,
  output [  0:0] \__mp_output271.A ,
  output [  0:0] \__mp_output271.Y ,
  output [  0:0] \__mp_output272.A ,
  output [  0:0] \__mp_output272.Y ,
  output [  0:0] \__mp_output273.A ,
  output [  0:0] \__mp_output273.Y ,
  output [  0:0] \__mp_output274.A ,
  output [  0:0] \__mp_output274.Y ,
  output [  0:0] \__mp_output275.A ,
  output [  0:0] \__mp_output275.Y ,
  output [  0:0] \__mp_output276.A ,
  output [  0:0] \__mp_output276.Y ,
  output [  0:0] \__mp_output277.A ,
  output [  0:0] \__mp_output277.Y ,
  output [  0:0] \__mp_output278.A ,
  output [  0:0] \__mp_output278.Y ,
  output [  0:0] \__mp_output279.A ,
  output [  0:0] \__mp_output279.Y ,
  output [  0:0] \__mp_output280.A ,
  output [  0:0] \__mp_output280.Y ,
  output [  0:0] \__mp_output281.A ,
  output [  0:0] \__mp_output281.Y ,
  output [  0:0] \__mp_output282.A ,
  output [  0:0] \__mp_output282.Y ,
  output [  0:0] \__mp_output283.A ,
  output [  0:0] \__mp_output283.Y ,
  output [  0:0] \__mp_output284.A ,
  output [  0:0] \__mp_output284.Y ,
  output [  0:0] \__mp_output285.A ,
  output [  0:0] \__mp_output285.Y ,
  output [  0:0] \__mp_output286.A ,
  output [  0:0] \__mp_output286.Y ,
  output [  0:0] \__mp_output287.A ,
  output [  0:0] \__mp_output287.Y ,
  output [  0:0] \__mp_output288.A ,
  output [  0:0] \__mp_output288.Y ,
  output [  0:0] \__mp_output289.A ,
  output [  0:0] \__mp_output289.Y ,
  output [  0:0] \__mp_output290.A ,
  output [  0:0] \__mp_output290.Y ,
  output [  0:0] \__mp_output291.A ,
  output [  0:0] \__mp_output291.Y ,
  output [  0:0] \__mp_output292.A ,
  output [  0:0] \__mp_output292.Y ,
  output [  0:0] \__mp_output293.A ,
  output [  0:0] \__mp_output293.Y ,
  output [  0:0] \__mp_output294.A ,
  output [  0:0] \__mp_output294.Y ,
  output [  0:0] \__mp_output295.A ,
  output [  0:0] \__mp_output295.Y ,
  output [  0:0] \__mp_output296.A ,
  output [  0:0] \__mp_output296.Y ,
  output [  0:0] \__mp_output297.A ,
  output [  0:0] \__mp_output297.Y ,
  output [  0:0] \__mp_output298.A ,
  output [  0:0] \__mp_output298.Y ,
  output [  0:0] \__mp_output299.A ,
  output [  0:0] \__mp_output299.Y ,
  output [  0:0] \__mp_output300.A ,
  output [  0:0] \__mp_output300.Y ,
  output [  0:0] \__mp_output301.A ,
  output [  0:0] \__mp_output301.Y ,
  output [  0:0] \__mp_output302.A ,
  output [  0:0] \__mp_output302.Y ,
  output [  0:0] \__mp_output303.A ,
  output [  0:0] \__mp_output303.Y ,
  output [  0:0] \__mp_output304.A ,
  output [  0:0] \__mp_output304.Y ,
  output [  0:0] \__mp_output305.A ,
  output [  0:0] \__mp_output305.Y ,
  output [  0:0] \__mp_output306.A ,
  output [  0:0] \__mp_output306.Y ,
  output [  0:0] \__mp_output307.A ,
  output [  0:0] \__mp_output307.Y ,
  output [  0:0] \__mp_output308.A ,
  output [  0:0] \__mp_output308.Y ,
  output [  0:0] \__mp_output309.A ,
  output [  0:0] \__mp_output309.Y ,
  output [  0:0] \__mp_output310.A ,
  output [  0:0] \__mp_output310.Y ,
  output [  0:0] \__mp_output311.A ,
  output [  0:0] \__mp_output311.Y ,
  output [  0:0] \__mp_output312.A ,
  output [  0:0] \__mp_output312.Y ,
  output [  0:0] \__mp_output313.A ,
  output [  0:0] \__mp_output313.Y ,
  output [  0:0] \__mp_output314.A ,
  output [  0:0] \__mp_output314.Y ,
  output [  0:0] \__mp_output315.A ,
  output [  0:0] \__mp_output315.Y ,
  output [  0:0] \__mp_output316.A ,
  output [  0:0] \__mp_output316.Y ,
  output [  0:0] \__mp_output317.A ,
  output [  0:0] \__mp_output317.Y ,
  output [  0:0] \__mp_output318.A ,
  output [  0:0] \__mp_output318.Y ,
  output [  0:0] \__mp_output319.A ,
  output [  0:0] \__mp_output319.Y ,
  output [  0:0] \__mp_output320.A ,
  output [  0:0] \__mp_output320.Y ,
  output [  0:0] \__mp_output321.A ,
  output [  0:0] \__mp_output321.Y ,
  output [  0:0] \__mp_output322.A ,
  output [  0:0] \__mp_output322.Y ,
  output [  0:0] \__mp_output323.A ,
  output [  0:0] \__mp_output323.Y ,
  output [  0:0] \__mp_output324.A ,
  output [  0:0] \__mp_output324.Y ,
  output [  0:0] \__mp_output325.A ,
  output [  0:0] \__mp_output325.Y ,
  output [  0:0] \__mp_output326.A ,
  output [  0:0] \__mp_output326.Y ,
  output [  0:0] \__mp_output327.A ,
  output [  0:0] \__mp_output327.Y ,
  output [  0:0] \__mp_output328.A ,
  output [  0:0] \__mp_output328.Y ,
  output [  0:0] \__mp_output329.A ,
  output [  0:0] \__mp_output329.Y ,
  output [  0:0] \__mp_output330.A ,
  output [  0:0] \__mp_output330.Y ,
  output [  0:0] \__mp_output331.A ,
  output [  0:0] \__mp_output331.Y ,
  output [  0:0] \__mp_output332.A ,
  output [  0:0] \__mp_output332.Y ,
  output [  0:0] \__mp_output333.A ,
  output [  0:0] \__mp_output333.Y ,
  output [  0:0] \__mp_output334.A ,
  output [  0:0] \__mp_output334.Y ,
  output [  0:0] \__mp_output335.A ,
  output [  0:0] \__mp_output335.Y ,
  output [  0:0] \__mp_output336.A ,
  output [  0:0] \__mp_output336.Y ,
  output [  0:0] \__mp_output337.A ,
  output [  0:0] \__mp_output337.Y ,
  output [  0:0] \__mp_output338.A ,
  output [  0:0] \__mp_output338.Y ,
  output [  0:0] \__mp_output339.A ,
  output [  0:0] \__mp_output339.Y ,
  output [  0:0] \__mp_output340.A ,
  output [  0:0] \__mp_output340.Y ,
  output [  0:0] \__mp_output341.A ,
  output [  0:0] \__mp_output341.Y ,
  output [  0:0] \__mp_output342.A ,
  output [  0:0] \__mp_output342.Y ,
  output [  0:0] \__mp_output343.A ,
  output [  0:0] \__mp_output343.Y ,
  output [  0:0] \__mp_output344.A ,
  output [  0:0] \__mp_output344.Y ,
  output [  0:0] \__mp_output345.A ,
  output [  0:0] \__mp_output345.Y ,
  output [  0:0] \__mp_output346.A ,
  output [  0:0] \__mp_output346.Y ,
  output [  0:0] \__mp_output347.A ,
  output [  0:0] \__mp_output347.Y ,
  output [  0:0] \__mp_output348.A ,
  output [  0:0] \__mp_output348.Y ,
  output [  0:0] \__mp_output349.A ,
  output [  0:0] \__mp_output349.Y ,
  output [  0:0] \__mp_output350.A ,
  output [  0:0] \__mp_output350.Y ,
  output [  0:0] \__mp_output351.A ,
  output [  0:0] \__mp_output351.Y ,
  output [  0:0] \__mp_output352.A ,
  output [  0:0] \__mp_output352.Y ,
  output [  0:0] \__mp_output353.A ,
  output [  0:0] \__mp_output353.Y ,
  output [  0:0] \__mp_output354.A ,
  output [  0:0] \__mp_output354.Y ,
  output [  0:0] \__mp_output355.A ,
  output [  0:0] \__mp_output355.Y ,
  output [  0:0] \__mp_output356.A ,
  output [  0:0] \__mp_output356.Y ,
  output [  0:0] \__mp_output357.A ,
  output [  0:0] \__mp_output357.Y ,
  output [  0:0] \__mp_output358.A ,
  output [  0:0] \__mp_output358.Y ,
  output [  0:0] \__mp_output359.A ,
  output [  0:0] \__mp_output359.Y ,
  output [  0:0] \__mp_output360.A ,
  output [  0:0] \__mp_output360.Y ,
  output [  0:0] \__mp_output361.A ,
  output [  0:0] \__mp_output361.Y ,
  output [  0:0] \__mp_output362.A ,
  output [  0:0] \__mp_output362.Y ,
  output [  0:0] \__mp_output363.A ,
  output [  0:0] \__mp_output363.Y ,
  output [  0:0] \__mp_output364.A ,
  output [  0:0] \__mp_output364.Y ,
  output [  0:0] \__mp_output365.A ,
  output [  0:0] \__mp_output365.Y ,
  output [  0:0] \__mp_output366.A ,
  output [  0:0] \__mp_output366.Y ,
  output [  0:0] \__mp_output367.A ,
  output [  0:0] \__mp_output367.Y ,
  output [  0:0] \__mp_output368.A ,
  output [  0:0] \__mp_output368.Y ,
  output [  0:0] \__mp_output369.A ,
  output [  0:0] \__mp_output369.Y ,
  output [  0:0] \__mp_output370.A ,
  output [  0:0] \__mp_output370.Y ,
  output [  0:0] \__mp_output371.A ,
  output [  0:0] \__mp_output371.Y ,
  output [  0:0] \__mp_output372.A ,
  output [  0:0] \__mp_output372.Y ,
  output [  0:0] \__mp_output373.A ,
  output [  0:0] \__mp_output373.Y ,
  output [  0:0] \__mp_output374.A ,
  output [  0:0] \__mp_output374.Y ,
  output [  0:0] \__mp_output375.A ,
  output [  0:0] \__mp_output375.Y ,
  output [  0:0] \__mp_output376.A ,
  output [  0:0] \__mp_output376.Y ,
  output [  0:0] \__mp_output377.A ,
  output [  0:0] \__mp_output377.Y ,
  output [  0:0] \__mp_output378.A ,
  output [  0:0] \__mp_output378.Y ,
  output [  0:0] \__mp_output379.A ,
  output [  0:0] \__mp_output379.Y ,
  output [  0:0] \__mp_output380.A ,
  output [  0:0] \__mp_output380.Y ,
  output [  0:0] \__mp_output381.A ,
  output [  0:0] \__mp_output381.Y ,
  output [  0:0] \__mp_output382.A ,
  output [  0:0] \__mp_output382.Y ,
  output [  0:0] \__mp_output383.A ,
  output [  0:0] \__mp_output383.Y ,
  output [  0:0] \__mp_output384.A ,
  output [  0:0] \__mp_output384.Y ,
  output [  0:0] \__mp_output385.A ,
  output [  0:0] \__mp_output385.Y ,
  output [  0:0] \__mp_output386.A ,
  output [  0:0] \__mp_output386.Y ,
  output [  0:0] \__mp_output387.A ,
  output [  0:0] \__mp_output387.Y ,
  output [  0:0] \__mp_sa00_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_in_r[0]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[100]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[101]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[102]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[103]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[104]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[105]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[106]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[107]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[108]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[109]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[10]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[110]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[111]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[112]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[113]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[114]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[115]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[116]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[117]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[118]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[119]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[11]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[120]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[121]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[122]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[123]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[124]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[125]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[126]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[127]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[12]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[13]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[14]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[15]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[16]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[17]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[18]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[19]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[1]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[20]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[21]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[22]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[23]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[24]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[25]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[26]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[27]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[28]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[29]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[2]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[30]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[31]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[32]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[33]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[34]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[35]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[36]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[37]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[38]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[39]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[3]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[40]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[41]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[42]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[43]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[44]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[45]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[46]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[47]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[48]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[49]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[4]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[50]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[51]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[52]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[53]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[54]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[55]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[56]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[57]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[58]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[59]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[5]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[60]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[61]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[62]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[63]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[64]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[65]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[66]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[67]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[68]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[69]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[6]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[70]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[71]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[72]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[73]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[74]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[75]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[76]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[77]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[78]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[79]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[7]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[80]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[81]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[82]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[83]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[84]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[85]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[86]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[87]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[88]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[89]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[8]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[90]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[91]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[92]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[93]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[94]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[95]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[96]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[97]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[98]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[99]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[9]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK ,
  output [  0:0] \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.u0.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][9]$_DFF_P_.CLK ,
  output [  0:0] \__po_done ,
  output [127:0] \__po_text_out
);
endmodule
module \gate.aes_cipher_top (
  input  [  0:0] \__pi_clk ,
  input  [127:0] \__pi_key ,
  input  [  0:0] \__pi_ld ,
  input  [  0:0] \__pi_rst ,
  input  [127:0] \__pi_text_in ,
  output [  0:0] \__mp_clkbuf_0_clk.A ,
  output [  0:0] \__mp_clkbuf_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_0_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_1_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_2_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.A ,
  output [  0:0] \__mp_clkbuf_2_3_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_0_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_10_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_11_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_12_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_13_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_14_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_15_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_16_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_17_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_18_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_19_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_1_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_20_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_21_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_22_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_23_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_24_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_25_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_26_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_27_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_28_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_29_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_2_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_30_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_31_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_32_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_33_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_3_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_4_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_5_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_6_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_7_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_8_clk.Y ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.A ,
  output [  0:0] \__mp_clkbuf_leaf_9_clk.Y ,
  output [  0:0] \__mp_clkload0.A ,
  output [  0:0] \__mp_clkload0.Y ,
  output [  0:0] \__mp_clkload1.A ,
  output [  0:0] \__mp_clkload10.A ,
  output [  0:0] \__mp_clkload11.A ,
  output [  0:0] \__mp_clkload12.A ,
  output [  0:0] \__mp_clkload13.A ,
  output [  0:0] \__mp_clkload14.A ,
  output [  0:0] \__mp_clkload15.A ,
  output [  0:0] \__mp_clkload16.A ,
  output [  0:0] \__mp_clkload17.A ,
  output [  0:0] \__mp_clkload18.A ,
  output [  0:0] \__mp_clkload18.Y ,
  output [  0:0] \__mp_clkload19.A ,
  output [  0:0] \__mp_clkload2.A ,
  output [  0:0] \__mp_clkload20.A ,
  output [  0:0] \__mp_clkload21.A ,
  output [  0:0] \__mp_clkload22.A ,
  output [  0:0] \__mp_clkload23.A ,
  output [  0:0] \__mp_clkload24.A ,
  output [  0:0] \__mp_clkload25.A ,
  output [  0:0] \__mp_clkload26.A ,
  output [  0:0] \__mp_clkload27.A ,
  output [  0:0] \__mp_clkload28.A ,
  output [  0:0] \__mp_clkload29.A ,
  output [  0:0] \__mp_clkload3.A ,
  output [  0:0] \__mp_clkload30.A ,
  output [  0:0] \__mp_clkload31.A ,
  output [  0:0] \__mp_clkload31.Y ,
  output [  0:0] \__mp_clkload32.A ,
  output [  0:0] \__mp_clkload4.A ,
  output [  0:0] \__mp_clkload5.A ,
  output [  0:0] \__mp_clkload6.A ,
  output [  0:0] \__mp_clkload7.A ,
  output [  0:0] \__mp_clkload8.A ,
  output [  0:0] \__mp_clkload9.A ,
  output [  0:0] \__mp_clknet_0_clk ,
  output [  0:0] \__mp_clknet_2_0_0_clk ,
  output [  0:0] \__mp_clknet_2_1_0_clk ,
  output [  0:0] \__mp_clknet_2_2_0_clk ,
  output [  0:0] \__mp_clknet_2_3_0_clk ,
  output [  0:0] \__mp_clknet_leaf_0_clk ,
  output [  0:0] \__mp_clknet_leaf_10_clk ,
  output [  0:0] \__mp_clknet_leaf_11_clk ,
  output [  0:0] \__mp_clknet_leaf_12_clk ,
  output [  0:0] \__mp_clknet_leaf_13_clk ,
  output [  0:0] \__mp_clknet_leaf_14_clk ,
  output [  0:0] \__mp_clknet_leaf_15_clk ,
  output [  0:0] \__mp_clknet_leaf_16_clk ,
  output [  0:0] \__mp_clknet_leaf_17_clk ,
  output [  0:0] \__mp_clknet_leaf_18_clk ,
  output [  0:0] \__mp_clknet_leaf_19_clk ,
  output [  0:0] \__mp_clknet_leaf_1_clk ,
  output [  0:0] \__mp_clknet_leaf_20_clk ,
  output [  0:0] \__mp_clknet_leaf_21_clk ,
  output [  0:0] \__mp_clknet_leaf_22_clk ,
  output [  0:0] \__mp_clknet_leaf_23_clk ,
  output [  0:0] \__mp_clknet_leaf_24_clk ,
  output [  0:0] \__mp_clknet_leaf_25_clk ,
  output [  0:0] \__mp_clknet_leaf_26_clk ,
  output [  0:0] \__mp_clknet_leaf_27_clk ,
  output [  0:0] \__mp_clknet_leaf_28_clk ,
  output [  0:0] \__mp_clknet_leaf_29_clk ,
  output [  0:0] \__mp_clknet_leaf_2_clk ,
  output [  0:0] \__mp_clknet_leaf_30_clk ,
  output [  0:0] \__mp_clknet_leaf_31_clk ,
  output [  0:0] \__mp_clknet_leaf_32_clk ,
  output [  0:0] \__mp_clknet_leaf_33_clk ,
  output [  0:0] \__mp_clknet_leaf_3_clk ,
  output [  0:0] \__mp_clknet_leaf_4_clk ,
  output [  0:0] \__mp_clknet_leaf_5_clk ,
  output [  0:0] \__mp_clknet_leaf_6_clk ,
  output [  0:0] \__mp_clknet_leaf_7_clk ,
  output [  0:0] \__mp_clknet_leaf_8_clk ,
  output [  0:0] \__mp_clknet_leaf_9_clk ,
  output [  0:0] \__mp_dcnt[0]$_SDFFE_PN0P_.CLK ,
  output [  0:0] \__mp_dcnt[1]$_SDFFE_PN0P_.CLK ,
  output [  0:0] \__mp_dcnt[2]$_SDFFE_PP0P_.CLK ,
  output [  0:0] \__mp_dcnt[3]$_SDFFE_PN0P_.CLK ,
  output [  0:0] \__mp_done$_DFF_P_.CLK ,
  output [  0:0] \__mp_done$_DFF_P_.QN ,
  output [  0:0] \__mp_done$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_input1.A ,
  output [  0:0] \__mp_input1.Y ,
  output [  0:0] \__mp_input10.A ,
  output [  0:0] \__mp_input10.Y ,
  output [  0:0] \__mp_input100.A ,
  output [  0:0] \__mp_input100.Y ,
  output [  0:0] \__mp_input101.A ,
  output [  0:0] \__mp_input101.Y ,
  output [  0:0] \__mp_input102.A ,
  output [  0:0] \__mp_input102.Y ,
  output [  0:0] \__mp_input103.A ,
  output [  0:0] \__mp_input103.Y ,
  output [  0:0] \__mp_input104.A ,
  output [  0:0] \__mp_input104.Y ,
  output [  0:0] \__mp_input105.A ,
  output [  0:0] \__mp_input105.Y ,
  output [  0:0] \__mp_input106.A ,
  output [  0:0] \__mp_input106.Y ,
  output [  0:0] \__mp_input107.A ,
  output [  0:0] \__mp_input107.Y ,
  output [  0:0] \__mp_input108.A ,
  output [  0:0] \__mp_input108.Y ,
  output [  0:0] \__mp_input109.A ,
  output [  0:0] \__mp_input109.Y ,
  output [  0:0] \__mp_input11.A ,
  output [  0:0] \__mp_input11.Y ,
  output [  0:0] \__mp_input110.A ,
  output [  0:0] \__mp_input110.Y ,
  output [  0:0] \__mp_input111.A ,
  output [  0:0] \__mp_input111.Y ,
  output [  0:0] \__mp_input112.A ,
  output [  0:0] \__mp_input112.Y ,
  output [  0:0] \__mp_input113.A ,
  output [  0:0] \__mp_input113.Y ,
  output [  0:0] \__mp_input114.A ,
  output [  0:0] \__mp_input114.Y ,
  output [  0:0] \__mp_input115.A ,
  output [  0:0] \__mp_input115.Y ,
  output [  0:0] \__mp_input116.A ,
  output [  0:0] \__mp_input116.Y ,
  output [  0:0] \__mp_input117.A ,
  output [  0:0] \__mp_input117.Y ,
  output [  0:0] \__mp_input118.A ,
  output [  0:0] \__mp_input118.Y ,
  output [  0:0] \__mp_input119.A ,
  output [  0:0] \__mp_input119.Y ,
  output [  0:0] \__mp_input12.A ,
  output [  0:0] \__mp_input12.Y ,
  output [  0:0] \__mp_input120.A ,
  output [  0:0] \__mp_input120.Y ,
  output [  0:0] \__mp_input121.A ,
  output [  0:0] \__mp_input121.Y ,
  output [  0:0] \__mp_input122.A ,
  output [  0:0] \__mp_input122.Y ,
  output [  0:0] \__mp_input123.A ,
  output [  0:0] \__mp_input123.Y ,
  output [  0:0] \__mp_input124.A ,
  output [  0:0] \__mp_input124.Y ,
  output [  0:0] \__mp_input125.A ,
  output [  0:0] \__mp_input125.Y ,
  output [  0:0] \__mp_input126.A ,
  output [  0:0] \__mp_input126.Y ,
  output [  0:0] \__mp_input127.A ,
  output [  0:0] \__mp_input127.Y ,
  output [  0:0] \__mp_input128.A ,
  output [  0:0] \__mp_input128.Y ,
  output [  0:0] \__mp_input129.A ,
  output [  0:0] \__mp_input129.Y ,
  output [  0:0] \__mp_input13.A ,
  output [  0:0] \__mp_input13.Y ,
  output [  0:0] \__mp_input130.A ,
  output [  0:0] \__mp_input130.Y ,
  output [  0:0] \__mp_input131.A ,
  output [  0:0] \__mp_input131.Y ,
  output [  0:0] \__mp_input132.A ,
  output [  0:0] \__mp_input132.Y ,
  output [  0:0] \__mp_input133.A ,
  output [  0:0] \__mp_input133.Y ,
  output [  0:0] \__mp_input134.A ,
  output [  0:0] \__mp_input134.Y ,
  output [  0:0] \__mp_input135.A ,
  output [  0:0] \__mp_input135.Y ,
  output [  0:0] \__mp_input136.A ,
  output [  0:0] \__mp_input136.Y ,
  output [  0:0] \__mp_input137.A ,
  output [  0:0] \__mp_input137.Y ,
  output [  0:0] \__mp_input138.A ,
  output [  0:0] \__mp_input138.Y ,
  output [  0:0] \__mp_input139.A ,
  output [  0:0] \__mp_input139.Y ,
  output [  0:0] \__mp_input14.A ,
  output [  0:0] \__mp_input14.Y ,
  output [  0:0] \__mp_input140.A ,
  output [  0:0] \__mp_input140.Y ,
  output [  0:0] \__mp_input141.A ,
  output [  0:0] \__mp_input141.Y ,
  output [  0:0] \__mp_input142.A ,
  output [  0:0] \__mp_input142.Y ,
  output [  0:0] \__mp_input143.A ,
  output [  0:0] \__mp_input143.Y ,
  output [  0:0] \__mp_input144.A ,
  output [  0:0] \__mp_input144.Y ,
  output [  0:0] \__mp_input145.A ,
  output [  0:0] \__mp_input145.Y ,
  output [  0:0] \__mp_input146.A ,
  output [  0:0] \__mp_input146.Y ,
  output [  0:0] \__mp_input147.A ,
  output [  0:0] \__mp_input147.Y ,
  output [  0:0] \__mp_input148.A ,
  output [  0:0] \__mp_input148.Y ,
  output [  0:0] \__mp_input149.A ,
  output [  0:0] \__mp_input149.Y ,
  output [  0:0] \__mp_input15.A ,
  output [  0:0] \__mp_input15.Y ,
  output [  0:0] \__mp_input150.A ,
  output [  0:0] \__mp_input150.Y ,
  output [  0:0] \__mp_input151.A ,
  output [  0:0] \__mp_input151.Y ,
  output [  0:0] \__mp_input152.A ,
  output [  0:0] \__mp_input152.Y ,
  output [  0:0] \__mp_input153.A ,
  output [  0:0] \__mp_input153.Y ,
  output [  0:0] \__mp_input154.A ,
  output [  0:0] \__mp_input154.Y ,
  output [  0:0] \__mp_input155.A ,
  output [  0:0] \__mp_input155.Y ,
  output [  0:0] \__mp_input156.A ,
  output [  0:0] \__mp_input156.Y ,
  output [  0:0] \__mp_input157.A ,
  output [  0:0] \__mp_input157.Y ,
  output [  0:0] \__mp_input158.A ,
  output [  0:0] \__mp_input158.Y ,
  output [  0:0] \__mp_input159.A ,
  output [  0:0] \__mp_input159.Y ,
  output [  0:0] \__mp_input16.A ,
  output [  0:0] \__mp_input16.Y ,
  output [  0:0] \__mp_input160.A ,
  output [  0:0] \__mp_input160.Y ,
  output [  0:0] \__mp_input161.A ,
  output [  0:0] \__mp_input161.Y ,
  output [  0:0] \__mp_input162.A ,
  output [  0:0] \__mp_input162.Y ,
  output [  0:0] \__mp_input163.A ,
  output [  0:0] \__mp_input163.Y ,
  output [  0:0] \__mp_input164.A ,
  output [  0:0] \__mp_input164.Y ,
  output [  0:0] \__mp_input165.A ,
  output [  0:0] \__mp_input165.Y ,
  output [  0:0] \__mp_input166.A ,
  output [  0:0] \__mp_input166.Y ,
  output [  0:0] \__mp_input167.A ,
  output [  0:0] \__mp_input167.Y ,
  output [  0:0] \__mp_input168.A ,
  output [  0:0] \__mp_input168.Y ,
  output [  0:0] \__mp_input169.A ,
  output [  0:0] \__mp_input169.Y ,
  output [  0:0] \__mp_input17.A ,
  output [  0:0] \__mp_input17.Y ,
  output [  0:0] \__mp_input170.A ,
  output [  0:0] \__mp_input170.Y ,
  output [  0:0] \__mp_input171.A ,
  output [  0:0] \__mp_input171.Y ,
  output [  0:0] \__mp_input172.A ,
  output [  0:0] \__mp_input172.Y ,
  output [  0:0] \__mp_input173.A ,
  output [  0:0] \__mp_input173.Y ,
  output [  0:0] \__mp_input174.A ,
  output [  0:0] \__mp_input174.Y ,
  output [  0:0] \__mp_input175.A ,
  output [  0:0] \__mp_input175.Y ,
  output [  0:0] \__mp_input176.A ,
  output [  0:0] \__mp_input176.Y ,
  output [  0:0] \__mp_input177.A ,
  output [  0:0] \__mp_input177.Y ,
  output [  0:0] \__mp_input178.A ,
  output [  0:0] \__mp_input178.Y ,
  output [  0:0] \__mp_input179.A ,
  output [  0:0] \__mp_input179.Y ,
  output [  0:0] \__mp_input18.A ,
  output [  0:0] \__mp_input18.Y ,
  output [  0:0] \__mp_input180.A ,
  output [  0:0] \__mp_input180.Y ,
  output [  0:0] \__mp_input181.A ,
  output [  0:0] \__mp_input181.Y ,
  output [  0:0] \__mp_input182.A ,
  output [  0:0] \__mp_input182.Y ,
  output [  0:0] \__mp_input183.A ,
  output [  0:0] \__mp_input183.Y ,
  output [  0:0] \__mp_input184.A ,
  output [  0:0] \__mp_input184.Y ,
  output [  0:0] \__mp_input185.A ,
  output [  0:0] \__mp_input185.Y ,
  output [  0:0] \__mp_input186.A ,
  output [  0:0] \__mp_input186.Y ,
  output [  0:0] \__mp_input187.A ,
  output [  0:0] \__mp_input187.Y ,
  output [  0:0] \__mp_input188.A ,
  output [  0:0] \__mp_input188.Y ,
  output [  0:0] \__mp_input189.A ,
  output [  0:0] \__mp_input189.Y ,
  output [  0:0] \__mp_input19.A ,
  output [  0:0] \__mp_input19.Y ,
  output [  0:0] \__mp_input190.A ,
  output [  0:0] \__mp_input190.Y ,
  output [  0:0] \__mp_input191.A ,
  output [  0:0] \__mp_input191.Y ,
  output [  0:0] \__mp_input192.A ,
  output [  0:0] \__mp_input192.Y ,
  output [  0:0] \__mp_input193.A ,
  output [  0:0] \__mp_input193.Y ,
  output [  0:0] \__mp_input194.A ,
  output [  0:0] \__mp_input194.Y ,
  output [  0:0] \__mp_input195.A ,
  output [  0:0] \__mp_input195.Y ,
  output [  0:0] \__mp_input196.A ,
  output [  0:0] \__mp_input196.Y ,
  output [  0:0] \__mp_input197.A ,
  output [  0:0] \__mp_input197.Y ,
  output [  0:0] \__mp_input198.A ,
  output [  0:0] \__mp_input198.Y ,
  output [  0:0] \__mp_input199.A ,
  output [  0:0] \__mp_input199.Y ,
  output [  0:0] \__mp_input2.A ,
  output [  0:0] \__mp_input2.Y ,
  output [  0:0] \__mp_input20.A ,
  output [  0:0] \__mp_input20.Y ,
  output [  0:0] \__mp_input200.A ,
  output [  0:0] \__mp_input200.Y ,
  output [  0:0] \__mp_input201.A ,
  output [  0:0] \__mp_input201.Y ,
  output [  0:0] \__mp_input202.A ,
  output [  0:0] \__mp_input202.Y ,
  output [  0:0] \__mp_input203.A ,
  output [  0:0] \__mp_input203.Y ,
  output [  0:0] \__mp_input204.A ,
  output [  0:0] \__mp_input204.Y ,
  output [  0:0] \__mp_input205.A ,
  output [  0:0] \__mp_input205.Y ,
  output [  0:0] \__mp_input206.A ,
  output [  0:0] \__mp_input206.Y ,
  output [  0:0] \__mp_input207.A ,
  output [  0:0] \__mp_input207.Y ,
  output [  0:0] \__mp_input208.A ,
  output [  0:0] \__mp_input208.Y ,
  output [  0:0] \__mp_input209.A ,
  output [  0:0] \__mp_input209.Y ,
  output [  0:0] \__mp_input21.A ,
  output [  0:0] \__mp_input21.Y ,
  output [  0:0] \__mp_input210.A ,
  output [  0:0] \__mp_input210.Y ,
  output [  0:0] \__mp_input211.A ,
  output [  0:0] \__mp_input211.Y ,
  output [  0:0] \__mp_input212.A ,
  output [  0:0] \__mp_input212.Y ,
  output [  0:0] \__mp_input213.A ,
  output [  0:0] \__mp_input213.Y ,
  output [  0:0] \__mp_input214.A ,
  output [  0:0] \__mp_input214.Y ,
  output [  0:0] \__mp_input215.A ,
  output [  0:0] \__mp_input215.Y ,
  output [  0:0] \__mp_input216.A ,
  output [  0:0] \__mp_input216.Y ,
  output [  0:0] \__mp_input217.A ,
  output [  0:0] \__mp_input217.Y ,
  output [  0:0] \__mp_input218.A ,
  output [  0:0] \__mp_input218.Y ,
  output [  0:0] \__mp_input219.A ,
  output [  0:0] \__mp_input219.Y ,
  output [  0:0] \__mp_input22.A ,
  output [  0:0] \__mp_input22.Y ,
  output [  0:0] \__mp_input220.A ,
  output [  0:0] \__mp_input220.Y ,
  output [  0:0] \__mp_input221.A ,
  output [  0:0] \__mp_input221.Y ,
  output [  0:0] \__mp_input222.A ,
  output [  0:0] \__mp_input222.Y ,
  output [  0:0] \__mp_input223.A ,
  output [  0:0] \__mp_input223.Y ,
  output [  0:0] \__mp_input224.A ,
  output [  0:0] \__mp_input224.Y ,
  output [  0:0] \__mp_input225.A ,
  output [  0:0] \__mp_input225.Y ,
  output [  0:0] \__mp_input226.A ,
  output [  0:0] \__mp_input226.Y ,
  output [  0:0] \__mp_input227.A ,
  output [  0:0] \__mp_input227.Y ,
  output [  0:0] \__mp_input228.A ,
  output [  0:0] \__mp_input228.Y ,
  output [  0:0] \__mp_input229.A ,
  output [  0:0] \__mp_input229.Y ,
  output [  0:0] \__mp_input23.A ,
  output [  0:0] \__mp_input23.Y ,
  output [  0:0] \__mp_input230.A ,
  output [  0:0] \__mp_input230.Y ,
  output [  0:0] \__mp_input231.A ,
  output [  0:0] \__mp_input231.Y ,
  output [  0:0] \__mp_input232.A ,
  output [  0:0] \__mp_input232.Y ,
  output [  0:0] \__mp_input233.A ,
  output [  0:0] \__mp_input233.Y ,
  output [  0:0] \__mp_input234.A ,
  output [  0:0] \__mp_input234.Y ,
  output [  0:0] \__mp_input235.A ,
  output [  0:0] \__mp_input235.Y ,
  output [  0:0] \__mp_input236.A ,
  output [  0:0] \__mp_input236.Y ,
  output [  0:0] \__mp_input237.A ,
  output [  0:0] \__mp_input237.Y ,
  output [  0:0] \__mp_input238.A ,
  output [  0:0] \__mp_input238.Y ,
  output [  0:0] \__mp_input239.A ,
  output [  0:0] \__mp_input239.Y ,
  output [  0:0] \__mp_input24.A ,
  output [  0:0] \__mp_input24.Y ,
  output [  0:0] \__mp_input240.A ,
  output [  0:0] \__mp_input240.Y ,
  output [  0:0] \__mp_input241.A ,
  output [  0:0] \__mp_input241.Y ,
  output [  0:0] \__mp_input242.A ,
  output [  0:0] \__mp_input242.Y ,
  output [  0:0] \__mp_input243.A ,
  output [  0:0] \__mp_input243.Y ,
  output [  0:0] \__mp_input244.A ,
  output [  0:0] \__mp_input244.Y ,
  output [  0:0] \__mp_input245.A ,
  output [  0:0] \__mp_input245.Y ,
  output [  0:0] \__mp_input246.A ,
  output [  0:0] \__mp_input246.Y ,
  output [  0:0] \__mp_input247.A ,
  output [  0:0] \__mp_input247.Y ,
  output [  0:0] \__mp_input248.A ,
  output [  0:0] \__mp_input248.Y ,
  output [  0:0] \__mp_input249.A ,
  output [  0:0] \__mp_input249.Y ,
  output [  0:0] \__mp_input25.A ,
  output [  0:0] \__mp_input25.Y ,
  output [  0:0] \__mp_input250.A ,
  output [  0:0] \__mp_input250.Y ,
  output [  0:0] \__mp_input251.A ,
  output [  0:0] \__mp_input251.Y ,
  output [  0:0] \__mp_input252.A ,
  output [  0:0] \__mp_input252.Y ,
  output [  0:0] \__mp_input253.A ,
  output [  0:0] \__mp_input253.Y ,
  output [  0:0] \__mp_input254.A ,
  output [  0:0] \__mp_input254.Y ,
  output [  0:0] \__mp_input255.A ,
  output [  0:0] \__mp_input255.Y ,
  output [  0:0] \__mp_input256.A ,
  output [  0:0] \__mp_input256.Y ,
  output [  0:0] \__mp_input257.A ,
  output [  0:0] \__mp_input257.Y ,
  output [  0:0] \__mp_input258.A ,
  output [  0:0] \__mp_input258.Y ,
  output [  0:0] \__mp_input26.A ,
  output [  0:0] \__mp_input26.Y ,
  output [  0:0] \__mp_input27.A ,
  output [  0:0] \__mp_input27.Y ,
  output [  0:0] \__mp_input28.A ,
  output [  0:0] \__mp_input28.Y ,
  output [  0:0] \__mp_input29.A ,
  output [  0:0] \__mp_input29.Y ,
  output [  0:0] \__mp_input3.A ,
  output [  0:0] \__mp_input3.Y ,
  output [  0:0] \__mp_input30.A ,
  output [  0:0] \__mp_input30.Y ,
  output [  0:0] \__mp_input31.A ,
  output [  0:0] \__mp_input31.Y ,
  output [  0:0] \__mp_input32.A ,
  output [  0:0] \__mp_input32.Y ,
  output [  0:0] \__mp_input33.A ,
  output [  0:0] \__mp_input33.Y ,
  output [  0:0] \__mp_input34.A ,
  output [  0:0] \__mp_input34.Y ,
  output [  0:0] \__mp_input35.A ,
  output [  0:0] \__mp_input35.Y ,
  output [  0:0] \__mp_input36.A ,
  output [  0:0] \__mp_input36.Y ,
  output [  0:0] \__mp_input37.A ,
  output [  0:0] \__mp_input37.Y ,
  output [  0:0] \__mp_input38.A ,
  output [  0:0] \__mp_input38.Y ,
  output [  0:0] \__mp_input39.A ,
  output [  0:0] \__mp_input39.Y ,
  output [  0:0] \__mp_input4.A ,
  output [  0:0] \__mp_input4.Y ,
  output [  0:0] \__mp_input40.A ,
  output [  0:0] \__mp_input40.Y ,
  output [  0:0] \__mp_input41.A ,
  output [  0:0] \__mp_input41.Y ,
  output [  0:0] \__mp_input42.A ,
  output [  0:0] \__mp_input42.Y ,
  output [  0:0] \__mp_input43.A ,
  output [  0:0] \__mp_input43.Y ,
  output [  0:0] \__mp_input44.A ,
  output [  0:0] \__mp_input44.Y ,
  output [  0:0] \__mp_input45.A ,
  output [  0:0] \__mp_input45.Y ,
  output [  0:0] \__mp_input46.A ,
  output [  0:0] \__mp_input46.Y ,
  output [  0:0] \__mp_input47.A ,
  output [  0:0] \__mp_input47.Y ,
  output [  0:0] \__mp_input48.A ,
  output [  0:0] \__mp_input48.Y ,
  output [  0:0] \__mp_input49.A ,
  output [  0:0] \__mp_input49.Y ,
  output [  0:0] \__mp_input5.A ,
  output [  0:0] \__mp_input5.Y ,
  output [  0:0] \__mp_input50.A ,
  output [  0:0] \__mp_input50.Y ,
  output [  0:0] \__mp_input51.A ,
  output [  0:0] \__mp_input51.Y ,
  output [  0:0] \__mp_input52.A ,
  output [  0:0] \__mp_input52.Y ,
  output [  0:0] \__mp_input53.A ,
  output [  0:0] \__mp_input53.Y ,
  output [  0:0] \__mp_input54.A ,
  output [  0:0] \__mp_input54.Y ,
  output [  0:0] \__mp_input55.A ,
  output [  0:0] \__mp_input55.Y ,
  output [  0:0] \__mp_input56.A ,
  output [  0:0] \__mp_input56.Y ,
  output [  0:0] \__mp_input57.A ,
  output [  0:0] \__mp_input57.Y ,
  output [  0:0] \__mp_input58.A ,
  output [  0:0] \__mp_input58.Y ,
  output [  0:0] \__mp_input59.A ,
  output [  0:0] \__mp_input59.Y ,
  output [  0:0] \__mp_input6.A ,
  output [  0:0] \__mp_input6.Y ,
  output [  0:0] \__mp_input60.A ,
  output [  0:0] \__mp_input60.Y ,
  output [  0:0] \__mp_input61.A ,
  output [  0:0] \__mp_input61.Y ,
  output [  0:0] \__mp_input62.A ,
  output [  0:0] \__mp_input62.Y ,
  output [  0:0] \__mp_input63.A ,
  output [  0:0] \__mp_input63.Y ,
  output [  0:0] \__mp_input64.A ,
  output [  0:0] \__mp_input64.Y ,
  output [  0:0] \__mp_input65.A ,
  output [  0:0] \__mp_input65.Y ,
  output [  0:0] \__mp_input66.A ,
  output [  0:0] \__mp_input66.Y ,
  output [  0:0] \__mp_input67.A ,
  output [  0:0] \__mp_input67.Y ,
  output [  0:0] \__mp_input68.A ,
  output [  0:0] \__mp_input68.Y ,
  output [  0:0] \__mp_input69.A ,
  output [  0:0] \__mp_input69.Y ,
  output [  0:0] \__mp_input7.A ,
  output [  0:0] \__mp_input7.Y ,
  output [  0:0] \__mp_input70.A ,
  output [  0:0] \__mp_input70.Y ,
  output [  0:0] \__mp_input71.A ,
  output [  0:0] \__mp_input71.Y ,
  output [  0:0] \__mp_input72.A ,
  output [  0:0] \__mp_input72.Y ,
  output [  0:0] \__mp_input73.A ,
  output [  0:0] \__mp_input73.Y ,
  output [  0:0] \__mp_input74.A ,
  output [  0:0] \__mp_input74.Y ,
  output [  0:0] \__mp_input75.A ,
  output [  0:0] \__mp_input75.Y ,
  output [  0:0] \__mp_input76.A ,
  output [  0:0] \__mp_input76.Y ,
  output [  0:0] \__mp_input77.A ,
  output [  0:0] \__mp_input77.Y ,
  output [  0:0] \__mp_input78.A ,
  output [  0:0] \__mp_input78.Y ,
  output [  0:0] \__mp_input79.A ,
  output [  0:0] \__mp_input79.Y ,
  output [  0:0] \__mp_input8.A ,
  output [  0:0] \__mp_input8.Y ,
  output [  0:0] \__mp_input80.A ,
  output [  0:0] \__mp_input80.Y ,
  output [  0:0] \__mp_input81.A ,
  output [  0:0] \__mp_input81.Y ,
  output [  0:0] \__mp_input82.A ,
  output [  0:0] \__mp_input82.Y ,
  output [  0:0] \__mp_input83.A ,
  output [  0:0] \__mp_input83.Y ,
  output [  0:0] \__mp_input84.A ,
  output [  0:0] \__mp_input84.Y ,
  output [  0:0] \__mp_input85.A ,
  output [  0:0] \__mp_input85.Y ,
  output [  0:0] \__mp_input86.A ,
  output [  0:0] \__mp_input86.Y ,
  output [  0:0] \__mp_input87.A ,
  output [  0:0] \__mp_input87.Y ,
  output [  0:0] \__mp_input88.A ,
  output [  0:0] \__mp_input88.Y ,
  output [  0:0] \__mp_input89.A ,
  output [  0:0] \__mp_input89.Y ,
  output [  0:0] \__mp_input9.A ,
  output [  0:0] \__mp_input9.Y ,
  output [  0:0] \__mp_input90.A ,
  output [  0:0] \__mp_input90.Y ,
  output [  0:0] \__mp_input91.A ,
  output [  0:0] \__mp_input91.Y ,
  output [  0:0] \__mp_input92.A ,
  output [  0:0] \__mp_input92.Y ,
  output [  0:0] \__mp_input93.A ,
  output [  0:0] \__mp_input93.Y ,
  output [  0:0] \__mp_input94.A ,
  output [  0:0] \__mp_input94.Y ,
  output [  0:0] \__mp_input95.A ,
  output [  0:0] \__mp_input95.Y ,
  output [  0:0] \__mp_input96.A ,
  output [  0:0] \__mp_input96.Y ,
  output [  0:0] \__mp_input97.A ,
  output [  0:0] \__mp_input97.Y ,
  output [  0:0] \__mp_input98.A ,
  output [  0:0] \__mp_input98.Y ,
  output [  0:0] \__mp_input99.A ,
  output [  0:0] \__mp_input99.Y ,
  output [  0:0] \__mp_ld_r$_DFF_P_.CLK ,
  output [  0:0] \__mp_ld_r$_DFF_P_.D ,
  output [  0:0] \__mp_output259.A ,
  output [  0:0] \__mp_output259.Y ,
  output [  0:0] \__mp_output260.A ,
  output [  0:0] \__mp_output260.Y ,
  output [  0:0] \__mp_output261.A ,
  output [  0:0] \__mp_output261.Y ,
  output [  0:0] \__mp_output262.A ,
  output [  0:0] \__mp_output262.Y ,
  output [  0:0] \__mp_output263.A ,
  output [  0:0] \__mp_output263.Y ,
  output [  0:0] \__mp_output264.A ,
  output [  0:0] \__mp_output264.Y ,
  output [  0:0] \__mp_output265.A ,
  output [  0:0] \__mp_output265.Y ,
  output [  0:0] \__mp_output266.A ,
  output [  0:0] \__mp_output266.Y ,
  output [  0:0] \__mp_output267.A ,
  output [  0:0] \__mp_output267.Y ,
  output [  0:0] \__mp_output268.A ,
  output [  0:0] \__mp_output268.Y ,
  output [  0:0] \__mp_output269.A ,
  output [  0:0] \__mp_output269.Y ,
  output [  0:0] \__mp_output270.A ,
  output [  0:0] \__mp_output270.Y ,
  output [  0:0] \__mp_output271.A ,
  output [  0:0] \__mp_output271.Y ,
  output [  0:0] \__mp_output272.A ,
  output [  0:0] \__mp_output272.Y ,
  output [  0:0] \__mp_output273.A ,
  output [  0:0] \__mp_output273.Y ,
  output [  0:0] \__mp_output274.A ,
  output [  0:0] \__mp_output274.Y ,
  output [  0:0] \__mp_output275.A ,
  output [  0:0] \__mp_output275.Y ,
  output [  0:0] \__mp_output276.A ,
  output [  0:0] \__mp_output276.Y ,
  output [  0:0] \__mp_output277.A ,
  output [  0:0] \__mp_output277.Y ,
  output [  0:0] \__mp_output278.A ,
  output [  0:0] \__mp_output278.Y ,
  output [  0:0] \__mp_output279.A ,
  output [  0:0] \__mp_output279.Y ,
  output [  0:0] \__mp_output280.A ,
  output [  0:0] \__mp_output280.Y ,
  output [  0:0] \__mp_output281.A ,
  output [  0:0] \__mp_output281.Y ,
  output [  0:0] \__mp_output282.A ,
  output [  0:0] \__mp_output282.Y ,
  output [  0:0] \__mp_output283.A ,
  output [  0:0] \__mp_output283.Y ,
  output [  0:0] \__mp_output284.A ,
  output [  0:0] \__mp_output284.Y ,
  output [  0:0] \__mp_output285.A ,
  output [  0:0] \__mp_output285.Y ,
  output [  0:0] \__mp_output286.A ,
  output [  0:0] \__mp_output286.Y ,
  output [  0:0] \__mp_output287.A ,
  output [  0:0] \__mp_output287.Y ,
  output [  0:0] \__mp_output288.A ,
  output [  0:0] \__mp_output288.Y ,
  output [  0:0] \__mp_output289.A ,
  output [  0:0] \__mp_output289.Y ,
  output [  0:0] \__mp_output290.A ,
  output [  0:0] \__mp_output290.Y ,
  output [  0:0] \__mp_output291.A ,
  output [  0:0] \__mp_output291.Y ,
  output [  0:0] \__mp_output292.A ,
  output [  0:0] \__mp_output292.Y ,
  output [  0:0] \__mp_output293.A ,
  output [  0:0] \__mp_output293.Y ,
  output [  0:0] \__mp_output294.A ,
  output [  0:0] \__mp_output294.Y ,
  output [  0:0] \__mp_output295.A ,
  output [  0:0] \__mp_output295.Y ,
  output [  0:0] \__mp_output296.A ,
  output [  0:0] \__mp_output296.Y ,
  output [  0:0] \__mp_output297.A ,
  output [  0:0] \__mp_output297.Y ,
  output [  0:0] \__mp_output298.A ,
  output [  0:0] \__mp_output298.Y ,
  output [  0:0] \__mp_output299.A ,
  output [  0:0] \__mp_output299.Y ,
  output [  0:0] \__mp_output300.A ,
  output [  0:0] \__mp_output300.Y ,
  output [  0:0] \__mp_output301.A ,
  output [  0:0] \__mp_output301.Y ,
  output [  0:0] \__mp_output302.A ,
  output [  0:0] \__mp_output302.Y ,
  output [  0:0] \__mp_output303.A ,
  output [  0:0] \__mp_output303.Y ,
  output [  0:0] \__mp_output304.A ,
  output [  0:0] \__mp_output304.Y ,
  output [  0:0] \__mp_output305.A ,
  output [  0:0] \__mp_output305.Y ,
  output [  0:0] \__mp_output306.A ,
  output [  0:0] \__mp_output306.Y ,
  output [  0:0] \__mp_output307.A ,
  output [  0:0] \__mp_output307.Y ,
  output [  0:0] \__mp_output308.A ,
  output [  0:0] \__mp_output308.Y ,
  output [  0:0] \__mp_output309.A ,
  output [  0:0] \__mp_output309.Y ,
  output [  0:0] \__mp_output310.A ,
  output [  0:0] \__mp_output310.Y ,
  output [  0:0] \__mp_output311.A ,
  output [  0:0] \__mp_output311.Y ,
  output [  0:0] \__mp_output312.A ,
  output [  0:0] \__mp_output312.Y ,
  output [  0:0] \__mp_output313.A ,
  output [  0:0] \__mp_output313.Y ,
  output [  0:0] \__mp_output314.A ,
  output [  0:0] \__mp_output314.Y ,
  output [  0:0] \__mp_output315.A ,
  output [  0:0] \__mp_output315.Y ,
  output [  0:0] \__mp_output316.A ,
  output [  0:0] \__mp_output316.Y ,
  output [  0:0] \__mp_output317.A ,
  output [  0:0] \__mp_output317.Y ,
  output [  0:0] \__mp_output318.A ,
  output [  0:0] \__mp_output318.Y ,
  output [  0:0] \__mp_output319.A ,
  output [  0:0] \__mp_output319.Y ,
  output [  0:0] \__mp_output320.A ,
  output [  0:0] \__mp_output320.Y ,
  output [  0:0] \__mp_output321.A ,
  output [  0:0] \__mp_output321.Y ,
  output [  0:0] \__mp_output322.A ,
  output [  0:0] \__mp_output322.Y ,
  output [  0:0] \__mp_output323.A ,
  output [  0:0] \__mp_output323.Y ,
  output [  0:0] \__mp_output324.A ,
  output [  0:0] \__mp_output324.Y ,
  output [  0:0] \__mp_output325.A ,
  output [  0:0] \__mp_output325.Y ,
  output [  0:0] \__mp_output326.A ,
  output [  0:0] \__mp_output326.Y ,
  output [  0:0] \__mp_output327.A ,
  output [  0:0] \__mp_output327.Y ,
  output [  0:0] \__mp_output328.A ,
  output [  0:0] \__mp_output328.Y ,
  output [  0:0] \__mp_output329.A ,
  output [  0:0] \__mp_output329.Y ,
  output [  0:0] \__mp_output330.A ,
  output [  0:0] \__mp_output330.Y ,
  output [  0:0] \__mp_output331.A ,
  output [  0:0] \__mp_output331.Y ,
  output [  0:0] \__mp_output332.A ,
  output [  0:0] \__mp_output332.Y ,
  output [  0:0] \__mp_output333.A ,
  output [  0:0] \__mp_output333.Y ,
  output [  0:0] \__mp_output334.A ,
  output [  0:0] \__mp_output334.Y ,
  output [  0:0] \__mp_output335.A ,
  output [  0:0] \__mp_output335.Y ,
  output [  0:0] \__mp_output336.A ,
  output [  0:0] \__mp_output336.Y ,
  output [  0:0] \__mp_output337.A ,
  output [  0:0] \__mp_output337.Y ,
  output [  0:0] \__mp_output338.A ,
  output [  0:0] \__mp_output338.Y ,
  output [  0:0] \__mp_output339.A ,
  output [  0:0] \__mp_output339.Y ,
  output [  0:0] \__mp_output340.A ,
  output [  0:0] \__mp_output340.Y ,
  output [  0:0] \__mp_output341.A ,
  output [  0:0] \__mp_output341.Y ,
  output [  0:0] \__mp_output342.A ,
  output [  0:0] \__mp_output342.Y ,
  output [  0:0] \__mp_output343.A ,
  output [  0:0] \__mp_output343.Y ,
  output [  0:0] \__mp_output344.A ,
  output [  0:0] \__mp_output344.Y ,
  output [  0:0] \__mp_output345.A ,
  output [  0:0] \__mp_output345.Y ,
  output [  0:0] \__mp_output346.A ,
  output [  0:0] \__mp_output346.Y ,
  output [  0:0] \__mp_output347.A ,
  output [  0:0] \__mp_output347.Y ,
  output [  0:0] \__mp_output348.A ,
  output [  0:0] \__mp_output348.Y ,
  output [  0:0] \__mp_output349.A ,
  output [  0:0] \__mp_output349.Y ,
  output [  0:0] \__mp_output350.A ,
  output [  0:0] \__mp_output350.Y ,
  output [  0:0] \__mp_output351.A ,
  output [  0:0] \__mp_output351.Y ,
  output [  0:0] \__mp_output352.A ,
  output [  0:0] \__mp_output352.Y ,
  output [  0:0] \__mp_output353.A ,
  output [  0:0] \__mp_output353.Y ,
  output [  0:0] \__mp_output354.A ,
  output [  0:0] \__mp_output354.Y ,
  output [  0:0] \__mp_output355.A ,
  output [  0:0] \__mp_output355.Y ,
  output [  0:0] \__mp_output356.A ,
  output [  0:0] \__mp_output356.Y ,
  output [  0:0] \__mp_output357.A ,
  output [  0:0] \__mp_output357.Y ,
  output [  0:0] \__mp_output358.A ,
  output [  0:0] \__mp_output358.Y ,
  output [  0:0] \__mp_output359.A ,
  output [  0:0] \__mp_output359.Y ,
  output [  0:0] \__mp_output360.A ,
  output [  0:0] \__mp_output360.Y ,
  output [  0:0] \__mp_output361.A ,
  output [  0:0] \__mp_output361.Y ,
  output [  0:0] \__mp_output362.A ,
  output [  0:0] \__mp_output362.Y ,
  output [  0:0] \__mp_output363.A ,
  output [  0:0] \__mp_output363.Y ,
  output [  0:0] \__mp_output364.A ,
  output [  0:0] \__mp_output364.Y ,
  output [  0:0] \__mp_output365.A ,
  output [  0:0] \__mp_output365.Y ,
  output [  0:0] \__mp_output366.A ,
  output [  0:0] \__mp_output366.Y ,
  output [  0:0] \__mp_output367.A ,
  output [  0:0] \__mp_output367.Y ,
  output [  0:0] \__mp_output368.A ,
  output [  0:0] \__mp_output368.Y ,
  output [  0:0] \__mp_output369.A ,
  output [  0:0] \__mp_output369.Y ,
  output [  0:0] \__mp_output370.A ,
  output [  0:0] \__mp_output370.Y ,
  output [  0:0] \__mp_output371.A ,
  output [  0:0] \__mp_output371.Y ,
  output [  0:0] \__mp_output372.A ,
  output [  0:0] \__mp_output372.Y ,
  output [  0:0] \__mp_output373.A ,
  output [  0:0] \__mp_output373.Y ,
  output [  0:0] \__mp_output374.A ,
  output [  0:0] \__mp_output374.Y ,
  output [  0:0] \__mp_output375.A ,
  output [  0:0] \__mp_output375.Y ,
  output [  0:0] \__mp_output376.A ,
  output [  0:0] \__mp_output376.Y ,
  output [  0:0] \__mp_output377.A ,
  output [  0:0] \__mp_output377.Y ,
  output [  0:0] \__mp_output378.A ,
  output [  0:0] \__mp_output378.Y ,
  output [  0:0] \__mp_output379.A ,
  output [  0:0] \__mp_output379.Y ,
  output [  0:0] \__mp_output380.A ,
  output [  0:0] \__mp_output380.Y ,
  output [  0:0] \__mp_output381.A ,
  output [  0:0] \__mp_output381.Y ,
  output [  0:0] \__mp_output382.A ,
  output [  0:0] \__mp_output382.Y ,
  output [  0:0] \__mp_output383.A ,
  output [  0:0] \__mp_output383.Y ,
  output [  0:0] \__mp_output384.A ,
  output [  0:0] \__mp_output384.Y ,
  output [  0:0] \__mp_output385.A ,
  output [  0:0] \__mp_output385.Y ,
  output [  0:0] \__mp_output386.A ,
  output [  0:0] \__mp_output386.Y ,
  output [  0:0] \__mp_output387.A ,
  output [  0:0] \__mp_output387.Y ,
  output [  0:0] \__mp_sa00_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa00_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa01_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa02_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa03_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa10_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa11_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa12_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa13_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa20_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa21_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa22_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa23_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa30_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa31_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa32_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_sa33_sr[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_in_r[0]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[100]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[101]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[102]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[103]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[104]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[105]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[106]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[107]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[108]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[109]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[10]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[110]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[111]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[112]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[113]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[114]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[115]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[116]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[117]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[118]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[119]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[11]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[120]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[121]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[122]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[123]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[124]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[125]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[126]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[127]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[12]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[13]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[14]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[15]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[16]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[17]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[18]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[19]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[1]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[20]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[21]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[22]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[23]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[24]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[25]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[26]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[27]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[28]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[29]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[2]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[30]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[31]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[32]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[33]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[34]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[35]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[36]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[37]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[38]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[39]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[3]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[40]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[41]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[42]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[43]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[44]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[45]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[46]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[47]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[48]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[49]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[4]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[50]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[51]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[52]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[53]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[54]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[55]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[56]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[57]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[58]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[59]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[5]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[60]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[61]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[62]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[63]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[64]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[65]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[66]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[67]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[68]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[69]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[6]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[70]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[71]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[72]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[73]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[74]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[75]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[76]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[77]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[78]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[79]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[7]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[80]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[81]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[82]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[83]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[84]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[85]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[86]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[87]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[88]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[89]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[8]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[90]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[91]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[92]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[93]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[94]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[95]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[96]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[97]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[98]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[99]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_in_r[9]$_DFFE_PP_.CLK ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[0]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[100]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[101]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[102]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[103]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[104]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[105]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[106]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[107]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[108]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[109]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[10]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[110]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[111]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[112]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[113]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[114]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[115]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[116]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[117]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[118]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[119]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[11]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[120]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[121]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[122]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[123]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[124]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[125]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[126]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[127]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[12]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[13]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[14]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[15]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[16]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[17]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[18]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[19]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[1]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[20]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[21]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[22]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[23]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[24]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[25]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[26]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[27]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[28]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[29]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[2]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[30]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[31]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[32]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[33]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[34]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[35]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[36]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[37]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[38]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[39]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[3]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[40]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[41]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[42]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[43]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[44]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[45]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[46]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[47]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[48]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[49]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[4]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[50]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[51]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[52]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[53]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[54]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[55]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[56]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[57]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[58]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[59]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[5]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[60]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[61]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[62]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[63]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[64]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[65]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[66]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[67]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[68]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[69]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[6]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[70]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[71]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[72]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[73]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[74]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[75]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[76]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[77]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[78]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[79]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[7]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[80]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[81]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[82]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[83]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[84]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[85]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[86]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[87]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[88]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[89]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[8]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[90]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[91]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[92]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[93]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[94]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[95]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[96]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[97]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[98]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[99]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.QN ,
  output [  0:0] \__mp_text_out[9]$_DFF_P_.int_fwire_IQN ,
  output [  0:0] \__mp_u0.r0.out[24]$_SDFF_PP1_.CLK ,
  output [  0:0] \__mp_u0.r0.out[25]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[26]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[27]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[28]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[29]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[30]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.out[31]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[0]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[1]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[2]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.r0.rcnt[3]$_SDFF_PP0_.CLK ,
  output [  0:0] \__mp_u0.u0.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u0.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u1.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u2.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.u3.d[7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[0][9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[1][9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[2][9]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][0]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][10]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][11]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][12]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][13]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][14]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][15]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][16]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][17]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][18]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][19]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][1]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][20]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][21]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][22]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][23]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][24]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][25]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][26]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][27]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][28]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][29]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][2]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][30]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][31]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][3]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][4]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][5]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][6]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][7]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][8]$_DFF_P_.CLK ,
  output [  0:0] \__mp_u0.w[3][9]$_DFF_P_.CLK ,
  output [  0:0] \__po_done ,
  output [127:0] \__po_text_out
);
endmodule
